

package model_weights;


logic signed [31:0] VT_0 [37][37] ='{
{32'h80000800 , 32'h00000070 , 32'hFFFFFFB3 , 32'h0000004A , 32'h00000006 , 32'hFFFFFFFA , 32'h00000019 , 32'hFFFFFFF4 , 32'h00000017 , 32'h00000007 , 32'hFFFFFFFF , 32'hFFFFFFFB , 32'h00000005 , 32'h00000000 , 32'hFFFFFFFD , 32'h00000004 , 32'hFFFFFFFF , 32'h00000002 , 32'h00000005 , 32'hFFFFFFF4 , 32'h00000000 , 32'hFFFFFFFB , 32'hFFFFFFFE , 32'h00000000 , 32'hFFFFFFFD , 32'h0000000A , 32'h00000003 , 32'hFFFFFFF3 , 32'h00000001 , 32'hFFFFFFF9 , 32'h00000005 , 32'h00000000 , 32'h00000005 , 32'h00000000 , 32'hFFFFFFFC , 32'h00000002 , 32'h00000000} , 
{32'h00000070 , 32'h7FFFF800 , 32'hFFFFFFF0 , 32'h0000000A , 32'h00000047 , 32'h00000029 , 32'h0000001B , 32'h00000005 , 32'hFFFFFFF0 , 32'h00000000 , 32'hFFFFFFFB , 32'hFFFFFFEC , 32'h00000000 , 32'h00000007 , 32'h00000009 , 32'h0000000A , 32'hFFFFFFFE , 32'h00000003 , 32'h00000009 , 32'h00000009 , 32'hFFFFFFFB , 32'h00000001 , 32'hFFFFFFFA , 32'hFFFFFFFE , 32'hFFFFFFFF , 32'hFFFFFFF6 , 32'hFFFFFFFC , 32'h00000000 , 32'h00000000 , 32'hFFFFFFFF , 32'h00000000 , 32'h00000005 , 32'hFFFFFFF9 , 32'hFFFFFFF3 , 32'hFFFFFFF8 , 32'h00000007 , 32'hFFFFFFFD} , 
{32'hFFFFFFB3 , 32'h0000000E , 32'h7FFFF800 , 32'h00000085 , 32'hFFFFFF88 , 32'h0000004F , 32'hFFFFFFF6 , 32'h0000000C , 32'hFFFFFFF9 , 32'h0000000A , 32'hFFFFFFEC , 32'h0000000B , 32'hFFFFFFF8 , 32'hFFFFFFFB , 32'h00000009 , 32'h00000012 , 32'h00000010 , 32'hFFFFFFEB , 32'hFFFFFFF0 , 32'hFFFFFFFD , 32'hFFFFFFF9 , 32'h00000003 , 32'h00000000 , 32'h00000000 , 32'h00000005 , 32'hFFFFFFF4 , 32'hFFFFFFF3 , 32'hFFFFFFFE , 32'h00000002 , 32'hFFFFFFF7 , 32'hFFFFFFFF , 32'h00000004 , 32'h00000008 , 32'hFFFFFFFD , 32'hFFFFFFFE , 32'hFFFFFFFC , 32'hFFFFFFFD} , 
{32'h0000004A , 32'hFFFFFFF4 , 32'hFFFFFF79 , 32'h7FFFF800 , 32'h000000B7 , 32'hFFFFFF76 , 32'hFFFFFFA3 , 32'hFFFFFFFF , 32'hFFFFFFF1 , 32'h0000001E , 32'h00000009 , 32'hFFFFFFEF , 32'h0000000A , 32'h00000005 , 32'hFFFFFFFB , 32'hFFFFFFE4 , 32'hFFFFFFFC , 32'hFFFFFFF4 , 32'hFFFFFFFD , 32'hFFFFFFFF , 32'h00000013 , 32'h00000003 , 32'h00000005 , 32'hFFFFFFF5 , 32'hFFFFFFF6 , 32'h00000004 , 32'h0000000A , 32'h00000004 , 32'h00000008 , 32'hFFFFFFFB , 32'h0000000B , 32'hFFFFFFFE , 32'h00000000 , 32'hFFFFFFFC , 32'hFFFFFFFB , 32'h00000000 , 32'hFFFFFFFC} , 
{32'hFFFFFFF8 , 32'h00000047 , 32'hFFFFFF88 , 32'h000000B7 , 32'h80000800 , 32'hFFFFFDDE , 32'hFFFFFFF7 , 32'hFFFFFFF9 , 32'h0000000A , 32'hFFFFFFE0 , 32'hFFFFFFE5 , 32'hFFFFFFE1 , 32'h00000000 , 32'h00000001 , 32'h00000001 , 32'hFFFFFFF0 , 32'h0000000C , 32'hFFFFFFFF , 32'hFFFFFFF7 , 32'hFFFFFFFD , 32'h00000002 , 32'hFFFFFFFA , 32'hFFFFFFFB , 32'hFFFFFFFD , 32'hFFFFFFF7 , 32'hFFFFFFFD , 32'h00000000 , 32'hFFFFFFFB , 32'hFFFFFFF9 , 32'h00000004 , 32'h00000000 , 32'hFFFFFFFE , 32'hFFFFFFFB , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'hFFFFFFF7} , 
{32'h00000004 , 32'h00000029 , 32'h0000004F , 32'hFFFFFF76 , 32'h00000220 , 32'h80000800 , 32'h0000000F , 32'hFFFFFFEC , 32'hFFFFFFF7 , 32'h00000006 , 32'hFFFFFFC8 , 32'hFFFFFFF1 , 32'hFFFFFFFD , 32'hFFFFFFF0 , 32'h00000009 , 32'h0000001F , 32'h0000000E , 32'hFFFFFFFE , 32'h00000006 , 32'h00000000 , 32'hFFFFFFFE , 32'hFFFFFFFB , 32'hFFFFFFFE , 32'h00000002 , 32'hFFFFFFFE , 32'hFFFFFFFA , 32'hFFFFFFFF , 32'h00000004 , 32'h00000001 , 32'hFFFFFFFB , 32'hFFFFFFFA , 32'hFFFFFFFF , 32'h00000000 , 32'h00000008 , 32'h00000003 , 32'h00000000 , 32'h00000001} , 
{32'hFFFFFFE5 , 32'h0000001B , 32'hFFFFFFF6 , 32'hFFFFFFA3 , 32'h00000007 , 32'hFFFFFFEF , 32'h80000800 , 32'h00000024 , 32'hFFFFFFEE , 32'h00000003 , 32'h00000000 , 32'h00000004 , 32'h00000000 , 32'hFFFFFFDD , 32'hFFFFFFE3 , 32'h00000003 , 32'hFFFFFFF1 , 32'h00000018 , 32'hFFFFFFFC , 32'hFFFFFFFB , 32'h00000006 , 32'hFFFFFFF8 , 32'hFFFFFFFD , 32'h00000006 , 32'h00000007 , 32'hFFFFFFFB , 32'hFFFFFFF7 , 32'h00000004 , 32'h0000000F , 32'h00000004 , 32'hFFFFFFF7 , 32'h00000000 , 32'hFFFFFFFE , 32'h00000002 , 32'hFFFFFFF3 , 32'h00000001 , 32'hFFFFFFFA} , 
{32'h0000000A , 32'h00000005 , 32'h0000000C , 32'hFFFFFFFF , 32'h00000005 , 32'h00000012 , 32'hFFFFFFDA , 32'h80000800 , 32'h00000015 , 32'h00000025 , 32'hFFFFFFC3 , 32'hFFFFFFF5 , 32'h00000014 , 32'hFFFFFFEF , 32'hFFFFFFD9 , 32'hFFFFFFF8 , 32'hFFFFFFEB , 32'h0000000D , 32'h00000004 , 32'hFFFFFFE6 , 32'hFFFFFFF1 , 32'hFFFFFFEE , 32'hFFFFFFF7 , 32'hFFFFFFEF , 32'h00000002 , 32'h00000016 , 32'hFFFFFFE7 , 32'h00000002 , 32'h00000008 , 32'h00000000 , 32'hFFFFFFFA , 32'hFFFFFFFB , 32'h00000004 , 32'h00000001 , 32'hFFFFFFF5 , 32'h0000000A , 32'h00000004} , 
{32'hFFFFFFE7 , 32'hFFFFFFF0 , 32'hFFFFFFF9 , 32'hFFFFFFF1 , 32'hFFFFFFF4 , 32'h00000007 , 32'h00000010 , 32'hFFFFFFE9 , 32'h80000800 , 32'h0000009A , 32'h00000090 , 32'h0000001E , 32'hFFFFFFF1 , 32'hFFFFFFEE , 32'h00000008 , 32'hFFFFFFE7 , 32'h00000014 , 32'hFFFFFFF7 , 32'h00000019 , 32'h0000000F , 32'h0000000A , 32'hFFFFFFFD , 32'hFFFFFFFB , 32'h00000015 , 32'h0000000B , 32'hFFFFFFFF , 32'h00000016 , 32'h0000000F , 32'h0000000C , 32'hFFFFFFF7 , 32'hFFFFFFFE , 32'h0000000A , 32'h00000000 , 32'hFFFFFFFC , 32'h00000000 , 32'hFFFFFFFC , 32'hFFFFFFFB} , 
{32'h00000007 , 32'hFFFFFFFF , 32'hFFFFFFF4 , 32'hFFFFFFE0 , 32'hFFFFFFE0 , 32'h00000006 , 32'h00000003 , 32'h00000025 , 32'h0000009A , 32'h7FFFF800 , 32'hFFFFFF12 , 32'hFFFFFFB2 , 32'h00000027 , 32'h00000053 , 32'hFFFFFFFD , 32'h00000001 , 32'hFFFFFFFE , 32'hFFFFFFFA , 32'hFFFFFFE9 , 32'hFFFFFFDE , 32'h00000014 , 32'hFFFFFFF8 , 32'h00000005 , 32'hFFFFFFD6 , 32'h00000000 , 32'hFFFFFFF6 , 32'hFFFFFFF5 , 32'h00000004 , 32'hFFFFFFFD , 32'hFFFFFFF4 , 32'h00000002 , 32'h00000008 , 32'hFFFFFFF3 , 32'hFFFFFFFC , 32'hFFFFFFF3 , 32'h00000000 , 32'h00000007} , 
{32'h00000000 , 32'hFFFFFFFB , 32'hFFFFFFEC , 32'h00000009 , 32'h00000019 , 32'h00000036 , 32'hFFFFFFFE , 32'h0000003B , 32'hFFFFFF6E , 32'hFFFFFF12 , 32'h80000800 , 32'hFFFFFFD7 , 32'hFFFFFFDB , 32'h00000028 , 32'h0000000E , 32'h00000001 , 32'h0000001E , 32'hFFFFFFFA , 32'hFFFFFFF2 , 32'hFFFFFFF7 , 32'h0000000C , 32'h00000015 , 32'h00000002 , 32'hFFFFFFF5 , 32'h00000008 , 32'hFFFFFFFE , 32'h00000012 , 32'h00000001 , 32'h00000002 , 32'hFFFFFFF8 , 32'hFFFFFFFE , 32'h00000000 , 32'hFFFFFFFE , 32'hFFFFFFEF , 32'hFFFFFFF9 , 32'hFFFFFFFD , 32'h00000004} , 
{32'hFFFFFFFB , 32'h00000012 , 32'hFFFFFFF3 , 32'h0000000F , 32'hFFFFFFE1 , 32'hFFFFFFF1 , 32'h00000004 , 32'hFFFFFFF5 , 32'h0000001E , 32'h0000004C , 32'hFFFFFFD7 , 32'h7FFFF800 , 32'hFFFFFFAE , 32'h00000000 , 32'h0000000E , 32'h0000002D , 32'h0000000C , 32'hFFFFFFE0 , 32'h00000020 , 32'hFFFFFFC2 , 32'h00000009 , 32'hFFFFFFEE , 32'h00000016 , 32'hFFFFFFF1 , 32'hFFFFFFFE , 32'hFFFFFFFD , 32'hFFFFFFFA , 32'hFFFFFFF1 , 32'h00000017 , 32'h00000004 , 32'h00000005 , 32'h00000004 , 32'hFFFFFFEB , 32'hFFFFFFFA , 32'hFFFFFFFE , 32'h00000006 , 32'hFFFFFFFF} , 
{32'hFFFFFFF9 , 32'h00000000 , 32'hFFFFFFF8 , 32'h0000000A , 32'hFFFFFFFF , 32'h00000001 , 32'hFFFFFFFE , 32'hFFFFFFEA , 32'h0000000D , 32'h00000027 , 32'h00000023 , 32'hFFFFFFAE , 32'h80000800 , 32'h00000114 , 32'h0000006C , 32'hFFFFFF8C , 32'h00000032 , 32'hFFFFFFF9 , 32'h00000001 , 32'h00000032 , 32'hFFFFFFEC , 32'h0000000A , 32'h00000000 , 32'hFFFFFFFB , 32'h00000000 , 32'h00000017 , 32'hFFFFFFE6 , 32'h0000000A , 32'hFFFFFFFA , 32'h00000004 , 32'hFFFFFFF7 , 32'hFFFFFFF2 , 32'h00000017 , 32'h00000006 , 32'h00000001 , 32'h0000000D , 32'hFFFFFFFC} , 
{32'hFFFFFFFE , 32'h00000007 , 32'hFFFFFFFB , 32'h00000005 , 32'hFFFFFFFD , 32'h0000000E , 32'h00000021 , 32'h0000000F , 32'h00000010 , 32'h00000053 , 32'hFFFFFFD6 , 32'h00000000 , 32'hFFFFFEEA , 32'h80000800 , 32'hFFFFFE80 , 32'h00000032 , 32'h00000049 , 32'h0000001D , 32'hFFFFFFF0 , 32'hFFFFFFBC , 32'h00000023 , 32'h0000001D , 32'h00000000 , 32'hFFFFFFF8 , 32'hFFFFFFFF , 32'h0000000E , 32'h00000007 , 32'hFFFFFFEB , 32'h00000014 , 32'h0000000A , 32'hFFFFFFED , 32'h00000018 , 32'h00000008 , 32'h00000001 , 32'h0000000A , 32'h0000000E , 32'hFFFFFFF6} , 
{32'h00000001 , 32'h00000009 , 32'h00000009 , 32'hFFFFFFFB , 32'hFFFFFFFD , 32'hFFFFFFF5 , 32'h0000001B , 32'h00000025 , 32'hFFFFFFF6 , 32'hFFFFFFFD , 32'hFFFFFFF0 , 32'h0000000E , 32'hFFFFFF92 , 32'h0000017E , 32'h80000800 , 32'hFFFFFFC8 , 32'h0000003A , 32'hFFFFFFE9 , 32'hFFFFFFE7 , 32'hFFFFFFF8 , 32'h0000000C , 32'hFFFFFFE6 , 32'hFFFFFFF3 , 32'hFFFFFFEF , 32'hFFFFFFE1 , 32'h00000006 , 32'hFFFFFFF9 , 32'h00000022 , 32'h00000019 , 32'h0000000C , 32'hFFFFFFFA , 32'hFFFFFFFB , 32'hFFFFFFF9 , 32'h00000000 , 32'hFFFFFFFD , 32'hFFFFFFFB , 32'hFFFFFFF1} , 
{32'h00000004 , 32'hFFFFFFF4 , 32'hFFFFFFEC , 32'h0000001A , 32'hFFFFFFF0 , 32'h0000001F , 32'h00000003 , 32'hFFFFFFF8 , 32'hFFFFFFE7 , 32'hFFFFFFFD , 32'h00000001 , 32'hFFFFFFD1 , 32'hFFFFFF8C , 32'h00000032 , 32'hFFFFFFC8 , 32'h7FFFF800 , 32'hFFFFFF88 , 32'hFFFFFFF8 , 32'hFFFFFFFA , 32'hFFFFFFB7 , 32'h0000001A , 32'hFFFFFFED , 32'hFFFFFFF4 , 32'h0000000B , 32'h00000014 , 32'h00000013 , 32'h00000011 , 32'h00000001 , 32'h00000000 , 32'h00000001 , 32'h00000007 , 32'h00000000 , 32'hFFFFFFF7 , 32'h0000000D , 32'hFFFFFFF5 , 32'hFFFFFFFB , 32'h00000000} , 
{32'h00000000 , 32'hFFFFFFFE , 32'h00000010 , 32'hFFFFFFFC , 32'hFFFFFFF2 , 32'hFFFFFFF0 , 32'h0000000D , 32'h00000013 , 32'hFFFFFFEA , 32'hFFFFFFFE , 32'hFFFFFFE0 , 32'h0000000C , 32'hFFFFFFCC , 32'hFFFFFFB5 , 32'hFFFFFFC4 , 32'hFFFFFF88 , 32'h80000800 , 32'h0000003B , 32'h00000023 , 32'hFFFFFFDD , 32'h0000003B , 32'hFFFFFFC8 , 32'hFFFFFFE1 , 32'h00000007 , 32'hFFFFFFE4 , 32'hFFFFFFED , 32'h0000001B , 32'hFFFFFFF8 , 32'h0000000A , 32'h00000000 , 32'h00000009 , 32'hFFFFFFED , 32'h00000001 , 32'h00000003 , 32'h00000008 , 32'hFFFFFFE9 , 32'h00000018} , 
{32'h00000002 , 32'hFFFFFFFB , 32'h00000013 , 32'h0000000A , 32'hFFFFFFFF , 32'hFFFFFFFE , 32'h00000018 , 32'h0000000D , 32'hFFFFFFF7 , 32'h00000004 , 32'hFFFFFFFA , 32'h0000001E , 32'hFFFFFFF9 , 32'h0000001D , 32'hFFFFFFE9 , 32'h00000006 , 32'h0000003B , 32'h7FFFF800 , 32'h0000007F , 32'hFFFFFFEF , 32'h00000011 , 32'h0000002F , 32'hFFFFFFF6 , 32'hFFFFFFE7 , 32'hFFFFFFF6 , 32'h00000004 , 32'hFFFFFFEB , 32'h00000000 , 32'hFFFFFFF3 , 32'h00000010 , 32'h00000009 , 32'hFFFFFFF9 , 32'h00000007 , 32'h00000000 , 32'hFFFFFFFF , 32'hFFFFFFFD , 32'h00000000} , 
{32'hFFFFFFF9 , 32'h00000009 , 32'hFFFFFFF0 , 32'hFFFFFFFD , 32'h00000007 , 32'hFFFFFFF8 , 32'h00000002 , 32'hFFFFFFFA , 32'hFFFFFFE5 , 32'hFFFFFFE9 , 32'h0000000C , 32'h00000020 , 32'hFFFFFFFD , 32'h0000000E , 32'h00000017 , 32'hFFFFFFFA , 32'hFFFFFFDB , 32'h0000007F , 32'h80000800 , 32'h00000136 , 32'hFFFFFF81 , 32'hFFFFFFE0 , 32'hFFFFFFD3 , 32'hFFFFFFEF , 32'h0000001B , 32'hFFFFFFF8 , 32'h00000007 , 32'h00000001 , 32'h00000009 , 32'h00000003 , 32'h00000002 , 32'hFFFFFFEE , 32'hFFFFFFF6 , 32'h0000001B , 32'hFFFFFFFD , 32'hFFFFFFFD , 32'h00000004} , 
{32'hFFFFFFF4 , 32'hFFFFFFF5 , 32'h00000001 , 32'h00000000 , 32'hFFFFFFFD , 32'h00000000 , 32'hFFFFFFFB , 32'hFFFFFFE6 , 32'h0000000F , 32'h00000020 , 32'hFFFFFFF7 , 32'h0000003C , 32'h00000032 , 32'hFFFFFFBC , 32'hFFFFFFF8 , 32'h00000047 , 32'hFFFFFFDD , 32'h0000000F , 32'h00000136 , 32'h7FFFF800 , 32'h00000121 , 32'hFFFFFFE2 , 32'hFFFFFFC4 , 32'h00000009 , 32'h0000000D , 32'h00000017 , 32'hFFFFFFFD , 32'h00000008 , 32'hFFFFFFDD , 32'h00000007 , 32'h00000007 , 32'h00000001 , 32'hFFFFFFF1 , 32'h00000013 , 32'h00000000 , 32'hFFFFFFF9 , 32'hFFFFFFF7} , 
{32'h00000000 , 32'h00000003 , 32'h00000005 , 32'hFFFFFFEB , 32'h00000002 , 32'hFFFFFFFE , 32'h00000006 , 32'hFFFFFFF1 , 32'h0000000A , 32'hFFFFFFEA , 32'h0000000C , 32'hFFFFFFF5 , 32'hFFFFFFEC , 32'h00000023 , 32'h0000000C , 32'hFFFFFFE4 , 32'h0000003B , 32'hFFFFFFED , 32'hFFFFFF81 , 32'hFFFFFEDD , 32'h7FFFF800 , 32'hFFFFFF78 , 32'h00000011 , 32'h00000027 , 32'hFFFFFFF1 , 32'h00000018 , 32'h00000008 , 32'h00000004 , 32'h00000007 , 32'h00000014 , 32'h00000012 , 32'hFFFFFFF2 , 32'h00000001 , 32'h00000000 , 32'h00000016 , 32'hFFFFFFFD , 32'h00000008} , 
{32'h00000003 , 32'h00000001 , 32'h00000003 , 32'h00000003 , 32'h00000004 , 32'h00000003 , 32'h00000006 , 32'h00000010 , 32'h00000001 , 32'hFFFFFFF8 , 32'hFFFFFFE9 , 32'hFFFFFFEE , 32'hFFFFFFF4 , 32'hFFFFFFE1 , 32'h00000018 , 32'hFFFFFFED , 32'h00000036 , 32'h0000002F , 32'h0000001E , 32'hFFFFFFE2 , 32'hFFFFFF78 , 32'h80000800 , 32'hFFFFFF1B , 32'h00000044 , 32'h0000000F , 32'hFFFFFFBB , 32'hFFFFFFE6 , 32'h00000006 , 32'h00000017 , 32'hFFFFFFFF , 32'h00000003 , 32'hFFFFFFF1 , 32'h00000006 , 32'hFFFFFFF9 , 32'hFFFFFFEB , 32'hFFFFFFF8 , 32'hFFFFFFF4} , 
{32'h00000000 , 32'hFFFFFFFA , 32'h00000000 , 32'h00000005 , 32'h00000003 , 32'h00000000 , 32'h00000001 , 32'h00000007 , 32'h00000003 , 32'h00000005 , 32'hFFFFFFFC , 32'h00000016 , 32'hFFFFFFFE , 32'hFFFFFFFE , 32'h0000000B , 32'hFFFFFFF4 , 32'h0000001D , 32'hFFFFFFF6 , 32'h0000002B , 32'hFFFFFFC4 , 32'h00000011 , 32'h000000E3 , 32'h80000800 , 32'hFFFFFE59 , 32'hFFFFFF83 , 32'hFFFFFFCA , 32'hFFFFFFBE , 32'hFFFFFFB3 , 32'hFFFFFFC9 , 32'h00000011 , 32'h0000000C , 32'h00000003 , 32'h00000014 , 32'hFFFFFFE1 , 32'h00000027 , 32'hFFFFFFD1 , 32'h00000010} , 
{32'h00000000 , 32'h00000000 , 32'hFFFFFFFF , 32'h00000009 , 32'hFFFFFFFD , 32'h00000002 , 32'h00000006 , 32'hFFFFFFEF , 32'h00000015 , 32'h00000028 , 32'hFFFFFFF5 , 32'h0000000D , 32'hFFFFFFFB , 32'hFFFFFFF8 , 32'hFFFFFFEF , 32'hFFFFFFF3 , 32'h00000007 , 32'h00000017 , 32'hFFFFFFEF , 32'hFFFFFFF5 , 32'hFFFFFFD7 , 32'h00000044 , 32'hFFFFFE59 , 32'h7FFFF800 , 32'h00000017 , 32'hFFFFFFAC , 32'h00000039 , 32'hFFFFFFDD , 32'hFFFFFFCB , 32'h00000000 , 32'h0000001E , 32'hFFFFFFFB , 32'hFFFFFFEE , 32'hFFFFFFBE , 32'hFFFFFFF6 , 32'h0000000D , 32'h00000007} , 
{32'h00000001 , 32'hFFFFFFFF , 32'h00000005 , 32'hFFFFFFF6 , 32'h00000007 , 32'h00000000 , 32'hFFFFFFF7 , 32'hFFFFFFFC , 32'hFFFFFFF3 , 32'h00000000 , 32'hFFFFFFF6 , 32'hFFFFFFFE , 32'hFFFFFFFE , 32'h00000000 , 32'h0000001D , 32'h00000014 , 32'h0000001A , 32'hFFFFFFF6 , 32'hFFFFFFE3 , 32'h0000000D , 32'hFFFFFFF1 , 32'hFFFFFFEF , 32'h0000007B , 32'h00000017 , 32'h80000800 , 32'hFFFFFF73 , 32'h0000009A , 32'hFFFFFF2A , 32'h00000059 , 32'h00000014 , 32'hFFFFFFED , 32'h0000002D , 32'hFFFFFFFF , 32'hFFFFFFF5 , 32'hFFFFFFD2 , 32'hFFFFFFDA , 32'hFFFFFFFF} , 
{32'hFFFFFFF4 , 32'hFFFFFFF6 , 32'hFFFFFFF4 , 32'h00000004 , 32'h00000001 , 32'h00000004 , 32'h00000003 , 32'hFFFFFFE8 , 32'h00000000 , 32'hFFFFFFF6 , 32'h00000000 , 32'hFFFFFFFD , 32'hFFFFFFE7 , 32'hFFFFFFF0 , 32'hFFFFFFF8 , 32'h00000013 , 32'h00000011 , 32'h00000004 , 32'h00000006 , 32'h00000017 , 32'h00000018 , 32'h00000043 , 32'h00000034 , 32'hFFFFFFAC , 32'h0000008B , 32'h80000800 , 32'hFFFFFF32 , 32'h00000182 , 32'hFFFFFFE1 , 32'hFFFFFFD6 , 32'hFFFFFFB9 , 32'hFFFFFFD8 , 32'h00000013 , 32'h00000024 , 32'hFFFFFFF1 , 32'h00000017 , 32'hFFFFFFFC} , 
{32'hFFFFFFFB , 32'hFFFFFFFC , 32'hFFFFFFF3 , 32'h0000000A , 32'hFFFFFFFF , 32'h00000000 , 32'h00000007 , 32'h00000017 , 32'hFFFFFFE8 , 32'hFFFFFFF5 , 32'hFFFFFFEC , 32'hFFFFFFFA , 32'h00000018 , 32'hFFFFFFF7 , 32'h00000005 , 32'h00000011 , 32'hFFFFFFE3 , 32'hFFFFFFEB , 32'hFFFFFFF7 , 32'hFFFFFFFD , 32'h00000008 , 32'h00000018 , 32'h00000040 , 32'h00000039 , 32'hFFFFFF64 , 32'h000000CC , 32'h80000800 , 32'h00000194 , 32'h00000014 , 32'h00000029 , 32'hFFFFFFAE , 32'h00000064 , 32'h00000021 , 32'h00000021 , 32'hFFFFFFF4 , 32'h00000007 , 32'hFFFFFFE8} , 
{32'h0000000B , 32'h00000000 , 32'hFFFFFFFE , 32'h00000004 , 32'h00000003 , 32'hFFFFFFFA , 32'hFFFFFFFA , 32'hFFFFFFFC , 32'hFFFFFFEF , 32'h00000004 , 32'hFFFFFFFD , 32'hFFFFFFF1 , 32'hFFFFFFF4 , 32'h00000013 , 32'hFFFFFFDC , 32'h00000001 , 32'h00000006 , 32'h00000000 , 32'hFFFFFFFD , 32'h00000008 , 32'h00000004 , 32'hFFFFFFF8 , 32'h0000004B , 32'hFFFFFFDD , 32'h000000D4 , 32'hFFFFFE7C , 32'hFFFFFE6A , 32'h80000800 , 32'h000000FB , 32'hFFFFFFA4 , 32'hFFFFFFAA , 32'hFFFFFFFC , 32'hFFFFFFDC , 32'h00000012 , 32'h0000000B , 32'hFFFFFFEF , 32'hFFFFFFD8} , 
{32'h00000001 , 32'hFFFFFFFF , 32'hFFFFFFFC , 32'hFFFFFFF6 , 32'hFFFFFFF9 , 32'h00000001 , 32'h0000000F , 32'h00000008 , 32'h0000000C , 32'h00000001 , 32'h00000002 , 32'hFFFFFFE7 , 32'hFFFFFFFA , 32'h00000014 , 32'h00000019 , 32'hFFFFFFFF , 32'h0000000A , 32'h0000000B , 32'h00000009 , 32'h00000021 , 32'hFFFFFFF7 , 32'h00000017 , 32'hFFFFFFC9 , 32'h00000033 , 32'h00000059 , 32'hFFFFFFE1 , 32'h00000014 , 32'h000000FB , 32'h7FFFF800 , 32'h000000B8 , 32'h00000041 , 32'hFFFFFF95 , 32'hFFFFFFED , 32'h0000000F , 32'h0000002E , 32'hFFFFFFEE , 32'h00000000} , 
{32'h00000005 , 32'hFFFFFFFF , 32'hFFFFFFF7 , 32'hFFFFFFFB , 32'hFFFFFFFA , 32'h00000003 , 32'hFFFFFFFA , 32'hFFFFFFFE , 32'h00000007 , 32'hFFFFFFF4 , 32'h00000006 , 32'h00000004 , 32'hFFFFFFFA , 32'hFFFFFFF4 , 32'hFFFFFFF2 , 32'h00000001 , 32'hFFFFFFFE , 32'h00000010 , 32'hFFFFFFFB , 32'h00000007 , 32'h00000014 , 32'h00000000 , 32'hFFFFFFED , 32'h00000000 , 32'hFFFFFFEA , 32'h00000028 , 32'hFFFFFFD5 , 32'h0000005A , 32'h000000B8 , 32'h80000800 , 32'h0000024A , 32'h00000000 , 32'hFFFFFF90 , 32'h0000007B , 32'hFFFFFFC0 , 32'hFFFFFFBD , 32'h00000021} , 
{32'hFFFFFFF9 , 32'h00000000 , 32'hFFFFFFFF , 32'h0000000B , 32'hFFFFFFFE , 32'h00000004 , 32'h00000007 , 32'h00000004 , 32'h00000000 , 32'h00000002 , 32'h00000000 , 32'h00000005 , 32'h00000007 , 32'h00000011 , 32'h00000004 , 32'h00000007 , 32'hFFFFFFF5 , 32'h00000009 , 32'hFFFFFFFC , 32'h00000007 , 32'h00000012 , 32'hFFFFFFFB , 32'hFFFFFFF2 , 32'h0000001E , 32'h00000011 , 32'h00000045 , 32'h00000050 , 32'h00000054 , 32'h00000041 , 32'hFFFFFDB4 , 32'h80000800 , 32'hFFFFFECB , 32'h000000A3 , 32'hFFFFFFCE , 32'h00000064 , 32'hFFFFFFB5 , 32'hFFFFFFF8} , 
{32'hFFFFFFFE , 32'h00000005 , 32'h00000004 , 32'hFFFFFFFE , 32'h00000000 , 32'h00000000 , 32'hFFFFFFFF , 32'h00000003 , 32'hFFFFFFF4 , 32'h00000008 , 32'hFFFFFFFF , 32'h00000004 , 32'h0000000C , 32'hFFFFFFE6 , 32'h00000003 , 32'h00000000 , 32'h00000011 , 32'hFFFFFFF9 , 32'h00000010 , 32'h00000001 , 32'hFFFFFFF2 , 32'h0000000D , 32'hFFFFFFFB , 32'hFFFFFFFB , 32'hFFFFFFD1 , 32'h00000026 , 32'hFFFFFF9A , 32'h00000002 , 32'hFFFFFF95 , 32'hFFFFFFFE , 32'h00000133 , 32'h80000800 , 32'hFFFFFFFA , 32'hFFFFFFB0 , 32'hFFFFFFAD , 32'hFFFFFFA3 , 32'hFFFFFFDB} , 
{32'hFFFFFFF9 , 32'hFFFFFFF9 , 32'h00000008 , 32'h00000000 , 32'h00000003 , 32'hFFFFFFFE , 32'h00000000 , 32'hFFFFFFFA , 32'hFFFFFFFF , 32'hFFFFFFF3 , 32'h00000000 , 32'hFFFFFFEB , 32'hFFFFFFE7 , 32'hFFFFFFF6 , 32'h00000005 , 32'hFFFFFFF7 , 32'hFFFFFFFD , 32'h00000007 , 32'h00000008 , 32'hFFFFFFF1 , 32'h00000001 , 32'hFFFFFFF8 , 32'hFFFFFFEA , 32'hFFFFFFEE , 32'h00000000 , 32'hFFFFFFEB , 32'hFFFFFFDD , 32'h00000022 , 32'hFFFFFFED , 32'h0000006E , 32'hFFFFFF5B , 32'h00000004 , 32'h80000800 , 32'h0000003E , 32'h00000022 , 32'hFFFFFFFD , 32'hFFFFFFD2} , 
{32'hFFFFFFFF , 32'hFFFFFFF3 , 32'hFFFFFFFD , 32'hFFFFFFFC , 32'hFFFFFFFF , 32'hFFFFFFF6 , 32'hFFFFFFFC , 32'hFFFFFFFD , 32'h00000002 , 32'hFFFFFFFC , 32'h0000000F , 32'hFFFFFFFA , 32'hFFFFFFF8 , 32'hFFFFFFFD , 32'hFFFFFFFF , 32'h0000000D , 32'hFFFFFFFB , 32'h00000000 , 32'hFFFFFFE3 , 32'h00000013 , 32'h00000000 , 32'h00000005 , 32'h0000001D , 32'hFFFFFFBE , 32'h00000009 , 32'hFFFFFFDA , 32'hFFFFFFDD , 32'hFFFFFFEC , 32'h0000000F , 32'hFFFFFF83 , 32'h00000030 , 32'h0000004E , 32'hFFFFFFC0 , 32'h80000800 , 32'h00000089 , 32'h00000063 , 32'h00000040} , 
{32'h00000002 , 32'hFFFFFFF8 , 32'hFFFFFFFE , 32'hFFFFFFFB , 32'hFFFFFFFE , 32'hFFFFFFFB , 32'h0000000B , 32'h00000009 , 32'hFFFFFFFE , 32'hFFFFFFF3 , 32'h00000005 , 32'hFFFFFFFE , 32'hFFFFFFFD , 32'hFFFFFFF4 , 32'h00000001 , 32'hFFFFFFF5 , 32'hFFFFFFF6 , 32'hFFFFFFFF , 32'h00000001 , 32'h00000000 , 32'h00000016 , 32'h00000013 , 32'hFFFFFFD7 , 32'hFFFFFFF6 , 32'h0000002C , 32'h0000000D , 32'h0000000A , 32'hFFFFFFF3 , 32'h0000002E , 32'h0000003E , 32'hFFFFFF9A , 32'h00000051 , 32'hFFFFFFDC , 32'hFFFFFF75 , 32'h80000800 , 32'h000003E8 , 32'h00000091} , 
{32'h00000002 , 32'hFFFFFFF7 , 32'h00000002 , 32'hFFFFFFFF , 32'h00000000 , 32'h00000000 , 32'h00000001 , 32'h0000000A , 32'hFFFFFFFC , 32'hFFFFFFFE , 32'hFFFFFFFD , 32'hFFFFFFF8 , 32'h0000000D , 32'h0000000E , 32'hFFFFFFFB , 32'h00000003 , 32'hFFFFFFE9 , 32'h00000001 , 32'hFFFFFFFD , 32'h00000005 , 32'h00000001 , 32'hFFFFFFF8 , 32'hFFFFFFD1 , 32'hFFFFFFF1 , 32'hFFFFFFDA , 32'h00000017 , 32'h00000007 , 32'hFFFFFFEF , 32'h00000010 , 32'hFFFFFFBD , 32'hFFFFFFB5 , 32'hFFFFFFA3 , 32'hFFFFFFFD , 32'h00000063 , 32'h000003E8 , 32'h7FFFF800 , 32'h00000029} , 
{32'hFFFFFFFE , 32'hFFFFFFFD , 32'hFFFFFFFD , 32'hFFFFFFFC , 32'h00000007 , 32'hFFFFFFFD , 32'h00000004 , 32'hFFFFFFFA , 32'h00000003 , 32'h00000007 , 32'hFFFFFFFA , 32'hFFFFFFFF , 32'h00000002 , 32'h00000008 , 32'h0000000D , 32'h00000000 , 32'hFFFFFFE6 , 32'h00000000 , 32'hFFFFFFFA , 32'hFFFFFFF7 , 32'h00000008 , 32'h0000000A , 32'hFFFFFFEE , 32'h00000007 , 32'h00000000 , 32'h00000002 , 32'h00000016 , 32'h00000026 , 32'h00000000 , 32'hFFFFFFDD , 32'h00000006 , 32'h00000023 , 32'h0000002C , 32'hFFFFFFBE , 32'hFFFFFF6D , 32'h00000029 , 32'h80000800}
};

logic signed [31:0] VT_1 [37][300] ='{
{32'hFD02A1DC , 32'hA3E68A00 , 32'h000015DA , 32'hEA0FADA0 , 32'hFFFE4AA0 , 32'h0889E4C0 , 32'hFFFF2E89 , 32'h0001952F , 32'hFFF8CFEC , 32'hFFFF429D , 32'h0ABDD950 , 32'hE8A9AC00 , 32'h1343E9E0 , 32'hFFFF1CB2 , 32'hFFF9FC43 , 32'hE9F20540 , 32'hFFFE9741 , 32'h01329B40 , 32'hF5E65930 , 32'h00013808 , 32'hFFFF93FB , 32'h004CE82C , 32'hF672CB20 , 32'hFB2E0EF0 , 32'h061D7B98 , 32'h00007855 , 32'hFC2B5FC0 , 32'hFF019849 , 32'hFFFD706A , 32'h0AA57480 , 32'hFFFED8BE , 32'h007269EF , 32'h00002C4C , 32'hFFFA13FF , 32'hFFFF23D4 , 32'hE4BD5120 , 32'h07135D40 , 32'h04CE97F0 , 32'h0002FAE1 , 32'h07B124D8 , 32'h1C675540 , 32'h00012C58 , 32'h00058023 , 32'hF9203BC0 , 32'h02FB1F44 , 32'h208B7D80 , 32'hF0FBEC30 , 32'hFFFE7645 , 32'h0B20AF60 , 32'hC1B23140 , 32'hFE9B8A60 , 32'h000064E7 , 32'h0727B1F0 , 32'h1F1649C0 , 32'h08A1E840 , 32'hFFFFE0E5 , 32'h07A39658 , 32'hFFFFC810 , 32'h0002623F , 32'h01BF4F58 , 32'hFFA1F5B5 , 32'h0E1D39B0 , 32'hC47F7880 , 32'h0001F36A , 32'hE4C51D20 , 32'hFFFEC781 , 32'hEED58880 , 32'h0120D604 , 32'hFFFFAD64 , 32'h0014A77B , 32'h05FE1CE8 , 32'hF4806D10 , 32'hFFFFCCA5 , 32'h0005A534 , 32'h0000135D , 32'hDEC5F400 , 32'hF571F7D0 , 32'h0000FD84 , 32'hD40FB7C0 , 32'h02A60E30 , 32'hFFFE04C0 , 32'hD44CD240 , 32'hEF394AA0 , 32'h0000042B , 32'h03CA46B0 , 32'h261A4BC0 , 32'hF3538680 , 32'h0001892B , 32'hFFFE180F , 32'h35B420C0 , 32'h0003D3AC , 32'hF54AC460 , 32'h0000A925 , 32'hF6AA31D0 , 32'hFE5C5714 , 32'h0004D7CC , 32'hFFFCA76C , 32'hFFFF6404 , 32'h00049120 , 32'hECE063A0 , 32'hFC67D5BC , 32'h0003178E , 32'h01C033F0 , 32'h057F1508 , 32'h05E51E68 , 32'h0002F7F3 , 32'h00A3A08A , 32'h0000E809 , 32'h0FD65A10 , 32'h55DC6700 , 32'hFFFF1EC4 , 32'h04D45298 , 32'hFFFDB49F , 32'h000129AD , 32'hEFD5CAA0 , 32'h05FAD3B0 , 32'hFF56F81D , 32'h000064F3 , 32'hF3BE8A20 , 32'h0003C813 , 32'hFFFC2815 , 32'hEFAA2E40 , 32'h00059647 , 32'h0000A431 , 32'hFF5B3A5C , 32'hECB9A140 , 32'h0000757E , 32'hFFFDEAFB , 32'h00031312 , 32'hFFFC030B , 32'hFFFEEFA9 , 32'h0270A8E8 , 32'hF3498780 , 32'h0002E721 , 32'hFFFE6B25 , 32'h6714E100 , 32'h1E6441A0 , 32'h00036A14 , 32'hFFFE0D36 , 32'hFF3B5337 , 32'h000023AB , 32'hFFFFB97D , 32'hFD118024 , 32'h09187100 , 32'h0158F088 , 32'hF9484708 , 32'hFFFDC01A , 32'hFFFDF3D8 , 32'h097EE1C0 , 32'hFFFF5ED9 , 32'hFFFBDBC6 , 32'hFE5840B0 , 32'hFFFE939D , 32'h0000904E , 32'h099C5340 , 32'hFFF748AC , 32'hE519C760 , 32'hFC2367E8 , 32'h00032EF1 , 32'h0003794A , 32'hFFFBD272 , 32'hE6342260 , 32'hFDBD6D64 , 32'h15F34680 , 32'h094CBBA0 , 32'hFFFE01A0 , 32'hE17E2F80 , 32'h0000D185 , 32'h0001C7A2 , 32'hD84C9100 , 32'h005DC028 , 32'h03E245CC , 32'hFFFCDD55 , 32'hDB5944C0 , 32'hFC7016EC , 32'hFB9D8260 , 32'hD363CC80 , 32'hF8DFF178 , 32'hFCB62034 , 32'hFE5F5CD4 , 32'h07859F80 , 32'h000070C5 , 32'hFFFD1D40 , 32'hFFFE0348 , 32'hF6216060 , 32'h0AC08050 , 32'h02432650 , 32'h02A0A374 , 32'hF2A41F60 , 32'h0624DB20 , 32'h00046A0C , 32'hEBE484A0 , 32'hEC0C8840 , 32'hFFFAC585 , 32'h00650BFC , 32'hFFFD8572 , 32'h1122FFE0 , 32'h03B42664 , 32'hFFFC6BA6 , 32'h00057C7D , 32'hFFFDEA8A , 32'h00095F1C , 32'h0005359D , 32'hFFFF7623 , 32'h085848D0 , 32'h02E15950 , 32'hEF85AD20 , 32'h0595DFC8 , 32'h1C21DAA0 , 32'h23D2B4C0 , 32'h00011D71 , 32'hFFFFE96E , 32'h00055E08 , 32'h00002658 , 32'hFFFE2D72 , 32'h01A46FB4 , 32'h0151EA00 , 32'h181BDF40 , 32'h0003D983 , 32'hFFFE6765 , 32'h0003BB7A , 32'hFFF6B005 , 32'hF8AA4450 , 32'h1D13A920 , 32'hFFFDE94E , 32'hFFFC4AA2 , 32'hFFFAD8CE , 32'hD8CFCD80 , 32'h05873888 , 32'h13550880 , 32'hFFFC469B , 32'hFFFBFCC3 , 32'h000578AF , 32'hFC89F01C , 32'h04FFFAD8 , 32'h1E1828A0 , 32'hFFFE199F , 32'hFE61B534 , 32'h00046A3F , 32'h0567A2D8 , 32'h0002D1C3 , 32'hF6222E40 , 32'h0001E366 , 32'hE2C40F40 , 32'hF8A4ADD0 , 32'h183B2840 , 32'hFB5EBDE8 , 32'hFFFE1EE5 , 32'h0A8906A0 , 32'hFC675F84 , 32'h0005804C , 32'hEF1D8880 , 32'h0002A9A0 , 32'h009E8442 , 32'hF1F56FD0 , 32'hFBEA3860 , 32'hFFFD681E , 32'hFFFCA26F , 32'hFE0F8CB4 , 32'h00006985 , 32'hFC746684 , 32'hFFFFB6EC , 32'h00F49CDB , 32'hFFFEFBD4 , 32'hF2DC23B0 , 32'hFFFF41A1 , 32'hFFFBAB7F , 32'h000109E4 , 32'hFEB9FC4C , 32'hF0B149A0 , 32'hFFFD6183 , 32'hFFF98050 , 32'hFFFEB1AA , 32'h00004F96 , 32'hF4E7BC70 , 32'hF6E25430 , 32'hFFC820D9 , 32'h4195C600 , 32'h0B1924C0 , 32'h00038853 , 32'h000187CC , 32'h0000E73B , 32'h09651230 , 32'hFFFE3B40 , 32'h0006AFE9 , 32'h075F1B58 , 32'h067691D0 , 32'h0001B32B , 32'h255D3040 , 32'hFF4AD714 , 32'h09DA9640 , 32'h003CAB61 , 32'h000172AB , 32'h03633864 , 32'hE53EAFA0 , 32'hF7E054C0 , 32'h00010BA8 , 32'hD4F9E540 , 32'hEFD45CE0 , 32'hE4740660} , 
{32'h0C985ED0 , 32'hCE8FCAC0 , 32'hFFFFE426 , 32'h0563C4F0 , 32'h000420EA , 32'h04097458 , 32'h00077ACE , 32'h00037B2E , 32'hFFFAD215 , 32'hFFFE621B , 32'h03267594 , 32'hE5A5AF60 , 32'hFEEA6FF4 , 32'h0003CC75 , 32'hFFFFD433 , 32'hDA074D00 , 32'hFFFA8717 , 32'h0F6E23B0 , 32'h0D789550 , 32'h00054542 , 32'h00012990 , 32'h03952298 , 32'hFAF8C610 , 32'hE0AB3BE0 , 32'hE21749A0 , 32'hFFF94EB6 , 32'hFEB94520 , 32'hFF741C7A , 32'h0004208D , 32'hE6CF0B60 , 32'hFFFC6709 , 32'h150F60C0 , 32'hFFFDEBE8 , 32'hFFFBE621 , 32'h0003965A , 32'hE9398840 , 32'hFF887313 , 32'h1DE3CD80 , 32'hFFFC2D45 , 32'hFC3D302C , 32'h01183824 , 32'hFFFEFF76 , 32'hFFFFBCF4 , 32'h0A344C10 , 32'h07B7B820 , 32'hF69ED790 , 32'hF8FC8A00 , 32'h000109B7 , 32'h1B782440 , 32'hD8E56D00 , 32'hFCA4A3EC , 32'h00069C13 , 32'hF7077EA0 , 32'h09636020 , 32'hFE64D9C0 , 32'hFFFE84DF , 32'hF78049B0 , 32'h0005563E , 32'h00036043 , 32'h03B325DC , 32'hFDE7632C , 32'hFF2AB0F0 , 32'h4A7BE780 , 32'h00041C9D , 32'hF446D090 , 32'hFFFE7D8F , 32'hFB7C4BC8 , 32'h019A3B48 , 32'hFFFFFBA6 , 32'hF2785C60 , 32'hFA082330 , 32'h0CB51FD0 , 32'h00063914 , 32'hFFFD75A2 , 32'hFFFB7FFE , 32'hED4AF840 , 32'h0635F1E0 , 32'hFFFC8301 , 32'hFE88C01C , 32'h034F5234 , 32'h0000F884 , 32'hF8A4B300 , 32'hF2BD1D00 , 32'hFFFCDE3E , 32'h0AE45700 , 32'hF492FE90 , 32'h0E3B1790 , 32'hFFFD337F , 32'hFFFEE206 , 32'hF7C8EAB0 , 32'h0004EE86 , 32'hEDE24100 , 32'hFFFE4E06 , 32'h17007D20 , 32'hFFDBDC96 , 32'h0000A5DB , 32'h00007035 , 32'hFFFB32CD , 32'h0001AC3F , 32'hEEBA4FA0 , 32'hFE067C98 , 32'h0000B84C , 32'h05AF1CF8 , 32'h0D9C9450 , 32'hFC1F65C8 , 32'hFFFA02E7 , 32'h00E0A1D8 , 32'hFFFACD56 , 32'hF71A65F0 , 32'hA5349B80 , 32'hFFFDD4B5 , 32'hE88434A0 , 32'h0003499B , 32'hFFFDE4F8 , 32'h09AA3060 , 32'hFFE1B3D2 , 32'hFD4CFF94 , 32'hFFF703FE , 32'h03E0E99C , 32'hFFFEB643 , 32'hFFFF48C4 , 32'hFC9270DC , 32'h0003BF1B , 32'hFFFF662C , 32'h085C7D10 , 32'hF1C818A0 , 32'hFFFD8279 , 32'hFFFE1B76 , 32'hFFFE399B , 32'hFFFF1400 , 32'h0002D03A , 32'hE609E6E0 , 32'h0C2E68B0 , 32'h000043ED , 32'h000214C1 , 32'h0CE2AE20 , 32'hFF7D4A50 , 32'h000104D3 , 32'h00048400 , 32'h114272E0 , 32'hFFFE0942 , 32'hFFF98CD1 , 32'h09F8D370 , 32'hFA46AA28 , 32'h043612B0 , 32'hFF37C5E3 , 32'hFFFEFDFD , 32'hFFFBDF11 , 32'h015C6974 , 32'hFFFF9422 , 32'hFFFFEEC4 , 32'hF8FD2308 , 32'hFFFEA80B , 32'h00022778 , 32'hF52B0B90 , 32'h00002725 , 32'h07034718 , 32'hFF5BC484 , 32'h000060F0 , 32'hFFFCF485 , 32'h0006EC9E , 32'hD23B9240 , 32'hF8FEE790 , 32'hE790F8A0 , 32'hF3D22CB0 , 32'h0001B69A , 32'h18E23420 , 32'h00045767 , 32'h0003DD38 , 32'h08243B40 , 32'hFD6AA414 , 32'h04127790 , 32'h0003497A , 32'hD7F5C900 , 32'h026CED30 , 32'hFFFCA2A1 , 32'hFE9E3E98 , 32'hFCF3C050 , 32'h4B820780 , 32'hFE2829E8 , 32'hFAE06370 , 32'h0002672F , 32'hFFFF89F2 , 32'hFFFECFC8 , 32'hF3554E10 , 32'hCE6FC080 , 32'h08AE1970 , 32'hFE9D5D30 , 32'hF8ED1500 , 32'hF42DD230 , 32'h0001A0BD , 32'hEBEC1220 , 32'hF56AFF90 , 32'hFFFBB765 , 32'hFDCE0F14 , 32'h00033282 , 32'hF8DA34D8 , 32'hCF128D40 , 32'h000850DD , 32'h0001DB12 , 32'hFFFDC378 , 32'hFFFD95B1 , 32'h00020FE0 , 32'hFFFDB001 , 32'h02438F50 , 32'h0FE09310 , 32'h0381EBF4 , 32'h17D70740 , 32'h0D09B2F0 , 32'hD5AB20C0 , 32'h0002AEC8 , 32'hFFFAE523 , 32'hFFFD7FDB , 32'h00021351 , 32'h000245E2 , 32'h03E49B40 , 32'h0DAAA880 , 32'h0BB5DC90 , 32'h0001466E , 32'hFFFD13EC , 32'h00007045 , 32'h0004E74D , 32'h18113120 , 32'hE18DE500 , 32'h00015460 , 32'h0004A70E , 32'h0000589C , 32'hE329AB20 , 32'h156DFDA0 , 32'hE92D5FE0 , 32'hFFFD104B , 32'hFFFDD759 , 32'hFFFF6403 , 32'h05795638 , 32'h01954E2C , 32'hDC535BC0 , 32'h00027A54 , 32'h026B1744 , 32'h0003751D , 32'h1219DE20 , 32'h00049919 , 32'hCB0ACEC0 , 32'h00062597 , 32'hD0E7C380 , 32'h09F6CCA0 , 32'h6CF08180 , 32'h1F6D0420 , 32'h00042A76 , 32'hFC5B5E5C , 32'hFBDF6158 , 32'hFFFD02D5 , 32'h150741A0 , 32'h00048558 , 32'hFDBA8C88 , 32'hF6541850 , 32'h007F1BB5 , 32'h0003A98A , 32'h0002B2F8 , 32'h21EF6640 , 32'h00030469 , 32'hEE3BAC60 , 32'h0001D330 , 32'h00FA2782 , 32'hFFFFE935 , 32'hFD362E90 , 32'hFFFF2F57 , 32'h0001AD1A , 32'h0000FB0F , 32'hFFFC4F5A , 32'h091A8DC0 , 32'hFFFC8DD4 , 32'h0000D668 , 32'hFFFE9178 , 32'h0000D2F1 , 32'hF0BBF880 , 32'h18C9DB20 , 32'hD71BE340 , 32'h161710E0 , 32'hEF0DDD80 , 32'h00019D3E , 32'hFFFFF515 , 32'hFFFF3B53 , 32'h039FB020 , 32'hFFFCF87A , 32'hFFFD5D50 , 32'hF96A05D0 , 32'h1519CEE0 , 32'hFFFD53AC , 32'hE0F04D00 , 32'h06956E70 , 32'hFE9D87B0 , 32'hE18CC860 , 32'hFFFE051F , 32'h05990700 , 32'h0543A638 , 32'hFC89B0C4 , 32'hFFFD6D6B , 32'hF78A65C0 , 32'h177AB580 , 32'h1E077F80} , 
{32'h0E978750 , 32'hC451B6C0 , 32'h00051D42 , 32'hF04FB740 , 32'h00027A27 , 32'hFEFE1D18 , 32'h000196A0 , 32'hFFFF592A , 32'h0005A33E , 32'h00026AB9 , 32'hFEE0FD7C , 32'hF6FAF6C0 , 32'hF9F01B70 , 32'h0000D2D0 , 32'h00040507 , 32'h19B581E0 , 32'hFFFC9D53 , 32'hCEE677C0 , 32'h009D5BD5 , 32'hFFFDFEBF , 32'hFFFFB89E , 32'h064C71B0 , 32'h08D36A00 , 32'h03D67278 , 32'hDAD20380 , 32'h00018055 , 32'h0A087910 , 32'hFCFC977C , 32'hFFFC549E , 32'hFC7C54B0 , 32'hFFFFE691 , 32'hF87E13F0 , 32'h0000FB2C , 32'hFFFFD3BE , 32'hFFFB1172 , 32'hEABC0520 , 32'hEAB70080 , 32'h117EE6A0 , 32'hFFFBD308 , 32'hE64A1820 , 32'h0DCAB1E0 , 32'h00004634 , 32'hFFFBB506 , 32'hF466F280 , 32'h2B5CE980 , 32'hCE120140 , 32'hFFFD366F , 32'hFFFEEC01 , 32'hF60D3360 , 32'h03350340 , 32'h015E5428 , 32'h0002EC24 , 32'hFC1FAE9C , 32'h025E0D78 , 32'hF986A0D8 , 32'h00041550 , 32'h009047F6 , 32'h0002BE94 , 32'h00013B61 , 32'h061F9C50 , 32'h023852D8 , 32'h036FD6EC , 32'hEE7FD760 , 32'h0000B6AB , 32'h1586A6E0 , 32'hFFFFCB33 , 32'hA7EEC600 , 32'hFA78E390 , 32'h0004215E , 32'h03DF363C , 32'h30658040 , 32'hE91ACB20 , 32'hFFFFE85F , 32'hFFFFC2CA , 32'hFFFBD3C3 , 32'hF8ACEE08 , 32'hF3792F70 , 32'h0002505E , 32'hF84E8DB8 , 32'hFC1DA0A0 , 32'hFFFE4F8F , 32'hDEDB3740 , 32'hF52F5C00 , 32'h00012139 , 32'hFDE3808C , 32'hDA17ED00 , 32'hF509BBF0 , 32'hFFFE186C , 32'hFFFEEEB5 , 32'h217D7380 , 32'hFFFFB418 , 32'hF9405170 , 32'h0001D50E , 32'hF8E8A260 , 32'h001914FA , 32'hFFFEE494 , 32'hFFFC4819 , 32'hFFFF7A24 , 32'hFFFEC862 , 32'hF8F5BB80 , 32'h0BF1D010 , 32'hFFFAC6B2 , 32'hF4E51650 , 32'hFDCC329C , 32'hFF359F76 , 32'h00030B82 , 32'hFF4B27A2 , 32'h0001A415 , 32'h08EBEBA0 , 32'h0652CFC0 , 32'hFFFC52FF , 32'h0D3E83C0 , 32'h00071C75 , 32'hFFFC677D , 32'h037993CC , 32'hFA5D63C0 , 32'h00C8F8F2 , 32'h0001C65A , 32'hF2530200 , 32'hFFFDF5DF , 32'h00001257 , 32'hFC5072C4 , 32'hFFFDB991 , 32'hFFFEE69E , 32'h17E18760 , 32'h05BC11E8 , 32'h0001D1A3 , 32'hFFFE451B , 32'h0004D26A , 32'h000151DE , 32'h0000A912 , 32'hFA062728 , 32'h11C234C0 , 32'h0002268F , 32'hFFFB688E , 32'hAC785C80 , 32'hFA40E618 , 32'hFFFF1860 , 32'hFFFF39D2 , 32'h06A3E020 , 32'hFFFE2374 , 32'h00018022 , 32'h0563ABE0 , 32'h06846F00 , 32'hFC961C90 , 32'h04A8BE58 , 32'h00090608 , 32'hFFFA0CEE , 32'hF9A9B6D0 , 32'h0006BF74 , 32'h0002D38A , 32'h0091B39F , 32'h0004C23B , 32'h0003E6D1 , 32'hF7C692A0 , 32'h0001EEE7 , 32'h132A14C0 , 32'h00367CAE , 32'hFFF9254C , 32'h0000D9DD , 32'hFFFE8C5D , 32'hF2C223B0 , 32'hFE85BA74 , 32'hFC833A6C , 32'hE74F9A20 , 32'h000052FD , 32'hE6341E00 , 32'h00068C75 , 32'hFFFC7D30 , 32'h011AB0C0 , 32'hF7BE1960 , 32'hED976C00 , 32'hFFFD099D , 32'h2F7613C0 , 32'hF95E3048 , 32'hF5A8D800 , 32'h3AF82340 , 32'hF5BA90F0 , 32'hF46BA180 , 32'h006F70CD , 32'hC2CC2680 , 32'hFFFE885F , 32'h0003A84B , 32'h00022F36 , 32'h0AA35FD0 , 32'hBB463E00 , 32'hFF637000 , 32'hFE636750 , 32'h04D51A98 , 32'hF3667380 , 32'hFFFB8D75 , 32'h001E818B , 32'hF67D2580 , 32'h00011F4B , 32'hE7272A80 , 32'hFFFD5D79 , 32'hF9D73040 , 32'h01823530 , 32'hFFFF4D1A , 32'h0001AE9F , 32'h0004836A , 32'h0000732A , 32'hFFFE0D43 , 32'h0000A1E8 , 32'h06520CE8 , 32'hD03DB800 , 32'h08316990 , 32'h1F4268C0 , 32'h107DDA60 , 32'hFD507C68 , 32'hFFFD1953 , 32'hFFFDC7A9 , 32'h00019BD8 , 32'hFFFA5BB1 , 32'h00051942 , 32'hFFD6C787 , 32'h0CFED890 , 32'h0AE60C80 , 32'hFFFE3483 , 32'h0004CE30 , 32'h00006EF3 , 32'h00044519 , 32'h157609A0 , 32'h53E90D00 , 32'h00075297 , 32'hFFFE8C42 , 32'hFFFE67E1 , 32'h1628DCA0 , 32'h3AB6F900 , 32'h1A440B80 , 32'h00003D00 , 32'hFFFE5EA2 , 32'h0001DCB1 , 32'hF3F49B90 , 32'hFFD98D29 , 32'h09BD2050 , 32'h00043CAF , 32'h00A3BA30 , 32'h00065A71 , 32'hEF105C20 , 32'h0009DF1D , 32'h09241510 , 32'h00067CE3 , 32'hE500C800 , 32'hF9164F20 , 32'hF761F260 , 32'h1656BF80 , 32'h00046523 , 32'hE756E0A0 , 32'hFEAD31A8 , 32'hFFFE79C3 , 32'hFD19F050 , 32'hFFFF9983 , 32'h022AF98C , 32'hDE645BC0 , 32'h0CBCF740 , 32'h00039C6A , 32'h0000DDF5 , 32'hF8833248 , 32'h0002ACFE , 32'h09661830 , 32'hFFFEFAFF , 32'hFB6B1AB8 , 32'hFFFFF3DA , 32'hFF7583D5 , 32'h00021AF1 , 32'h000921CF , 32'hFFF9167D , 32'hFA6E9180 , 32'hE8903860 , 32'hFFFA00E6 , 32'h0005BBA5 , 32'hFFFE9D2C , 32'h00006655 , 32'hE902E7E0 , 32'hFC4C5DB8 , 32'h1CD970A0 , 32'h15626CC0 , 32'h1B414660 , 32'hFFFC7477 , 32'h0000DFF1 , 32'hFFFEE441 , 32'h00A4639D , 32'h0001D86C , 32'hFFFEA1C8 , 32'hFF47E907 , 32'h0D9F0660 , 32'hFFFEA6FE , 32'hE5D24EA0 , 32'hFF1DBC4C , 32'hF638CEE0 , 32'h165B0D00 , 32'h00016B54 , 32'h0E920040 , 32'hF2CE5E30 , 32'hFE4174E4 , 32'h0000393F , 32'h1BE0BFC0 , 32'h07E19F90 , 32'hF8E1AF40} , 
{32'h076A96E8 , 32'hD9B66D80 , 32'h0000C036 , 32'hFA97AD40 , 32'hFFFC381D , 32'h04BCC848 , 32'h00015F2C , 32'hFFFEA57C , 32'hFFFBDBFA , 32'h000102C3 , 32'hEEA26500 , 32'hE4149280 , 32'hFF28C35F , 32'h00025814 , 32'h0000CC6C , 32'hFADF4868 , 32'h000336DD , 32'h016668BC , 32'hFC2ED4F0 , 32'hFFFDDEB4 , 32'h0006E86C , 32'h06A00010 , 32'hFEB98E98 , 32'hFD488064 , 32'hFDECB69C , 32'h0002C014 , 32'h03D0901C , 32'hFA9A62E8 , 32'hFFFDA3E7 , 32'h282A4F40 , 32'h0004C4C3 , 32'hF1B85D60 , 32'hFFF9B8DF , 32'h0002338A , 32'hFFFFD3A8 , 32'h061104A8 , 32'h224E6700 , 32'h1957EF60 , 32'h0002790B , 32'h15B55D80 , 32'h039A10D0 , 32'h0000C294 , 32'h00017347 , 32'hF31A2090 , 32'h06530B48 , 32'h165DAD20 , 32'h1F3DF200 , 32'h0006C3CB , 32'h0548CB60 , 32'h044405F8 , 32'h047F6558 , 32'h0002AA92 , 32'hFDC2D868 , 32'h163BCF60 , 32'h12D1B960 , 32'hFFFF98CA , 32'h00B34757 , 32'h00005807 , 32'h0005E162 , 32'hF38DE920 , 32'h042A5B68 , 32'hFCFCD65C , 32'h09E766A0 , 32'h0000B518 , 32'hE460D5C0 , 32'hFFFDE5FF , 32'h48292300 , 32'h0083B032 , 32'h00038918 , 32'hE547A7E0 , 32'hF24244D0 , 32'h031CA96C , 32'h0003265C , 32'h00008A80 , 32'hFFFDC597 , 32'h062B0278 , 32'hFC07C7E0 , 32'h00008DE4 , 32'h078DB888 , 32'h0071A893 , 32'h000746A0 , 32'h15F4F4E0 , 32'h01AFBC40 , 32'hFFFE88DA , 32'h089CF890 , 32'h0AA8A5F0 , 32'h09F148C0 , 32'hFFFFE180 , 32'hFFFF1161 , 32'hDD10E980 , 32'h0000D5DE , 32'h1083A600 , 32'h000084C2 , 32'h0D6074A0 , 32'hFDCBE080 , 32'h00021FF5 , 32'h00007DF7 , 32'hFFFFBB35 , 32'hFFFE884C , 32'hFE80B8F8 , 32'h16DC90E0 , 32'hFFFAA441 , 32'hFD80E468 , 32'h247D6640 , 32'h0BE06080 , 32'hFFFEE3F6 , 32'h00048FC1 , 32'hFFFF2F69 , 32'hFEA26C14 , 32'h0B077BC0 , 32'h0002EF0B , 32'hFA65AC58 , 32'h0000F607 , 32'h00053DD9 , 32'h17C10140 , 32'h13B75380 , 32'h048406C0 , 32'h00002CE3 , 32'hF7FE3D60 , 32'h0000E7E0 , 32'h0000F63A , 32'hF9206F40 , 32'hFFFEBBF6 , 32'h000078C8 , 32'hE8AE64A0 , 32'h05683940 , 32'h000413BF , 32'hFFFFAA6E , 32'h0001EB66 , 32'hFFFD7ECD , 32'hFFFF776B , 32'h000B501E , 32'h14434AC0 , 32'h00026857 , 32'h0001DB59 , 32'h26FB1D40 , 32'h0280BED4 , 32'hFFFA530F , 32'hFFFE2B9F , 32'h005215AC , 32'h0001B23A , 32'hFFFFE4AE , 32'hFF226EDA , 32'h190C35E0 , 32'h0C0C45A0 , 32'h01BB802C , 32'hFFFE3571 , 32'h0004773E , 32'h0254DA44 , 32'h0005287A , 32'hFFFDBCAA , 32'hFF0A4457 , 32'h00014A29 , 32'hFFFD143E , 32'hFB017988 , 32'hFFFF07BC , 32'h1F3F52C0 , 32'hFFB72FC2 , 32'h0003DD79 , 32'h0001B2BA , 32'hFFFDF68E , 32'hEA8760A0 , 32'h12EB5080 , 32'h011E1BF4 , 32'h0F3C6250 , 32'h0002C806 , 32'hE3E39780 , 32'h0000FCC0 , 32'hFFFDDC00 , 32'hEA845560 , 32'h133D5A60 , 32'hFEA6E010 , 32'hFFFBB6F7 , 32'h00C96623 , 32'hF64A27E0 , 32'hF73483D0 , 32'h7FFFF800 , 32'hFC84CC14 , 32'hFCF808C8 , 32'h07CF64D0 , 32'h01404720 , 32'h0000F37B , 32'h0001697F , 32'hFFFF9236 , 32'h1943B400 , 32'hE10C0E80 , 32'hFF529DAB , 32'h05F376C8 , 32'hF907D488 , 32'h06D84470 , 32'hFFF930A0 , 32'hF30A6EA0 , 32'hF01E7F10 , 32'hFFFBEE4B , 32'hFAC07C78 , 32'hFFFB36A4 , 32'h0CF84D60 , 32'h18F4D400 , 32'hFFFF91BE , 32'h00040302 , 32'hFFFF0BDA , 32'h0001E418 , 32'h00006297 , 32'h0004394E , 32'h0C2D5B80 , 32'hED5BC6A0 , 32'hF4E7A210 , 32'h13BBFB80 , 32'hFFA8B7DE , 32'h0C8F82C0 , 32'h0001792E , 32'hFFFE7ECF , 32'h00030E92 , 32'h00032B44 , 32'hFFFEEAD4 , 32'hFF46D7C8 , 32'h0059A08A , 32'h09E405C0 , 32'h00033675 , 32'hFFFDC534 , 32'hFFFDE43B , 32'h0000DF5C , 32'h03ADE40C , 32'hD6A09900 , 32'h000488FD , 32'hFFFE2D92 , 32'h0004E9C7 , 32'hC3EB3600 , 32'h2E953CC0 , 32'h0264DA04 , 32'hFFFE104B , 32'h00056EAD , 32'h000146B7 , 32'hFB74CFA8 , 32'h071B47D8 , 32'hBE1CE200 , 32'h000081CC , 32'hFFEA76BB , 32'hFFFA6FF1 , 32'hEAE1DE00 , 32'hFFFAAF4B , 32'h43581900 , 32'h0002BD53 , 32'h2B6AE4C0 , 32'h27B06640 , 32'h045D9300 , 32'h2012C100 , 32'h0003F795 , 32'hF228BFA0 , 32'hFE2A76E4 , 32'h00003058 , 32'hFFE876C1 , 32'hFFFE7BEB , 32'h04116968 , 32'h150F7640 , 32'h12BED0C0 , 32'hFFFCD352 , 32'hFFFA2305 , 32'hE91291C0 , 32'h0004C4FD , 32'h1DD373E0 , 32'h00006829 , 32'hFE818870 , 32'h0004F5B1 , 32'h18BD0B40 , 32'h0001F518 , 32'h000085B5 , 32'hFFFA8397 , 32'h31383840 , 32'hF1BCE390 , 32'hFFFD563B , 32'hFFFE4AC0 , 32'h00004A26 , 32'hFFFDB13B , 32'h10EF1380 , 32'hEFCE02E0 , 32'h40D3B580 , 32'hFD553CFC , 32'h16DB5C80 , 32'hFFFCEE2F , 32'hFFFF3164 , 32'h00077F38 , 32'h04D49D20 , 32'hFFFE66E2 , 32'h000156CA , 32'h0CF33140 , 32'hFAA56160 , 32'h0001CF39 , 32'hFA71C000 , 32'h042106F0 , 32'h0731BCE0 , 32'h09458F40 , 32'h000285FB , 32'h05E09788 , 32'h025A9AEC , 32'hFF291274 , 32'hFFFD43EF , 32'hF94C08D0 , 32'hEFEE0940 , 32'h1E4A2700} , 
{32'h10367E80 , 32'h2F0F02C0 , 32'hFFFADAF7 , 32'hFC6D69A8 , 32'hFFF6D2BE , 32'h00EB3EB9 , 32'hFFFCCCB0 , 32'hFFFDC4B4 , 32'hFFFAF2E0 , 32'hFFFF1BF5 , 32'hFBD880D0 , 32'hFAB359A0 , 32'h059476A8 , 32'hFFFA75B8 , 32'hFFFC87B4 , 32'h1313D1C0 , 32'h00005B30 , 32'hD0F020C0 , 32'hEAB2EAC0 , 32'hFFFFC143 , 32'h00009481 , 32'h00768109 , 32'h1057FAA0 , 32'hF76A2AB0 , 32'h09BFD590 , 32'h000104C5 , 32'hFCADD024 , 32'hFB31E958 , 32'hFFFBD9BF , 32'h17296A20 , 32'h0000A483 , 32'hE24815C0 , 32'hFFFB166E , 32'h00021306 , 32'h000069BC , 32'h0FE964A0 , 32'hE4D46640 , 32'hF37EB5C0 , 32'h0002C08B , 32'h1A814B60 , 32'h0D2A35C0 , 32'h00034A06 , 32'h00038EB6 , 32'h04FEF630 , 32'h0933B840 , 32'h1D4DEDE0 , 32'hE5937880 , 32'h0001C747 , 32'hFEDC8994 , 32'h3CA38B00 , 32'hFF626308 , 32'h000A7253 , 32'hFB025C48 , 32'h02C4F4B8 , 32'hF2E7A560 , 32'hFFFE8355 , 32'hFF1BE585 , 32'h000250EB , 32'hFFFF4741 , 32'h02115108 , 32'hFCA9C508 , 32'h07ABC0C8 , 32'hF7C44110 , 32'h0001F73F , 32'hB6309C00 , 32'h0002F931 , 32'hCA3C01C0 , 32'hFD9076C4 , 32'h000247F7 , 32'hE5A2E360 , 32'h01C1032C , 32'h1E510140 , 32'hFFFD9DBF , 32'hFFF9E5F8 , 32'hFFFE3D85 , 32'h099EF4F0 , 32'h08028280 , 32'h00000078 , 32'h24F6A580 , 32'hFFCE02B3 , 32'h00025643 , 32'h189A3CE0 , 32'hF9659940 , 32'h00046653 , 32'hFE7FE3C8 , 32'hFF5CC6E3 , 32'h004D3D9B , 32'h00011F4E , 32'hFFFE2D5A , 32'hFFB3049E , 32'h000067CB , 32'h0E936510 , 32'hFFFDED62 , 32'hE093F340 , 32'hFD5BCF9C , 32'hFFFB0598 , 32'hFFFF3C10 , 32'h00027D85 , 32'h00053829 , 32'h111C1B40 , 32'h0975C4C0 , 32'h00073D5C , 32'hF5CB4560 , 32'hEA6FFB40 , 32'h0B11F350 , 32'hFFFEF45C , 32'h01A287AC , 32'h0001DF36 , 32'h0786C4E8 , 32'h31499740 , 32'hFFF7A15B , 32'h0B0827B0 , 32'hFFF87795 , 32'hFFFDBC12 , 32'hEFD26F80 , 32'h0B505800 , 32'hFCD9CC1C , 32'hFFFF8C9E , 32'hD9FC3240 , 32'h00013C2E , 32'h0004A8D7 , 32'hFBE63460 , 32'h00045EA2 , 32'h00021018 , 32'hE4E55140 , 32'h0BAEC8F0 , 32'h0001F6D8 , 32'hFFFD5D31 , 32'hFFFFBBF8 , 32'hFFFCDBD8 , 32'hFFFBE64C , 32'h0FADDEB0 , 32'h020F7CCC , 32'hFFFCEE07 , 32'hFFFE126C , 32'h06EEB7C8 , 32'h12BE78A0 , 32'h00083353 , 32'hFFFF20F2 , 32'h07D026D8 , 32'hFFF82A92 , 32'hFFFA1953 , 32'hFB40C4D0 , 32'hFA189F60 , 32'h035F22C8 , 32'hFB356C90 , 32'hFFFE58A8 , 32'h0002B626 , 32'hFFF2BDFF , 32'hFFFDC62B , 32'h000232AF , 32'h01FDF1E4 , 32'hFFFEB31F , 32'h00018C7E , 32'h037A46F4 , 32'hFFFE5CC9 , 32'h09594E00 , 32'h025CBB1C , 32'h0003074A , 32'hFFFF72F1 , 32'hFFFD09F2 , 32'h34CB6E80 , 32'h05237A90 , 32'hFA48E138 , 32'h052458A0 , 32'hFFFFA084 , 32'hFC543A98 , 32'hFFFEE69D , 32'hFFFF629C , 32'h080EDDA0 , 32'h01799A78 , 32'h04E72CC0 , 32'h00027018 , 32'hD5EE79C0 , 32'h03673F10 , 32'h074D7E20 , 32'h327F9BC0 , 32'hF6121840 , 32'h547CD280 , 32'h00F257FD , 32'hF4D84930 , 32'hFFFC6AC8 , 32'h00040227 , 32'h0000C6EF , 32'hFE08CD7C , 32'h16E3ED60 , 32'hFBF2F918 , 32'h00363084 , 32'hFD9BC410 , 32'hFA8AFA90 , 32'hFFF824A3 , 32'hF1C24610 , 32'hFF467555 , 32'h00051F9B , 32'h1288B440 , 32'h0002D3C8 , 32'h1BCF4EE0 , 32'hFF259579 , 32'h00032095 , 32'h000233EB , 32'hFFFEFA9E , 32'h00029E4F , 32'hFFFFCA49 , 32'h0000ECA1 , 32'hFBB0CDE0 , 32'hF0A09100 , 32'h14701380 , 32'hE85089A0 , 32'hF705EE00 , 32'hFCD7F0EC , 32'h0003EFE3 , 32'h000373CD , 32'h00030069 , 32'h000312EB , 32'hFFFC6BAF , 32'h042D76D0 , 32'h17311260 , 32'hD1CC14C0 , 32'hFFFE2EA1 , 32'hFFFFAC2D , 32'h0000A39F , 32'h0000088D , 32'h16682FA0 , 32'h24C5BA40 , 32'h0001A332 , 32'h000381A7 , 32'h0002D344 , 32'hDE7383C0 , 32'h1BB686E0 , 32'hD0436080 , 32'hFFFDDC64 , 32'h00027847 , 32'h00000FA6 , 32'hFA4E2BA8 , 32'h03A06078 , 32'hFFB68C88 , 32'hFFFD8589 , 32'h00317ECD , 32'hFFFBCFD2 , 32'hFB491FD8 , 32'h0001A41D , 32'hD966A900 , 32'h000531B3 , 32'hD0F4AA00 , 32'h0031374B , 32'h21E4C600 , 32'hC416B1C0 , 32'h00050BD9 , 32'h0EC75470 , 32'h050F4868 , 32'h0002CC60 , 32'hF029D9F0 , 32'hFFFC8FD9 , 32'hFF4741AE , 32'h1AF04040 , 32'h214623C0 , 32'h0002BA55 , 32'hFFFBEBAC , 32'h12397660 , 32'h00032B01 , 32'hEE116A20 , 32'hFFFFAAB7 , 32'hFC771B60 , 32'hFFFCD7CD , 32'hF9925AD0 , 32'h00014FC7 , 32'h0002353A , 32'hFFFD8E64 , 32'hF9355E90 , 32'hFD5EFCC4 , 32'hFFFE8FB8 , 32'hFFFCB646 , 32'hFFFEFE9D , 32'h0000F4E4 , 32'hF3E368F0 , 32'hF30C44F0 , 32'h090CDB30 , 32'h0CEF3AA0 , 32'h041E8078 , 32'hFFFE18D4 , 32'hFFFD363B , 32'hFFFE98D8 , 32'hFE8F8CAC , 32'h000194C9 , 32'h00013AD8 , 32'hFDE63E54 , 32'h36DE4440 , 32'hFFFAB997 , 32'hFF7ABF9E , 32'h00843F05 , 32'h071C8AA0 , 32'h1824A960 , 32'h000117AF , 32'hE69EBD00 , 32'h2AFC7BC0 , 32'hF8F08150 , 32'hFFFE1248 , 32'hE26CECA0 , 32'h2853F540 , 32'h1F2997E0} , 
{32'hF311DA00 , 32'h2A9A1480 , 32'h00028B66 , 32'hDBE5B580 , 32'h0001F58A , 32'hFC909714 , 32'hFFF70AB2 , 32'h0003391D , 32'h0000C879 , 32'hFFFFB6A5 , 32'h0F893B50 , 32'h310509C0 , 32'hFB880FD8 , 32'hFFFDABB5 , 32'h000254D5 , 32'hE2100160 , 32'hFFF9D400 , 32'h389984C0 , 32'h03DA54FC , 32'hFFFBBBE1 , 32'h0001B120 , 32'h04558078 , 32'hECA233E0 , 32'hF2B96690 , 32'hFCE2D4F8 , 32'hFFFC38E8 , 32'h059E3840 , 32'h072865E8 , 32'h0002615E , 32'h0D85C900 , 32'h0001E045 , 32'hFAD0CB08 , 32'h0004FC80 , 32'h00018D46 , 32'hFFFA86E8 , 32'hF9D624F0 , 32'h230FF6C0 , 32'hE1AF40A0 , 32'hFFFD3EC3 , 32'hE508A360 , 32'hFF5513D3 , 32'h00022EC7 , 32'h0004C535 , 32'hFED886C4 , 32'hE28794C0 , 32'hD1116C40 , 32'h1CBE2720 , 32'h0001C9B8 , 32'hF31A0620 , 32'hEC188C80 , 32'h01FB9E04 , 32'hFFFFD47B , 32'h063625C0 , 32'h1D86D3A0 , 32'h10B60E80 , 32'h00039F2A , 32'hFED6E4E8 , 32'hFFFB1E86 , 32'h00021C7A , 32'hF5CF6BE0 , 32'h041472F0 , 32'hF06D3720 , 32'h20074840 , 32'hFFFB432E , 32'hF5BA2CC0 , 32'hFFFEB692 , 32'hCB016280 , 32'hFFC33158 , 32'h00048D24 , 32'h01AEDF14 , 32'h0D80E280 , 32'h0C571D20 , 32'h00021F3B , 32'h0002FB9A , 32'hFFFE999A , 32'h0C167390 , 32'hFF399471 , 32'h0000C5F9 , 32'h0196B680 , 32'h00BC6ED1 , 32'hFFFD3645 , 32'hCE5BC980 , 32'hF9F7E418 , 32'h00046EDC , 32'h0213604C , 32'hE9644BC0 , 32'h00425A7B , 32'hFFFA3D37 , 32'h00018F5F , 32'hFECCCB1C , 32'hFFFEB133 , 32'h1019EC00 , 32'hFFFC0A97 , 32'h07B537D8 , 32'hFFB70F54 , 32'h00014A84 , 32'hFFFCED40 , 32'hFFFD2254 , 32'h000220CF , 32'hEDB6AF20 , 32'h00237F30 , 32'hFFFF370D , 32'hC7330EC0 , 32'hE0F9E320 , 32'h0CD3C750 , 32'hFFFE7F82 , 32'h00A2EB8E , 32'h00024D9D , 32'hF7F10950 , 32'hF7FD45F0 , 32'hFFFF366C , 32'h02894424 , 32'h00014AA6 , 32'hFFFF24D9 , 32'h12F3C500 , 32'h0C4FFE20 , 32'hFE43E11C , 32'hFFFD7233 , 32'h045054C0 , 32'hFFFF4530 , 32'hFFF921AA , 32'hFC9C2294 , 32'hFFFF5B7A , 32'hFFFD5DC0 , 32'hF54405E0 , 32'h00AE462D , 32'h0002706B , 32'hFFFDB9A1 , 32'hFFFFDEAA , 32'h0005B934 , 32'hFFFE1E81 , 32'hFC5AEBC8 , 32'h0994ACD0 , 32'h00011D38 , 32'hFFFDABEB , 32'h2EEAFF00 , 32'hF3F95A20 , 32'hFFFAB318 , 32'hFFFF408F , 32'h18F9E940 , 32'h000518D2 , 32'hFFFE5CAD , 32'h04558E50 , 32'h05C1EFF0 , 32'h0BDF6DC0 , 32'h03B4911C , 32'hFFF9C8B4 , 32'h0000F79B , 32'h013FF8D4 , 32'h0000FCFD , 32'h0006B44B , 32'hFD83E9A0 , 32'h0002BC26 , 32'h00046DA2 , 32'hE0615D60 , 32'hFFFFB2EF , 32'h00CBA06E , 32'h0383CAA4 , 32'hFFFFC4B9 , 32'h00020E3B , 32'h0000C35C , 32'hE49C7EA0 , 32'h0E319210 , 32'hF6E36560 , 32'hED0EBA40 , 32'hFFFC70AF , 32'hE6D54C60 , 32'hFFFC9C2F , 32'hFFF96F13 , 32'h2B90D840 , 32'h008D0F79 , 32'h099C30F0 , 32'h00025FBE , 32'h02B22B68 , 32'hFF28A8D6 , 32'hFD3F6D64 , 32'h1185E220 , 32'hF9B4EA40 , 32'hF6EE6930 , 32'h064359C8 , 32'hFCB755D8 , 32'hFFFF1D51 , 32'hFFFF569C , 32'h00018EEA , 32'hF3103F50 , 32'hDA868D00 , 32'h00DEE942 , 32'hFDF2BCF0 , 32'hF7026490 , 32'h07F302D0 , 32'hFFFDBFB8 , 32'hF77BD8C0 , 32'h17619080 , 32'hFFFCC162 , 32'hF12CD3E0 , 32'hFFFBD211 , 32'hFA7EE040 , 32'hDA19C2C0 , 32'h00003CA0 , 32'h00010D2C , 32'hFFFF79A3 , 32'hFFFD345D , 32'hFFFF9F26 , 32'h00036627 , 32'hF3B14560 , 32'hDB834C40 , 32'h0BEFAB20 , 32'hFCCC2030 , 32'hF0BBF680 , 32'h0AB27AA0 , 32'hFFFCF7E5 , 32'h0000FCF2 , 32'h0004166B , 32'h00029994 , 32'hFFF89E2D , 32'hFD72EF34 , 32'hF45C6400 , 32'hFC3A304C , 32'h00044B07 , 32'h0004A3F9 , 32'hFFFF2FD0 , 32'hFFFE10B0 , 32'h09432160 , 32'h2C6C0980 , 32'h00044AE3 , 32'hFFFFBA5E , 32'h00004700 , 32'hBE518880 , 32'hAD6A7E80 , 32'h278603C0 , 32'hFFFB40D0 , 32'h00012C06 , 32'hFFFC2F92 , 32'hFD006EC0 , 32'h04E965E8 , 32'h2481FD80 , 32'hFFFF27BE , 32'h00EE2BF7 , 32'hFFF9F8BD , 32'h3E097A80 , 32'h00000B0F , 32'h38A9CCC0 , 32'h000258A7 , 32'h19CA1400 , 32'hE6250080 , 32'hF89CFE58 , 32'hE7C1E420 , 32'h0003EB99 , 32'hF9161288 , 32'h00EDF059 , 32'h000428E7 , 32'h0A949EA0 , 32'h00047B6F , 32'h09B40030 , 32'h2FEEA880 , 32'h07FB68B8 , 32'hFFFFCEBA , 32'h0002992F , 32'hF7317740 , 32'h0004A596 , 32'hEBBDB340 , 32'h0001804B , 32'h0091F10B , 32'h00010016 , 32'h06BA7720 , 32'hFFFD950B , 32'hFFFE4EB8 , 32'hFFFF5929 , 32'h12CEBBC0 , 32'h03E8524C , 32'hFFFBFFE4 , 32'h00009231 , 32'h000043F1 , 32'h000541E6 , 32'h0D80B780 , 32'hF432E580 , 32'hFF357B6C , 32'h012BB2C4 , 32'hF7433B60 , 32'h0001C880 , 32'h0000E1B0 , 32'h0000E2C3 , 32'h05E71CB0 , 32'h0000026E , 32'hFFFF0210 , 32'hF93F62C0 , 32'h414A5E80 , 32'hFFFF8483 , 32'h07588B20 , 32'h09DDA7E0 , 32'h00B32483 , 32'h0639BCC8 , 32'h00018E8C , 32'h10A550A0 , 32'h297C5A80 , 32'hFE5E8DFC , 32'h0001E8DD , 32'hF6348AF0 , 32'hF8B48738 , 32'h16C87840} , 
{32'hED7FC4C0 , 32'h1E2E5BE0 , 32'h00058165 , 32'h113A2C80 , 32'h0001C058 , 32'hF881F328 , 32'h0003F4C0 , 32'h0001A6DD , 32'h000072F7 , 32'h0003ED72 , 32'hEF558B80 , 32'h0EF09DA0 , 32'h028404AC , 32'h0001E283 , 32'hFFFC82B3 , 32'h49BC4500 , 32'h000419D1 , 32'h1A836D20 , 32'hF63E0ED0 , 32'hFFFC41C4 , 32'hFFFC9E57 , 32'h06F55C30 , 32'h275A3B80 , 32'h100DAFE0 , 32'hFAE1A6B8 , 32'h0002F36E , 32'h06B15460 , 32'h026B95F0 , 32'h0006CA28 , 32'h1FE754A0 , 32'hFFFCCECF , 32'h11935AE0 , 32'h0001354E , 32'h00015A51 , 32'hFFFC6F57 , 32'hE97BD540 , 32'hF739C240 , 32'hF7D97480 , 32'hFFF97067 , 32'h2D2164C0 , 32'h1C6B9A20 , 32'h0002A8F6 , 32'hFFFC2562 , 32'h01E41A00 , 32'h15B79F00 , 32'h0F757FB0 , 32'h1D0DE360 , 32'hFFFC35CC , 32'hE8C8BD40 , 32'hDD5C2680 , 32'h00979BA6 , 32'hFFFF7657 , 32'h0CBE9A40 , 32'h0A253340 , 32'hFB582A70 , 32'hFFFA3C6D , 32'hFFF705D7 , 32'hFFFEB346 , 32'h000212CC , 32'h0A703580 , 32'h00FCDBAD , 32'hFEDE6B34 , 32'h01408DC8 , 32'h00030EF9 , 32'hEBADCC80 , 32'hFFFC44AC , 32'h231264C0 , 32'hFA1B4470 , 32'h0001EC96 , 32'h07101210 , 32'h0D204C10 , 32'hF27C74E0 , 32'h00031FEB , 32'hFFF8B2B7 , 32'hFFFE37C4 , 32'h095A9830 , 32'hFABD6898 , 32'h00031A3D , 32'h2A35DD40 , 32'hFC7F0AC8 , 32'h0000352E , 32'hE6551240 , 32'hF94A5E90 , 32'hFFFE0809 , 32'h0405E500 , 32'h05132608 , 32'h0B07E920 , 32'hFFFC8899 , 32'h00025AE5 , 32'hE9D5DA80 , 32'h0006B616 , 32'hE75B7740 , 32'h000181C8 , 32'h0BB6C320 , 32'h003AE20A , 32'hFFFE1F59 , 32'hFFFDD23E , 32'h000007BC , 32'h000520D5 , 32'h0B4182F0 , 32'h0662C390 , 32'hFFFE7A96 , 32'hF9923AA0 , 32'h1DD1CFA0 , 32'hF52A24A0 , 32'h00002696 , 32'h000B0AAA , 32'h000228B2 , 32'h0D01E450 , 32'h012A3BCC , 32'hFFFD175A , 32'h0315B908 , 32'h00032A64 , 32'h000386A0 , 32'h0BE42340 , 32'h083C1D50 , 32'hF9D297B8 , 32'hFFFC8783 , 32'hF02DEC40 , 32'h00033A27 , 32'hFFFB066D , 32'h06A4F7C0 , 32'h00004627 , 32'hFFFED0BD , 32'h1ED3DF80 , 32'h0854A870 , 32'h0004E559 , 32'hFFFED514 , 32'h00025791 , 32'hFFFCF85E , 32'h0004396C , 32'h1775BA00 , 32'h044DF7A8 , 32'h000146FA , 32'h0003D6B9 , 32'hFE047FDC , 32'h0E3D9BF0 , 32'h000070FD , 32'hFFFC2C6B , 32'h1100F880 , 32'hFFFF4133 , 32'h0001B6CB , 32'h00D6FA9F , 32'hE05C4540 , 32'h036AD8B4 , 32'h0009A120 , 32'h0005AB7F , 32'h0004219A , 32'hF91E22D0 , 32'hFFFE7A73 , 32'hFFFD091F , 32'h078B46F8 , 32'h0004B4F0 , 32'h0003A08D , 32'hFE125430 , 32'h00063469 , 32'h09E06040 , 32'h02BC8490 , 32'h00026C18 , 32'h00035965 , 32'hFFFC7357 , 32'h12196B40 , 32'hFE5D1B54 , 32'h0A04C8C0 , 32'hFF9E23EB , 32'h0001E0D7 , 32'h235543C0 , 32'h00015F22 , 32'h0002B54F , 32'hF195E4C0 , 32'h05D76B50 , 32'hF06E6450 , 32'h00007D5B , 32'h0D50D770 , 32'hF381B8C0 , 32'h0C2B9480 , 32'hDD98EE00 , 32'hFEA56DB0 , 32'hF2073F00 , 32'hFDD9882C , 32'hE93194E0 , 32'h000129A2 , 32'h00021940 , 32'h00019BAB , 32'h0C68E800 , 32'h8239DF80 , 32'hFC365644 , 32'hFE98BB20 , 32'h178EB880 , 32'hEA6A6880 , 32'hFFFA3E6D , 32'h19F8FEE0 , 32'hFEAE3D2C , 32'h000418DC , 32'h08FE0990 , 32'hFFFE2216 , 32'h0C624E00 , 32'hF9A599E8 , 32'h0001F446 , 32'hFFFE304A , 32'h00023D3C , 32'h0008168A , 32'hFFFFF627 , 32'h000047BF , 32'hF6823810 , 32'h187EB880 , 32'hFA3C7B20 , 32'h04BEA800 , 32'h09956FF0 , 32'h0BDC6300 , 32'hFFFE33AD , 32'hFFFB815D , 32'h000768F3 , 32'h000002CE , 32'hFFFC6423 , 32'h092E6970 , 32'h1B5320C0 , 32'h0463E940 , 32'h00007C16 , 32'h0000CE3A , 32'hFFFE5AB6 , 32'h0004AEA5 , 32'h01539D40 , 32'hD593D8C0 , 32'h0001B30F , 32'hFFFD77E4 , 32'hFFFFDB19 , 32'hCB87EBC0 , 32'hDE8E8740 , 32'hD42C0200 , 32'hFFFD53F8 , 32'hFFFF615B , 32'h0000CB88 , 32'hFBE7E1C0 , 32'hFE756214 , 32'hF76BB6F0 , 32'hFFFE7EBD , 32'hFC754D70 , 32'h0005127D , 32'h060845D8 , 32'h0003032C , 32'hF79816F0 , 32'hFFFD00D5 , 32'hC9F74240 , 32'hF4176900 , 32'hDE1663C0 , 32'hD9E00FC0 , 32'h00001451 , 32'h067F38D8 , 32'hFFA85D8A , 32'hFFF64534 , 32'hF3C3B060 , 32'h0003A05B , 32'h02644518 , 32'hEFA163E0 , 32'h045E31F8 , 32'h00006349 , 32'hFFFD9E46 , 32'hF338B770 , 32'hFFF92175 , 32'h006A8E96 , 32'hFFFBC520 , 32'h0161EF3C , 32'hFFFD76FB , 32'h007FC007 , 32'h00019DA1 , 32'h000B55A2 , 32'hFFFE3210 , 32'hF94D6D70 , 32'hE01AA580 , 32'hFFFDD59B , 32'hFFFD85BA , 32'hFFFF908E , 32'h0002BFFB , 32'hF735ABC0 , 32'h1FDCE240 , 32'hEE4A8E00 , 32'h30F38340 , 32'h24C5F700 , 32'hFFFDED84 , 32'h0004A476 , 32'h0004654F , 32'hF8A4A2F0 , 32'hFFFB19E4 , 32'hFFFD7864 , 32'h011A0618 , 32'hFF323085 , 32'h000453D3 , 32'h44D25680 , 32'hFFC16F8F , 32'hF5F21A70 , 32'h084C5BF0 , 32'h00012CBE , 32'h0586DDE0 , 32'h1D3E2720 , 32'h063B0980 , 32'hFFFF2DFD , 32'h381CF840 , 32'hE8FA5B60 , 32'hFFE3BED7} , 
{32'h1DEF22A0 , 32'h06C2A838 , 32'h00014969 , 32'hF5C1C9A0 , 32'h00018DC7 , 32'hF648CEC0 , 32'h0004F670 , 32'hFFFFB959 , 32'h0000174B , 32'h00073F4B , 32'h1A48DBC0 , 32'hD4AAAE80 , 32'hEC0956A0 , 32'h00000220 , 32'hFFFA7FF0 , 32'h04E2C9B8 , 32'hFFFB8D84 , 32'h08437DB0 , 32'hFCC337DC , 32'hFFFF99C1 , 32'h0001DE4B , 32'h0024FFF1 , 32'hD7CDBE40 , 32'h0637FD18 , 32'h0D32C5D0 , 32'h0000E86C , 32'hFEF6BE48 , 32'hF66E07C0 , 32'h00037366 , 32'hF2DCA5C0 , 32'hFFFDC431 , 32'hE4C7FF80 , 32'h0001CB0E , 32'h0001A3BE , 32'hFFFCD9AA , 32'h238A4280 , 32'hE7478780 , 32'hE24EBD40 , 32'h00002D72 , 32'hE7D3AE60 , 32'hE5D279A0 , 32'hFFFFDD70 , 32'h0001D58C , 32'hF25139F0 , 32'hDFB21180 , 32'hE8636E20 , 32'hF0BCA550 , 32'hFFFF34FA , 32'h01E9E9CC , 32'h2B11D580 , 32'hFE5E8338 , 32'hFFFA3EA1 , 32'hF7C8D450 , 32'hEB6D52A0 , 32'h03CD8184 , 32'h000269F9 , 32'hFEFA0874 , 32'h000122A3 , 32'hFFFDBA2B , 32'h0BFEF3E0 , 32'h03FE7C3C , 32'hEDDB66C0 , 32'h2599D2C0 , 32'h00051C93 , 32'h8E403200 , 32'h000216B3 , 32'hFDC4FF64 , 32'hFDD067D0 , 32'h00026EB4 , 32'hFD4072B0 , 32'h2A060540 , 32'hFDF8428C , 32'hFFFCB5A2 , 32'hFFFF3303 , 32'hFFFD8429 , 32'hEF60F260 , 32'hF72DCA60 , 32'h00022F00 , 32'hF4FABFA0 , 32'hFE516F04 , 32'h0000C651 , 32'hD03BBE00 , 32'h06C8F368 , 32'hFFFF7348 , 32'hFA63B6A0 , 32'hF8FA5D20 , 32'h03A94F08 , 32'h0000D20B , 32'hFFFFF756 , 32'h26A57B00 , 32'h00049B00 , 32'h0D6E6170 , 32'h00057F41 , 32'hFD0014D8 , 32'h03361624 , 32'h000208C9 , 32'hFFFBFC65 , 32'hFFFBC13E , 32'h0004C264 , 32'h2773E480 , 32'hFCA88DF8 , 32'hFFFD5A11 , 32'h0D4A0F80 , 32'h21A42D40 , 32'h0186712C , 32'hFFF920D9 , 32'h0078B499 , 32'h00020717 , 32'h06D75580 , 32'hF8CB4AB0 , 32'hFFFEB7F4 , 32'h09279A00 , 32'hFFFFC443 , 32'h000212A5 , 32'hFC4611B4 , 32'h083A38B0 , 32'h03F719F8 , 32'hFFFCAACC , 32'hE1D22020 , 32'hFFF9FAA7 , 32'hFFFD4A55 , 32'h07DB38B0 , 32'h0001B981 , 32'h00042CCA , 32'hAD1B3380 , 32'hFED74068 , 32'h0002B8AC , 32'h00023C2E , 32'h00022534 , 32'hFFFEA784 , 32'h00028EF5 , 32'h023901E0 , 32'hEB3371C0 , 32'hFFFFDC14 , 32'h00043F01 , 32'h0C37E470 , 32'hE933C3A0 , 32'h000346B2 , 32'hFFFF6790 , 32'h0A49C530 , 32'h000500AB , 32'h0003D2D9 , 32'hFEC6FD78 , 32'h001C0E82 , 32'h00AA8524 , 32'hFF4C5734 , 32'h0007587D , 32'h00012750 , 32'h008EA806 , 32'hFFFE5031 , 32'h00004DE3 , 32'h0651DF38 , 32'h0003D299 , 32'h00080A23 , 32'hEE5E34A0 , 32'hFFFBF28F , 32'h029AC0F8 , 32'h00B26514 , 32'hFFFFBFCA , 32'hFFFBECE4 , 32'h0000634B , 32'h045AA058 , 32'h088B2150 , 32'h07D61420 , 32'hF7F349C0 , 32'h0001B405 , 32'hFEB05268 , 32'h0002689B , 32'h0003C3E6 , 32'hF5E2D970 , 32'h066FDA18 , 32'h0A274030 , 32'hFFFDA6A7 , 32'hE7C90440 , 32'h06150788 , 32'hF031DFD0 , 32'hEBA4F5C0 , 32'hF8441408 , 32'hFA1FF548 , 32'hFBA89C08 , 32'h0107AE74 , 32'hFFFEBB2C , 32'h0007CABD , 32'h00040E53 , 32'h12C4A1A0 , 32'hEDC27700 , 32'h0A2A2E80 , 32'hFBDC4CD0 , 32'hFD45CEF0 , 32'hFC023208 , 32'h00062A16 , 32'hE74481E0 , 32'hED913C00 , 32'hFFFF0C2C , 32'hEFA5FD60 , 32'h00008D3F , 32'hED1C8DC0 , 32'hD768A900 , 32'h000479C3 , 32'h00030E6C , 32'h00099A50 , 32'h0000D507 , 32'hFFF9CA20 , 32'h00007918 , 32'hF74AF000 , 32'h09EEA030 , 32'h3909F4C0 , 32'h097908A0 , 32'hEDD03EE0 , 32'hE96E2CA0 , 32'h000211F7 , 32'hFFFF3EB5 , 32'h00034935 , 32'h000222EE , 32'h0007CCDF , 32'hFAF72778 , 32'h0F4BCDC0 , 32'h1AA98F60 , 32'h0000B97C , 32'h0000F5EB , 32'h00000C5A , 32'hFFFFC8EE , 32'h05D016C8 , 32'hE1F90E80 , 32'hFFFDBD48 , 32'hFFFDDF44 , 32'h00037E82 , 32'hF8098218 , 32'h225D0BC0 , 32'h351A6500 , 32'h00011F44 , 32'h000231D9 , 32'h0005914E , 32'hFF696FC0 , 32'hFDC66FA0 , 32'hF122FF70 , 32'h00064587 , 32'hFF7241C1 , 32'h0001ABCF , 32'hF68F9500 , 32'h0000A415 , 32'hE474FB00 , 32'hFFFFEF79 , 32'hFBA48058 , 32'hF6D2CEE0 , 32'hB5DCAB00 , 32'h241EE340 , 32'hFFFEEDE7 , 32'h16CA58A0 , 32'h0233FA54 , 32'h0003F960 , 32'hFB9E08C0 , 32'hFFFBB8BD , 32'hFC88D148 , 32'hE2BBCC40 , 32'hE901C540 , 32'h00020654 , 32'h0003C0B9 , 32'hF72BDDE0 , 32'h00059D34 , 32'h0BA67B80 , 32'hFFFA5E3F , 32'hFD68B6C4 , 32'hFFFE61DE , 32'hDF8ABC40 , 32'h0004C0ED , 32'h0000F002 , 32'h00021C1D , 32'h26DC7800 , 32'h0F99E860 , 32'h000159B3 , 32'hFFFB7CFB , 32'h00022BB0 , 32'hFFFEB054 , 32'h04006228 , 32'h12585260 , 32'hED2E3760 , 32'hE85A4B00 , 32'h1B8BDD00 , 32'h000072CC , 32'h000609C2 , 32'hFFFEA372 , 32'hF931D010 , 32'h000371F3 , 32'h000166BE , 32'hFED8FEB4 , 32'hFB808258 , 32'h0004D33F , 32'h2609A800 , 32'hF8D28CF0 , 32'h0017CC9F , 32'hE7B163E0 , 32'hFFFD17F8 , 32'h030646B4 , 32'hFA168C98 , 32'h05BE0820 , 32'h00031E9C , 32'h1E8E04E0 , 32'hEBCC9080 , 32'hEDCAB120} , 
{32'h128FDAE0 , 32'h13A39D40 , 32'hFFFCF074 , 32'hEB09D640 , 32'hFFFE7052 , 32'h049325A8 , 32'h0002D795 , 32'hFFFF1E4E , 32'hFFFC14D0 , 32'h00075882 , 32'h03596158 , 32'hC9F68680 , 32'hF09D9160 , 32'hFFFE430E , 32'hFFFDA4B3 , 32'h3B5CF6C0 , 32'h0002F55B , 32'h073F5478 , 32'h0B454BD0 , 32'hFFFE4BA1 , 32'hFFFEEC9C , 32'h004C00E9 , 32'h1F786660 , 32'h0FCD4180 , 32'hFDEDC614 , 32'h00063302 , 32'hFD71DF90 , 32'h00213689 , 32'hFFFCC19F , 32'hC7886A80 , 32'h00047E61 , 32'h02E3B4C4 , 32'h00087873 , 32'h000256EB , 32'hFFFC5D12 , 32'h39CBD4C0 , 32'h22223440 , 32'hDCAA8E40 , 32'hFFFC3687 , 32'h0E85FA00 , 32'h002DACE7 , 32'hFFFC5860 , 32'hFFFB69A2 , 32'h04A57BF0 , 32'hD4C4AAC0 , 32'hFB57F9A8 , 32'hFDEF9764 , 32'hFFFE0F1D , 32'h18DAF7E0 , 32'h01C1FABC , 32'hFEA74370 , 32'h0000F7B5 , 32'hFFC59DD3 , 32'h2CA3EA00 , 32'h05E22CC8 , 32'h00029752 , 32'h00A7C43E , 32'hFFFBF1C0 , 32'hFFFED1FB , 32'h03496D38 , 32'hFCAB35E8 , 32'h00555ADE , 32'hE66BF220 , 32'h000084AB , 32'h0867E6C0 , 32'h00029972 , 32'hE050E200 , 32'h05DD6430 , 32'hFFFE965D , 32'hC8C32A40 , 32'h0D1BABC0 , 32'h0BEC9EC0 , 32'h00011DCA , 32'h00058445 , 32'hFFFE97D5 , 32'hFF13155B , 32'h0A794A90 , 32'h00039D58 , 32'hF2F3A3B0 , 32'hFD808728 , 32'hFFFE14F9 , 32'h2252E7C0 , 32'h06A14E40 , 32'hFFFC0C3E , 32'h0D73B080 , 32'h18E891E0 , 32'h007B44EB , 32'h0001AD2E , 32'hFFFF03DF , 32'h2AAB6B80 , 32'h00006A8B , 32'hE1745880 , 32'h0003422D , 32'h147CF440 , 32'h0051B875 , 32'h00058BD5 , 32'h0004858E , 32'hFFFE6164 , 32'h0002B82F , 32'h105A3260 , 32'h05D80818 , 32'hFFFC097D , 32'h0963CFF0 , 32'hEDC1FC40 , 32'h0312B9F8 , 32'h00017AA7 , 32'hFFFE89FE , 32'hFFFAAAB7 , 32'hF84C4800 , 32'hD1607700 , 32'h00017666 , 32'h1E13C560 , 32'hFFFAD196 , 32'hFFFD7518 , 32'h1708AB20 , 32'h0D0EFB30 , 32'h021B0D80 , 32'hFFFA079B , 32'h0F2CDCF0 , 32'hFFFBD7FB , 32'h000247DB , 32'hFFA5A758 , 32'hFFFE6FAF , 32'h00053987 , 32'h260E4EC0 , 32'hD34352C0 , 32'h000190A6 , 32'hFFF89C9B , 32'h0005354B , 32'h00036616 , 32'h0000425D , 32'h06E71E18 , 32'h0E17E5B0 , 32'h00021EFB , 32'hFFFC8254 , 32'h3343DD40 , 32'h0095F4BF , 32'hFFFC7ED7 , 32'h00006A75 , 32'h027D9098 , 32'h0004AA99 , 32'hFFFD8B6C , 32'hFEBB7240 , 32'h0A729B20 , 32'hFF0318C8 , 32'hFA8BA9A0 , 32'hFFFF10D7 , 32'hFFFC4986 , 32'hFDC2A270 , 32'hFFF6E90E , 32'hFFF9E619 , 32'h10AC5940 , 32'hFFFB18BA , 32'h00005661 , 32'hF6C63980 , 32'hFFFFA81E , 32'h026FF348 , 32'h044B7F00 , 32'hFFFB6DD4 , 32'hFFFD5C2C , 32'h00013251 , 32'hFAAF5BA8 , 32'h0BF53170 , 32'hF5F8E4A0 , 32'h0C935570 , 32'hFFFE78A3 , 32'h1A43A340 , 32'h00011E19 , 32'h000263CA , 32'h2EC6FCC0 , 32'h0C49DDC0 , 32'hEDBCC660 , 32'hFFF8EDD5 , 32'hFAFDAD00 , 32'hF6D477C0 , 32'h02262D5C , 32'hDE3EE080 , 32'h0EBABDE0 , 32'hFA1F2E98 , 32'hFEE160D0 , 32'hEA418B20 , 32'hFFFFB4E5 , 32'hFFFF9F45 , 32'h00035A2C , 32'hF9FB6E38 , 32'hDFEACAC0 , 32'h16054C60 , 32'hFEDDD62C , 32'hEABF5EA0 , 32'h1555C640 , 32'hFFF95825 , 32'hECAC9300 , 32'h0CE535A0 , 32'h0003C431 , 32'hFFBEC11A , 32'h000312EA , 32'hF8BDB9B0 , 32'h1EC178C0 , 32'h00027393 , 32'h000A47B2 , 32'hFFFA6A01 , 32'hFFFD7E96 , 32'h00030F37 , 32'hFFFDBA47 , 32'hFF0859B2 , 32'hEE9DEC20 , 32'h1666F520 , 32'hF3CCBCA0 , 32'hE6D32A00 , 32'hF9A6C0A8 , 32'h00000960 , 32'h0003FD35 , 32'hFFF96523 , 32'hFFFBB542 , 32'hFFFC70DD , 32'h01DC4850 , 32'hF71CE680 , 32'hF4ACB7B0 , 32'h00024F98 , 32'hFFF9A4EE , 32'h00046848 , 32'hFFFDA1A9 , 32'hFA763FD8 , 32'h12BC9B20 , 32'hFFF9CD92 , 32'hFFFF52E3 , 32'h00033A71 , 32'hFF0D74B3 , 32'h1CA6A820 , 32'hCEB01940 , 32'hFFFC8D6B , 32'h00019379 , 32'h0000AC6B , 32'h0391D3D4 , 32'h03F29710 , 32'h01BDFC44 , 32'h00028347 , 32'hFFD32E58 , 32'h000518F1 , 32'hDB441F80 , 32'h000747F8 , 32'h0C531BA0 , 32'h000033BA , 32'h0A65B2B0 , 32'hF424C910 , 32'hCC591DC0 , 32'h0E729F70 , 32'h0003A491 , 32'h0AAD8AB0 , 32'h0061F693 , 32'h00037E78 , 32'h1233C220 , 32'hFFFD7084 , 32'hF8B65B90 , 32'h00BE5566 , 32'hF70EC0C0 , 32'hFFFB3A46 , 32'h0004C05E , 32'hFA0A0850 , 32'h0006B451 , 32'h0FA97BA0 , 32'h000157B8 , 32'h0033A055 , 32'hFFFF2E4C , 32'h1DB956E0 , 32'hFFFDA658 , 32'hFFF9D8F4 , 32'h0000C5B7 , 32'h1D147CC0 , 32'h0C585E10 , 32'hFFFF045D , 32'h0001933E , 32'hFFFF9D87 , 32'hFFFAA26E , 32'h17C81700 , 32'hEB7F1EC0 , 32'hE73D0AC0 , 32'h4EB7D200 , 32'hF62884A0 , 32'h00026824 , 32'hFFFD82EC , 32'h0001A857 , 32'hFF032D84 , 32'h0000FA83 , 32'h0001B4E2 , 32'h08E35770 , 32'hE2BCCC80 , 32'hFFFDC3EC , 32'hCAC7E140 , 32'hF2C0BF30 , 32'hE0AC4E00 , 32'h1FCF3000 , 32'h000073D8 , 32'hFD4B0A6C , 32'hF4755E90 , 32'hFE851C50 , 32'h00026320 , 32'hE1CB9E20 , 32'hFCD1DF3C , 32'h26C58F00} , 
{32'hEA759300 , 32'h45FCFB80 , 32'hFFFE897D , 32'hFE644A84 , 32'hFFF71A0C , 32'h0348EF70 , 32'h0004E637 , 32'hFFFEFB8F , 32'hFFFD4884 , 32'hFFFBD42C , 32'hEA5FE6E0 , 32'hEFF64600 , 32'hF66144F0 , 32'h00055647 , 32'h0006D706 , 32'hD81A3640 , 32'hFFFD36F3 , 32'hF87DBB18 , 32'hFE93C9E8 , 32'hFFF8F2B7 , 32'h0001524A , 32'hF8C6F5A8 , 32'h0B0B5A20 , 32'hECE95700 , 32'h11BFB0A0 , 32'h000598D0 , 32'hFEDCE6B4 , 32'h08B626F0 , 32'hFFFE0C2F , 32'h05A0F540 , 32'hFFFCB241 , 32'hFA1FB5E8 , 32'hFFFD1F20 , 32'hFFFE7812 , 32'h0005DA2B , 32'hEDAA4580 , 32'hEF4C5640 , 32'h1089E540 , 32'h000234BF , 32'h0822B050 , 32'hE2233D00 , 32'h0002BC0D , 32'h0000BCE1 , 32'h0A16B000 , 32'h07CF2B60 , 32'hE8071DC0 , 32'hDE13C880 , 32'h0003BB3E , 32'hF8129DB8 , 32'hCCDDC8C0 , 32'h0143C374 , 32'hFFFB3730 , 32'h0083405C , 32'hDE540AC0 , 32'h0E281510 , 32'hFFFFF238 , 32'hFB8458B8 , 32'h0007C39A , 32'h0001DC88 , 32'h0208F3AC , 32'hFB336D00 , 32'hF597CFA0 , 32'h1AB2F420 , 32'hFFFEB282 , 32'h21395D40 , 32'hFFFFD496 , 32'hD095B640 , 32'h02EE26C0 , 32'hFFFC2796 , 32'h0AAC2980 , 32'hEE264260 , 32'h27DDF9C0 , 32'hFFFC8582 , 32'h0000CC00 , 32'hFFFDC0AB , 32'hE70D0FA0 , 32'h023C4588 , 32'h000195B8 , 32'h2831D3C0 , 32'hFDB53B48 , 32'hFFFD0ECD , 32'hE8D662A0 , 32'hFF71D9E7 , 32'h00003E4C , 32'hEDE947A0 , 32'h3FF9C800 , 32'h0AB612A0 , 32'h00001A8C , 32'h0007261E , 32'hD7ECB3C0 , 32'h00030CAD , 32'h010E2C38 , 32'hFFFE04B0 , 32'h018676A4 , 32'h010ECD2C , 32'h00082F68 , 32'h0005E712 , 32'hFFFEA413 , 32'h0004AB24 , 32'h047C5D40 , 32'hF5FBD700 , 32'h0000BD84 , 32'hF5524910 , 32'h03F4949C , 32'h077AEA68 , 32'h0000861D , 32'h01CE051C , 32'h0000AE33 , 32'hEB5CB9A0 , 32'h0E36C570 , 32'hFFFF3EE6 , 32'h1BA449A0 , 32'hFFFEA38B , 32'hFFFD2B05 , 32'hF52CCF20 , 32'hFFF2A8C3 , 32'hFBEC6090 , 32'hFFFE6C38 , 32'hF9A4A2D8 , 32'h0001DC29 , 32'h00035B61 , 32'h0176F9E4 , 32'h00048134 , 32'hFFF6CA2C , 32'hD54E04C0 , 32'hE61E2020 , 32'hFFFDEBF3 , 32'h0006E983 , 32'h0006A000 , 32'hFFFC82B8 , 32'hFFFE045A , 32'hE596DCE0 , 32'hF58D0BD0 , 32'hFFFE1605 , 32'hFFFCEA15 , 32'h0686CE38 , 32'hF9126968 , 32'h00014976 , 32'h00054BFE , 32'hF83BFDF8 , 32'h0000C6AF , 32'h0003347F , 32'hF1289920 , 32'hFF482299 , 32'h01AB05D8 , 32'h0146B958 , 32'h000060E2 , 32'hFFFDF0F8 , 32'h06C0B110 , 32'hFFFEDE9B , 32'h00043EE3 , 32'hFC9761F4 , 32'h0001EFFA , 32'h00062347 , 32'h08140E00 , 32'h0000C97D , 32'hD6FFAE00 , 32'hFD03D704 , 32'h00028DB8 , 32'hFFFEB199 , 32'hFFFE3BD3 , 32'h14E40140 , 32'h0275233C , 32'hEC5A6120 , 32'h1A7D5EE0 , 32'hFFFFCA83 , 32'hCE2E5B00 , 32'h0001289F , 32'hFFFFF35A , 32'hDD442C80 , 32'h06409BD0 , 32'h090D33B0 , 32'hFFFEAB35 , 32'h3EBCADC0 , 32'h04073AC8 , 32'hFBD9C5E0 , 32'hC94B74C0 , 32'h41EEC080 , 32'h08E65DA0 , 32'hFB5A0080 , 32'hF8DC7EF8 , 32'hFFFE67D8 , 32'h0000164B , 32'h0002E55F , 32'hFC807950 , 32'hE358AD00 , 32'hFFDA7BC9 , 32'hFA819A88 , 32'hFE38E7CC , 32'h0230BA04 , 32'hFFFFFB76 , 32'h0B3EBA20 , 32'hFE96A4FC , 32'h00015547 , 32'hDB325400 , 32'hFFF96983 , 32'h0E112A00 , 32'h18F29180 , 32'hFFFE00BA , 32'h000251F9 , 32'hFFFF50A4 , 32'h0006BD83 , 32'hFFFF5BF8 , 32'hFFFBB804 , 32'hFCDDF5D8 , 32'hF870F990 , 32'h0C832A70 , 32'h07487E70 , 32'h03B83DF8 , 32'h1FEF9540 , 32'h0003A671 , 32'h00022054 , 32'hFFFCF287 , 32'h0000652F , 32'hFFFB0671 , 32'h0CE0D5A0 , 32'h2C2756C0 , 32'h0428F170 , 32'h00002C26 , 32'h0000A8A2 , 32'hFFFC6C25 , 32'hFFFDD67F , 32'h0D69BE90 , 32'h0DE16A70 , 32'hFFF7F81B , 32'hFFFB6DF6 , 32'hFFFE6146 , 32'hD410C7C0 , 32'h424DB300 , 32'h094529A0 , 32'hFFFC3C99 , 32'h00039DC7 , 32'hFFFCFECF , 32'hFC325230 , 32'h02FBB294 , 32'hFC629B28 , 32'h00026160 , 32'hFF5CEF85 , 32'h0005EC7D , 32'hCCA20A80 , 32'h000A7812 , 32'h11A06AE0 , 32'h00036165 , 32'h1CF32100 , 32'h061323D0 , 32'h1536EA20 , 32'h0EB382B0 , 32'hFFFF1FA5 , 32'hFF7D783C , 32'hFB8B8528 , 32'hFFFABF1F , 32'hF65819D0 , 32'h00015EDC , 32'h0854C240 , 32'h196ADF80 , 32'hEAEAE020 , 32'h00024A69 , 32'hFFFD390F , 32'h0462F2F8 , 32'h00003B84 , 32'h1625AD00 , 32'h0005B560 , 32'h034C44D4 , 32'hFFFB0FCC , 32'h029A4678 , 32'hFFFABB63 , 32'hFFFAD1CB , 32'hFFFD99FE , 32'h01D19BD8 , 32'hE1C5F800 , 32'h0003E11A , 32'hFFFE7E7A , 32'h00011165 , 32'h0002E5C9 , 32'h202B3D00 , 32'hEDB08560 , 32'hE13C6B80 , 32'h08D53DA0 , 32'h121E0900 , 32'hFFFF718D , 32'h00013DC1 , 32'hFFFFEC28 , 32'h02222480 , 32'hFFFEEF1A , 32'h000514FE , 32'h0E5060B0 , 32'hE8495400 , 32'h0001CBBB , 32'hEF6F4A20 , 32'hFF70B03A , 32'hFC261870 , 32'hD58F7400 , 32'hFFFF138D , 32'hF95F8208 , 32'h15AF9180 , 32'h01777820 , 32'h00038075 , 32'h120DBE20 , 32'h2496CD40 , 32'h06062BB8} , 
{32'h061F8418 , 32'h37353240 , 32'h00027434 , 32'hEF980DC0 , 32'h0003D63E , 32'h03B68FE0 , 32'hFFF4E9AA , 32'hFFFE4A6C , 32'h0000C72B , 32'hFFF62B9B , 32'h090AECA0 , 32'h1B064440 , 32'h09AF3530 , 32'hFFFEF10E , 32'hFFFC9E69 , 32'hF2FC45A0 , 32'hFFFC0BEC , 32'hF3322560 , 32'hF343EF00 , 32'hFFFE1258 , 32'h0004232E , 32'h06E39170 , 32'h1A3E5840 , 32'h04C6F778 , 32'hF4EC9050 , 32'h0005D0CF , 32'h0A46D690 , 32'hFD96F4E0 , 32'h0005B13E , 32'hE5020260 , 32'h00034735 , 32'h0FCD6F50 , 32'h0002CE82 , 32'hFFFB9D63 , 32'hFFFDA542 , 32'hD19B6E80 , 32'hF7E6F5F0 , 32'hEDFE5B80 , 32'h0001909B , 32'h04917050 , 32'h322EC8C0 , 32'h00040A4B , 32'hFFFEAD64 , 32'h04704280 , 32'h03491664 , 32'hDA7B4340 , 32'h26A7C400 , 32'h00064C3F , 32'h1B026B20 , 32'h054429A8 , 32'hFE45AFB4 , 32'h000685CD , 32'hF2B954E0 , 32'h1DE82300 , 32'hF56A4A70 , 32'h000362F3 , 32'h065D8420 , 32'h0004EA4A , 32'h00011490 , 32'h0D5D1980 , 32'h02F9E900 , 32'h02CE2254 , 32'hF9EDDE98 , 32'hFFFF936E , 32'hFEC5FB88 , 32'hFFFD35A5 , 32'h3A03B2C0 , 32'h04A09E88 , 32'hFFFE54AD , 32'hF8733C68 , 32'hF4DB9020 , 32'hDF068640 , 32'hFFFD8FEF , 32'hFFFEFBAC , 32'hFFFFC72C , 32'h0859B800 , 32'hFDCCC6C4 , 32'hFFFF7D77 , 32'h172A7060 , 32'hFB5F63D8 , 32'h0001FED4 , 32'h33C66A00 , 32'hEFD85C40 , 32'h0002C06F , 32'h09337C70 , 32'hDC81C580 , 32'h09DB0BB0 , 32'h00001F6E , 32'hFFF9DD85 , 32'h33800E40 , 32'h00036FFE , 32'h123A3880 , 32'hFFFE904D , 32'hED8FE120 , 32'h025AD2B4 , 32'hFFFC56DC , 32'hFFFF606C , 32'h00015504 , 32'hFFFEA46F , 32'hEBFF1A80 , 32'h08AEE240 , 32'h0000BE95 , 32'h24B8C880 , 32'h1883FAC0 , 32'h07B16988 , 32'h0000F0E0 , 32'hFEF0B500 , 32'h0000DA60 , 32'hFFDBE6A7 , 32'h1B7F60C0 , 32'h00029438 , 32'hF20104D0 , 32'h000711DD , 32'hFFFEADB6 , 32'hFDDAFC24 , 32'h0D55EF90 , 32'hFD04BD68 , 32'hFFFFD1E9 , 32'hEB262D60 , 32'hFFFE6C22 , 32'hFFFDC553 , 32'hF697F9F0 , 32'hFFFCD37F , 32'h00051295 , 32'hE8E294E0 , 32'h1CB6EAC0 , 32'hFFFDB942 , 32'hFFFD58CA , 32'hFFFC83A1 , 32'h00034730 , 32'h0002C7FE , 32'h00BBCD28 , 32'hFFCFD48F , 32'h0001C81D , 32'h0000FA55 , 32'h193B20C0 , 32'hFD8A9384 , 32'hFFFB9C14 , 32'hFFFEB6E1 , 32'h03F99988 , 32'h00025A3A , 32'h00019D4B , 32'h03FA79BC , 32'h09180EE0 , 32'h04964D40 , 32'h05201B70 , 32'hFFFC85F1 , 32'hFFFF83AB , 32'hF5A3F800 , 32'h000476A7 , 32'hFFFAC8D2 , 32'h015F904C , 32'h0001031B , 32'hFFF5FD9D , 32'hFC681350 , 32'hFFFE3089 , 32'hFCBA624C , 32'h01CDD9CC , 32'hFFFBBC6C , 32'h0002D04C , 32'h0000F266 , 32'hFB0282B8 , 32'hE887CC40 , 32'hFFE273CF , 32'h135DB1A0 , 32'h0000505E , 32'hEBE25880 , 32'hFFFC555B , 32'h000200C9 , 32'h1202B180 , 32'hFADA3DB0 , 32'h01F3F3EC , 32'hFFFE2754 , 32'h1935BC80 , 32'h05DB2940 , 32'h083C5D00 , 32'hF0C75F50 , 32'hF4E6F800 , 32'h009FE812 , 32'hFAEDD770 , 32'hEE3815E0 , 32'h00005C68 , 32'hFFFAFF0A , 32'hFFFA45DA , 32'h07A43F40 , 32'hDDA9B640 , 32'hFDCDA068 , 32'hFEC0355C , 32'hF92CBDC0 , 32'h035D400C , 32'h0000760A , 32'h011CC2E8 , 32'h356F9D00 , 32'h00004130 , 32'h0C162A20 , 32'hFFFF0E14 , 32'h042CA068 , 32'h02D70F90 , 32'hFFFBD4FD , 32'h0005BF89 , 32'hFFF85B0B , 32'hFFFE8B6F , 32'h00007042 , 32'h00040B12 , 32'h05412230 , 32'hF665FA10 , 32'hE7A23520 , 32'hEC84EC80 , 32'hF0EAA0E0 , 32'hF9604480 , 32'hFFFBC2A5 , 32'h0000089A , 32'h0001A34C , 32'hFFFAF9D4 , 32'h0001EB39 , 32'hF7A76B20 , 32'hE7FEC5A0 , 32'hF5B1A1E0 , 32'h0001E8BB , 32'h000629E8 , 32'h000200C5 , 32'h00000A05 , 32'h0224B440 , 32'hF389E530 , 32'h00018FC7 , 32'hFFFB84B4 , 32'hFFFE4E10 , 32'hE94495E0 , 32'h58E7C800 , 32'h0A973640 , 32'hFFFC34B6 , 32'hFFFECC92 , 32'h0002C90A , 32'h04964D28 , 32'h0E95D310 , 32'h69091380 , 32'h00043BAE , 32'hFFF36505 , 32'hFFFD4C8B , 32'h0778EF70 , 32'hFFFF8001 , 32'hD094D700 , 32'hFFFE9E20 , 32'h21F73EC0 , 32'hE16B3200 , 32'h153929C0 , 32'h40618A80 , 32'h000688B6 , 32'h16D5A240 , 32'hFEE06C00 , 32'h00004AF9 , 32'hF5EA6440 , 32'hFFFE2D65 , 32'h027AA664 , 32'h03A99724 , 32'h01349040 , 32'hFFFDE941 , 32'hFFFD7EAB , 32'hFD41974C , 32'h000158B9 , 32'h01D1A3FC , 32'h0001A1F5 , 32'hFE1D3874 , 32'h00044B55 , 32'h0B7D7950 , 32'hFFFC78C5 , 32'h00004AAC , 32'hFFFF86A7 , 32'hFCC4B940 , 32'hEECDAA60 , 32'h0002A803 , 32'hFFFF0F55 , 32'h000163B8 , 32'hFFFCFD59 , 32'hDC778EC0 , 32'h12A3DA40 , 32'hFBB58E80 , 32'hDFCB2940 , 32'hF80D7270 , 32'hFFFF0C49 , 32'hFFFE3FC0 , 32'h00040BD4 , 32'hFF994F24 , 32'hFFFDDD8B , 32'h0003D901 , 32'hEC5FEDE0 , 32'hF6DA1F30 , 32'hFFFD63DF , 32'hF1D9F600 , 32'hFEEDDEF0 , 32'h047FCD70 , 32'hDCAF31C0 , 32'hFFFDCFD0 , 32'h108FFE80 , 32'h25908480 , 32'h08561140 , 32'h0005BA0B , 32'hE768AE40 , 32'hDC414440 , 32'h04837290} , 
{32'hF31DD4E0 , 32'hF5D7C660 , 32'hFFFF33FE , 32'h19E85AA0 , 32'hFFFE5BC9 , 32'hFF318D1B , 32'hFFFC6603 , 32'hFFFD4746 , 32'h0001D92B , 32'hFFFD984B , 32'hDD5B3D00 , 32'h1A09CCA0 , 32'h042B0ED0 , 32'hFFFF6B99 , 32'hFFF9CAD1 , 32'hE52C9520 , 32'h00011763 , 32'h28EAD4C0 , 32'h00D9F59B , 32'h00009D64 , 32'hFFFC9B97 , 32'h01C61790 , 32'h01A7DCDC , 32'hF14B5BE0 , 32'hFE2FC408 , 32'h0003B70B , 32'h022C11F8 , 32'hF8331D48 , 32'hFFFC60AE , 32'hFF637405 , 32'hFFFD506C , 32'h01A00BEC , 32'h0006D26B , 32'h0001F938 , 32'hFFFE7AA7 , 32'h152DC2A0 , 32'hCFD2D940 , 32'hFDCE9074 , 32'h00037B62 , 32'hDCB0CA80 , 32'hF307B0C0 , 32'hFFFF3E53 , 32'hFFFFFDF3 , 32'h081B6760 , 32'hE95DE340 , 32'hFD060DEC , 32'h12CB9A80 , 32'hFFFDBB51 , 32'h12EF5CA0 , 32'h0E2039F0 , 32'hFEBFA968 , 32'h000290CC , 32'hFE7A9D00 , 32'h304DF000 , 32'h0CB944F0 , 32'h0005B8FC , 32'h07EEF6A8 , 32'h00001BA7 , 32'h000074B9 , 32'h0813D9A0 , 32'hF87C7398 , 32'h068946A8 , 32'hBA944300 , 32'hFFFD676E , 32'h0CEE9E00 , 32'h00058462 , 32'h07586968 , 32'h0A612250 , 32'hFFFC0E7A , 32'h11111E60 , 32'h128FD960 , 32'hE4260060 , 32'h00061BD5 , 32'h00047BA3 , 32'h0005C3C5 , 32'h0C3BB2B0 , 32'hEFEB3BE0 , 32'h00019304 , 32'hEDC1F580 , 32'hFEF416F4 , 32'hFFFCA509 , 32'hF1684270 , 32'h018CE104 , 32'h0001070E , 32'hFA0A2008 , 32'hEDD4C1C0 , 32'hFE979438 , 32'hFFFB0F76 , 32'hFFFF8240 , 32'h38BB53C0 , 32'h000554E1 , 32'hFEF42534 , 32'hFFFF96EF , 32'hFEA33344 , 32'h0185A4F8 , 32'h00092346 , 32'hFFFFB30D , 32'h0000634D , 32'hFFFC87B1 , 32'hFA346FC0 , 32'hF6FEC400 , 32'h00016752 , 32'hD9F1ED80 , 32'h2CEC8580 , 32'hF707AFB0 , 32'h0004B1E0 , 32'hFF50D487 , 32'h000173A2 , 32'hE9AEF7A0 , 32'h1008CDA0 , 32'hFFFBC201 , 32'hF2F80E70 , 32'h0002CA02 , 32'hFFFEC2D9 , 32'hE6488160 , 32'h14170600 , 32'h000C965B , 32'h000259B2 , 32'h01B6AC9C , 32'hFFFCA52D , 32'hFFFD281E , 32'h1320F060 , 32'h000516EB , 32'h0000BD1E , 32'hE2AF73A0 , 32'hEABF1560 , 32'hFFFB3987 , 32'h00054A13 , 32'h0004494A , 32'hFFFDEDF7 , 32'h0000481F , 32'hF57723A0 , 32'h1638AEC0 , 32'hFFFE57FA , 32'hFFF7DA0C , 32'hEAFCED40 , 32'hE278F100 , 32'h00057328 , 32'hFFFF87B0 , 32'h0B1A7A80 , 32'hFFFF7757 , 32'hFFFDCF75 , 32'h04CE50D0 , 32'hF235BA90 , 32'h08E6B280 , 32'h0A2DD0D0 , 32'hFFF80F01 , 32'hFFFD0FD6 , 32'hF8045338 , 32'h00025F41 , 32'hFFF49417 , 32'hF3E72630 , 32'hFFFE0751 , 32'hFFFAC745 , 32'hFDFA6D2C , 32'hFFFF7B9D , 32'hF4228A10 , 32'hFFA05C6C , 32'h00068F9C , 32'hFFFAC764 , 32'h000526CE , 32'hF15BAB90 , 32'hFFE32450 , 32'hF89DF208 , 32'hEF7EE9E0 , 32'h0001980D , 32'h36A7D640 , 32'h00002521 , 32'hFFFDFE22 , 32'h11EADB00 , 32'h03A0CBC8 , 32'hF7A1D730 , 32'hFFFE8FFA , 32'h392AD880 , 32'hF979F988 , 32'hF777E4B0 , 32'h0BD3FF40 , 32'h1B587A80 , 32'h57556B80 , 32'hFEFA1F40 , 32'h24D4F300 , 32'hFFFFDB72 , 32'hFFFC6B87 , 32'hFFFF66D7 , 32'hFD8D0D78 , 32'h13209240 , 32'h06C8FDA8 , 32'h01949AB8 , 32'h204A9EC0 , 32'h0B86B790 , 32'hFFFDED0F , 32'h1003E7A0 , 32'hFF235C50 , 32'hFFFCE914 , 32'hF5063EA0 , 32'hFFFF8A2A , 32'h0688FEA8 , 32'h2540B7C0 , 32'h00021433 , 32'hFFFDEC80 , 32'hFFFD9723 , 32'hFFFC9EA4 , 32'hFFFE047F , 32'h000348BC , 32'hFD8DE5BC , 32'hE4BDC960 , 32'hD548A240 , 32'h01A870F8 , 32'hF1FC2710 , 32'h1DD9E100 , 32'hFFFD97B8 , 32'h00018B66 , 32'h0000E8B4 , 32'h00042843 , 32'h00057888 , 32'hF9FD5740 , 32'hFA3540D0 , 32'h10C8A860 , 32'h0001454B , 32'h0003BA0E , 32'hFFFE1713 , 32'hFFFDEC08 , 32'hE2D54A80 , 32'hE4747020 , 32'hFFFFC17C , 32'hFFFE460A , 32'hFFFBD7A9 , 32'hDC0ACD00 , 32'h36148700 , 32'hFBD26A18 , 32'h00017E2C , 32'h0001E3A3 , 32'h00001AD9 , 32'hF68E1B20 , 32'h09D5DDE0 , 32'hD78F7380 , 32'hFFFB907D , 32'h02D688EC , 32'hFFFA0778 , 32'h012211B8 , 32'h0002D81A , 32'hFB251990 , 32'h00035901 , 32'h003357D1 , 32'hF54C95B0 , 32'hFD108064 , 32'hC8DCED80 , 32'hFFFD12AA , 32'h0531B590 , 32'hFEEB1A74 , 32'hFFFC6DDB , 32'h023D90A8 , 32'hFFF8E86F , 32'h07194FB8 , 32'h25D29E80 , 32'h105D9F60 , 32'h0003D4E1 , 32'h00039BF8 , 32'h09D77920 , 32'hFFFE6070 , 32'hE0B5C040 , 32'h0004CF0F , 32'h004D6CF6 , 32'hFFFD9A46 , 32'hF46DCE90 , 32'h00004AB8 , 32'h0001D45B , 32'hFFFF9922 , 32'h0C82FD20 , 32'h2DABC600 , 32'h0003D55E , 32'h00066D34 , 32'h0001AD17 , 32'hFFFD86BE , 32'h116C58C0 , 32'h0BDB82B0 , 32'hC8CCDD00 , 32'h02C52BFC , 32'h116A1960 , 32'h00017F14 , 32'hFFF8CB76 , 32'h000514DE , 32'h04276380 , 32'h00003D45 , 32'h00043F64 , 32'h03ECA63C , 32'h0B7BB300 , 32'hFFF71070 , 32'hF0337840 , 32'h02832AEC , 32'hED9D9CC0 , 32'h17C64B60 , 32'hFFFE29E9 , 32'h0D0922A0 , 32'hE52CDB40 , 32'h044DE9F0 , 32'h00084E37 , 32'h2A8485C0 , 32'hE949EDA0 , 32'hF3A55370} , 
{32'h19055DA0 , 32'hCD877740 , 32'h0003738B , 32'hF477D340 , 32'h00027661 , 32'h11577C80 , 32'hFFFA1001 , 32'hFFFE8DF8 , 32'hFFFFB3AB , 32'h0000EE74 , 32'h0A7EF3F0 , 32'h15542D20 , 32'h055F02B0 , 32'hFFFB6944 , 32'hFFF5DA2D , 32'hE2A80100 , 32'h00098D4F , 32'h1A850F00 , 32'hF46469B0 , 32'hFFFE3251 , 32'h0000B461 , 32'hFBFD6690 , 32'h0BF44D70 , 32'hE1563280 , 32'h026AD9FC , 32'hFFFB6CE6 , 32'h08361400 , 32'hFD13F1D8 , 32'h00026642 , 32'h1DA81AC0 , 32'h000285FC , 32'h07142198 , 32'hFFFFCA1D , 32'hFFFE5E3D , 32'hFFFD2E33 , 32'h00F41D83 , 32'h1A9785C0 , 32'hE8EA72E0 , 32'hFFFB7210 , 32'h0CB693A0 , 32'hEF0DBBC0 , 32'hFFFEE31B , 32'hFFF9FB23 , 32'hFBBEBA50 , 32'h13D30BC0 , 32'h00BCF3A5 , 32'h07D48140 , 32'h00055451 , 32'hD53B8400 , 32'hEE15FB20 , 32'h028E864C , 32'hFFF90C83 , 32'h0B141CA0 , 32'hE9FAF200 , 32'hEC175760 , 32'hFFFF8497 , 32'h0063B000 , 32'hFFFF4E22 , 32'hFFFC130E , 32'hF6F1F890 , 32'h00D2644E , 32'hE39F4020 , 32'hF5E67120 , 32'hFFFF7A2F , 32'hB965CE80 , 32'h0006360D , 32'hE3FDF9E0 , 32'h01D3D6E0 , 32'hFFFB57BF , 32'h24730E40 , 32'h028F6CF4 , 32'h06289F10 , 32'h00002B84 , 32'h0001E867 , 32'h00019978 , 32'h0BE36490 , 32'h0B3DEC10 , 32'hFFF7FB37 , 32'hDACE9F40 , 32'h04A76070 , 32'hFFFCE5E8 , 32'h4F39B700 , 32'h0C3176A0 , 32'h0000D152 , 32'hF8B69698 , 32'hE1B27640 , 32'hFB679370 , 32'h00099FA1 , 32'h00019ED1 , 32'hC04EFC00 , 32'h0000D531 , 32'hFDB19F30 , 32'h0000450E , 32'hFDF16EA8 , 32'h00CEA39C , 32'hFFFBA5E6 , 32'h00006B2F , 32'h000065ED , 32'hFFFF0461 , 32'hF21336B0 , 32'hF40363A0 , 32'hFFFF1BC5 , 32'hE9AE1320 , 32'h1A9F8700 , 32'h07A0AA70 , 32'hFFFDBEA6 , 32'hFF824CBD , 32'hFFFE7F93 , 32'h0C8808A0 , 32'h01447DB8 , 32'hFFFECF30 , 32'hD9731680 , 32'h00004788 , 32'hFFFE5D7C , 32'h06E92B60 , 32'hF634FC90 , 32'h021B3D64 , 32'h000185CC , 32'hFE3809D0 , 32'h0000DBBE , 32'h00058736 , 32'h02255688 , 32'hFFFED9B6 , 32'h0006187E , 32'hD53C9FC0 , 32'h09906BB0 , 32'hFFFCB01E , 32'hFFF73387 , 32'h0003B5ED , 32'h0000A36C , 32'h0002E3F5 , 32'h08C88400 , 32'h1AB66EE0 , 32'hFFFB37F7 , 32'hFFF9E590 , 32'hED194200 , 32'hF056C1B0 , 32'hFFFE4370 , 32'h000144C0 , 32'hFB9569E8 , 32'h0002FED3 , 32'h0001C5F8 , 32'h0CAEF5B0 , 32'h10F26160 , 32'hF92E7BB0 , 32'h018C4700 , 32'hFFFCE4F0 , 32'hFFFA5586 , 32'hF64C0680 , 32'h000166D2 , 32'h0002A83A , 32'h07C06600 , 32'hFFFFAEDB , 32'hFFFF90AC , 32'h0108CF34 , 32'h00018F10 , 32'hF13E06A0 , 32'h0345FBB8 , 32'hFFF8C8CD , 32'h00029DEE , 32'hFFFD5E2D , 32'h0D44A5A0 , 32'h0FDC7120 , 32'h0876C2A0 , 32'h25362740 , 32'hFFFC79B6 , 32'hF391E900 , 32'h0001087B , 32'h0002CDA5 , 32'hFF882D28 , 32'h00822BEF , 32'hEB7A3C80 , 32'hFFFC1A38 , 32'h1EACA1A0 , 32'hF926DA48 , 32'h06711F38 , 32'hDE5F21C0 , 32'hD1A70E80 , 32'h4EC30500 , 32'hFFBED0B5 , 32'h0DAB2A60 , 32'hFFFD24A9 , 32'h0002AA29 , 32'hFFFE6079 , 32'hFBF806A0 , 32'hE4336DA0 , 32'hF47D29F0 , 32'h018FE794 , 32'hE912C7A0 , 32'h0267D794 , 32'h0002622C , 32'h0FBD4EA0 , 32'h192BB6A0 , 32'h0001F9B6 , 32'h00C0044F , 32'h00042CA1 , 32'h00A441FF , 32'hE8AB0DC0 , 32'hFFFE5C8A , 32'h0005EF07 , 32'hFFFE49B8 , 32'hFFFFFA99 , 32'hFFFB24A0 , 32'h0003E388 , 32'h061106D8 , 32'h1361A5E0 , 32'h1B539220 , 32'h09C44450 , 32'hFF72A7D2 , 32'h0DAD7A40 , 32'h00034438 , 32'h00003174 , 32'h0001BA31 , 32'hFFFF68E7 , 32'h000110BF , 32'hF11ECCB0 , 32'h125D1A60 , 32'hE9BF2640 , 32'h0005E20F , 32'h00010489 , 32'hFFFB867F , 32'hFFFCE679 , 32'hF5177DF0 , 32'hE89EFA00 , 32'hFFFFC76A , 32'h0000003E , 32'hFFFAC749 , 32'h1B6608E0 , 32'hF675B170 , 32'h00EE0D01 , 32'hFFFCDEEE , 32'hFFF7B77A , 32'hFFFEB1C8 , 32'h04404FC0 , 32'h01246074 , 32'h27B4E440 , 32'hFFFB8162 , 32'h00A3DCCD , 32'hFFFE7BE0 , 32'hE5561600 , 32'h0001429B , 32'h1DDF6F60 , 32'h00042F57 , 32'h164F0D60 , 32'hED5397C0 , 32'hE6365E40 , 32'hFD7697A8 , 32'h0000235C , 32'hF317DA30 , 32'h00E785B7 , 32'h00021EB4 , 32'h036273EC , 32'hFFFDD830 , 32'hFE1A84E8 , 32'hF9B14020 , 32'hE352A580 , 32'hFFFFA935 , 32'hFFF81BF6 , 32'h2157F9C0 , 32'h00031A2F , 32'h061E9B70 , 32'hFFFF6142 , 32'hFD8F5714 , 32'h000344A2 , 32'hF715AB10 , 32'hFFFA7702 , 32'hFFF7B2AA , 32'h00036F52 , 32'hE2F33EE0 , 32'hF88EBA08 , 32'h0002D827 , 32'hFFFDD53E , 32'hFFFC4F46 , 32'hFFFFA19D , 32'hFD1276E4 , 32'hEAA36660 , 32'h084B8080 , 32'h47FB4D80 , 32'hF2284370 , 32'h00022632 , 32'hFFFCB0FB , 32'hFFFBB230 , 32'hF769E000 , 32'hFFFDF453 , 32'h00003651 , 32'h0C562230 , 32'hE4234F40 , 32'hFFFF6859 , 32'hC0C17B00 , 32'hF92316E8 , 32'h0660CC18 , 32'h188239E0 , 32'h000445D6 , 32'hF82F6FD8 , 32'h00E09C85 , 32'h05F60258 , 32'h0003DA34 , 32'h05592870 , 32'hD3BB4E00 , 32'hE93A6A00} , 
{32'h418DB780 , 32'hF32D83E0 , 32'h0000ACD4 , 32'h098D4770 , 32'h00041813 , 32'h0C45E800 , 32'h000079BD , 32'hFFFFC664 , 32'hFFFFE1BE , 32'h00025816 , 32'h02A10740 , 32'hF4D3A210 , 32'hE07EA360 , 32'hFFFE3222 , 32'hFFFE7301 , 32'hFD86DB38 , 32'hFFFFFC0F , 32'hEEEDB3E0 , 32'hFA0350D8 , 32'hFFFC7FFA , 32'h0004E0CA , 32'h00D3B82C , 32'hEE462520 , 32'h18331DA0 , 32'hFBCA4AA0 , 32'hFFFC4F07 , 32'h07635980 , 32'h05169E00 , 32'h0002611B , 32'hFA66F0C0 , 32'h00010BE3 , 32'h14950760 , 32'h0001373E , 32'hFFFA0133 , 32'hFFF9EBB9 , 32'h17580120 , 32'hFA798908 , 32'hF36D5A50 , 32'hFFFEB5B2 , 32'hD37BECC0 , 32'hE2706120 , 32'h000416F2 , 32'hFFFF48B0 , 32'hFD080A64 , 32'hE62FB8C0 , 32'h0198E14C , 32'h0F483A40 , 32'hFFF96EFE , 32'h008ACEEA , 32'h165C1D80 , 32'hFE68414C , 32'hFFFE50EC , 32'h00070EE3 , 32'h0378B4CC , 32'h11D4AD80 , 32'hFFFDE7C7 , 32'h0134A90C , 32'hFFFC3921 , 32'h0004871F , 32'hFC19DAD4 , 32'hFE31EFB0 , 32'hFC830780 , 32'h28825B00 , 32'hFFFF44F8 , 32'hF7FBAD30 , 32'h000243C4 , 32'h1DFCF000 , 32'h06746BA8 , 32'h0004E3F4 , 32'h1B6D49C0 , 32'hF5956CB0 , 32'h245E7840 , 32'h0000405A , 32'hFFFD0E9D , 32'h0001FD8B , 32'h25579380 , 32'h11FD55A0 , 32'hFFFF5EDC , 32'hCCA8F400 , 32'h0590D8E0 , 32'hFFFE60E5 , 32'hE6FB6DC0 , 32'h0DFDDBD0 , 32'h0001320B , 32'h114589A0 , 32'hEC282440 , 32'hFFD2E4B7 , 32'hFFF9750B , 32'h00016CC9 , 32'hE2775740 , 32'h00030722 , 32'h15D25000 , 32'h0001C77F , 32'hF60C9340 , 32'h00F71594 , 32'h0003BD36 , 32'h000436C0 , 32'hFFF92C5E , 32'hFFFC9487 , 32'hF3CAE590 , 32'hFCED75B4 , 32'h0000BE96 , 32'h0C245080 , 32'hF6646A90 , 32'h093FD300 , 32'hFFFE6CC6 , 32'hFFA4D352 , 32'h00014258 , 32'h05ACB998 , 32'h30C9FD40 , 32'h0001E1B4 , 32'hF6AACE60 , 32'h00009B00 , 32'h000530C8 , 32'hF0549FC0 , 32'h071E9C08 , 32'hFDB6E9E8 , 32'hFFFEFFE0 , 32'hE7E333C0 , 32'hFFFF45AF , 32'hFFFE22B0 , 32'hF956DD28 , 32'h00032701 , 32'hFFFC8760 , 32'h40947E00 , 32'hEC2F7BA0 , 32'hFFFE02AC , 32'h00038540 , 32'h0000C6F2 , 32'hFFFB56AE , 32'h00025941 , 32'hF9B66480 , 32'hFA2AF810 , 32'hFFFE2109 , 32'hFFFE4C1B , 32'h0F387100 , 32'hDA532140 , 32'hFFFE3D0A , 32'h0001A946 , 32'hF0CE0CB0 , 32'h0001CA77 , 32'hFFFF840A , 32'hFBF3AEF0 , 32'h02053AF0 , 32'h040F4540 , 32'h05C14508 , 32'h0004A92C , 32'hFFFAEBFB , 32'hF8D217E8 , 32'hFFFEE838 , 32'h0000A853 , 32'h0721E848 , 32'hFFFD65FB , 32'h000403E3 , 32'h010E4404 , 32'h0001E1AC , 32'hFC8DF17C , 32'h01897F48 , 32'h00019A77 , 32'hFFFF7B78 , 32'hFFFC01C8 , 32'h355E5B00 , 32'h0D63B7D0 , 32'hFE893A28 , 32'h0D3531A0 , 32'h00013A16 , 32'h10A0EDA0 , 32'h00005500 , 32'hFFF741DA , 32'hFF1218FC , 32'hF38C6C60 , 32'h072F22B8 , 32'hFFFE7ADE , 32'h39860240 , 32'h01A507C0 , 32'h10F091E0 , 32'h116AC620 , 32'h07B38E58 , 32'hDD022F80 , 32'hFD3F4410 , 32'h084CBF70 , 32'h00037AE6 , 32'h00040E81 , 32'h00017C95 , 32'hED1FF680 , 32'hF8A998A8 , 32'h03B7FD6C , 32'hFF6E2906 , 32'hE4689CE0 , 32'hFF27896B , 32'hFFFFD218 , 32'hE1BB4E80 , 32'h19782B80 , 32'h000236CC , 32'hF3130E70 , 32'hFFF84913 , 32'hFAF32890 , 32'hF3E39290 , 32'hFFFAA802 , 32'hFFFF2546 , 32'hFFFB244D , 32'h000348B0 , 32'hFFF92AD4 , 32'hFFFC49BD , 32'h0C004B50 , 32'hDF5312C0 , 32'hEF05AD00 , 32'hF90D6CC8 , 32'h0C31E3B0 , 32'hECF3D980 , 32'hFFFF8CB1 , 32'hFFF81D82 , 32'h00001B60 , 32'h00008FA9 , 32'h0006D037 , 32'hFC817430 , 32'h28EDF300 , 32'h1B0E3E80 , 32'h00022798 , 32'h0000EB51 , 32'hFFFCA9CE , 32'h000125DC , 32'h172544E0 , 32'hE248A4E0 , 32'hFFFE16A6 , 32'h0004EC7D , 32'h00036C92 , 32'h0BF24F40 , 32'hF61B1F50 , 32'hE9C4EB60 , 32'hFFFE5DC9 , 32'h00051076 , 32'hFFFE4D47 , 32'hF2D26020 , 32'h083FB500 , 32'h0F1C16C0 , 32'h00060772 , 32'h01D58490 , 32'h0003AF1B , 32'hEC2C14A0 , 32'h00007AA1 , 32'h06E920F8 , 32'hFFFFE2DD , 32'hB5FE3C80 , 32'hF1F0E050 , 32'h0A866130 , 32'h13CB2680 , 32'hFFFF9CE8 , 32'hFE144720 , 32'hFF4C31AC , 32'h0001B1A7 , 32'hF26B8370 , 32'hFFFC5287 , 32'h0B5860C0 , 32'h5FC94800 , 32'h13527360 , 32'h0000E988 , 32'h0005A5C2 , 32'hF4816C30 , 32'h00001E66 , 32'hF2C61630 , 32'hFFFFD667 , 32'hFFCFAB25 , 32'h000A0293 , 32'h11607560 , 32'hFFFE8DAA , 32'hFFFD4103 , 32'hFFFD816E , 32'hC9C8F880 , 32'hED3B6A60 , 32'h00007A21 , 32'hFFFEBE3A , 32'h0004402C , 32'h000146D4 , 32'hF2F43780 , 32'hFC1A7AF4 , 32'hE09ED080 , 32'h11330E80 , 32'h377DF100 , 32'h00008C74 , 32'hFFFBDA86 , 32'h0002CE9D , 32'h03A8CC84 , 32'hFFFEE521 , 32'h00026697 , 32'hF853BCB8 , 32'hF98C6E30 , 32'h00003CC4 , 32'h02EF8598 , 32'hFC3BC4D8 , 32'h02756750 , 32'hDA469480 , 32'h000082AB , 32'h0DC7AD90 , 32'hDB0B3E00 , 32'h0469F168 , 32'hFFFCFC0E , 32'hDF5CA100 , 32'hF1C30260 , 32'h0B451B80} , 
{32'h1197CD60 , 32'h127631E0 , 32'hFFFE4656 , 32'hD102D940 , 32'hFFFDF643 , 32'hFC564A5C , 32'h0001C4BA , 32'hFFFE2EEC , 32'h000072A6 , 32'hFFFCD8E7 , 32'hDC74A380 , 32'h01ACFAD0 , 32'h1474B3E0 , 32'h00030606 , 32'hFFF7EF12 , 32'hFE089548 , 32'h0001B010 , 32'hF138DF40 , 32'h01BBB1A4 , 32'hFFFB1994 , 32'hFFFEB35F , 32'h04A9D548 , 32'h029F3BA8 , 32'h01A35B7C , 32'h17EFD380 , 32'hFFF81D55 , 32'hF6DF74F0 , 32'hFBA19C58 , 32'h0000C50F , 32'h2146F0C0 , 32'hFFFE4B67 , 32'h0B092780 , 32'h0001520D , 32'h000253A7 , 32'h00008D9F , 32'h09EB9FD0 , 32'h0DC20CE0 , 32'hFA875A98 , 32'hFFFF0DFE , 32'hDF5E6100 , 32'h28CCCAC0 , 32'h00003936 , 32'h00034326 , 32'hFFEF9A67 , 32'hF4E31EC0 , 32'h1B6823C0 , 32'hEFFAE4C0 , 32'h00033B37 , 32'h1AFBC020 , 32'hF2ABDD90 , 32'hFD764218 , 32'h00024A2D , 32'hFA94C580 , 32'h1D1C8120 , 32'h04F0CCF8 , 32'hFFFBA6A3 , 32'hFEE47E38 , 32'h0003940F , 32'h0004A63F , 32'h0CDF4D30 , 32'h076D2698 , 32'h0C3639F0 , 32'h26047580 , 32'h0003B9AD , 32'hDBD82980 , 32'hFFFAA186 , 32'hDFC10940 , 32'hFF0F2F84 , 32'hFFFEC0E4 , 32'h392F0C40 , 32'hE71E09E0 , 32'hF7996690 , 32'h000B33BC , 32'h00012AD5 , 32'hFFFD138C , 32'h316F25C0 , 32'hF84DF890 , 32'hFFFD8086 , 32'hF85F01A8 , 32'h029F1F88 , 32'hFFFD5C29 , 32'h22122580 , 32'hF188C680 , 32'h0001EF7D , 32'h015B9E7C , 32'h0D31DF80 , 32'h07B96678 , 32'hFFF4FB05 , 32'hFFF8AC5C , 32'h05A09F08 , 32'hFFFEC96B , 32'h05D94A38 , 32'h0000B4A2 , 32'h133C4740 , 32'hFCC330D8 , 32'hFFFAD648 , 32'hFFFEE9A2 , 32'h000013E7 , 32'h00038ED6 , 32'hFD7AB854 , 32'hF8A0C178 , 32'h000434E2 , 32'hF3852EA0 , 32'h0FFB4BC0 , 32'hF8ED8FE0 , 32'hFFFC9DD0 , 32'hFE71AF08 , 32'hFFFE73AB , 32'h0B754F70 , 32'hEC432500 , 32'hFFFEFCC3 , 32'h05E18EF8 , 32'hFFFA8566 , 32'h00013DEE , 32'h1D081020 , 32'hF7C8EC00 , 32'h03EFFD90 , 32'h00010D74 , 32'h0E043C30 , 32'h00033915 , 32'h0001B954 , 32'hE8109460 , 32'h00024B77 , 32'h0002A919 , 32'hE3996AE0 , 32'h0AB0B700 , 32'hFFFD215D , 32'h00028258 , 32'hFFFF1AEA , 32'hFFFBA29C , 32'hFFFCBCEE , 32'h0BA57AF0 , 32'hEE562DA0 , 32'h0001B6EF , 32'h0000214F , 32'hD25E0D80 , 32'hF9CC42C8 , 32'h0000E50F , 32'h0000C37D , 32'hFA793E70 , 32'h00041187 , 32'hFFFF031A , 32'hF7CCF9C0 , 32'hF28C5570 , 32'hFB97D9F8 , 32'hFB2F8530 , 32'hFFFD84CF , 32'hFFFFDB3A , 32'h060FD9C8 , 32'hFFFC6C22 , 32'hFFF8325F , 32'hFD430B54 , 32'hFFFE49A2 , 32'hFFFC192F , 32'hE85B6C60 , 32'h000266F2 , 32'hEADDD460 , 32'h020080D8 , 32'hFFFE05C8 , 32'hFFFFE0BA , 32'hFFFEFAD2 , 32'hE14C8540 , 32'hE2DA5A40 , 32'h04FDA658 , 32'hF2824860 , 32'h00012BEF , 32'hA761B680 , 32'h000205FB , 32'hFFFA40FC , 32'h1576A680 , 32'hF70DF560 , 32'hFF903BD7 , 32'h00056354 , 32'hCF79F880 , 32'hFBF25678 , 32'h15E34660 , 32'hF13C8BE0 , 32'h12EC8740 , 32'hE0897040 , 32'hFDCB4300 , 32'h2BFFB780 , 32'h0003F3C7 , 32'h0000CB08 , 32'hFFFF8522 , 32'hE947D7C0 , 32'hD9783C80 , 32'hFE761010 , 32'h026D2058 , 32'hFA5C4A30 , 32'hFA719500 , 32'hFFFD6EB0 , 32'hD8FDBF00 , 32'hD8735EC0 , 32'hFFFE2133 , 32'hE5A45CA0 , 32'h0003BAC9 , 32'hFFCAF9E0 , 32'h3AAC40C0 , 32'hFFFDF346 , 32'h00023E36 , 32'hFFFD6ADC , 32'h00024C88 , 32'h00005A02 , 32'hFFFE1D3E , 32'h036C1B00 , 32'h046686B0 , 32'hDE1515C0 , 32'hFCC41098 , 32'hD20695C0 , 32'hF758C390 , 32'h0000126B , 32'hFFFDE1D9 , 32'h00054B4E , 32'hFFFD241C , 32'h0006A5E0 , 32'hFDC23634 , 32'hD67670C0 , 32'h0F60FA60 , 32'hFFFB945F , 32'hFFFE28C1 , 32'hFFF711B1 , 32'h0003516E , 32'hE5F36840 , 32'h04449370 , 32'h000017A3 , 32'h00040319 , 32'h0000A829 , 32'h33A2C280 , 32'h2391B140 , 32'hF2E80B30 , 32'h00026908 , 32'hFFFD966E , 32'h0000225F , 32'h02C33548 , 32'h00B87E80 , 32'hDAE1CF00 , 32'h00032D0A , 32'h00E95F6D , 32'hFFFB1E32 , 32'h1F7DD6E0 , 32'hFFFC96EE , 32'h09A2D1A0 , 32'hFFFF08FD , 32'hE9E7D9C0 , 32'h0870DF60 , 32'hF1BB3500 , 32'hE8DB0F80 , 32'hFFFB4B46 , 32'h094CBFC0 , 32'hFF353EE6 , 32'h0004AD34 , 32'h0F188910 , 32'h00011B3C , 32'hFD071B00 , 32'h14479CC0 , 32'h21388B40 , 32'h0004E121 , 32'h0001CB09 , 32'h028024A0 , 32'h0003D9FC , 32'hC356AE00 , 32'hFFF6A5F2 , 32'h0511FDD0 , 32'hFFFFFDBC , 32'h077A0C70 , 32'hFFFCFCD1 , 32'h000265A8 , 32'hFFF9BD3F , 32'hEE270040 , 32'hCF6AF200 , 32'h00065234 , 32'hFFFFCE23 , 32'h00009539 , 32'h0000BB98 , 32'hF5920C20 , 32'hFC6C6454 , 32'hEBCC70C0 , 32'h0EE6EC00 , 32'h09028CA0 , 32'hFFFF64E7 , 32'hFFFDBA56 , 32'h00008F9E , 32'h0150DF68 , 32'hFFFF94C4 , 32'hFFFEF308 , 32'hF23CCB40 , 32'hE2A45960 , 32'hFFFD9576 , 32'h08CF0260 , 32'hF670DB00 , 32'h1052D240 , 32'hF73F7410 , 32'h0000D7B1 , 32'hEF752880 , 32'h0280CF18 , 32'hF89B3E00 , 32'hFFFD8D0A , 32'h0A935A90 , 32'hF21D4960 , 32'h031309F0} , 
{32'hD2186C80 , 32'hD0E8A380 , 32'hFFFC8BFC , 32'hE9E386A0 , 32'h0001CC1F , 32'h1474FE00 , 32'hFFFEE7A4 , 32'h00005FA0 , 32'hFFFE5DAC , 32'h0007C580 , 32'h05291A60 , 32'h1D71BF40 , 32'hFFEBFD0E , 32'h00043A33 , 32'hFFFE96FD , 32'h4BB6F100 , 32'h00018BDA , 32'hF4B9B2B0 , 32'hEE570DA0 , 32'h000379A8 , 32'hFFFEB856 , 32'h03E81858 , 32'h0C3CA470 , 32'h1CD94980 , 32'h1708C060 , 32'hFFFC074C , 32'hFF2A5B39 , 32'h0194B1B4 , 32'hFFFE8BF0 , 32'hD8D33500 , 32'hFFFC4225 , 32'hEEA7DFE0 , 32'hFFF9AEFB , 32'hFFFDB772 , 32'hFFFDF67E , 32'h02001474 , 32'hCE7C6100 , 32'h09AF0720 , 32'h0001C385 , 32'h1176A4A0 , 32'h10DB0840 , 32'h00052170 , 32'h00011C7F , 32'hF68C88A0 , 32'hFC049210 , 32'h17BBB360 , 32'hE5C16220 , 32'hFFFA0D87 , 32'hFCA3B6A4 , 32'h0D528890 , 32'hFF515728 , 32'hFFFC32C8 , 32'h0115DBAC , 32'h0615BC78 , 32'hFE1BF004 , 32'h00029B84 , 32'hFDF17704 , 32'h00043005 , 32'hFFFC7B01 , 32'h01C1403C , 32'hFDABAD84 , 32'hF78B7A80 , 32'h1F12BCE0 , 32'h00083C0B , 32'h14786F00 , 32'hFFFC8790 , 32'hBF7DF000 , 32'hFFB82CC5 , 32'h0001AF1D , 32'h2ED96AC0 , 32'h22DE7F80 , 32'h13FE4E00 , 32'h0000763D , 32'h00021E2F , 32'h00041F7C , 32'hF1FC4640 , 32'h0A31F1C0 , 32'h0000BCC3 , 32'hF74D0840 , 32'hF9C12308 , 32'hFFF9240E , 32'h0402BC88 , 32'hFEA2D658 , 32'hFFFBD584 , 32'h1825E780 , 32'hDCFB2CC0 , 32'hF1035900 , 32'hFFFE8AFC , 32'hFFFF97C1 , 32'h155D3EE0 , 32'hFFFB9A4F , 32'hEE3BF180 , 32'hFFFDFE5A , 32'hFDF8E74C , 32'hFE657D4C , 32'h00015BCC , 32'h00013B7C , 32'h0001E363 , 32'hFFFF4354 , 32'hE2A4D500 , 32'hF9015840 , 32'h00001A0B , 32'hDCC46180 , 32'h129692E0 , 32'h07654810 , 32'h000506DB , 32'h00665B5F , 32'hFFFF55FB , 32'h0D6171A0 , 32'hF3EF52B0 , 32'hFFFD9698 , 32'h0CADFB30 , 32'h0000A879 , 32'hFFFD21BE , 32'hEABA4B00 , 32'hE6C05F40 , 32'hFD8F9CA8 , 32'hFFFEEC3A , 32'h03E5D420 , 32'h0002B166 , 32'hFFF8C525 , 32'hFD2F64B0 , 32'hFFFE77CE , 32'hFFFE6C40 , 32'hF5C327A0 , 32'h03BCB358 , 32'h0000641D , 32'hFFFEC65E , 32'hFFFE08DD , 32'h000439A0 , 32'h0000BAB4 , 32'h14B5BAA0 , 32'h0A809CB0 , 32'hFFFCD6CD , 32'hFFFD252A , 32'h07C26518 , 32'hEBCC5A80 , 32'hFFFF6982 , 32'h00030A97 , 32'h2087CE40 , 32'h000021B4 , 32'hFFF92522 , 32'h15B18820 , 32'h00FDC5F5 , 32'h0634A4D0 , 32'h0020276A , 32'h00073189 , 32'hFFFC08DE , 32'h0A312740 , 32'hFFFCF693 , 32'hFFFFAB55 , 32'h02D9AB00 , 32'h0006F013 , 32'h0002F8CA , 32'hE783F5C0 , 32'h0004891E , 32'hFF48B50F , 32'h01D25E10 , 32'hFFFC205A , 32'h00018982 , 32'hFFFE4A21 , 32'h2D3A7140 , 32'h01A600D0 , 32'h077F8BD8 , 32'h270260C0 , 32'hFFFE537C , 32'hF7201C40 , 32'h00016E8E , 32'h00013261 , 32'h11CC3480 , 32'hF43663F0 , 32'h047CC518 , 32'hFFFEC626 , 32'hFC0A4C04 , 32'hFCB6B324 , 32'hCD598340 , 32'h00E3F490 , 32'h0F3950C0 , 32'hFF8742DF , 32'hFE23E578 , 32'h148427A0 , 32'h0001A448 , 32'h0004530D , 32'hFFFE569D , 32'h100AC960 , 32'h0201D548 , 32'h077EAAA0 , 32'h003ACDD3 , 32'h06B87148 , 32'hF5A89E20 , 32'h000176A1 , 32'hD0638400 , 32'hF8F919B0 , 32'hFFFBB552 , 32'h33C66AC0 , 32'hFFFB9F89 , 32'hF9638D78 , 32'hF644BF50 , 32'h00023C79 , 32'hFFFE74BC , 32'h0000151D , 32'hFFFECB7B , 32'hFFF85820 , 32'h0002EFC5 , 32'h04FDEC10 , 32'h2785A880 , 32'hE3425540 , 32'hF5455AB0 , 32'h18EB9260 , 32'hF3E67C30 , 32'h0005DE57 , 32'hFFFFB69C , 32'h000004C8 , 32'hFFFA7EBF , 32'h00022378 , 32'hF5F7FE70 , 32'h0E351AE0 , 32'hEDFC2820 , 32'h0000DC08 , 32'hFFFF8D4C , 32'h0003C6A0 , 32'h0000DA75 , 32'h0CC2F0C0 , 32'hBB8F0080 , 32'h0001A076 , 32'hFFF73E40 , 32'hFFFA95D5 , 32'hE7AB0880 , 32'h1CE885C0 , 32'hF88DF0B0 , 32'h0001B385 , 32'hFFFB6E30 , 32'hFFFCC13C , 32'h0436D938 , 32'h030BA0C0 , 32'hF8310158 , 32'hFFFF6610 , 32'h001D0552 , 32'h00004CC0 , 32'h33411280 , 32'hFFFF6B3F , 32'h1BCD9500 , 32'h0000473D , 32'h4204A880 , 32'hFAD8A7F8 , 32'h0FBBFB60 , 32'h13AA4380 , 32'h0000EC14 , 32'hDFBD4780 , 32'h032A6AB8 , 32'h0001AF4E , 32'hFEDFB1EC , 32'h0000A2C9 , 32'h08926790 , 32'h18A9D4E0 , 32'hF4AF16A0 , 32'hFFFE061C , 32'h0000A13C , 32'hD8DD4800 , 32'h0000AF3B , 32'h20825B40 , 32'h0006F5B6 , 32'hFEAECD28 , 32'hFFFEFF03 , 32'h2BA738C0 , 32'hFFFF5E69 , 32'hFFFF2D88 , 32'h00056397 , 32'hE22BE8C0 , 32'hEE352400 , 32'hFFFACB9E , 32'hFFFDB798 , 32'h000058AA , 32'h00001165 , 32'h198BB500 , 32'hF5BE8DB0 , 32'hEC247020 , 32'hF242C2D0 , 32'hEC3177A0 , 32'h00043018 , 32'h0001E890 , 32'h00007892 , 32'hFA3627B0 , 32'hFFFC6A8E , 32'hFFFC4A39 , 32'h027A2660 , 32'h065C65F8 , 32'h00039580 , 32'h17D609E0 , 32'hE8B5B660 , 32'hFB25DB18 , 32'hF794E7B0 , 32'hFFFA2AFB , 32'hF8ACB8E0 , 32'hF74E0DE0 , 32'hFD96FD5C , 32'h0003E2FA , 32'hEE228A20 , 32'h143A77A0 , 32'hE999A8C0} , 
{32'h12B7F3E0 , 32'h03008304 , 32'h00003022 , 32'h0EA158E0 , 32'hFFFFE9E6 , 32'hF3A61180 , 32'h00036806 , 32'h0002E8CD , 32'h0000DB08 , 32'h00002A82 , 32'hE36B8760 , 32'h1F4E0A80 , 32'hF8E34038 , 32'h00008B95 , 32'h0000A8FD , 32'hE82681E0 , 32'h00019890 , 32'hFC7B1838 , 32'h12DC5EE0 , 32'hFFFB92BD , 32'h00018F0D , 32'h00DF5952 , 32'h0B37E530 , 32'h08989310 , 32'hF20DD3B0 , 32'h0004660B , 32'hF9456288 , 32'h03ED90AC , 32'h0000BFE7 , 32'hFA71D060 , 32'h00002B90 , 32'hE3D1B700 , 32'h000193D2 , 32'hFFFD1ADB , 32'h00012ABC , 32'h2094A880 , 32'h35ECCF00 , 32'hFD04B59C , 32'h000002E9 , 32'h15BEDCE0 , 32'hDF81A040 , 32'h000460AF , 32'h000188E2 , 32'h02742208 , 32'hFD8A6E6C , 32'hF837C798 , 32'hFC0B4A58 , 32'h00036084 , 32'h05FD8AD8 , 32'hD049CA00 , 32'hFFE9A2AD , 32'h00020F69 , 32'h05AD0030 , 32'hEF7E9FE0 , 32'h09C586D0 , 32'h00002486 , 32'h06D41170 , 32'hFFFE0484 , 32'hFFFB645F , 32'hF162E680 , 32'hFBE1C6D8 , 32'hF9FF9AD0 , 32'hF1100150 , 32'hFFFE2D16 , 32'hE2E8E200 , 32'h0000F0D2 , 32'hC628EA40 , 32'h01C4D004 , 32'h0006FDAB , 32'hF3FCA120 , 32'hC119CF40 , 32'h0F2262B0 , 32'h000109A4 , 32'hFFFC171E , 32'hFFFD353E , 32'hDAAF3540 , 32'h0762B5A0 , 32'hFFFFD8F5 , 32'h25926840 , 32'h00DEC7C6 , 32'hFFF37146 , 32'h184DA1C0 , 32'h06C26788 , 32'h00057FB0 , 32'h053487B8 , 32'hC760FF40 , 32'hF5569C60 , 32'hFFFDF67E , 32'h0003C3E5 , 32'hE51234A0 , 32'h00012346 , 32'hF7D56AF0 , 32'hFFFEC6C6 , 32'h03658334 , 32'h009B426C , 32'h00029C56 , 32'hFFFCE944 , 32'hFFFDB248 , 32'hFFFEDD8F , 32'h0AC51ED0 , 32'hF4ABA690 , 32'hFFFB873A , 32'hEB549860 , 32'h076851D8 , 32'hFA0D8250 , 32'hFFF969B0 , 32'hFF0F445A , 32'hFFF9F1D5 , 32'h05D12CE0 , 32'h59E03480 , 32'h0000D2AF , 32'h0F17FE70 , 32'h000064C5 , 32'hFFFB9AF0 , 32'hEDF9E760 , 32'h0F8C6650 , 32'h026370E0 , 32'h000377EC , 32'h195ABC80 , 32'h000287D4 , 32'h00018BE6 , 32'h07501F80 , 32'h00044603 , 32'h00038649 , 32'h111962C0 , 32'h0234F0FC , 32'h00021204 , 32'hFFFA77BF , 32'hFFFF18BC , 32'h0001232D , 32'hFFFF52E9 , 32'hF8288140 , 32'hEFA50340 , 32'h000377C4 , 32'hFFFCD51C , 32'hD20454C0 , 32'hF0749440 , 32'h0001DA04 , 32'h00003D00 , 32'h1C7980C0 , 32'hFFFE96BD , 32'h0002DC2C , 32'h0A90EAD0 , 32'h068AD630 , 32'hF6EE54D0 , 32'h02F632C8 , 32'hFFFCE213 , 32'hFFF8709F , 32'hFD09BC48 , 32'hFFFB9B7F , 32'h0004F657 , 32'hFE22B928 , 32'h0004F6F9 , 32'h0000C685 , 32'hF351AA30 , 32'h0009D8D0 , 32'hFC474994 , 32'h0179A90C , 32'hFFFEF856 , 32'hFFFF2E62 , 32'hFFFA5294 , 32'hEA5EB700 , 32'h05DA8400 , 32'h0D46C320 , 32'h0297A354 , 32'hFFFB3DA2 , 32'h1CC5A8C0 , 32'h0002B23D , 32'hFFFD26BF , 32'h2200CBC0 , 32'h02BCAFE4 , 32'hF48DB340 , 32'h000226C3 , 32'hAE1C8C80 , 32'hFF9CE15F , 32'hF1C3D240 , 32'hDEB1CE40 , 32'h13A16440 , 32'hCF8BE200 , 32'h054A20E0 , 32'hFC54BE1C , 32'h0000C762 , 32'hFFFD3529 , 32'hFFFCB11A , 32'h0E1C3B80 , 32'hF483A4A0 , 32'hFF3C639A , 32'hFDE26D08 , 32'h13AD10C0 , 32'h0F3B1900 , 32'hFFFE893E , 32'h1A9ECA00 , 32'h09B39760 , 32'hFFFF5116 , 32'h056232E8 , 32'hFFFDF8D6 , 32'h188472C0 , 32'h05183330 , 32'hFFFBB35D , 32'h0003E397 , 32'h00038626 , 32'h00022CDD , 32'hFFFE5466 , 32'h0001A511 , 32'hFAB68058 , 32'hFB763A38 , 32'hF03B25B0 , 32'h0781D280 , 32'h02ECFE54 , 32'hF55084D0 , 32'hFFFC1974 , 32'h0002BCEC , 32'h0000987C , 32'h00038713 , 32'hFFFE6BF0 , 32'hF57E1570 , 32'h136D29E0 , 32'h28F08500 , 32'h00028399 , 32'h0004A042 , 32'hFFFCF664 , 32'h0004AC1A , 32'h05232BD0 , 32'hE26A1A00 , 32'h00003A7C , 32'h0002D2EE , 32'h00022397 , 32'hE9E79220 , 32'h1C7115A0 , 32'hE3EA37A0 , 32'h0000998D , 32'h0004ACF3 , 32'hFFFE9F59 , 32'hF74EB520 , 32'hFFD3698A , 32'hF5C15030 , 32'h0001BDBC , 32'hFE66861C , 32'hFFFD3855 , 32'hF6E94FD0 , 32'hFFFFE1E4 , 32'h0EB4D660 , 32'hFFFFD675 , 32'hFD9B8304 , 32'h0A72DF00 , 32'hF6CE6550 , 32'h283C7FC0 , 32'h00022040 , 32'h0330102C , 32'h01A456E4 , 32'hFFFBE7AA , 32'h0DF6A880 , 32'h00036BF1 , 32'hFAA8C148 , 32'hDF9AE040 , 32'h3182BCC0 , 32'hFFFFD1C3 , 32'h00003C60 , 32'hEDD9D320 , 32'hFFFD93B5 , 32'h04A5AFA0 , 32'hFFFF5BAC , 32'h0572A9B0 , 32'hFFFDF57D , 32'h0ABF65B0 , 32'hFFFC5C62 , 32'h00014F48 , 32'hFFFFA850 , 32'hF34C71E0 , 32'h301161C0 , 32'hFFFF1AF2 , 32'h0006090A , 32'hFFFDB5CA , 32'hFFFB8E6F , 32'hF37CF730 , 32'h1F16D600 , 32'hF467F470 , 32'hE1331220 , 32'h154B60C0 , 32'hFFF978D6 , 32'hFFFB2C40 , 32'h0001CC8B , 32'h0C4D2D40 , 32'h00025BFC , 32'hFFFF0D35 , 32'h04B01C18 , 32'h33E55940 , 32'hFFF86998 , 32'hE037BC20 , 32'h0A3BE040 , 32'hF72E7BB0 , 32'hF1F73570 , 32'hFFFE099F , 32'h032702A8 , 32'hF2B91070 , 32'hFE96DB74 , 32'h000997DA , 32'hE4A95280 , 32'hE33F3AA0 , 32'hE65E3860} , 
{32'h294EFB80 , 32'h088424D0 , 32'hFFFABD4B , 32'hFAC34AF0 , 32'hFFFC5DDF , 32'h0F396AF0 , 32'hFFFCEDB7 , 32'hFFFAEAC6 , 32'h0003A3AE , 32'h00015F32 , 32'h0DC0B350 , 32'hF0BEBAD0 , 32'hF47869E0 , 32'h0001486D , 32'h00020485 , 32'h10C56BA0 , 32'hFFFFF3B3 , 32'h13756080 , 32'hF7FF47F0 , 32'hFFFEE01C , 32'hFFFA1243 , 32'hFFC115B8 , 32'hEE25A3E0 , 32'h131B7480 , 32'h11F806C0 , 32'h000098E8 , 32'h012B46B8 , 32'hFF9D48DC , 32'h00000431 , 32'h2FA98080 , 32'hFFFBCD49 , 32'h0471DBD0 , 32'hFFFC5E20 , 32'h0000611B , 32'h00059126 , 32'hDE0D0DC0 , 32'hCCE86500 , 32'hD7464740 , 32'hFFFE17AD , 32'h13C58B60 , 32'hDE598B00 , 32'h000049C7 , 32'hFFFF17BE , 32'h0D0BA870 , 32'h39139940 , 32'hCCBABE00 , 32'h0291918C , 32'h00012A1B , 32'h10BD35C0 , 32'h0E03E470 , 32'hFE311CD8 , 32'hFFFDD598 , 32'hF57993C0 , 32'h033C8A74 , 32'hED5D1FE0 , 32'h0004EA21 , 32'h00B8A98B , 32'hFFFE0BF6 , 32'hFFFEEB6B , 32'h06A764C0 , 32'hFC235774 , 32'h1677FBA0 , 32'hE9F50F20 , 32'hFFFDB1D2 , 32'h1B153AC0 , 32'h000027CB , 32'hD28CDE00 , 32'h012F0610 , 32'hFFFBC183 , 32'hF9164F18 , 32'hC72BD080 , 32'hE38C86C0 , 32'hFFFFA97A , 32'h0001C71C , 32'hFFFE3CDC , 32'h115DDEA0 , 32'hF4951F60 , 32'hFFFD27CA , 32'hEF0BCE80 , 32'h05E55760 , 32'h0000CCD3 , 32'h295EB600 , 32'h04126F10 , 32'h000105A1 , 32'h0FF32CB0 , 32'h078ED200 , 32'h0B66DE90 , 32'hFFFF6C13 , 32'hFFFFF298 , 32'h0CDB04D0 , 32'hFFFD0E68 , 32'h02716CF0 , 32'hFFFEC60C , 32'hEB6DE300 , 32'h00AD7A71 , 32'h0001FE21 , 32'hFFFEFA40 , 32'hFFFBF614 , 32'hFFFF7FE4 , 32'hE5450D20 , 32'hFFD13806 , 32'h0004AD8D , 32'hEA5762C0 , 32'h06C68358 , 32'h042BC870 , 32'hFFFE33FB , 32'h0065FB1E , 32'h000363C7 , 32'h0E715130 , 32'hE4606FC0 , 32'hFFFE7363 , 32'h17ADB760 , 32'h0001887D , 32'h00026FD1 , 32'hF436B380 , 32'hF2DDA020 , 32'h026F4B44 , 32'hFFFC2AD0 , 32'h0E2B1990 , 32'h00012BEF , 32'h0003C0D9 , 32'h07CA1968 , 32'h0004CE4E , 32'hFFFB3B02 , 32'hEF902B20 , 32'hEFD4C480 , 32'hFFFB52E9 , 32'h0006BE98 , 32'hFFFB53DF , 32'hFFFA35DB , 32'h0002934A , 32'h077DEFC0 , 32'hED8CB560 , 32'hFFFD7377 , 32'hFFFE1CFF , 32'h178D53A0 , 32'hF9365E90 , 32'hFFFF82F8 , 32'h0000D124 , 32'h1A68DCE0 , 32'h000001A5 , 32'hFFF89123 , 32'h03D50764 , 32'h074A3E80 , 32'hFE79C400 , 32'hFBA32FF8 , 32'h0000599B , 32'hFFFFDC95 , 32'h009E244F , 32'hFFFD54B4 , 32'hFFFD7A4A , 32'hFADD1910 , 32'h000094FA , 32'h0005E33F , 32'h17926940 , 32'hFFFE5F14 , 32'hF32E5270 , 32'h027FDBF8 , 32'hFFFFF8EA , 32'h000043F3 , 32'hFFFE0671 , 32'hF80645F0 , 32'h0502D728 , 32'h08085A70 , 32'h084B21F0 , 32'h00007C6F , 32'hEB7B8640 , 32'hFFFA71CB , 32'h0003A652 , 32'hF5334CC0 , 32'h05EBE7E0 , 32'h002165A7 , 32'h0002B737 , 32'h0B3D0670 , 32'h016B28E0 , 32'h01C40D28 , 32'h0848E8B0 , 32'hF0B955B0 , 32'hA9216080 , 32'h01413818 , 32'hF84ED720 , 32'h0003F2AE , 32'h00014D72 , 32'hFFFEA4BF , 32'hFC6FAA8C , 32'h2AF48700 , 32'hF80C0BE8 , 32'hFE467DC0 , 32'h047FFF88 , 32'hF3072710 , 32'h0008CE55 , 32'h12452C60 , 32'hF3128580 , 32'hFFFEB71C , 32'hDFD7E040 , 32'h00025B78 , 32'hF59962E0 , 32'hE90E2420 , 32'h00031067 , 32'h0000C901 , 32'h00010DF7 , 32'hFFFAEBB2 , 32'h0006A8C7 , 32'hFFFCEEC6 , 32'h188E1440 , 32'hF5982750 , 32'h440FE700 , 32'h002F21ED , 32'hF511D890 , 32'hF63D5080 , 32'h000263E7 , 32'h00013416 , 32'hFFFF42CC , 32'h0002B3CB , 32'hFFFD83DE , 32'hFCDBB860 , 32'hEAC68680 , 32'hE5F806E0 , 32'h0001C97E , 32'h00042057 , 32'hFFFFC442 , 32'hFFFDC5D4 , 32'hFEC1E4B4 , 32'hD4021B80 , 32'hFFF952D9 , 32'hFFFE11D4 , 32'hFFF82E38 , 32'hDA940D40 , 32'hF72BB780 , 32'hEA0BBD60 , 32'h0002FC53 , 32'hFFFE64BE , 32'hFFFD4526 , 32'h09D2AB60 , 32'hF1AFA600 , 32'hCE92CA40 , 32'h0001FF90 , 32'hFDFE103C , 32'h000060C9 , 32'h06BB3870 , 32'hFFFACC9C , 32'hD143BBC0 , 32'h00047AE1 , 32'h076C0EC8 , 32'hFBB5DC98 , 32'h2E0FC480 , 32'hE0651AC0 , 32'hFFFBB50A , 32'hF1968C90 , 32'hFE8018CC , 32'hFFFEA734 , 32'hF4C142E0 , 32'h0004238C , 32'h05FA6748 , 32'h0F4D4890 , 32'h015F9FFC , 32'hFFFEBBF8 , 32'hFFFE08C4 , 32'hDF5C3A00 , 32'hFFFDB0C5 , 32'h2260AB00 , 32'hFFFF187F , 32'hFFE6FFFD , 32'hFFFF05CB , 32'hFD08EACC , 32'h0003674F , 32'h00006381 , 32'hFFFE51CC , 32'h11AEDF80 , 32'hF61EE3F0 , 32'h0002C50E , 32'h000132F6 , 32'hFFFFE5EB , 32'hFFFC5F2D , 32'hDB86A000 , 32'h0A968AB0 , 32'hE99050A0 , 32'h1E3CDF40 , 32'h06B81EF8 , 32'hFFFFDA49 , 32'h0002BA2B , 32'hFFFCF56C , 32'hFF1D8750 , 32'h0002ED87 , 32'h0004E45C , 32'hF2CCBD70 , 32'h1A820E40 , 32'hFFFF8AA3 , 32'hDDA48A80 , 32'h03ECC870 , 32'h0DC1DD90 , 32'h07340940 , 32'h0003FC82 , 32'hFD7E1964 , 32'hEED5F7E0 , 32'hFECFCAF0 , 32'h0000808B , 32'h1A7D1700 , 32'hBCC63800 , 32'h057370D8} , 
{32'h03730728 , 32'h0E47E440 , 32'h00031E89 , 32'h0D8498D0 , 32'hFFFF0B7C , 32'h052E2D50 , 32'hFFFB9C28 , 32'h000092E1 , 32'h00026D1F , 32'hFFFD136C , 32'hF174DB00 , 32'hFDDE6620 , 32'h126C9FE0 , 32'h0001F84B , 32'hFFFF9485 , 32'hFF17A556 , 32'h0001AD2A , 32'h0E78A5E0 , 32'hFC962FC4 , 32'hFFFD2114 , 32'hFFFF2DFE , 32'hF7F87000 , 32'h00EA52F7 , 32'h131CE5E0 , 32'h275A7B40 , 32'h0000E895 , 32'h00D5C883 , 32'h00EEDACF , 32'hFFFCA973 , 32'h1A1AD800 , 32'h0006A493 , 32'h2C800280 , 32'hFFF7A6BA , 32'hFFFFAB5B , 32'hFFFDCA6A , 32'hEA7AA2C0 , 32'h385F1240 , 32'hC7CE1800 , 32'h00002752 , 32'hCFE580C0 , 32'hFDDE606C , 32'h000016FD , 32'h000026D7 , 32'h09A0A010 , 32'h30D4F200 , 32'hE3FC2040 , 32'hE68C0740 , 32'hFFF92BFF , 32'hFEF134C4 , 32'hDF0CCA00 , 32'h00BF6D24 , 32'h0001C931 , 32'h02A80D94 , 32'h18DCC300 , 32'hE6E5CDE0 , 32'hFFFBA071 , 32'h022191BC , 32'hFFFFFB3B , 32'h000330A0 , 32'hFA4D8BB0 , 32'hFD4BCA60 , 32'hF0A8F070 , 32'hDF429E00 , 32'hFFFFB23B , 32'hEDAD6560 , 32'hFFFE06B2 , 32'hEB8E0300 , 32'h007A5CE9 , 32'h000194F8 , 32'h02A74F90 , 32'hF10576C0 , 32'hF33CEF30 , 32'h00047DA9 , 32'h0002CDC7 , 32'h0000C1AC , 32'hFDE7666C , 32'h0A78C5E0 , 32'h00029A63 , 32'h068CB298 , 32'h03DBEF4C , 32'hFFFD4D51 , 32'hF8B3AF48 , 32'hEAE26720 , 32'h00013DCD , 32'h23D15BC0 , 32'hF820A2B0 , 32'h0CEDC660 , 32'h00050A85 , 32'h00003900 , 32'h125F3300 , 32'hFFFCDA4C , 32'h16616640 , 32'h0000DF42 , 32'h1239EC80 , 32'hFEF99364 , 32'hFFFD597F , 32'h0001F371 , 32'h000002C1 , 32'h000323F8 , 32'hF18E8DF0 , 32'hFD90F99C , 32'hFFFDA2E0 , 32'hFA74D938 , 32'h0F414DA0 , 32'h02A38650 , 32'h0000F6C1 , 32'h006DCB99 , 32'hFFFB7B58 , 32'h24DE7F40 , 32'h0F4627E0 , 32'h00002C71 , 32'hE2DC4E80 , 32'h0002593B , 32'h00040E17 , 32'h0951D830 , 32'h054C2BA8 , 32'hF9F476D8 , 32'h00059F6A , 32'h02BCF328 , 32'h0001265E , 32'h000487F4 , 32'h01D01AD4 , 32'hFFFC40C4 , 32'hFFFD282F , 32'h1A8CDD80 , 32'h05D28BB8 , 32'hFFFE0EA1 , 32'hFFFBEE29 , 32'h0004647E , 32'h0001AC2A , 32'hFFFE5534 , 32'h130EB0E0 , 32'h0A9513A0 , 32'h00001F4A , 32'hFFFD2DC1 , 32'hEFC198E0 , 32'hEBDF9100 , 32'hFFFDD50C , 32'h00056ECB , 32'h013092A0 , 32'h00019F48 , 32'hFFFF983F , 32'hFD603C74 , 32'h01426860 , 32'h0318F750 , 32'hF7CDCFC0 , 32'hFFFF8F5A , 32'hFFFAB8E2 , 32'hFBA41000 , 32'h0003FD90 , 32'hFFFFA69E , 32'h0416D260 , 32'hFFFE9E98 , 32'h00010FD8 , 32'h07A4AE98 , 32'h00025DDB , 32'h04CC5260 , 32'hFF7CB2E5 , 32'hFFFA7108 , 32'h00068FEC , 32'h00008B9E , 32'hF225E5D0 , 32'h079C1260 , 32'h0F0D40E0 , 32'h0DF93830 , 32'h0002556F , 32'h2F7BBE40 , 32'h0001C931 , 32'h0001087A , 32'hE2287C00 , 32'hFFEBA218 , 32'hFE19D884 , 32'h0000932D , 32'hFFBC4580 , 32'h05228D78 , 32'h17C85480 , 32'h03D45ACC , 32'hE1F353E0 , 32'hE0439A40 , 32'h03E59AB8 , 32'hFF84BCCD , 32'hFFFF9C6C , 32'h0000669D , 32'h00023F21 , 32'hEB4FDBE0 , 32'h06F77D88 , 32'hF85994B0 , 32'hFDCDEA74 , 32'hFC16AAA8 , 32'h09B78DE0 , 32'hFFFB6806 , 32'h06503188 , 32'h06130578 , 32'hFFFE54CB , 32'h4B53DC80 , 32'h000081D9 , 32'hFAA8EB18 , 32'hF5EB4E30 , 32'h00022DD2 , 32'h0000E37A , 32'hFFFEF171 , 32'hFFFF9BA7 , 32'hFFFBAF6A , 32'h0000B259 , 32'hF2F1D4C0 , 32'h1F3F10E0 , 32'h2D3C4480 , 32'h16E82260 , 32'h0063D978 , 32'hF5511C00 , 32'h0000E343 , 32'h00006C18 , 32'h00016AFA , 32'hFFFDA649 , 32'h00047429 , 32'h040FA840 , 32'h05F6C178 , 32'hF0C99FC0 , 32'h0006B0F7 , 32'hFFFF00B0 , 32'hFFFA16C6 , 32'hFFFFCC7E , 32'h03273BA4 , 32'hF6564F60 , 32'hFFFC1DD6 , 32'h000110C6 , 32'h00032F3A , 32'h19D3B0C0 , 32'h3C9D2240 , 32'h273196C0 , 32'h000062AB , 32'h00044047 , 32'hFFF8D0C4 , 32'h0D12C170 , 32'h09044D20 , 32'hFCDD4DF8 , 32'h0000FBEB , 32'h02E36848 , 32'h00013210 , 32'hF910BF88 , 32'h0003985F , 32'hFC111408 , 32'h00043753 , 32'hEA43C140 , 32'h08043EB0 , 32'h167D3B80 , 32'h19EF7EE0 , 32'hFFFF5D51 , 32'h06AD0920 , 32'hFE946C84 , 32'h000127CD , 32'h12EA2FA0 , 32'hFFFE000D , 32'h08A9F240 , 32'h35210340 , 32'h03CF2800 , 32'hFFFFCD9A , 32'h0000AB56 , 32'hECDEE840 , 32'hFFFE2FF6 , 32'hEBF06FC0 , 32'h00005B5C , 32'h0213F008 , 32'hFFFCE538 , 32'hEFE92340 , 32'hFFFB0EA4 , 32'hFFFEC875 , 32'hFFFFE50F , 32'h1B708DA0 , 32'h0C6FBD70 , 32'hFFFD1A32 , 32'hFFFEE9D1 , 32'hFFFE41DC , 32'hFFFDAAD0 , 32'h68464F00 , 32'hEC8F37E0 , 32'hFC70F618 , 32'hF8FF8300 , 32'hF67132F0 , 32'h00001347 , 32'h00007AFC , 32'h000338ED , 32'h04ED4A88 , 32'hFFFCF611 , 32'h00025FE5 , 32'h056D4AB8 , 32'hF534EDD0 , 32'hFFFEC06A , 32'h22A82980 , 32'h02A79C88 , 32'h01FFAA64 , 32'h1EEDB000 , 32'h0000AAF7 , 32'hF3C01520 , 32'h0BBAD520 , 32'h010761FC , 32'h000151AE , 32'h12C78120 , 32'h5419C680 , 32'h13F8E940} , 
{32'h008380FB , 32'h08D6ACC0 , 32'h00002499 , 32'hF6145290 , 32'h00061708 , 32'h01A041AC , 32'hFFFB0293 , 32'h000091DF , 32'hFFF99F06 , 32'h000821AD , 32'h0CD65600 , 32'h1235DFC0 , 32'h1387ACC0 , 32'h00030128 , 32'h00010A6E , 32'hEE744880 , 32'hFFFF9D3C , 32'h0A5E6F00 , 32'h08D33850 , 32'hFFFDFD0D , 32'hFFFFCD17 , 32'h03FF4634 , 32'h1B9C4EC0 , 32'hFBCEAB68 , 32'hD60DD300 , 32'hFFFFA999 , 32'h026BB8EC , 32'h08FBE9D0 , 32'h000402CB , 32'hD3DB9AC0 , 32'h000169FB , 32'h1500E580 , 32'hFFFFED42 , 32'h0006ABC7 , 32'h00010802 , 32'hF89F27E0 , 32'hC1194EC0 , 32'h092E0030 , 32'h0002F764 , 32'hF4B402A0 , 32'h047F06F8 , 32'h0000976F , 32'hFFFE4CEA , 32'hFD5D6BD8 , 32'hFB232548 , 32'hDAF68E80 , 32'hFDA5BEB8 , 32'h0002620A , 32'hFBC4E5B8 , 32'hF875BE50 , 32'h04325CB0 , 32'hFFFCB4F7 , 32'h0ED92B60 , 32'hF337A450 , 32'h22176240 , 32'h0002D631 , 32'h026053E0 , 32'hFFFF90B5 , 32'h000462E6 , 32'hFDE50320 , 32'h04169870 , 32'hF8F9DB20 , 32'hD6C740C0 , 32'hFFFE8A43 , 32'hE67F9160 , 32'h000234AC , 32'h0C236380 , 32'hFFFF72C2 , 32'h000517EB , 32'hE7489220 , 32'hFD0759E0 , 32'hF9BAC2C8 , 32'h0000E9C6 , 32'h00005F87 , 32'hFFFD4129 , 32'h0B1706D0 , 32'h06382BB0 , 32'h00023F1E , 32'h27110C80 , 32'hFD9D5E3C , 32'h00033485 , 32'h421E4080 , 32'hE90114A0 , 32'hFFF78677 , 32'h016727C4 , 32'hF4A70760 , 32'h03EF7CE0 , 32'h0001141D , 32'h00023079 , 32'hF46427E0 , 32'hFFFD9354 , 32'h0B2FCC20 , 32'hFFFF6AF0 , 32'hFE65AFD0 , 32'h0066D7F4 , 32'h0001C2E2 , 32'h00003B7D , 32'hFFFF1B65 , 32'h0005FF50 , 32'h017AE950 , 32'hFBD054F8 , 32'h0008AAB2 , 32'hDA8232C0 , 32'hE1E76BA0 , 32'h0C299E10 , 32'h0000ABB0 , 32'hFEB3F7B4 , 32'h0002E9C0 , 32'hF0BAA100 , 32'h0DD916C0 , 32'hFFFD04EE , 32'h042C0320 , 32'h0001DE94 , 32'hFFFBBE2B , 32'hEE70FAA0 , 32'hF22EE720 , 32'h0241E5B8 , 32'hFFFD6B96 , 32'hFEED8E84 , 32'hFFFE9802 , 32'h0000D83D , 32'hFBD19830 , 32'hFFFEE5AC , 32'hFFFFD0AF , 32'h0D03C2A0 , 32'h26F89540 , 32'h00001B2C , 32'hFFFF15DF , 32'hFFFBE562 , 32'h0002FB1A , 32'hFFFEE961 , 32'hE744FB40 , 32'hF9808F78 , 32'h00003578 , 32'h000301FC , 32'h42ED2500 , 32'h110603E0 , 32'hFFFA6E92 , 32'h00030DC1 , 32'h0A7BA720 , 32'hFFFFB0B0 , 32'hFFFC7672 , 32'hFDCA6708 , 32'hF8435AE8 , 32'h02FB2DA4 , 32'hFC97B08C , 32'hFFFD643F , 32'hFFFF05BA , 32'hFDD2048C , 32'hFFFDB3C3 , 32'h00035724 , 32'hF4E984B0 , 32'hFFFD2CB0 , 32'h0000F9B3 , 32'hD8E4F940 , 32'h0001C53F , 32'hFFA89B0A , 32'h029F1C6C , 32'hFFFCB2F9 , 32'h000323CF , 32'h0003A518 , 32'h0FB7E170 , 32'hEE3445E0 , 32'hEFFE5EE0 , 32'h051B44F0 , 32'h0002DA58 , 32'h1591FF20 , 32'h0001CFB2 , 32'h00054BB3 , 32'hF019F010 , 32'hF769DF90 , 32'hF66325F0 , 32'hFFFDCBB6 , 32'hD8DE25C0 , 32'hF7C4D8E0 , 32'h15C653C0 , 32'h165B1460 , 32'h31DB69C0 , 32'hFE9A9A48 , 32'h026C2E28 , 32'hE39ABE80 , 32'hFFFBF9E3 , 32'h0001E9F2 , 32'h00026F0B , 32'hF0A131A0 , 32'h26E5BF40 , 32'h0CCC7A60 , 32'hFD4276C4 , 32'hFEBEC03C , 32'hF43904E0 , 32'h0001461A , 32'hDFBB2000 , 32'hF7034C40 , 32'hFFFED470 , 32'hF6C3AA20 , 32'hFFFF5BAF , 32'hF94E90D0 , 32'hF14255B0 , 32'h00005FEA , 32'hFFFEEF64 , 32'hFFFDAAFE , 32'h0000E670 , 32'h000292A8 , 32'h00008B86 , 32'h07DC1528 , 32'h076010C8 , 32'h17D7FF60 , 32'h00180C49 , 32'h10AFF040 , 32'h02823F04 , 32'hFFFDAF7C , 32'hFFFCCBAD , 32'hFFFDCBC4 , 32'h00058962 , 32'hFFFF9C05 , 32'hF8434CF0 , 32'hFDDEF7A4 , 32'h16212C60 , 32'h0001075E , 32'hFFFFCD50 , 32'h0000BCE2 , 32'hFFFE1D5A , 32'h07FEAEF0 , 32'h1764E720 , 32'hFFFF41F9 , 32'h0004C1E5 , 32'hFFFDC939 , 32'h302DBD80 , 32'h06A84D70 , 32'hE5EE35C0 , 32'h0001F2C6 , 32'hFFFE6964 , 32'hFFFED4DC , 32'hE276EA40 , 32'hFBD27FE0 , 32'hD7A998C0 , 32'h00012B80 , 32'h02B30DBC , 32'hFFFE9E46 , 32'h093A9E70 , 32'hFFFD74E7 , 32'h34D0A1C0 , 32'h000520DF , 32'hF2715510 , 32'hFDB644E8 , 32'hF4B247A0 , 32'h47DB6D80 , 32'hFFFFA4BA , 32'hE71081A0 , 32'hFFE6B3DD , 32'h0000E0ED , 32'h0EEEA490 , 32'hFFFFA17B , 32'h020ACC8C , 32'h28B00740 , 32'hF357D820 , 32'hFFFAA62F , 32'hFFFDB1B1 , 32'h0BDEB490 , 32'hFFFA0A0C , 32'hEBEF9260 , 32'hFFFD6CA5 , 32'h031B97D4 , 32'hFFFF0C95 , 32'hE8D72C20 , 32'h0000918D , 32'hFFFBC71E , 32'h0002BA8F , 32'hF32D6A40 , 32'hF9536538 , 32'hFFFFBC39 , 32'hFFFBF993 , 32'hFFFADE6E , 32'hFFFE80C6 , 32'hFBB90B38 , 32'h00E967AA , 32'h03DE87A0 , 32'h2BA9F8C0 , 32'hE690DCC0 , 32'h0002052C , 32'hFFFD3EB9 , 32'h00010ABA , 32'hFD05C1BC , 32'hFFFB0F38 , 32'hFFF96CC9 , 32'h041DE690 , 32'hFA7DBBE8 , 32'h0000346C , 32'h28AD92C0 , 32'h02BA2E38 , 32'h006220BB , 32'hFA1AAE20 , 32'hFFFA9130 , 32'h086BC6C0 , 32'h144C0CE0 , 32'hFB755AE8 , 32'h00010D03 , 32'h631B6580 , 32'hF37113E0 , 32'hD4970880} , 
{32'hF21F0190 , 32'h0AE83C60 , 32'h00044657 , 32'hC2069F00 , 32'h000092D4 , 32'hF4EDF0F0 , 32'h00025DA5 , 32'h00024E7D , 32'h00036B95 , 32'h0000854E , 32'hE9DD0CC0 , 32'h1C8142A0 , 32'hF1F04D60 , 32'hFFFE46A1 , 32'hFFFD66FB , 32'h019B1DDC , 32'h0000EEFA , 32'h52191980 , 32'h0183B388 , 32'h0007449B , 32'hFFFFD1DC , 32'h0BA47470 , 32'hFC47E518 , 32'hFD2D51B4 , 32'hF00A0120 , 32'h0002F51C , 32'h05270748 , 32'hFCCD3A64 , 32'h000455E9 , 32'hF4242890 , 32'hFFFFA68E , 32'h0EACD520 , 32'h000155BF , 32'h0003EEC5 , 32'hFFFD4009 , 32'h18A957E0 , 32'hF55787C0 , 32'hE9B97760 , 32'hFFFEF70A , 32'h17AB0BA0 , 32'hFB4F1F58 , 32'h00020533 , 32'hFFFFCD37 , 32'h01BE81AC , 32'h03B21768 , 32'h29A1CC00 , 32'h0702E3B8 , 32'h0001E824 , 32'h07E6A7A0 , 32'h101F6A60 , 32'h003D30F5 , 32'h0007CC33 , 32'h025D35EC , 32'h08399550 , 32'hEF915D60 , 32'h000359E4 , 32'h0224694C , 32'hFFFD05BE , 32'hFFFFD957 , 32'hF5E2EDA0 , 32'h01080660 , 32'hF6815B10 , 32'hF69BB600 , 32'h0000DA63 , 32'hEEDE4580 , 32'h000015F4 , 32'hC69A8780 , 32'h04B3D860 , 32'h00001A04 , 32'h01A16BC8 , 32'hEB4065E0 , 32'hFDA8BA24 , 32'h0003475D , 32'hFFFF699E , 32'hFFFE04A2 , 32'hD86EB200 , 32'hFB9F9E50 , 32'h0008D864 , 32'h14E0A700 , 32'h03B6B688 , 32'h00003B10 , 32'hDD66A200 , 32'h096AC520 , 32'h000022AF , 32'h02A409E8 , 32'h1585FD40 , 32'h01E85204 , 32'h00068DE1 , 32'h0001973E , 32'hE9190320 , 32'h0000D68D , 32'h03C521AC , 32'h0001C84C , 32'hF839C970 , 32'h01941010 , 32'hFFFB58E7 , 32'h0004037E , 32'h00012EF5 , 32'hFFFD771E , 32'h0DDBA9E0 , 32'h0D3C8940 , 32'hFFFE4F69 , 32'h10F1BA00 , 32'hFEB8CC34 , 32'h07114860 , 32'h000281D6 , 32'h00171916 , 32'h0000994C , 32'hFD32658C , 32'h004ADEE8 , 32'h00032BD2 , 32'h076C4BA8 , 32'hFFFF5621 , 32'hFFFEA1AC , 32'hF1D26AA0 , 32'h15C452A0 , 32'h03DF4824 , 32'h000468F6 , 32'h065B6580 , 32'hFFFC8976 , 32'hFFFF815E , 32'h0160E3C8 , 32'hFFFD5FCE , 32'h00029DFE , 32'h45BCBB80 , 32'h2B49C540 , 32'hFFFEA84F , 32'hFFFFF5EE , 32'hFFF8BE4F , 32'h0004E9C1 , 32'hFFFFEE7F , 32'h00BFAE78 , 32'h0E1DBED0 , 32'hFFFE9268 , 32'h00010C81 , 32'hFFC1426D , 32'h0634A348 , 32'hFFFDCC24 , 32'hFFFEE7FF , 32'h10478FC0 , 32'h00031C54 , 32'h000453DC , 32'hFE2791B0 , 32'hF57A4620 , 32'h02973FE8 , 32'hFEA2FED8 , 32'hFFFF0199 , 32'hFFFE8EA0 , 32'hF8620A40 , 32'h00043F6D , 32'h0002D7DB , 32'hFD85F2B8 , 32'hFFFA65E7 , 32'hFFF74F09 , 32'hFEB820A0 , 32'h000739D3 , 32'h1E798380 , 32'hFE0E0A28 , 32'hFFFFE9DD , 32'h0001A0A3 , 32'hFFFDA0F8 , 32'h0719C790 , 32'hFE047068 , 32'h06E03FF0 , 32'h1AD0AEC0 , 32'hFFFFC45A , 32'hA2D44280 , 32'hFFFF0D68 , 32'h0000F32E , 32'h169C4840 , 32'h13DDAA60 , 32'hFFFE7B22 , 32'hFFFEF7DB , 32'h441D4F00 , 32'h003985C2 , 32'h160929E0 , 32'h19D34E60 , 32'hE7570B60 , 32'h07715738 , 32'hFB165508 , 32'h08E39CF0 , 32'h0008AB62 , 32'hFFFBE1DB , 32'hFFFFE5BF , 32'h0F12EC20 , 32'h3CC7AEC0 , 32'h04BF40B0 , 32'hFFDCA5AE , 32'h029B3D98 , 32'h0C44D840 , 32'h0000A3AD , 32'hE94D20C0 , 32'h218E3FC0 , 32'h0000E0EC , 32'h1F15CDC0 , 32'h000536D2 , 32'h08DDD1A0 , 32'hF8F75CA0 , 32'hFFFF70C8 , 32'h0004916A , 32'h00032C94 , 32'hFFFCB2BE , 32'h0000712E , 32'h00053AFF , 32'hF6B9C950 , 32'hFB6326A8 , 32'h0225E988 , 32'hFC330604 , 32'h01567064 , 32'hFBF5F518 , 32'hFFFE164E , 32'h0006BBEC , 32'h000121B7 , 32'h00021A3B , 32'h0003332E , 32'h08F00DB0 , 32'h08D63B30 , 32'h51F35F80 , 32'hFFFEDFEC , 32'h00011526 , 32'hFFFE9BD7 , 32'h0005E9D0 , 32'hF04FAA30 , 32'hDE2083C0 , 32'hFFFFD776 , 32'hFFFC28F4 , 32'h0003FD9B , 32'hF4057DE0 , 32'h0CC21660 , 32'hE7D37660 , 32'h000555CE , 32'h00005011 , 32'hFFFF539C , 32'h00FA085D , 32'hFFE27AF0 , 32'hFF0F8A76 , 32'hFFFFC7C9 , 32'hFB7633D0 , 32'hFFF8D3CA , 32'h14F46880 , 32'hFFFE2D9E , 32'hE61008C0 , 32'hFFFDFC6E , 32'hD31A8500 , 32'hFDDFF538 , 32'h0E7D0BC0 , 32'h11D428C0 , 32'hFFFEFC9B , 32'h0D16B050 , 32'h00253DD7 , 32'hFFFCB458 , 32'h15E29960 , 32'h00009A88 , 32'hF6DD8460 , 32'hCF5C8980 , 32'hD6398480 , 32'hFFFFF1C5 , 32'h0001A825 , 32'h02724B04 , 32'hFFFBF997 , 32'hDF485E40 , 32'hFFFCF606 , 32'hFD9D564C , 32'h000670E7 , 32'hEEF8C9E0 , 32'h0001C13A , 32'h0001F224 , 32'h0002B8A0 , 32'h1F85DC20 , 32'hFF78C71B , 32'h00052E4E , 32'hFFFFA0EB , 32'h0003C03C , 32'hFFFF2B84 , 32'hF4169BF0 , 32'hF5FF9040 , 32'h16263560 , 32'hF4223320 , 32'hFFFF6F85 , 32'hFFFE6CD2 , 32'h000181A5 , 32'h0001B97E , 32'hF95E91F8 , 32'hFFFDFCAF , 32'h00035818 , 32'hFECA90E4 , 32'hD4D61BC0 , 32'hFFFCFA1F , 32'hF0605D30 , 32'hF88A36B8 , 32'hF7D7AF10 , 32'hFC9AA888 , 32'h0001BCD6 , 32'h0BB57C30 , 32'hFABE8B10 , 32'h04AA2A70 , 32'hFFFF1493 , 32'h1B66A780 , 32'h051ED4E8 , 32'h09066A30} , 
{32'h038E021C , 32'h122F51A0 , 32'h0000C5C7 , 32'hEE6C6240 , 32'h00021D9C , 32'hF664A2A0 , 32'h000555CD , 32'h0003F6B7 , 32'h00054CF0 , 32'h00021905 , 32'h0FC5BF50 , 32'hE3F9EC80 , 32'hF6235750 , 32'hFFFDAA4D , 32'hFFFEFE96 , 32'hC5168340 , 32'h00029A53 , 32'hB9C21C80 , 32'h1A4F7120 , 32'hFFFE89A0 , 32'hFFFAD3EF , 32'h02933CF4 , 32'hEFB15360 , 32'hF3B82400 , 32'hD0A40B00 , 32'hFFFE8010 , 32'h01597E64 , 32'h0033433D , 32'hFFFF821D , 32'hE6DDDF60 , 32'hFFFB8B0C , 32'hF8F83358 , 32'hFFFAF3F6 , 32'hFFFEB0B2 , 32'hFFFAE131 , 32'h0DFC8EB0 , 32'h2D7D4540 , 32'h11D02500 , 32'h00053651 , 32'h0A2EAFF0 , 32'hEDD09FA0 , 32'h00042BE5 , 32'h0000E2A6 , 32'hFE61531C , 32'h287D4C40 , 32'hE8246240 , 32'hFA852D18 , 32'h000052C3 , 32'hE76B01C0 , 32'hF986DAA0 , 32'h018524CC , 32'hFFFDF218 , 32'h0906A320 , 32'hE3C11EA0 , 32'hFD0B2F50 , 32'hFFFF9439 , 32'h01D370A4 , 32'hFFFF666F , 32'h0002DEED , 32'h06F086B0 , 32'hFC09E618 , 32'hF738CDB0 , 32'hD0CDCA40 , 32'h0001FA70 , 32'hE3957AE0 , 32'hFFFC8EA2 , 32'hE11323A0 , 32'hFCF51680 , 32'h0004E12A , 32'h4FBC6E00 , 32'hFF29A49E , 32'hEB823600 , 32'h0000E78F , 32'hFFFFDC44 , 32'h00014855 , 32'hFEB02C94 , 32'h02C225FC , 32'h00024D2C , 32'h1D0E7280 , 32'hFCDAEE10 , 32'h0002784C , 32'h099BD240 , 32'h125B6F00 , 32'h000182DC , 32'hFFCFFE1D , 32'h04C327C8 , 32'hFD95C590 , 32'h0001C4B3 , 32'hFFFDC5A8 , 32'h415CC400 , 32'h0003A05D , 32'h00EB04FA , 32'hFFFAD78F , 32'h0625AD28 , 32'h0087587E , 32'h00048706 , 32'h000482B6 , 32'hFFFD2509 , 32'hFFFF4328 , 32'h0B2B5290 , 32'h02BC7CE8 , 32'h0001D4E9 , 32'h10052880 , 32'h27CED5C0 , 32'h0AEC9240 , 32'h0000DF3E , 32'h00268020 , 32'hFFFC8626 , 32'hF2DE42C0 , 32'h045A33C8 , 32'h0000B534 , 32'h51045E00 , 32'hFFFEB3E6 , 32'h0002EE09 , 32'h12C81E80 , 32'h0155B24C , 32'hF93DE568 , 32'h000013A0 , 32'h17F79F40 , 32'h0001F2D8 , 32'h0003EA9F , 32'h04547B88 , 32'h0002B229 , 32'h00049901 , 32'h08952D80 , 32'hE6E044C0 , 32'hFFFFB612 , 32'hFFF8603C , 32'h0000069E , 32'hFFFB214E , 32'h0002CD42 , 32'hEB220F80 , 32'h0B1FAD20 , 32'hFFFDB9B0 , 32'h0002966F , 32'h220CE800 , 32'h04C482C0 , 32'h00000E51 , 32'h00034356 , 32'hF8611B28 , 32'hFFFAC852 , 32'h0000BDD6 , 32'hFFAE3DDC , 32'hF8025180 , 32'h01CE5010 , 32'hFEB374D0 , 32'hFFFFA6CA , 32'hFFFF64F6 , 32'hF5813400 , 32'hFFFF6B65 , 32'h0002153B , 32'h05DECE30 , 32'hFFFCD9A5 , 32'h0002BF1A , 32'h18042520 , 32'h0001CFE4 , 32'h1236E6A0 , 32'hFE7D19D4 , 32'h000297EF , 32'h0002CE8F , 32'h00000E8E , 32'hEF074600 , 32'h14638B60 , 32'hF39150E0 , 32'h044AFDF8 , 32'hFFFD23B1 , 32'hFCD37E98 , 32'hFFFC52E0 , 32'h0003BF2C , 32'h1A362BA0 , 32'hF9956AE0 , 32'h08509A00 , 32'hFFFDCE67 , 32'h18CFE4C0 , 32'h02B02B98 , 32'h0597CDD0 , 32'h0E4A8610 , 32'h10504FC0 , 32'h1070C320 , 32'hFF81CCB6 , 32'h1BD87BA0 , 32'hFFFE05DE , 32'hFFFEAA8C , 32'hFFFF01F2 , 32'h10ACF720 , 32'hE7F83CE0 , 32'h036BA2F0 , 32'hFFA178F3 , 32'h02EDE82C , 32'hFD8898D8 , 32'hFFFF3A90 , 32'hFF178B2B , 32'hFCB2A74C , 32'hFFFBB036 , 32'h14F67E00 , 32'hFFF8F80D , 32'hE5DB17E0 , 32'hF54ECBE0 , 32'h00019F85 , 32'hFFFD0DE1 , 32'h00041588 , 32'hFFFE5FA8 , 32'hFFFA8ABC , 32'hFFFE415B , 32'hEA5DB620 , 32'h24499740 , 32'h06D5E518 , 32'h04217C58 , 32'h28A06500 , 32'hD3A383C0 , 32'h00009ABB , 32'hFFFBFD1A , 32'hFFFC3579 , 32'hFFFF15E9 , 32'hFFFF0353 , 32'hFC0406DC , 32'hF374DD70 , 32'hECE5D940 , 32'h000011BA , 32'h00016304 , 32'h00022C74 , 32'h00000A67 , 32'hEDC46B20 , 32'hE97A6860 , 32'h00002983 , 32'hFFFDF087 , 32'hFFFE4EF0 , 32'hF7D9AE60 , 32'hD2A2D140 , 32'hD41028C0 , 32'h0004FD1B , 32'hFFFBF5C6 , 32'h0002C04D , 32'hF413E950 , 32'hF688C530 , 32'h024822C4 , 32'h0005CB77 , 32'hFE806C90 , 32'h000A2F45 , 32'h0ECB9FC0 , 32'hFFFCE05E , 32'hFBF9CD88 , 32'hFFF6A6C6 , 32'hF50D42A0 , 32'h00D05876 , 32'h0EE66FF0 , 32'hF1917290 , 32'h00009140 , 32'h04883D70 , 32'hF9C293B8 , 32'h0004A43C , 32'hFA396F50 , 32'h00055238 , 32'h064B82B0 , 32'h2CF6C800 , 32'h13D1D0E0 , 32'hFFFCA63F , 32'h00026752 , 32'h222BD800 , 32'hFFF88217 , 32'h0E4E8AE0 , 32'hFFFD042C , 32'hFE0EA6B0 , 32'h0002E057 , 32'h09F54C80 , 32'hFFFD7CAE , 32'hFFFA304A , 32'h00005C82 , 32'h039502FC , 32'hE6916920 , 32'h00014FA5 , 32'hFFFA0DF6 , 32'hFFF92999 , 32'hFFFFAA56 , 32'h07C01650 , 32'hF2E41AE0 , 32'h1798ECE0 , 32'hCC1D24C0 , 32'h07E150E0 , 32'h0000CF83 , 32'h0001ECA0 , 32'h0004AE65 , 32'h06B49018 , 32'h0002041C , 32'h0003E768 , 32'hF58462A0 , 32'hC9933000 , 32'hFFFF18A6 , 32'h1A7E32A0 , 32'hFDA83328 , 32'hE73AEE00 , 32'h21A50580 , 32'hFFFDBC50 , 32'h168E44E0 , 32'h06A78730 , 32'h02B303D0 , 32'hFFFF6344 , 32'h036DA0C0 , 32'hE13D60A0 , 32'hFB6CDAB8} , 
{32'h065261A8 , 32'hF3AA7B70 , 32'h0002B642 , 32'hFA343CA8 , 32'h00012049 , 32'h02ED936C , 32'hFFFBFE1D , 32'h00013859 , 32'hFFFCBC59 , 32'h0002B6C0 , 32'hF63166A0 , 32'h216289C0 , 32'hFA490168 , 32'hFFFCB53A , 32'hFFFF0962 , 32'hEA5B4E40 , 32'h0001F674 , 32'h22CA7F80 , 32'hFBE71198 , 32'h0001EC0B , 32'hFFFD86A8 , 32'h09F53260 , 32'hF592B520 , 32'hFBEEC2A8 , 32'hEC0CC4A0 , 32'h00024E99 , 32'h04572AA0 , 32'hFB542F78 , 32'h00005378 , 32'hF3D71610 , 32'h00005429 , 32'hD4D9EC80 , 32'h00019519 , 32'hFFFFC009 , 32'h000125CE , 32'h196FB4C0 , 32'hEAA1FD40 , 32'h00C47232 , 32'hFFFB285B , 32'h15107960 , 32'h0F80C630 , 32'h0000661E , 32'h000480A6 , 32'h0040A725 , 32'h168AFB60 , 32'hD4F2CF80 , 32'h149DCEC0 , 32'h000429A7 , 32'hEDCF3AA0 , 32'h01B6341C , 32'hFF516DE4 , 32'hFFFF3D95 , 32'h04BD94D0 , 32'hD9264000 , 32'hF5EFBCE0 , 32'h0003D467 , 32'hFC27ECB0 , 32'hFFF816F5 , 32'h0006A1EC , 32'h08F4B5A0 , 32'hFDF7F290 , 32'hEBD7E200 , 32'h3B987600 , 32'hFFFF7C54 , 32'hF44ED230 , 32'h000320A6 , 32'hEEDAF020 , 32'h04DCEDD0 , 32'h0007168E , 32'hBD998800 , 32'hF546F5E0 , 32'hEE3FE7E0 , 32'hFFFEE9CA , 32'h0000C462 , 32'hFFFFDCBE , 32'hFD824280 , 32'h0463ED18 , 32'hFFFFE055 , 32'hE3C70BC0 , 32'h0048D9ED , 32'h000098B7 , 32'hF0BB3710 , 32'h01951C30 , 32'h00012FF4 , 32'h0CBD9040 , 32'h06E07340 , 32'h0D42F0A0 , 32'hFFFF879F , 32'hFFFE3244 , 32'hF69D3860 , 32'hFFFF3365 , 32'h03E9AA14 , 32'h00039335 , 32'h04D26680 , 32'h0010489C , 32'h00002833 , 32'h00003E67 , 32'hFFFD1195 , 32'hFFFCFF0A , 32'hE22ECB40 , 32'hF492C810 , 32'h000073CF , 32'hDEE952C0 , 32'h22657C00 , 32'hFFC7B9F7 , 32'hFFFE8270 , 32'hFE040BC8 , 32'h00009A2B , 32'h06816130 , 32'h0573FDA8 , 32'hFFFE594F , 32'hFD0C090C , 32'hFFFF67F7 , 32'h00011B54 , 32'hFBBD7AF8 , 32'hF74F47D0 , 32'hFD55A2EC , 32'h0000E07C , 32'hF3212C70 , 32'hFFFE9B9C , 32'hFFFE4D96 , 32'h0CCDFD20 , 32'h000414BB , 32'h0005E087 , 32'hBBA45A80 , 32'hED8E9CE0 , 32'hFFFE2359 , 32'hFFFE4F49 , 32'h0002BEF4 , 32'hFFFFC2E9 , 32'hFFFCCDB5 , 32'hFA7B1CB8 , 32'h0B144D10 , 32'h00002B0D , 32'h0001DF5A , 32'h400DA200 , 32'h1440C000 , 32'hFFF9E29A , 32'h000130D6 , 32'h1F32BAC0 , 32'h0001C9FF , 32'h000279C2 , 32'hFBE74FD0 , 32'h00199C00 , 32'h00FCB210 , 32'h00D58020 , 32'h00078E59 , 32'h0002C009 , 32'hF1DF0FF0 , 32'h00011EFE , 32'hFFFF5E0D , 32'h04A292E0 , 32'hFFFBC89A , 32'h00064763 , 32'h002115EC , 32'hFFFD38A7 , 32'hFF317257 , 32'hFF4CE5F0 , 32'h00084772 , 32'h00005597 , 32'h0002F278 , 32'h11AF83E0 , 32'h163AE520 , 32'h01DCD188 , 32'h185BFF00 , 32'hFFFA6DE9 , 32'h16B23060 , 32'h00022A26 , 32'hFFFB1A82 , 32'h00F34689 , 32'hFF51FE08 , 32'h052CFC08 , 32'hFFFB9723 , 32'hF95FABA0 , 32'h01605B44 , 32'hF69C4180 , 32'h116B3780 , 32'hF819FEC0 , 32'hD7C4DD40 , 32'h0151D6B8 , 32'hFFD99279 , 32'hFFFDB46C , 32'hFFFE4812 , 32'h0001BD84 , 32'h043CD9E8 , 32'hE1B42A20 , 32'hF93AC338 , 32'h00A3976B , 32'h12D62D00 , 32'hF3264A60 , 32'h00047F44 , 32'h03CC52D8 , 32'h16F0AE80 , 32'hFFFD7165 , 32'h23867980 , 32'h000146D2 , 32'hF0157480 , 32'h6A8B6A80 , 32'hFFFA79C2 , 32'h00004508 , 32'hFFFC6AF5 , 32'hFFFBE6FF , 32'h00055E91 , 32'h0005491B , 32'h0F321FE0 , 32'hE9C22240 , 32'hE5EACE40 , 32'h0534D630 , 32'h03087AEC , 32'hFB5220D0 , 32'h00007A40 , 32'hFFFFEB79 , 32'h0002FE72 , 32'h00018B36 , 32'h000062E1 , 32'h04CDE350 , 32'h1C79BCA0 , 32'h1DAB3E20 , 32'hFFFBC12E , 32'h000709EF , 32'h00002903 , 32'hFFF9410F , 32'hFD70A570 , 32'h227BB600 , 32'h0001B11F , 32'hFFF71580 , 32'h0003F9F2 , 32'h52EED580 , 32'hEF50D340 , 32'hE69E1FA0 , 32'h0005FB36 , 32'hFFFE7201 , 32'h0000E874 , 32'hFFAE8F1B , 32'h01C25994 , 32'h14ABAD00 , 32'hFFFC6329 , 32'h00B91A17 , 32'hFFF824BD , 32'h03391620 , 32'hFFFD47E3 , 32'hDC075740 , 32'h00012421 , 32'hFF7C82E5 , 32'hF70319F0 , 32'h2920B780 , 32'hD3C5E280 , 32'hFFFAD7A5 , 32'h09C177D0 , 32'hFB7E0400 , 32'hFFFD772F , 32'h094A00A0 , 32'h00018C1D , 32'hFC44FBF0 , 32'hFAA4DD00 , 32'h14A5C300 , 32'h0001B002 , 32'hFFFF05AC , 32'hEDE229E0 , 32'h000697CB , 32'h01C2BB68 , 32'h00024582 , 32'hFD66158C , 32'h0002E94B , 32'h02D1FC10 , 32'hFFFD470F , 32'h00043557 , 32'h0005ED91 , 32'hF40C0A00 , 32'h14907E80 , 32'h0000DB87 , 32'h0002E251 , 32'hFFFFCEA9 , 32'h0005FE2C , 32'h16AFDDC0 , 32'h28455280 , 32'h0DD7F590 , 32'hF49DD130 , 32'hFDC51734 , 32'h00000131 , 32'hFFFF3F25 , 32'h00001DBF , 32'hFCDC5F70 , 32'hFFFA202C , 32'h00028B83 , 32'hFD44622C , 32'hBFADC180 , 32'hFFFE7716 , 32'h085BB680 , 32'h06443518 , 32'hF8026708 , 32'h159487A0 , 32'h0001E004 , 32'h0479B4D0 , 32'hF0E18260 , 32'hFB799078 , 32'h00050B6B , 32'h05CDE518 , 32'h1449C8C0 , 32'h0E466EF0} , 
{32'hFF81C5A2 , 32'h0F14B3A0 , 32'hFFFD1069 , 32'h22227980 , 32'h0000FB40 , 32'h02E9D188 , 32'h000214FF , 32'h00009CB6 , 32'h00000BA2 , 32'hFFFC0AF6 , 32'hF5DDAC90 , 32'h150777E0 , 32'hEE2F7160 , 32'h00022EDB , 32'hFFFF0D53 , 32'h0C9C43E0 , 32'h0001C992 , 32'hE40C2940 , 32'hFE82CC68 , 32'hFFFCBBE8 , 32'h00024168 , 32'hFBDB1D00 , 32'hF2AC14E0 , 32'hFF2FB119 , 32'hE85971C0 , 32'hFFFD4C3D , 32'h02EFD07C , 32'hFF9432FA , 32'hFFFEF9E7 , 32'h12293D40 , 32'h00030C9D , 32'hEBD54540 , 32'hFFFE39A5 , 32'hFFFE7406 , 32'hFFFF73FD , 32'h1A7CA360 , 32'hFAAB4380 , 32'hDDE433C0 , 32'hFFFCF833 , 32'h4681DE80 , 32'hE2EEC480 , 32'hFFFBEEEB , 32'hFFFB3E1C , 32'h09378C90 , 32'hF59AC900 , 32'h065A3838 , 32'hEF2FA6E0 , 32'hFFFF74B7 , 32'h0473D068 , 32'h0AC810B0 , 32'h0222ADA0 , 32'h00030A57 , 32'hF9C2A950 , 32'h337267C0 , 32'h0311E61C , 32'hFFFD4103 , 32'h013AC840 , 32'hFFFF9505 , 32'hFFFD553B , 32'hFA6B4F10 , 32'h02FF771C , 32'h077C2F88 , 32'hF0280720 , 32'hFFFE5007 , 32'hC068E580 , 32'hFFFDB058 , 32'h0253DE24 , 32'hFEDFC014 , 32'hFFFA441C , 32'h2EE13A00 , 32'hEBD26BC0 , 32'hDFB06040 , 32'h00020670 , 32'h0001C332 , 32'hFFFF69CB , 32'hFE40F3BC , 32'h047E6968 , 32'hFFFD0872 , 32'hF7D06AB0 , 32'h00C2BC08 , 32'h0002652E , 32'hC9AD6240 , 32'h1BA3B820 , 32'hFFFE993B , 32'h152FFB20 , 32'h206F0E80 , 32'hEBD7B020 , 32'hFFFB33F2 , 32'hFFFC3384 , 32'h2AB339C0 , 32'h000268D8 , 32'hF981E778 , 32'hFFFD4975 , 32'hF1B63180 , 32'hFF2623CB , 32'h000A04C3 , 32'h00027D88 , 32'hFFFD3524 , 32'hFFFD71FD , 32'hF6778950 , 32'hFC5E0CEC , 32'h0006CEC1 , 32'h09E33230 , 32'hEB493C40 , 32'hFE67FE18 , 32'hFFFC27A5 , 32'hFEF0BCC4 , 32'h0004A77B , 32'hFB0F1E48 , 32'h03038A20 , 32'h0003B18E , 32'hCCC5F0C0 , 32'hFFFDA9DE , 32'h00003533 , 32'hFA8ECBB8 , 32'h027ABD1C , 32'h05A42B90 , 32'hFFFAA407 , 32'h03C4C05C , 32'hFFFE444D , 32'hFFFDE299 , 32'hF26151D0 , 32'hFFFF5BF2 , 32'hFFFC040B , 32'hF31741F0 , 32'h041A26D0 , 32'hFFFF48B2 , 32'h000A1764 , 32'h0002D8EC , 32'hFFFF6F80 , 32'h0001DD2F , 32'hFA3D32E8 , 32'h126A2440 , 32'h00022F49 , 32'h0002BE1D , 32'hE9DFA080 , 32'h085361E0 , 32'h000184A8 , 32'h0001127E , 32'hF9A70448 , 32'h00023BA8 , 32'h000261E2 , 32'hFE15862C , 32'hF407A810 , 32'hFE8D9824 , 32'hFF302D15 , 32'hFFFF7F82 , 32'hFFFB007F , 32'hFEAFD494 , 32'hFFFD6F4F , 32'hFFFE3589 , 32'hEC9AEE80 , 32'h0001BC98 , 32'h00008A41 , 32'hF5FDCFB0 , 32'h0001852B , 32'hF09E67B0 , 32'h02B53450 , 32'hFFF91C5D , 32'hFFFBB45B , 32'h00012539 , 32'hE5B83A20 , 32'h08974560 , 32'hEFF86B80 , 32'hE51C1240 , 32'hFFFFD641 , 32'h12C94380 , 32'h0002147A , 32'hFFFB68E1 , 32'hE88AFA00 , 32'hF503EA40 , 32'hF6FE6800 , 32'hFFFBEDB5 , 32'hFF3C9B61 , 32'hF9ABB0E0 , 32'hFA660D40 , 32'h08C0EF20 , 32'hF51EB2B0 , 32'h0B587EA0 , 32'h00A45A62 , 32'hF50F9D00 , 32'h0002ECF5 , 32'h000170DC , 32'h0002C852 , 32'hF839D050 , 32'h0958D9E0 , 32'h0329688C , 32'h02C08C94 , 32'hFDDEDAD0 , 32'h067D64D8 , 32'hFFF77A0E , 32'h163BEBE0 , 32'h0B2539E0 , 32'hFFFFC387 , 32'hDC6B3340 , 32'hFFFD1713 , 32'hEE7B1320 , 32'h1BE2B080 , 32'h00053ED2 , 32'hFFFFFA22 , 32'h0004E32E , 32'h000300FD , 32'h0001B9E6 , 32'h0002289F , 32'h0875D740 , 32'hFFD8C114 , 32'h241BB480 , 32'hEEF313E0 , 32'hEF0D46E0 , 32'h0064271F , 32'hFFFA573E , 32'h0003DB6E , 32'h0001D900 , 32'h0000B1D7 , 32'h00000532 , 32'h05DA7EE0 , 32'hDB2B3F40 , 32'h31057800 , 32'hFFFE1DD9 , 32'hFFFD5775 , 32'hFFFE4062 , 32'h00005855 , 32'hFA9C9000 , 32'hEAD4E3E0 , 32'hFFFFFA51 , 32'hFFFC396F , 32'hFFFC30AE , 32'h2F88DE40 , 32'hE4CD7880 , 32'hDA8D51C0 , 32'h00028582 , 32'hFFFF7326 , 32'h0003EB5C , 32'hFE714334 , 32'hFDEF8108 , 32'h1C10C460 , 32'hFFFE1B69 , 32'hFCE412E0 , 32'h0003727A , 32'hE8EF1C20 , 32'hFFFFE1F5 , 32'h349D6E00 , 32'hFFFE2440 , 32'h307EFF80 , 32'hDA6A3FC0 , 32'h4C18DC80 , 32'h2A8F0F00 , 32'hFFFEF37A , 32'hDCF05940 , 32'hFDF02D58 , 32'h0002EEC3 , 32'h086DAE70 , 32'h0002F4F9 , 32'hFAE7F180 , 32'hE24D07E0 , 32'hF6020CE0 , 32'h0000361A , 32'hFFFD4D33 , 32'hFE9E02B0 , 32'h0001350A , 32'h18EB5460 , 32'hFFFB5BDD , 32'hFE8C12D8 , 32'hFFF7622F , 32'h38ACC780 , 32'h0002419C , 32'hFFFFD85C , 32'hFFF9292F , 32'hEBBFF080 , 32'hE7AE1DA0 , 32'h0005E404 , 32'h000101EB , 32'h0000A641 , 32'h000211A2 , 32'hFC647144 , 32'hF6304410 , 32'hEACE1160 , 32'h124F5720 , 32'h1C03E680 , 32'hFFFF6681 , 32'hFFFE6018 , 32'h000206A5 , 32'h03C13D08 , 32'hFFFFFD81 , 32'hFFFF7EE1 , 32'hF4B4D180 , 32'h0FDD36A0 , 32'h00024769 , 32'h1844C0E0 , 32'h0687DAA0 , 32'h03D99A44 , 32'hEF1C00A0 , 32'h00003170 , 32'h00A6C540 , 32'h1E5BBC60 , 32'h087ADDD0 , 32'hFFFBC25A , 32'h1771A1A0 , 32'h2B5BCBC0 , 32'h1F4C90C0} , 
{32'h0B352DF0 , 32'h1F6CB380 , 32'h00031D0F , 32'h171FD560 , 32'hFFFD6D08 , 32'hF8970148 , 32'hFFFFA1F0 , 32'h000183BF , 32'hFFFB0B1C , 32'h0002C9A4 , 32'hDF702480 , 32'h14766500 , 32'h0347AB08 , 32'hFFFFF66A , 32'h000277B1 , 32'hFC7B3140 , 32'h00027249 , 32'hD5CC6BC0 , 32'hF72033B0 , 32'h00001648 , 32'h0000CB53 , 32'h070D6718 , 32'hEF37A500 , 32'h0022607B , 32'h164F11A0 , 32'hFFFB096C , 32'hF9CA1B28 , 32'hFE42D588 , 32'hFFFF4CEA , 32'h15F417A0 , 32'h0004A367 , 32'h056AA980 , 32'hFFFF1BE2 , 32'h000373E3 , 32'hFFFD90BB , 32'hDF2331C0 , 32'hFCA50628 , 32'hE2CA5500 , 32'hFFFBCCB8 , 32'hE11479C0 , 32'hD4DC8080 , 32'hFFFF594E , 32'hFFFAEC1A , 32'h010866BC , 32'h06B210D0 , 32'hD33BEA00 , 32'h0B37ABE0 , 32'h00089FB8 , 32'hDC782F40 , 32'h123AFF60 , 32'h00274522 , 32'h00044A61 , 32'hFD58286C , 32'hFBC1E2D8 , 32'hF3EC1FE0 , 32'hFFFDEEE1 , 32'hFF683DFF , 32'h0001910F , 32'hFFFD6FB3 , 32'hFF3E6AD0 , 32'hFE5964DC , 32'h0AFDFD70 , 32'hF9612480 , 32'hFFFE9930 , 32'h461EDD00 , 32'hFFFEBE92 , 32'h090F4480 , 32'h02A14BD4 , 32'hFFFD4F2D , 32'h19367320 , 32'hF3BD3570 , 32'h1088C940 , 32'h000000AD , 32'h0002BC0C , 32'h00019D8B , 32'h8323AB00 , 32'hFAAC1EA8 , 32'h00050A48 , 32'hED6DBF40 , 32'h00E56203 , 32'h0000DB77 , 32'h02EC2030 , 32'hF52B06D0 , 32'h0001413F , 32'hF805C6D0 , 32'h1D937480 , 32'hDD90FC80 , 32'h00021E48 , 32'h0001F636 , 32'h07A32740 , 32'hFFFF9D2D , 32'h0374599C , 32'hFFFE7C9A , 32'h0943FD70 , 32'hFCB16F5C , 32'h000311C3 , 32'h00036F6F , 32'h00041F96 , 32'h0001577C , 32'h043824A8 , 32'h05FBAF10 , 32'h0002F4FB , 32'hF0FFFD80 , 32'h195B3C20 , 32'hF941F0F8 , 32'hFFFF85EC , 32'hFE48354C , 32'hFFFD6B2E , 32'h02C02A4C , 32'hE566B2E0 , 32'hFFFC51E8 , 32'h0E016610 , 32'h00021E66 , 32'h00053F54 , 32'h0FB6AB30 , 32'hF7A514E0 , 32'hFF321028 , 32'h00057DC3 , 32'h1915D9C0 , 32'hFFFE5081 , 32'hFFFBDD25 , 32'h04BC6C60 , 32'h0003030F , 32'h0005DEC6 , 32'h14AA1EA0 , 32'h140F9BA0 , 32'hFFFFB12D , 32'h00018177 , 32'hFFFF6A56 , 32'hFFFB4BDE , 32'hFFFCD60A , 32'h09AB74D0 , 32'h1E425A20 , 32'h0003AF0A , 32'h00034FD2 , 32'h2B336240 , 32'h061B6D58 , 32'hFFFF344B , 32'h00034849 , 32'hF61C2310 , 32'h000171D3 , 32'h0002A65A , 32'hF3A9BE40 , 32'h008D630C , 32'hFC61A5DC , 32'hFED8BC44 , 32'hFFFFCA41 , 32'hFFFEAD64 , 32'h06CEDA88 , 32'hFFFF829D , 32'hFFFF4D1B , 32'h064B0AB8 , 32'hFFFE06BC , 32'hFFFD15C5 , 32'hD97ED540 , 32'h00017A63 , 32'h10A88260 , 32'h0031C684 , 32'hFFFF9612 , 32'h000310DA , 32'hFFFF72DA , 32'h0EEE1F10 , 32'h08AE28F0 , 32'hFE5860EC , 32'h0AF10F60 , 32'hFFFCBB0E , 32'h04AD4338 , 32'hFFFC81E5 , 32'hFFFE4DF0 , 32'h17787040 , 32'hFEA34664 , 32'hF86B3800 , 32'h00049AF3 , 32'hCB578080 , 32'hF7E4B2F0 , 32'hEE9BECC0 , 32'h27B08EC0 , 32'hE00FF700 , 32'h1DF1A7E0 , 32'h03586104 , 32'h08FFADC0 , 32'h00042891 , 32'hFFFCB900 , 32'hFFFAC574 , 32'h00469866 , 32'hF1B704F0 , 32'h026159DC , 32'h0390B9C8 , 32'h15A87AE0 , 32'h024E7ECC , 32'hFFFAD7DB , 32'hE98EF5C0 , 32'hFDA60F78 , 32'h00049848 , 32'hDE38BE00 , 32'hFFFF6421 , 32'h233657C0 , 32'h0D003350 , 32'hFFFEDCDE , 32'hFFFFCD41 , 32'h0001E260 , 32'h00023C01 , 32'h000047F9 , 32'hFFFC723D , 32'hEE5CE780 , 32'hFE54420C , 32'h0088A9A1 , 32'hFA244028 , 32'hE7FD1900 , 32'hFA62E308 , 32'h000210E7 , 32'h00059130 , 32'h00001980 , 32'h0000E873 , 32'hFFFF3F58 , 32'h0A3CD0C0 , 32'h109776E0 , 32'h0CE0B010 , 32'hFFFF7566 , 32'hFFFD9C95 , 32'h00038F5B , 32'hFFFDF9A3 , 32'hF56A6BE0 , 32'hDD634E80 , 32'h000474CC , 32'h00022619 , 32'hFFFA3AD5 , 32'h345F4D00 , 32'h20EEE140 , 32'h08271000 , 32'hFFFD04C8 , 32'h00025A88 , 32'hFFFCA6DC , 32'h0025BD5D , 32'h04C63438 , 32'h06311A90 , 32'h0004845C , 32'h00BA9637 , 32'h0002412A , 32'h044EBE60 , 32'h000607F3 , 32'h135FB400 , 32'hFFF857AB , 32'hEB5D4320 , 32'hE49E9DE0 , 32'hF2842290 , 32'hEB355200 , 32'hFFFE854A , 32'hFC4BC5B8 , 32'hFF011947 , 32'hFFFD93DD , 32'h15697DA0 , 32'h00008DEC , 32'h020A48CC , 32'h0333EEF8 , 32'hC358F280 , 32'h0001DEE6 , 32'hFFFD1370 , 32'h0BFE1B70 , 32'hFFFC6890 , 32'hF76A81A0 , 32'h0001A13B , 32'hFFDFCFAA , 32'hFFFA128B , 32'hF2515600 , 32'h00029756 , 32'h0003D16C , 32'h0003A4CB , 32'hFBE0C780 , 32'h09B15DC0 , 32'hFFFF8EB6 , 32'h00059BD9 , 32'hFFFE3E5A , 32'h0005B746 , 32'hECAFB480 , 32'h176F67E0 , 32'h0DC6DD50 , 32'h1C6F1BC0 , 32'h2F254540 , 32'hFFF9CB86 , 32'hFFFBABA5 , 32'h0003FDA2 , 32'hF4E31370 , 32'hFFFC241F , 32'hFFFFE66F , 32'hFF1053D9 , 32'h05C82410 , 32'hFFFEDF11 , 32'h1CE9BD00 , 32'h064B1150 , 32'h05999348 , 32'hFA5177D0 , 32'hFFFB6CF8 , 32'hEAEBB600 , 32'h252CE6C0 , 32'hFE451FC0 , 32'h00037F31 , 32'hCAFBC2C0 , 32'hE64275A0 , 32'hF18FC2B0} , 
{32'h34366000 , 32'hFD1AAEF0 , 32'h00062B01 , 32'hDF592240 , 32'h0002A4D7 , 32'hFA5DDCD0 , 32'h00030CA1 , 32'h00030912 , 32'hFFFF357A , 32'hFFFEE7BF , 32'h1317C2A0 , 32'h1C76FEA0 , 32'hF1189B90 , 32'hFFFD3280 , 32'hFFFBD645 , 32'hEEE47440 , 32'h0003F02D , 32'h37A62100 , 32'hF9D3F7A0 , 32'hFFFA341F , 32'h0005287E , 32'h04386458 , 32'h0D21AB40 , 32'hF9317248 , 32'h11883660 , 32'hFFFF552C , 32'hFA7FC410 , 32'hFDA96238 , 32'h0002A6AD , 32'h05A86240 , 32'hFFFE6F2D , 32'hED422320 , 32'h00069F54 , 32'hFFFCA178 , 32'h00004538 , 32'h05CDDC90 , 32'h0C9B0820 , 32'hDF677AC0 , 32'hFFFDC691 , 32'hFF860B8F , 32'hF68EE540 , 32'h0001593E , 32'h0001FD3D , 32'h045040F8 , 32'h1B0D4360 , 32'hEC2BFE40 , 32'hE0FAA840 , 32'h00065779 , 32'hE90EB380 , 32'h03B57764 , 32'h00183BC0 , 32'hFFFC743C , 32'hFBA5E4E0 , 32'h0508ADA0 , 32'h0FFF0D30 , 32'hFFFE15F8 , 32'h01D47274 , 32'hFFFCFE20 , 32'h0000A0F3 , 32'hF53DF8C0 , 32'h094AF750 , 32'h062187C0 , 32'hED1A6160 , 32'hFFFE9AEC , 32'h527D3980 , 32'h000491B5 , 32'h12D58380 , 32'hFE6BA930 , 32'hFFFBDBAD , 32'hD9BA3EC0 , 32'hEBC22EE0 , 32'hFF8B0A2B , 32'h00005110 , 32'h0000C654 , 32'h00016CD0 , 32'h4F25CE00 , 32'hFC7624B8 , 32'hFFFEBF82 , 32'hE6355240 , 32'h01013848 , 32'h0001887D , 32'hF278A180 , 32'h12948760 , 32'hFFFFFB42 , 32'h00034590 , 32'h0DACEAA0 , 32'h0DB2DAB0 , 32'h0003214F , 32'h00077CB9 , 32'h1ABB51A0 , 32'h00009796 , 32'hF9F08BF0 , 32'h00010699 , 32'h183F3500 , 32'hFD23FF14 , 32'hFFFD944A , 32'h00052D51 , 32'hFFFE2D66 , 32'h0002233E , 32'hFFDEDCFC , 32'hFD487A38 , 32'hFFFB11F7 , 32'hD3FFC1C0 , 32'h143F0080 , 32'hEEF18E00 , 32'hFFFAA1A7 , 32'h0072A8F0 , 32'h00016F0C , 32'hF281B840 , 32'h27DB1680 , 32'h0001451D , 32'h04049250 , 32'hFFFF9F8C , 32'h00039366 , 32'hF3F0A0E0 , 32'hE6850100 , 32'h042C62A8 , 32'h0003C369 , 32'hE82A2300 , 32'h0002DA07 , 32'hFFF6BA00 , 32'hED47D240 , 32'h00002F85 , 32'h00049154 , 32'h27E6B100 , 32'hD9B66780 , 32'h0002ADA4 , 32'h00016245 , 32'h000127AB , 32'h00016A04 , 32'hFFFC76D5 , 32'h00FFDCE4 , 32'h18D37D40 , 32'h0001B085 , 32'h0001B7BA , 32'hF3B1B410 , 32'h01B80FC0 , 32'hFFFE9569 , 32'hFFFCF800 , 32'h05B8BC98 , 32'hFFFD1FA5 , 32'h0004A653 , 32'hFFAC97E3 , 32'h08235700 , 32'hF9708198 , 32'hFAC2F0E8 , 32'hFFF85DBD , 32'h0000412F , 32'h0D9D3AA0 , 32'hFFFDCBBC , 32'h0000C0D8 , 32'h088C4000 , 32'hFFFF934F , 32'hFFFD8F3D , 32'h0AF0BF00 , 32'hFFFF6134 , 32'hFE8374F4 , 32'h02563838 , 32'h0002AF82 , 32'h000267E3 , 32'hFFFBE9B2 , 32'h0B1B4340 , 32'h02D09EBC , 32'hFCE9D008 , 32'hF9ADE6E0 , 32'hFFFDB019 , 32'hDD1792C0 , 32'hFFFE141C , 32'h00030193 , 32'h0018E8AA , 32'hFF338F19 , 32'hF71D0C90 , 32'h000563ED , 32'hB4F7C700 , 32'hFAED93A0 , 32'hEF4FEF60 , 32'hFE38B314 , 32'h14A76F60 , 32'h45789400 , 32'h0672CE78 , 32'hE1231EC0 , 32'hFFFF0FF1 , 32'hFFFFA3EB , 32'h0004A459 , 32'h086702F0 , 32'hF37D1E70 , 32'h01C4E28C , 32'h05ECDAF8 , 32'hEACD0280 , 32'hF43C97D0 , 32'hFFF9CE1E , 32'hDD1A7180 , 32'h0FA4CF60 , 32'h0002229C , 32'hFE7CC5C4 , 32'hFFFFE234 , 32'hE80C0DE0 , 32'h0BD47BC0 , 32'hFFF970F7 , 32'hFFFE4B27 , 32'hFFFE8A60 , 32'hFFFE4FB0 , 32'hFFFFBB1E , 32'hFFFFB150 , 32'h0EE093C0 , 32'h03B5BCA4 , 32'h046ADA30 , 32'hE9F32A00 , 32'hE7182D80 , 32'hE0D2CE00 , 32'hFFFE45D1 , 32'h000228F6 , 32'hFFFF692B , 32'hFFFD2CC4 , 32'h0003F450 , 32'hF37EC1D0 , 32'h10C16C40 , 32'hE28BF8C0 , 32'h00009BAD , 32'hFFFDE0F0 , 32'hFFFFEAC0 , 32'hFFFE5E53 , 32'h07100AB0 , 32'hCEB05A40 , 32'h00019FFA , 32'hFFFE729D , 32'h00013D68 , 32'hF856EE70 , 32'hF440D810 , 32'h1595D100 , 32'h00005117 , 32'h0002935A , 32'hFFFF9C38 , 32'h00902470 , 32'h0869B3F0 , 32'h0311F2E4 , 32'hFFFF95B6 , 32'h007E2EEA , 32'hFFFE71E0 , 32'hEC1C32A0 , 32'hFFFB5942 , 32'hFD54ADCC , 32'hFFFCC25F , 32'hF4F65210 , 32'hE377E9E0 , 32'hF8BE9BF0 , 32'h0D1F22B0 , 32'hFFFEB1B4 , 32'h01811764 , 32'h0255B3F0 , 32'hFFFDD7EA , 32'h014FBB58 , 32'h00050152 , 32'hF5A143F0 , 32'hC938B300 , 32'h0FE38D60 , 32'hFFFFC3F1 , 32'hFFFDACB2 , 32'h2D6091C0 , 32'hFFFD203C , 32'h17606C20 , 32'h00014845 , 32'h0188AB34 , 32'hFFFE35F9 , 32'hFF9C0DF1 , 32'hFFFD4064 , 32'h00002BBB , 32'hFFFDFD8E , 32'h05B94028 , 32'hD2769380 , 32'hFFFB1E15 , 32'hFFFE9F81 , 32'h00026E2F , 32'hFFFAC276 , 32'h048889B0 , 32'hDD4C75C0 , 32'h0DC6A6B0 , 32'hCE71DD80 , 32'h20B71980 , 32'hFFFA6177 , 32'hFFFE52EB , 32'h00027DD2 , 32'hFFB9698B , 32'h0000AA5D , 32'h00054764 , 32'h00A91FB4 , 32'hFA341F88 , 32'h000453AC , 32'h18289760 , 32'hF9CE7708 , 32'hF5AED130 , 32'hF13573B0 , 32'h0003A718 , 32'hF9D787B8 , 32'hFBD33378 , 32'h002C1430 , 32'h00055E4A , 32'h21516F80 , 32'h17E47D00 , 32'hF0A52550} , 
{32'hDBE32B00 , 32'hE656D0C0 , 32'h0005A185 , 32'h0267FF94 , 32'hFFFDBEA5 , 32'hF99F6C58 , 32'hFFFBEB85 , 32'hFFFC841C , 32'hFFFED496 , 32'hFFFFDF47 , 32'h1E2142A0 , 32'h3E918200 , 32'hF7B67D40 , 32'h000096E6 , 32'h00002A70 , 32'hEAB75C80 , 32'hFFFDB140 , 32'hFCEB8DA0 , 32'h14A83460 , 32'hFFFCE7AE , 32'h0002EB1A , 32'h01AB4860 , 32'h143BD9A0 , 32'h00A7E24C , 32'hE0571CE0 , 32'h00024305 , 32'h013EF8DC , 32'h02FA5754 , 32'h00000E7F , 32'h2EEFDF40 , 32'hFFFF2D84 , 32'hFB687BD0 , 32'hFFFE2912 , 32'hFFFE76A1 , 32'h0002ECD9 , 32'h11EDAEC0 , 32'h089BB9D0 , 32'hE412F540 , 32'h00064A14 , 32'h0E9D9C80 , 32'h27D2C040 , 32'hFFFFAAAC , 32'hFFFF96BA , 32'hFDF9D9AC , 32'h1D65E1A0 , 32'hF71CA780 , 32'h16791F60 , 32'h00002929 , 32'h0C310B60 , 32'h05E27588 , 32'hFE6C64DC , 32'hFFFFAB2E , 32'hFAAC0A78 , 32'h0E707F60 , 32'hE0E06FA0 , 32'hFFFB1866 , 32'hFE97C7E4 , 32'h00013406 , 32'hFFFF7EF9 , 32'hF4760490 , 32'h0112B94C , 32'h0840D650 , 32'h0704F0C8 , 32'h000256C8 , 32'h04978D70 , 32'h00047DE7 , 32'hE86C9FC0 , 32'hFCB53D90 , 32'h00009723 , 32'h01C78E54 , 32'h0BBA4E50 , 32'hFD8CEC50 , 32'h00007BB6 , 32'hFFFABEE7 , 32'hFFFF7CEA , 32'h1F4CDC40 , 32'h034404A4 , 32'hFFFC7D7D , 32'hC56E1BC0 , 32'h0293F600 , 32'h0001066A , 32'h0675BC08 , 32'hFDED8850 , 32'h00005841 , 32'hEEC91380 , 32'h027C7CB0 , 32'h07CDC670 , 32'hFFFF880F , 32'hFFFEC4C2 , 32'hBCEB1000 , 32'hFFFF4CE3 , 32'h047E88F0 , 32'h000143F2 , 32'hEE715620 , 32'h0021C920 , 32'hFFFFF003 , 32'h0003CF93 , 32'h00020842 , 32'hFFFC939E , 32'h0ED84D10 , 32'h0120BD94 , 32'h0002FC57 , 32'h0B1D8220 , 32'hE0B86A00 , 32'h088783D0 , 32'hFFFF5531 , 32'h00953F93 , 32'h00013EAE , 32'hF670FC00 , 32'hF2619700 , 32'h0001909D , 32'h14D37840 , 32'hFFFF2555 , 32'hFFFB7C98 , 32'h024F9D20 , 32'h00513A95 , 32'hFEAB5628 , 32'hFFFE8A70 , 32'hFE41EF30 , 32'hFFFB6506 , 32'hFFFF3155 , 32'h0233D4A4 , 32'hFFFE6EFA , 32'hFFFFA5EE , 32'h0E4848F0 , 32'hE021B580 , 32'hFFFAB52D , 32'hFFFC4239 , 32'hFFFEF4ED , 32'h00017C91 , 32'hFFFF2986 , 32'hF82135B8 , 32'h0CD16870 , 32'hFFFF49BB , 32'hFFFF423C , 32'h31F02380 , 32'h11BB8420 , 32'h000096E0 , 32'h0000DACD , 32'hF34188B0 , 32'h00014548 , 32'h0000B211 , 32'h03B2E168 , 32'hE9C496A0 , 32'h035F3A38 , 32'h033134CC , 32'hFFFD4C97 , 32'hFFFB6860 , 32'hF0992E30 , 32'hFFFF8D29 , 32'hFFFCA38F , 32'h02C00D88 , 32'h0001F05D , 32'hFFFE1A51 , 32'hFBD97CD8 , 32'h0008EE0D , 32'hFB191538 , 32'hFE1EBFE8 , 32'hFFFE52FE , 32'h0001BDD9 , 32'hFFFE832F , 32'hF19416B0 , 32'h023B76C0 , 32'hFA36D8E0 , 32'hF28D53F0 , 32'hFFFE7BFD , 32'h23324780 , 32'h000327E2 , 32'hFFFFD92B , 32'h3583FB80 , 32'hF18C5AD0 , 32'h0C5BE150 , 32'hFFFCC2AF , 32'h0C29AEE0 , 32'h0AFAFFD0 , 32'h120BEA20 , 32'hEAD68E60 , 32'hE61FA460 , 32'h08F95FF0 , 32'h00081C6B , 32'hF6F88B90 , 32'h0000D8EF , 32'h00030C3A , 32'hFFFE3ABB , 32'hF486CF20 , 32'h0D2F5920 , 32'hFB85AA08 , 32'hFFDC3EFF , 32'hEAAFC280 , 32'h0A51CE60 , 32'h00018E49 , 32'h19505700 , 32'hF169FDF0 , 32'hFFFC74D0 , 32'hCB02BDC0 , 32'hFFFCC41D , 32'hEBE6A6C0 , 32'hF0C1C370 , 32'h0002F15C , 32'hFFFD2B39 , 32'h0005960C , 32'hFFFF07BD , 32'h000023F4 , 32'hFFFDEBBA , 32'hF0F762D0 , 32'h1B80D280 , 32'h2A5A64C0 , 32'h15652640 , 32'h0B86BA20 , 32'h181F87E0 , 32'hFFFAD4E6 , 32'h00019C52 , 32'h0000E11F , 32'h0004F76E , 32'hFFFF435C , 32'h04094830 , 32'h049B0EC0 , 32'h10ED7D40 , 32'hFFFC4C92 , 32'h0003A172 , 32'h00009AA9 , 32'hFFFDCF98 , 32'h0B60D450 , 32'h0E9C0340 , 32'h0000D229 , 32'hFFFF9567 , 32'hFFFFBF51 , 32'h00142A1C , 32'h61799480 , 32'hDE19AAC0 , 32'hFFFE2ABE , 32'hFFFF456C , 32'hFFFCFBF7 , 32'h05EE0438 , 32'h052F29C8 , 32'hDC1C20C0 , 32'h00007655 , 32'hFC9F388C , 32'h00049FFA , 32'hFE996B90 , 32'h0001098C , 32'hEB7C8200 , 32'hFFFDB58B , 32'h20BFFCC0 , 32'h128BCB40 , 32'hD9F4B9C0 , 32'hF6DBA5A0 , 32'hFFFB1657 , 32'h0B26BE00 , 32'h0042DA10 , 32'h000159C6 , 32'h1234AE60 , 32'h00017AB5 , 32'h020A86DC , 32'hFB024480 , 32'hF4417210 , 32'h0000EF3D , 32'hFFFCFC62 , 32'hFFF19F86 , 32'hFFFCC4B1 , 32'hF5FB4440 , 32'h0000ED8C , 32'hFA229970 , 32'h0002C0AD , 32'h18AEC640 , 32'h00032B5C , 32'hFFFC050C , 32'hFFFE9ADF , 32'hE2226700 , 32'hF1AA4580 , 32'h00023B73 , 32'h000060E1 , 32'h00041B45 , 32'h00000C3B , 32'hF10D4AC0 , 32'hEBF40440 , 32'h03194170 , 32'hC267DEC0 , 32'h0C672BD0 , 32'hFFFD9CD9 , 32'h0001FBB8 , 32'hFFFF87B4 , 32'hFE9E91A4 , 32'hFFFF5C2E , 32'h0001B7F6 , 32'h01499A60 , 32'h0D1C8570 , 32'hFFFEBABD , 32'h56369A80 , 32'hFCC4E6CC , 32'hE4C57EE0 , 32'hF1302E50 , 32'h0002906A , 32'hF671CC00 , 32'hE60E1FC0 , 32'h0296BF0C , 32'hFFFF490D , 32'hE5E8D3E0 , 32'h01DBECEC , 32'h0966EDF0} , 
{32'hE8EC4D60 , 32'h23E73F00 , 32'h00000148 , 32'hF07E4CB0 , 32'hFFFEE0D2 , 32'hFA306410 , 32'h0001CC48 , 32'hFFFF0DA1 , 32'h00049836 , 32'hFFF6AE00 , 32'hFA649128 , 32'hF8A212A8 , 32'hD9B95280 , 32'h0003CB54 , 32'h0000DDE1 , 32'h34B1BB40 , 32'hFFFD1F8C , 32'hEA5B4DE0 , 32'hFF8E0632 , 32'h0004A8A2 , 32'hFFFE82CC , 32'hFBEC81E8 , 32'h0EEBE1A0 , 32'h1000B8A0 , 32'h0143E89C , 32'h0006A57C , 32'hFFFB51AC , 32'h05AC41C0 , 32'hFFFEBEC4 , 32'h122B2BA0 , 32'h00033FD4 , 32'h00009264 , 32'h0006E026 , 32'hFFFEA872 , 32'h000174CD , 32'h1BEF56A0 , 32'h0F9C80E0 , 32'h334EA880 , 32'hFFFEFA1C , 32'hDA131540 , 32'hB11D9980 , 32'h0001013B , 32'h0002D646 , 32'h052D1580 , 32'h248DD740 , 32'hF394F600 , 32'h0EE2BD20 , 32'hFFFE783A , 32'h07DA0968 , 32'h01F60450 , 32'h025B6000 , 32'h0003A0E6 , 32'h01496EF0 , 32'hFB260AB8 , 32'h0B1A1C40 , 32'hFFF9F645 , 32'h02A9E504 , 32'h000005F1 , 32'hFFFB646B , 32'hFD922FC8 , 32'h00A73799 , 32'h01E2B86C , 32'hE44D5540 , 32'hFFFFE6F3 , 32'hDF5B4E00 , 32'h0005A7A8 , 32'hE514E440 , 32'h107A2C00 , 32'hFFFE590B , 32'hDE326940 , 32'hF1F88C60 , 32'hF3C7B4F0 , 32'h00034B11 , 32'h0006895D , 32'hFFFC9949 , 32'h16E05160 , 32'h009E8E9B , 32'hFFFEDD6F , 32'h1E574300 , 32'h0290A408 , 32'hFFFD4245 , 32'hE38CA900 , 32'h15E8A240 , 32'h00054F43 , 32'h0278F9BC , 32'hDD291900 , 32'h02A3653C , 32'hFFFE7A22 , 32'h0004B96D , 32'hE8D20DE0 , 32'h00029546 , 32'h06AB4AA0 , 32'hFFFEB802 , 32'h0D6F83E0 , 32'h004C84E8 , 32'hFFF936D8 , 32'h000006A6 , 32'h00008CA1 , 32'hFFFC72B0 , 32'hEEDF68E0 , 32'hF9654D90 , 32'h0002E824 , 32'hF5EC1C10 , 32'h00DDCA56 , 32'hF90B6C88 , 32'h00002C73 , 32'hFFB5D06F , 32'hFFF71695 , 32'h0EC28EA0 , 32'hD60BEC00 , 32'hFFFBBE26 , 32'hE5BE8A00 , 32'h000096B1 , 32'h00016989 , 32'hED189920 , 32'h070C3300 , 32'h04842EA0 , 32'h00036E98 , 32'h074E4D70 , 32'hFFFE8B69 , 32'h00013921 , 32'hF7DEE9C0 , 32'h00015F28 , 32'hFFFF402F , 32'hE59145A0 , 32'hF1208E70 , 32'hFFFE4DD5 , 32'h0006C688 , 32'h000120FB , 32'hFFFD7029 , 32'hFFFD652B , 32'h07916038 , 32'h0FCD8110 , 32'hFFFB7D2A , 32'hFFFD6FB7 , 32'h24689740 , 32'hECD466C0 , 32'h0001DCCA , 32'hFFFF55B4 , 32'hDC891D00 , 32'hFFFFC3A4 , 32'hFFFBB77B , 32'hFDAE24C0 , 32'hEFB60660 , 32'hFAC29D78 , 32'h04746A80 , 32'h00021063 , 32'h00003F90 , 32'hF7DC4A70 , 32'hFFFEF819 , 32'hFFFFCB8A , 32'hF4FC8B70 , 32'hFFFC3EC3 , 32'hFFFB16C1 , 32'h1C70FBE0 , 32'h0003661F , 32'hF6F5DF60 , 32'hF695E0D0 , 32'h0003C572 , 32'hFFFB15D1 , 32'hFFFDA5C8 , 32'hF14344A0 , 32'h0BE64BC0 , 32'h01C47154 , 32'hF192AF90 , 32'h00012C44 , 32'hF1D9DCE0 , 32'h000066C9 , 32'hFFFFAE7E , 32'hF165EE00 , 32'hF9D220F8 , 32'hF7270DC0 , 32'hFFFF58DD , 32'hD4281700 , 32'h018B1EE4 , 32'hFAEBF4D8 , 32'h0CE234C0 , 32'h0E268800 , 32'h0C104A80 , 32'h06D36A38 , 32'hD98BF980 , 32'hFFFE51C1 , 32'hFFFB5E9C , 32'hFFFFF896 , 32'hE6DCF8E0 , 32'h00AD4ABC , 32'hF286FA00 , 32'hF8732D40 , 32'hDA5EB240 , 32'h06049F58 , 32'h00065F20 , 32'h1E89AA20 , 32'h1FD76DA0 , 32'h00020F62 , 32'h16A888A0 , 32'hFFFFFC79 , 32'h0F6FFCB0 , 32'hE5EB47A0 , 32'h000037A9 , 32'hFFFDC0A2 , 32'h00035433 , 32'hFFF9CFEF , 32'h00034F3E , 32'h000036BC , 32'hF42A1D80 , 32'hF7DB7150 , 32'h9849C980 , 32'h047922C0 , 32'hF68BDC00 , 32'hF2500B40 , 32'hFFFD5A26 , 32'h0001132C , 32'h0001ACF0 , 32'hFFFFD145 , 32'hFFFE06D0 , 32'hF3DEFA00 , 32'hEFAED780 , 32'hF984BDE0 , 32'h0000B1D1 , 32'h000063C2 , 32'hFFFD135A , 32'hFFFB1E2C , 32'hEF4C1D80 , 32'h0B632560 , 32'h0000192E , 32'h00046046 , 32'h0001AC3C , 32'hF8D5B090 , 32'h095E0D30 , 32'h09B19C80 , 32'hFFFACE83 , 32'hFFFA2135 , 32'h0003333F , 32'h02ABF4D4 , 32'hFD0C7B80 , 32'h03C92C40 , 32'hFFFF05E8 , 32'hFFFE07EC , 32'h00053ADF , 32'hE6385560 , 32'hFFF97885 , 32'hF1E6D430 , 32'hFFFD6F44 , 32'h0A3794E0 , 32'h01C3DA28 , 32'h1A4502A0 , 32'h06952DF0 , 32'h000180B1 , 32'h062D6BF8 , 32'hFCCCBA8C , 32'hFFF93919 , 32'h011022AC , 32'h000068AA , 32'hFD0D84FC , 32'hFA8D1880 , 32'hA7BE1C80 , 32'h0000DAF0 , 32'h000104D7 , 32'hDFD034C0 , 32'h000216C6 , 32'hDB2D36C0 , 32'hFFFD0BB5 , 32'h02FB0D64 , 32'h00000EDD , 32'hF972B218 , 32'hFFFB175D , 32'hFFFDE1FF , 32'hFFFD9EBC , 32'hE8B99BE0 , 32'hE2374A60 , 32'hFFFFE46E , 32'h00064025 , 32'hFFFC3C41 , 32'hFFFD4A20 , 32'hE9993060 , 32'hD976D440 , 32'hF1A0A540 , 32'hF9987580 , 32'hFEC9BEA4 , 32'h0001A162 , 32'h0000D59A , 32'h00003A85 , 32'hFAFE7A48 , 32'h0002D88C , 32'h000AA8A0 , 32'h01BD6898 , 32'hF4B725D0 , 32'hFFF935A9 , 32'h281718C0 , 32'h00ECFA41 , 32'h033C4F08 , 32'h1D2FDD00 , 32'hFFFCCF49 , 32'hF6B43200 , 32'hD249E900 , 32'h081E38E0 , 32'hFFFE02DF , 32'hFDA1B8F0 , 32'hDF00A280 , 32'hF5D56CE0} , 
{32'hF8F5E4F8 , 32'hE8376400 , 32'hFFFFD209 , 32'hF43AB190 , 32'h00017820 , 32'h02E3AAB0 , 32'h0000B40B , 32'h00012CCB , 32'h00012A34 , 32'hFFFA029B , 32'h04254138 , 32'hF0918300 , 32'h057BF888 , 32'h00067198 , 32'hFFFF2739 , 32'hDA1DC580 , 32'h00004AAE , 32'hA436F780 , 32'hF20BBC10 , 32'hFFFB80A9 , 32'hFFFC6404 , 32'hF3373070 , 32'h21DE31C0 , 32'hFEFFA7FC , 32'hE63FD0E0 , 32'hFFFCED99 , 32'hFFF4051C , 32'hFEC4C8F0 , 32'h0001F13D , 32'h20BE5F00 , 32'hFFFD96C6 , 32'hF844D390 , 32'hFFFE0716 , 32'h00022C2C , 32'h000535C8 , 32'h2EF64740 , 32'hEEA5EFE0 , 32'hD20D0F00 , 32'h00014ABA , 32'h03A6ED30 , 32'h18730C40 , 32'h0002D51D , 32'h0004681C , 32'h064AFBD8 , 32'hD72694C0 , 32'h225C3940 , 32'hFC38D2F4 , 32'hFFFCEFB6 , 32'h1CEF8BC0 , 32'hDDCBF340 , 32'hFF94DD33 , 32'h0006DA5C , 32'hFF401A07 , 32'hE15AD060 , 32'hEB7A1CE0 , 32'hFFFCE684 , 32'hF9EAA460 , 32'h00002F03 , 32'hFFFCD3D2 , 32'h04412828 , 32'h00280E5E , 32'h00DF42DF , 32'h06544298 , 32'h0003CADB , 32'h2041C440 , 32'h00017803 , 32'hE803AD20 , 32'hFA04DA60 , 32'hFFF99E6B , 32'hE3075120 , 32'hD4FB71C0 , 32'h13285BA0 , 32'hFFFAF066 , 32'hFFFED7E2 , 32'hFFFE3DC3 , 32'h09DB52B0 , 32'h04BD5C00 , 32'h00033647 , 32'hD1E5F000 , 32'h07C86498 , 32'hFFFE217D , 32'hE5F92080 , 32'hFEF08E34 , 32'h0004BDE7 , 32'h03869CCC , 32'hC508D080 , 32'hF63DAF00 , 32'hFFFC4779 , 32'h00050824 , 32'h20B44F80 , 32'hFFFA3729 , 32'h0533AFA0 , 32'hFFFE0CC1 , 32'hECE83060 , 32'h01AEF4E4 , 32'hFFFCF5CF , 32'hFFFADBD3 , 32'hFFFBF5E0 , 32'h0000CE4C , 32'h0D5C3AA0 , 32'h0C0FA140 , 32'hFFFDE992 , 32'hF5CC1400 , 32'hEFB9C520 , 32'h11106680 , 32'hFFFD446A , 32'hFFAD254D , 32'h0001AFFC , 32'hFB1208B0 , 32'hE6D8B640 , 32'hFFFCE82A , 32'hE5F532E0 , 32'hFFFC1C6C , 32'h0003822A , 32'h1F877B60 , 32'hFCA74D38 , 32'h0639D5D0 , 32'hFFFA8E2F , 32'hF3CB6C20 , 32'h0001038F , 32'h00012B02 , 32'h16C029A0 , 32'hFFFFB379 , 32'hFFF7EF12 , 32'h0C86DC20 , 32'h26BCFDC0 , 32'hFFFCD205 , 32'h00005AA1 , 32'h000347A6 , 32'hFFFFD960 , 32'hFFFEC140 , 32'hF8BC2A60 , 32'h0EF2EF60 , 32'hFFFF764D , 32'h00085C48 , 32'h0843BFF0 , 32'h132F2180 , 32'h00004D07 , 32'h000636C9 , 32'hE3558320 , 32'hFFFE72F6 , 32'hFFFC7EB5 , 32'h075402D0 , 32'h011752F0 , 32'h04EF8B98 , 32'h03A88F9C , 32'h00032C6D , 32'h0000AA4B , 32'hFFCBDB99 , 32'h0003F0C5 , 32'hFFFD54C2 , 32'h0655BC70 , 32'hFFFD6EE6 , 32'h00011080 , 32'h0EDCD150 , 32'hFFFE1D78 , 32'hE7E38B80 , 32'h0152564C , 32'hFFFF2298 , 32'h00012E70 , 32'hFFFF7FB7 , 32'h1DED13E0 , 32'hE4F92B80 , 32'h08308150 , 32'h2EDDE000 , 32'hFFFD305D , 32'hF45B5470 , 32'hFFFE792F , 32'hFFFE883A , 32'hE05D2D20 , 32'h1422F920 , 32'hFA4479F8 , 32'hFFFE4E37 , 32'hEFF38520 , 32'hF4CCC9E0 , 32'hFFF5A27A , 32'hF766CB90 , 32'hE8FF9200 , 32'hEF3AFBA0 , 32'hFF9AF2E5 , 32'h053038E0 , 32'h0004ACA5 , 32'hFFFBF19D , 32'h0000393D , 32'hF1516B70 , 32'hE284CD20 , 32'hFE58A48C , 32'hFE1C91E4 , 32'h0737DE00 , 32'hEF804020 , 32'hFFFF3A33 , 32'h214685C0 , 32'h12759E80 , 32'hFFFB367B , 32'hE0B42920 , 32'hFFFD830E , 32'h1B2406C0 , 32'hF8C9D4A8 , 32'h000261E5 , 32'hFFFC4D33 , 32'hFFFFE344 , 32'h00005776 , 32'hFFF96CB2 , 32'hFFFCEEF8 , 32'h01186204 , 32'hF8BFE7D8 , 32'hEC254A20 , 32'hEDABCE40 , 32'hF857A168 , 32'hE3499660 , 32'h00008334 , 32'h0003A0BD , 32'h0003A702 , 32'hFFFE2E28 , 32'h0002166C , 32'hF20B7C70 , 32'h08895920 , 32'hE43C1000 , 32'hFFF63C1A , 32'hFFFEA96B , 32'h000183CC , 32'h00010BAB , 32'hF54E42F0 , 32'hF6A68F40 , 32'hFFFE6EB9 , 32'hFFFE2932 , 32'hFFFB2BA6 , 32'hE37A9780 , 32'h004CD12F , 32'hE154BCC0 , 32'hFFFBFAC1 , 32'h000311D3 , 32'hFFFE1180 , 32'h03FFE0B4 , 32'hF92CBAA0 , 32'h01E65D64 , 32'h0002AA2D , 32'hFE37BE54 , 32'hFFFCA40A , 32'h203D7740 , 32'hFFFFB6F3 , 32'h1A936380 , 32'hFFFE0937 , 32'h0A8E45B0 , 32'hE6F2E460 , 32'h06821CA0 , 32'hF9080BA0 , 32'h0004F3E7 , 32'h04408CB0 , 32'hFBE0B870 , 32'h00013C85 , 32'hE8E3E820 , 32'h0000FE2C , 32'hFB989EB0 , 32'h07639A30 , 32'hD83864C0 , 32'hFFFECEF5 , 32'h000179E8 , 32'h0F8B0BF0 , 32'hFFFE2AC5 , 32'hEC3AFE20 , 32'h00082554 , 32'hFCD04968 , 32'h0004539A , 32'hEDDA9320 , 32'h0000C009 , 32'hFFFFFAC5 , 32'hFFFDAD11 , 32'h346747C0 , 32'h3B725500 , 32'h00066232 , 32'h0003DDB6 , 32'h0000C425 , 32'h00058D54 , 32'h22A7E0C0 , 32'hF8629A50 , 32'h12A01F80 , 32'hEC8CF400 , 32'h13A74680 , 32'hFFFE632C , 32'h0001EBAD , 32'h00044475 , 32'hEFD11E60 , 32'hFFFBF8D1 , 32'hFFFD57BC , 32'hF1577D00 , 32'hEF6FBE80 , 32'hFFFBB2F2 , 32'h03B31FE8 , 32'h093AA110 , 32'h048F2300 , 32'hE5F84D40 , 32'hFFFAB86F , 32'h0DA9CC10 , 32'hEF192040 , 32'h0158D9C8 , 32'hFFFAD33B , 32'h47037580 , 32'h03BCEE40 , 32'h0785CCC0} , 
{32'hE867FE80 , 32'hF0853650 , 32'hFFF8F790 , 32'h024420D0 , 32'hFFFD2D19 , 32'hFBC2C548 , 32'h0000A5D9 , 32'hFFFB3A89 , 32'h00003A54 , 32'hFFFFEEDF , 32'hF9453F00 , 32'hDD039C80 , 32'h0F1AE5B0 , 32'hFFFE0C64 , 32'h00084488 , 32'h22011B80 , 32'hFFFFC23B , 32'h3A45CDC0 , 32'hEFC58E60 , 32'h0000B24D , 32'hFFF7923B , 32'hFE8AD0F0 , 32'hFA8FD948 , 32'h10DB93E0 , 32'hFA26D028 , 32'hFFFF3DD4 , 32'hFF639BDB , 32'hFF8BE9E1 , 32'h0003A2CE , 32'h20251740 , 32'h00003304 , 32'hEC609E60 , 32'h00018A97 , 32'h00052B6D , 32'hFFF6CD8F , 32'h025A2188 , 32'h0ACC5FE0 , 32'h0A318E30 , 32'h0001B099 , 32'h0A7EA3F0 , 32'hF162E2D0 , 32'h0003B239 , 32'hFFFFFB06 , 32'hFE540D1C , 32'h2740AA00 , 32'hC98B9340 , 32'hFA87FBA8 , 32'hFFFDF23A , 32'hF9321F68 , 32'h19C70880 , 32'hFFD068B5 , 32'hFFFFD490 , 32'hF36F5610 , 32'hEE57F2A0 , 32'hEE58BEE0 , 32'h0000FBCB , 32'h01D02FC4 , 32'h00027F9E , 32'hFFFE96B2 , 32'hF675CC30 , 32'hFB6809C8 , 32'h0B999C30 , 32'h07BEDE18 , 32'h0003C348 , 32'h077FDBB0 , 32'hFFF732FA , 32'hE4536540 , 32'hFEFEA5A4 , 32'h000B3734 , 32'h4C5C5600 , 32'hF5014B30 , 32'h0ED7B610 , 32'h000226D3 , 32'hFFFD7A9B , 32'hFFFC48E9 , 32'h155B7580 , 32'h08A10B80 , 32'h00021D3A , 32'hF1FB7370 , 32'hFD6F64B4 , 32'hFFFFFE0C , 32'h11C79160 , 32'h08D2B650 , 32'h0000650E , 32'hF3F8D9A0 , 32'h243CCE40 , 32'hFF5A0335 , 32'h0003EB49 , 32'hFFF7F43E , 32'h0884B410 , 32'hFFFDD4D3 , 32'h242BA480 , 32'hFFFB7968 , 32'hF0C11590 , 32'h00560FEA , 32'h00024A07 , 32'hFFFBA6E3 , 32'h00018A90 , 32'h0001BBE1 , 32'h13B24360 , 32'hFB257B70 , 32'hFFFF4441 , 32'h28F13F80 , 32'h004CFB20 , 32'h002F89AA , 32'h00027172 , 32'h0019B7D8 , 32'h000293CB , 32'h0A158260 , 32'h088BF1C0 , 32'hFFFF31FB , 32'hFF215DB0 , 32'h00016F4F , 32'hFFFF0481 , 32'hFC923B40 , 32'hFF494F3F , 32'hFC8713EC , 32'h0001CD24 , 32'h0B5B56B0 , 32'h00009B16 , 32'hFFFD1C84 , 32'h0E780D40 , 32'h00027604 , 32'h0004BEBA , 32'h0AACBCF0 , 32'hF9C99730 , 32'h0001255C , 32'hFFFC7088 , 32'h000304C7 , 32'h00036185 , 32'hFFFF9BF7 , 32'hFD181E94 , 32'h1A9355A0 , 32'h000047BB , 32'hFFFEB60A , 32'h151FF2C0 , 32'h04A5F388 , 32'hFFFD951D , 32'hFFFA62C2 , 32'h1C123580 , 32'h0006E3DF , 32'h00018151 , 32'h04508B70 , 32'h0462FEA8 , 32'h0598F8F0 , 32'h0CB342F0 , 32'hFFFFF9F8 , 32'h0007D51B , 32'hFBE131A0 , 32'hFFFF7F83 , 32'hFFFEB065 , 32'hF52169F0 , 32'h0008B940 , 32'h0004022E , 32'h105DC9A0 , 32'h00028CDC , 32'h080B7780 , 32'h00FC6AD2 , 32'h0006A722 , 32'h0004F5A7 , 32'hFFFDDF4E , 32'h1391D3C0 , 32'hF9E29980 , 32'hFD9C4C28 , 32'hE7FA91A0 , 32'hFFFA8221 , 32'h15D4B6A0 , 32'hFFFF06CE , 32'hFFFDC8B5 , 32'hF9C88D30 , 32'h0A2569A0 , 32'hFDF8C744 , 32'hFFFF1561 , 32'hDAA5CF40 , 32'hF7219830 , 32'h05CFF838 , 32'h140DC820 , 32'hCBBD9D00 , 32'h0E38E590 , 32'hFCD01600 , 32'h281B4740 , 32'hFFFEA6FA , 32'hFFFD9FF4 , 32'hFFFBDA46 , 32'h05D297D0 , 32'hFB40B4B0 , 32'hFB80B610 , 32'h0B5A3B30 , 32'h0BB05280 , 32'hF6856CB0 , 32'hFFFB86B8 , 32'h0705A0E8 , 32'hFD13F9F0 , 32'hFFFD132A , 32'hB71E6880 , 32'hFFFD5319 , 32'hFEEEC230 , 32'h1F3E6B60 , 32'hFFFB18ED , 32'hFFFF43B4 , 32'h0000BD16 , 32'h0000FD85 , 32'hFFFE6517 , 32'hFFFDB3BB , 32'hF9ACFE98 , 32'h0B1F1660 , 32'hA7D7F480 , 32'hF04A1DB0 , 32'hFB1B4BB8 , 32'h1E83CDA0 , 32'h0002A101 , 32'h00020524 , 32'hFFFA34CC , 32'h0005C08E , 32'hFFFF4EA6 , 32'hF9419C20 , 32'h0BEE65A0 , 32'hEDF57300 , 32'h0002AC4A , 32'h0000F7FB , 32'hFFFE49D0 , 32'h000172B3 , 32'h0871B0F0 , 32'h263A56C0 , 32'h0006AF74 , 32'h000093B4 , 32'hFFFDDD6C , 32'hE305E140 , 32'hE18A7560 , 32'hDDB559C0 , 32'hFFFB9D6B , 32'hFFFB744D , 32'h000102D9 , 32'hFFDB6A54 , 32'hFE7D6F28 , 32'h10A50660 , 32'hFFF94E97 , 32'h0041EE3A , 32'hFFFF888E , 32'h11532E60 , 32'h000311D3 , 32'hD780CDC0 , 32'hFFFD30CB , 32'hFBBD35A8 , 32'h01368E20 , 32'hDB3B7840 , 32'h7041C580 , 32'hFFFEFA6F , 32'h0FD83CF0 , 32'hFE845744 , 32'hFFFABA69 , 32'hF83753C8 , 32'hFFFC43A3 , 32'h06861958 , 32'h14037240 , 32'h0684B980 , 32'h00067A67 , 32'h00005643 , 32'hF7C5ADB0 , 32'hFFFD2AE7 , 32'hF8A3EEE8 , 32'h0002196D , 32'hFDBDAA7C , 32'hFFFDA5C1 , 32'hF4D786C0 , 32'hFFFF035C , 32'h00000387 , 32'h000028E3 , 32'h15A1ABA0 , 32'h107D6860 , 32'hFFFDC614 , 32'hFFFE7C0B , 32'hFFFECFEB , 32'h0002384E , 32'h1C569120 , 32'h08261FC0 , 32'hF3AFD2E0 , 32'h0871B2E0 , 32'hEFC86DC0 , 32'h00058AFC , 32'hFFFDBE8E , 32'h0005BE46 , 32'hF44CFA30 , 32'hFFFDD72A , 32'hFFFBC4CB , 32'hFE6B8A00 , 32'h067C6678 , 32'h0001734B , 32'hE5C9B920 , 32'hFDC5389C , 32'hFB778150 , 32'hE82AD340 , 32'h00009571 , 32'hF69C16D0 , 32'h01E24124 , 32'hF9E75548 , 32'h0001C531 , 32'h1B7337A0 , 32'h230F9FC0 , 32'hF929C220} , 
{32'hED16D240 , 32'hECC62300 , 32'hFFFEC90A , 32'h039CA72C , 32'hFFFF43B4 , 32'hFEEEEE3C , 32'hFFFEEDE1 , 32'hFFFEEB28 , 32'h00007A62 , 32'h0005DB9B , 32'hFEB70150 , 32'hDFF1A540 , 32'h069C1C90 , 32'h00039286 , 32'h00028882 , 32'hC72DDCC0 , 32'h00000523 , 32'h1C5E17C0 , 32'h0258DDF4 , 32'hFFFBFDF6 , 32'h00011081 , 32'hFC457480 , 32'hE4C20180 , 32'hF25FD100 , 32'hF7DCDA40 , 32'hFFFE9BB7 , 32'h017516A0 , 32'hFE567DDC , 32'hFFFF939C , 32'h120648E0 , 32'hFFFFAA19 , 32'h04F906D8 , 32'h00037E78 , 32'h00023A8D , 32'hFFFF7E07 , 32'h20602C00 , 32'hFBFAA0D8 , 32'h02E24024 , 32'hFFFFF2C1 , 32'h0A7450F0 , 32'hF50F8740 , 32'h000304CA , 32'hFFFFFD69 , 32'h0ABF4BC0 , 32'h1BBBA900 , 32'h3ABB9080 , 32'h009D57F3 , 32'hFFFD41D3 , 32'hEAA2FBE0 , 32'hFEEA8F1C , 32'h013B0700 , 32'hFFF89FBA , 32'hFCBED898 , 32'h081AD4E0 , 32'hED70A220 , 32'hFFFDA737 , 32'hFA57DB40 , 32'hFFFC3395 , 32'h0003BD36 , 32'hF934BAE0 , 32'hFE450C2C , 32'h04E4C428 , 32'h3595DF80 , 32'hFFF96CB9 , 32'h1EE53F00 , 32'hFFF73644 , 32'hE871AB60 , 32'hFA9FC368 , 32'h000755BA , 32'h0223A57C , 32'h2AE4D740 , 32'h037D91C4 , 32'h0002E8BD , 32'hFFFF360F , 32'hFFFEEF58 , 32'h2864E640 , 32'h01D0506C , 32'hFFF73F8C , 32'h6A995D00 , 32'hF95BDC50 , 32'hFFFB316A , 32'hD9873740 , 32'hFF4C0ADA , 32'h00005E28 , 32'h09D5F700 , 32'hED36BBE0 , 32'h15999660 , 32'hFFFE9320 , 32'hFFFF57BE , 32'h15EE2480 , 32'hFFFE1767 , 32'hF6DDE290 , 32'h0002753C , 32'h02381E48 , 32'h007DB429 , 32'h00018415 , 32'hFFFEA827 , 32'hFFFD3448 , 32'h0005A525 , 32'h04276BA0 , 32'h04EFD300 , 32'h0001C351 , 32'hEAC40540 , 32'h0CF1E3E0 , 32'hFFE38EEC , 32'h000162C9 , 32'h0062E363 , 32'h0002F734 , 32'h1A9DF640 , 32'hED50FF40 , 32'hFFFF06FA , 32'h06F325F0 , 32'h00045990 , 32'h00027108 , 32'hEFB8AB00 , 32'hF3364D80 , 32'hF35BE580 , 32'hFFFBFCE4 , 32'hF9D8F4D0 , 32'hFFFAC4B9 , 32'h0004F1E1 , 32'h02B61EE4 , 32'h00050C68 , 32'h00016375 , 32'h323C3580 , 32'hDF2FE900 , 32'hFFFF5B4A , 32'hFFFC0CBB , 32'h000373E5 , 32'h000490E2 , 32'h00014B4E , 32'hF4130DC0 , 32'hE219B740 , 32'hFFFF3820 , 32'hFFFFC6D4 , 32'hFF4C4895 , 32'hFD2163D0 , 32'hFFFFB76F , 32'h0000992C , 32'h0FA76E70 , 32'h0001C2B6 , 32'hFFFED434 , 32'h04A53F78 , 32'hF15F45E0 , 32'hFCF813D4 , 32'hFA5B55D0 , 32'h00002B9A , 32'h0000AF18 , 32'hFA31DC48 , 32'hFFFEBDF1 , 32'h0000DFDC , 32'hFDD0323C , 32'h0001839C , 32'h0000217A , 32'h23FB9A00 , 32'h000052F5 , 32'h0609B450 , 32'h04B26000 , 32'h0001B613 , 32'hFFFC6857 , 32'h000356A1 , 32'hFE530DE4 , 32'h0597BB38 , 32'h0D247D10 , 32'h1636D540 , 32'hFFFFEDB5 , 32'h2BAC6780 , 32'h000219F8 , 32'hFFFADF20 , 32'hF1BB2190 , 32'h08F7A430 , 32'h0CE05460 , 32'hFFFEFE4E , 32'hD886ED80 , 32'h1417F1E0 , 32'hE4E2B1C0 , 32'h173A6500 , 32'hE40EC3C0 , 32'hECCDA840 , 32'h02D972DC , 32'h11B2E820 , 32'hFFFE4DD7 , 32'h0002F55B , 32'hFFFEE209 , 32'h043B3F98 , 32'h2F5CDA40 , 32'hF94F4508 , 32'hFBF0EFC0 , 32'hEBCD3240 , 32'hF2CF30E0 , 32'h0004E218 , 32'h098739B0 , 32'hF9A66538 , 32'h00003D16 , 32'hDF79ADC0 , 32'hFFF99152 , 32'hF5631CE0 , 32'hF9DF9EB8 , 32'hFFF94D1A , 32'hFFFF62AE , 32'hFFFE9396 , 32'h0008BDB8 , 32'hFFFEA898 , 32'h00029F6A , 32'hFF474D56 , 32'hFD512ED0 , 32'hEEC8D660 , 32'hFF678A72 , 32'hF744E700 , 32'hFCACAED0 , 32'hFFFF7B5C , 32'hFFFD64C1 , 32'h0002F378 , 32'hFFFE837F , 32'h0004E44C , 32'hFC848A90 , 32'hFBD2AD30 , 32'h10561F00 , 32'hFFFFD1AC , 32'h00018DEC , 32'hFFFDF6A9 , 32'h0001594F , 32'h063DC640 , 32'hF8F7B740 , 32'h00029654 , 32'hFFF9DD37 , 32'hFFFF9499 , 32'h1B228220 , 32'h44944500 , 32'h07F38398 , 32'hFFFDA4F5 , 32'h0002B235 , 32'hFFFD3552 , 32'h0CD43CC0 , 32'hFDA2E9A0 , 32'h40CA8480 , 32'hFFFD0F00 , 32'h00C6F7CF , 32'h0001E112 , 32'hE8DB5180 , 32'h0001D741 , 32'h15327960 , 32'h000618F0 , 32'h0FA40720 , 32'hDE679500 , 32'hE2ED8220 , 32'hE4C57BC0 , 32'h0001F206 , 32'h029FFDA0 , 32'hFEA2A9FC , 32'hFFF922D2 , 32'hFCB55F04 , 32'hFFFF07D3 , 32'hFBE9F538 , 32'h174F93E0 , 32'h0A866E70 , 32'h0001A266 , 32'hFFFD223B , 32'h0D83FD80 , 32'h00025FA0 , 32'h065B2228 , 32'hFFFC4AD6 , 32'h07528BA8 , 32'h00002A30 , 32'h136E3120 , 32'h0003926C , 32'h00013B17 , 32'hFFFF9B08 , 32'h012B1DB8 , 32'h02F64768 , 32'hFFFEBFD5 , 32'h000414BD , 32'h0001949D , 32'h000180B9 , 32'hF2B75470 , 32'h03FD2158 , 32'h0AF60CA0 , 32'h31EE2C40 , 32'hE9BD3A80 , 32'h00000CE7 , 32'hFFFFBA40 , 32'h0000938C , 32'h041C6D58 , 32'h000224D3 , 32'hFFFFBC49 , 32'hFEC32408 , 32'hF3A39880 , 32'h000505DD , 32'h0AFC2EC0 , 32'hFF2DF1E8 , 32'h16B8F9E0 , 32'hF3C9ADC0 , 32'hFFFEEBA2 , 32'hFF0D5C32 , 32'h355FF480 , 32'hFD4D1550 , 32'hFFFA546C , 32'h11BAC640 , 32'hC40D1F00 , 32'h12567180} , 
{32'h992DDC00 , 32'hEA1F0DE0 , 32'h00031E6E , 32'hF654DA20 , 32'h0000FF0A , 32'hFC93E904 , 32'h0004468C , 32'hFFFE195F , 32'hFFFDF089 , 32'h000328E8 , 32'hFBD8AF68 , 32'hE5074200 , 32'h12110BC0 , 32'h000405E1 , 32'hFFFAD822 , 32'hFE626838 , 32'h00020F86 , 32'hF8BE59E8 , 32'hFD816C78 , 32'hFFFB3B67 , 32'h0004E413 , 32'hFC9C1FAC , 32'hFB79C910 , 32'h012D0A48 , 32'h02E202E0 , 32'h000178D9 , 32'hFA30BFC0 , 32'hFFC8AC79 , 32'h00015EC6 , 32'hF0C16DF0 , 32'h0001F8E5 , 32'h08E59750 , 32'h00017834 , 32'hFFFF033B , 32'hFFFEB074 , 32'hD814AEC0 , 32'h1CD3B8C0 , 32'hEE7BD340 , 32'h000351DD , 32'h1D7B1320 , 32'h01A6D698 , 32'h0000DC5F , 32'h0001A0A5 , 32'hF77D47F0 , 32'hF2243E10 , 32'hA921A700 , 32'hFDFAAE30 , 32'h0000FF09 , 32'hEB14E460 , 32'h13137740 , 32'h01BC19EC , 32'h00081700 , 32'h04289380 , 32'hE626F220 , 32'h1356DBA0 , 32'hFFFE2ADE , 32'h005359EA , 32'h0007AFBD , 32'hFFFA7C06 , 32'hFDA30E40 , 32'h088E2A80 , 32'hF69E3B20 , 32'hFA0D5C08 , 32'hFFF9E1F9 , 32'hE1DB6C20 , 32'h0002158D , 32'h39F20940 , 32'h03957B88 , 32'h0000559D , 32'hF691D370 , 32'hDC7E1A40 , 32'h0F1412A0 , 32'hFFFD6324 , 32'h00037C95 , 32'h0001B4C6 , 32'h0F96CA40 , 32'h017B9398 , 32'h00031E61 , 32'hCD803640 , 32'h039F24CC , 32'h0002E669 , 32'hA080A700 , 32'hF671DBF0 , 32'hFFFE6A79 , 32'h0D6763E0 , 32'h006DE3A2 , 32'hFB8A9A08 , 32'h00050B2E , 32'h00020596 , 32'h081E7300 , 32'hFFFF16D6 , 32'hF9E64120 , 32'h0000D159 , 32'h1011FF00 , 32'hFEAC7DAC , 32'hFFFCC314 , 32'h000274E3 , 32'hFFFE73A6 , 32'h0002582D , 32'hF503A3D0 , 32'h04357250 , 32'hFFFD8003 , 32'hECD36960 , 32'hE1878060 , 32'hF4EEF9B0 , 32'h00017525 , 32'h00C02EF0 , 32'h00024BB4 , 32'h0706E218 , 32'h1B302220 , 32'h0002FB9E , 32'h18B97E00 , 32'h00053187 , 32'hFFFEE321 , 32'hF9ADF6D8 , 32'hFE3BB3D4 , 32'h020AB99C , 32'h00034A56 , 32'h041F9EF0 , 32'h0005D8D0 , 32'hFFFBFA7C , 32'hFBAFD350 , 32'hFFFE9E15 , 32'hFFFC5D32 , 32'hFF072F50 , 32'hEF472600 , 32'h00059157 , 32'h00017388 , 32'h0003EEE9 , 32'hFFFC3C80 , 32'hFFFD75A7 , 32'hFFDA30C4 , 32'h102F1980 , 32'hFFFECABC , 32'hFFFC6E93 , 32'hE1507720 , 32'hFB5C0E38 , 32'hFFFE99E4 , 32'h00066F17 , 32'hF8804DB8 , 32'h00044F7B , 32'h0004A215 , 32'h041D9638 , 32'hD321AD40 , 32'hF7E00190 , 32'hFF5228EE , 32'hFFFE8001 , 32'hFFFD4D18 , 32'h04AA0EB0 , 32'hFFFF50BB , 32'hFFF88B20 , 32'h07093E58 , 32'hFFFFE590 , 32'h00033357 , 32'hF9E75310 , 32'hFFFFBF05 , 32'h10270BE0 , 32'h0557E178 , 32'h0003CE4F , 32'hFFFC1196 , 32'h0000235E , 32'h1AE55A60 , 32'hFF3DA855 , 32'hFFD1E770 , 32'hFEF3CAB0 , 32'hFFFE3F7E , 32'hF1150C50 , 32'hFFF81B41 , 32'h000047ED , 32'hFB3E3188 , 32'hF9CE42B0 , 32'h00138580 , 32'hFFFE1158 , 32'hF0E79A80 , 32'hFEE09200 , 32'h0ABE8DE0 , 32'h13E66A60 , 32'h0FAD5E90 , 32'hEDAC06E0 , 32'h01AF4F64 , 32'h13EFDCE0 , 32'hFFFD4755 , 32'hFFFF1426 , 32'h0002B245 , 32'hF7525A70 , 32'hFE3008A4 , 32'h0435BC78 , 32'h0251D38C , 32'hF57B38B0 , 32'h02414A3C , 32'h000045DD , 32'hE50B1EA0 , 32'h163AC600 , 32'h0003BA57 , 32'hFA4D6670 , 32'h00006754 , 32'h06E4B748 , 32'hD8002240 , 32'h0000835A , 32'hFFFD67DE , 32'h0000D4B5 , 32'h00026AE1 , 32'hFFFCECD5 , 32'hFFFCE6D0 , 32'hDFA42E00 , 32'h1B2956C0 , 32'h078583A8 , 32'hEA110FA0 , 32'hE6893C00 , 32'hF99DE8D8 , 32'hFFFF8464 , 32'hFFFFB213 , 32'hFFFAF0CC , 32'hFFFF6120 , 32'h00058691 , 32'hFA862338 , 32'h0997B310 , 32'hF9D4D080 , 32'hFFFFA3FC , 32'hFFFD776C , 32'h0002D0BB , 32'h000176A0 , 32'hFCB95110 , 32'hF03A0D90 , 32'h000255E1 , 32'hFFFDA00F , 32'h0001CF55 , 32'h0A206F50 , 32'h2CEC1400 , 32'hC9751840 , 32'hFFFB9842 , 32'h00034A1C , 32'hFFFD3B53 , 32'hF61B3770 , 32'h01B784F0 , 32'hF7659040 , 32'h0002F860 , 32'h016DA548 , 32'hFFF733EF , 32'hDF3CF680 , 32'h0000B20C , 32'hF44BD570 , 32'h0000662C , 32'h0F496500 , 32'hFA2277A8 , 32'h0512FF68 , 32'hD6B59BC0 , 32'h00019D9D , 32'hFD63E6D8 , 32'h01083CF4 , 32'hFFFE4AD8 , 32'hFDE56A0C , 32'h0002D246 , 32'hF98739A0 , 32'hF44BC450 , 32'h180E0380 , 32'hFFF9B3D9 , 32'h0000A7D3 , 32'hEA5382C0 , 32'hFFFECD67 , 32'hD0700180 , 32'h0000084D , 32'hFD51B89C , 32'h0001539C , 32'h01F47E28 , 32'h00020A5F , 32'hFFFE90B3 , 32'hFFFE279D , 32'hF7EEF5F0 , 32'hFA053300 , 32'h0000B1C0 , 32'h0005DD32 , 32'h00007638 , 32'h00017088 , 32'h0038E54F , 32'hF0CF7B90 , 32'h1582C6A0 , 32'h11FE3660 , 32'hBF076C80 , 32'h000195ED , 32'hFFFFB1CF , 32'h000203A7 , 32'h0395AD64 , 32'h0002E305 , 32'h0002536F , 32'hFFE9FDFA , 32'hFD243654 , 32'h00049610 , 32'hC394B7C0 , 32'hFF0D18F4 , 32'hF5181FE0 , 32'hF7BAF080 , 32'hFFFDE5BA , 32'hF942D1A0 , 32'h125CDC40 , 32'hFBB77A50 , 32'h00048CBE , 32'h0B6CADD0 , 32'hDEA8B740 , 32'hE807BCC0} , 
{32'h3639B880 , 32'h1D6C9080 , 32'hFFFEC925 , 32'h11C39840 , 32'hFFFD5C5F , 32'hFEF36D78 , 32'hFFFED217 , 32'hFFFD2137 , 32'h00025A83 , 32'h0000C259 , 32'h1EAF86C0 , 32'hFDE975E0 , 32'h0EA4CA50 , 32'h0001D6FF , 32'h000582FD , 32'h0F7D9730 , 32'hFFFDB3CF , 32'h31DEFBC0 , 32'hFFA37A7E , 32'hFFFD61BD , 32'h0003EDCD , 32'hFB22B778 , 32'hE878D280 , 32'h0CDB8540 , 32'hF6248890 , 32'hFFFD307A , 32'hFE5BEC68 , 32'hFB896A48 , 32'h0004639C , 32'hEE0238C0 , 32'hFFFE311C , 32'hF64D1BB0 , 32'hFFFED6F5 , 32'h00021538 , 32'h0006E9CA , 32'hF1C7DA00 , 32'h18A65440 , 32'h2B3D2FC0 , 32'hFFFD729E , 32'hF6345CD0 , 32'h22FACA40 , 32'h0003FBF6 , 32'h000237C4 , 32'hFC1CA7C0 , 32'hF22D37C0 , 32'h1E4BA1E0 , 32'hFA6EE098 , 32'h0005E1BA , 32'hEB6707E0 , 32'h14658040 , 32'h00303E8D , 32'h000193DE , 32'h006447FF , 32'hC9B82E40 , 32'hFDDF9ED4 , 32'h00016B47 , 32'hF60FE070 , 32'h0000CA7D , 32'hFFFD388B , 32'hFFD1E2DA , 32'h04910740 , 32'hFFE8CE5F , 32'hFF4EAA12 , 32'h0001762F , 32'hEEEE14C0 , 32'h0002683B , 32'hFB908000 , 32'hF8602E00 , 32'hFFFE8203 , 32'h0DF30A70 , 32'hE23483C0 , 32'h07704BA8 , 32'h0003A970 , 32'hFFFFD89F , 32'hFFFB2435 , 32'h1A8D5500 , 32'hF0462A20 , 32'hFFFA134B , 32'hCA6067C0 , 32'h0330F054 , 32'hFFFEB286 , 32'h1B7F4900 , 32'hF70F7B80 , 32'h000458FC , 32'h08E190B0 , 32'h2B16AC00 , 32'h05A126E8 , 32'hFFFF7FF9 , 32'h00015508 , 32'h1F40E900 , 32'h00069D8C , 32'h0E855340 , 32'hFFFD99FA , 32'hF9B93820 , 32'h0055A2F5 , 32'h00002740 , 32'h00012B47 , 32'h00038E85 , 32'h0000548A , 32'hFBD1B1B0 , 32'hF952B880 , 32'hFFFFC6C5 , 32'hF005E700 , 32'hDF420E80 , 32'hF9CDAE70 , 32'h0000324E , 32'h016045E4 , 32'h0002E40B , 32'hFC52DDAC , 32'hD4B0FFC0 , 32'hFFF8EA99 , 32'h32C78F80 , 32'h0002DFBE , 32'hFFFFB57C , 32'h27967A00 , 32'hF67B3980 , 32'h053F8100 , 32'h0003AF3B , 32'h1500BF80 , 32'hFFFF5EE8 , 32'h00031F75 , 32'h153E68C0 , 32'hFFFF388F , 32'h0002A596 , 32'hF72169E0 , 32'hE1209BA0 , 32'h000134A1 , 32'h0004A7D6 , 32'h000297C9 , 32'h00052FBC , 32'hFFFA9036 , 32'h043F1660 , 32'h0AAEF930 , 32'h0005EDE9 , 32'hFFFEE908 , 32'hDCCD0DC0 , 32'h05C5CDB0 , 32'h00000C61 , 32'h0000F238 , 32'hF4154790 , 32'h0001A6D8 , 32'h0002D181 , 32'hFA29AAF0 , 32'h10076400 , 32'hFA36BCB8 , 32'h0351B8CC , 32'h00001FE2 , 32'hFFFD3B24 , 32'hFADBEC48 , 32'hFFFE9089 , 32'h00034788 , 32'h03A83754 , 32'hFFFB06AA , 32'h0002C848 , 32'hD4D42840 , 32'hFFF39CD9 , 32'h02B456A8 , 32'hFB9F92D0 , 32'hFFFE49FB , 32'h00014F1F , 32'hFFFCE7A3 , 32'h12F34120 , 32'hF5E1B960 , 32'hFED35730 , 32'hF4F17460 , 32'hFFFDB0EA , 32'h0DEE3700 , 32'hFFFACD78 , 32'hFFFFD95C , 32'h0243CCA8 , 32'h0AE512F0 , 32'h0153036C , 32'hFFFF55BC , 32'hFFC2684C , 32'hFF7B101F , 32'hF5850AD0 , 32'hFA69C498 , 32'hE4A18BC0 , 32'hF07558F0 , 32'hFEB3A044 , 32'hF8737CE8 , 32'hFFFC74AB , 32'h000025DE , 32'hFFFE0519 , 32'h0240D344 , 32'hFF787FAB , 32'h09328DE0 , 32'h0739BAB0 , 32'hFD2B6790 , 32'h019C054C , 32'hFFF566B3 , 32'h1BFCB720 , 32'h0F530200 , 32'h00007813 , 32'h2EDA19C0 , 32'hFFFDE7C8 , 32'hED00E500 , 32'hEB97FBA0 , 32'h0002EA5F , 32'hFFFB880B , 32'h0001E762 , 32'h000159FF , 32'h00005F5E , 32'hFFFEB8E7 , 32'h0A324DC0 , 32'h1C0B7260 , 32'hCED03440 , 32'hE4B8C4C0 , 32'h12892A20 , 32'h0FA1F820 , 32'h000022F7 , 32'h0002B571 , 32'hFFFDF858 , 32'h0000EB1B , 32'hFFFF7B03 , 32'h08A98680 , 32'h000684AF , 32'h36268980 , 32'hFFFCC148 , 32'h0002DDD4 , 32'h0002D0F7 , 32'h00026F6A , 32'h04357B40 , 32'h0D17C160 , 32'h000063AB , 32'h0006E53D , 32'hFFFFB670 , 32'hE7C06A20 , 32'h3AA77AC0 , 32'hF38B32F0 , 32'hFFFA6F07 , 32'hFFFB42D7 , 32'h00002B44 , 32'hFE5FB9D0 , 32'hEF0BFB40 , 32'h3244AAC0 , 32'hFFFF14EC , 32'hFE4B34D4 , 32'h0002E818 , 32'hDA171140 , 32'h000197E4 , 32'h34CE8E80 , 32'h00014177 , 32'hFD52BF94 , 32'h0F6A6850 , 32'h3F346840 , 32'hDDE1DBC0 , 32'hFFFBA15C , 32'h00C42768 , 32'h027ED0E4 , 32'hFFFC519D , 32'h10FAF920 , 32'hFFFABF5F , 32'h063D7F90 , 32'h0B7B7A70 , 32'hF960EFB8 , 32'hFFFEDBBF , 32'hFFFD77A0 , 32'hFFF2B9D2 , 32'h00021EAD , 32'h0D6F5CB0 , 32'hFFFA6988 , 32'h01C50FA8 , 32'h00032264 , 32'hE71AB280 , 32'h000426DC , 32'h000216C3 , 32'h0001784A , 32'h2AC5BDC0 , 32'h17FEFDE0 , 32'hFFFD2968 , 32'hFFFFEEAF , 32'h00040C01 , 32'hFFFCCC9D , 32'hEDF84FA0 , 32'hEE9C2280 , 32'h126D2640 , 32'h0FFC0DE0 , 32'h1EEA9460 , 32'hFFFBE024 , 32'h0003A6FA , 32'h00006493 , 32'hFA878908 , 32'h000440CB , 32'h00039D99 , 32'hF7E5BFA0 , 32'h2D05F440 , 32'h0003099E , 32'h200DCC80 , 32'hF8A66360 , 32'hF836FB98 , 32'hF3F9BF90 , 32'hFFFEFC0F , 32'hF06EAB50 , 32'h02FAF54C , 32'h03BCD568 , 32'h0006B3E7 , 32'h1B9111C0 , 32'hF78A9070 , 32'hD0D7DA00} , 
{32'hD1C9C280 , 32'hE95C2F60 , 32'h0000F13B , 32'hEA95B700 , 32'h000265CE , 32'h0248BAF0 , 32'h00064FEF , 32'hFFF867B1 , 32'h0000B9F9 , 32'hFFFF0954 , 32'hFDFE9E88 , 32'hF102E410 , 32'hE98852A0 , 32'hFFF6B50F , 32'hFFFB2FB1 , 32'hEED17AE0 , 32'hFFFAB17D , 32'h117CB580 , 32'hEF7FA740 , 32'h0001B94A , 32'hFFFF41CD , 32'h04373F00 , 32'hE861A8C0 , 32'hF2D3F760 , 32'h1D7035C0 , 32'h000053F8 , 32'h0430EDB0 , 32'h00BF274A , 32'hFFFD835C , 32'h18BDCA00 , 32'h0003ECF6 , 32'h177DCFC0 , 32'hFFFFFEB4 , 32'h000090C0 , 32'hFFFEC558 , 32'h07675D48 , 32'h12890A60 , 32'h0B0395E0 , 32'hFFFFF25D , 32'hFD2E4F8C , 32'hFF100D71 , 32'h00017EB2 , 32'hFFFF39D8 , 32'hFAF93390 , 32'h0612B8E8 , 32'h29ECFE80 , 32'h04863A58 , 32'h00034F0D , 32'hF8B6F530 , 32'h11AD2880 , 32'hFE0A34D8 , 32'hFFF6523F , 32'hF47D4840 , 32'hFBE2C1D8 , 32'hFCAC7B54 , 32'h0000ABEE , 32'h06092988 , 32'h0005F6B3 , 32'h0001448B , 32'h091C3640 , 32'h01AB7DDC , 32'h05C7E6B8 , 32'hE8B135C0 , 32'hFFFDAAC6 , 32'h14A42660 , 32'h00017D89 , 32'hE9346BC0 , 32'h049BE348 , 32'hFFFFBB3D , 32'h9E237480 , 32'hF76CF450 , 32'h02C50540 , 32'hFFFE10BD , 32'h0008C457 , 32'hFFF9C897 , 32'hDDD0EA00 , 32'h078908E8 , 32'h0003072F , 32'hFFD84401 , 32'h01D23220 , 32'h0000E4C0 , 32'h09D94180 , 32'h0FDA9790 , 32'h00016166 , 32'hF0EDCE50 , 32'hFC9EBBD8 , 32'h00470BB8 , 32'h0004201D , 32'h0000BAE4 , 32'h1A4D9900 , 32'hFFF6DCDC , 32'h092FFF40 , 32'h0001F28F , 32'hFC77E8F4 , 32'h006D76E8 , 32'hFFFA7837 , 32'hFFFDEA2A , 32'hFFFE1107 , 32'h0001AFBD , 32'h06CFCE40 , 32'hF89590F8 , 32'h0001F4D6 , 32'hE80DC080 , 32'hB6F82780 , 32'h038E11A4 , 32'h00019139 , 32'hFECCCF88 , 32'hFFFFD68F , 32'h04E3DF30 , 32'h1B787F60 , 32'h00020F6A , 32'h17BAB900 , 32'hFFFFA298 , 32'h00036FB0 , 32'h19A83F40 , 32'hFF1D4D92 , 32'h05F8C6C8 , 32'h0001FC8C , 32'h07020B50 , 32'h0001B561 , 32'h00074D9E , 32'h016A9700 , 32'h00011ACF , 32'hFFF9C932 , 32'hD9C4A080 , 32'hFA553AD8 , 32'h0003F4DB , 32'hFFFCF4E5 , 32'h00002035 , 32'hFFFBB717 , 32'hFFFD4D9C , 32'h012D1464 , 32'hF6C0BAB0 , 32'h0002D9B3 , 32'h00054BDC , 32'hD0040840 , 32'hE05725E0 , 32'hFFFD242D , 32'h0000096C , 32'h0D133B40 , 32'hFFFF93C1 , 32'hFFF9D8E0 , 32'h04340EF0 , 32'hF86104C8 , 32'hFF019411 , 32'h082AB5B0 , 32'h00005870 , 32'h00015D4E , 32'h006D738E , 32'h000256E2 , 32'h0006B6C9 , 32'h040DB478 , 32'h0001F452 , 32'h000172C0 , 32'hE1C3EE80 , 32'h0002E031 , 32'hFCC63D14 , 32'h03C83A5C , 32'hFFFA675F , 32'h0003968F , 32'h000433C3 , 32'hF9F87668 , 32'h041F0CC0 , 32'h04C3C360 , 32'hFC4CCEB8 , 32'hFFFAFEB5 , 32'hE5D740E0 , 32'hFFFB908A , 32'hFFFD55D2 , 32'h01AAC1B0 , 32'h07495F68 , 32'hEFE49AC0 , 32'hFFFFE897 , 32'h33ACF680 , 32'hF9B7AD90 , 32'h110D3900 , 32'h0BD9CBC0 , 32'hDFD8A840 , 32'h110824A0 , 32'h043F5038 , 32'hD51446C0 , 32'hFFFF2125 , 32'h000270F8 , 32'h0000BFF0 , 32'h08EA9A00 , 32'hDB184AC0 , 32'hFAD422F8 , 32'h01AF0904 , 32'h091FF700 , 32'h012D4234 , 32'h00084039 , 32'hF79588A0 , 32'hF9C3E030 , 32'h0000647A , 32'hCC70E0C0 , 32'hFFFF2C79 , 32'h019AAB44 , 32'h22FCF300 , 32'hFFFCFC1D , 32'hFFFDC8E8 , 32'hFFFFD40B , 32'h0000B6FE , 32'h0001DCF2 , 32'h00025267 , 32'h03FA56E4 , 32'h364362C0 , 32'hF4EA2550 , 32'hFE3F2A78 , 32'h03F2DDE4 , 32'hD55E03C0 , 32'h00008A5D , 32'hFFFF12F6 , 32'hFFFF7CE7 , 32'h0003DB68 , 32'hFFFE05C8 , 32'h0071E0CF , 32'hE840FEC0 , 32'h01A2A318 , 32'hFFFFBE6C , 32'h00016318 , 32'hFFFD718F , 32'h0002935A , 32'h08F3C050 , 32'hD14C63C0 , 32'hFFFF2F7D , 32'hFFF8EAA8 , 32'h0006049F , 32'h111A6FE0 , 32'hDE711580 , 32'hF3C30720 , 32'h0000FCAD , 32'hFFFF042B , 32'h000061D3 , 32'h035C1CFC , 32'h01D21338 , 32'h022511B4 , 32'h0000A6E4 , 32'h006028E7 , 32'hFFFBF214 , 32'hD54D6B80 , 32'hFFFF63A2 , 32'hE97CCBE0 , 32'h0002AA53 , 32'h037E85C8 , 32'hFD896854 , 32'h07ADEDD8 , 32'h331AEC00 , 32'h0005C1D9 , 32'h06D966B0 , 32'hFC51D068 , 32'h0000B9B4 , 32'hFBA4F2F8 , 32'hFFFF65D8 , 32'h0A180F30 , 32'h3F3292C0 , 32'h10B157C0 , 32'h000240BE , 32'hFFFD389A , 32'h17C496C0 , 32'h00000481 , 32'h06BFB570 , 32'h0000DF08 , 32'h02D9EFE8 , 32'h0001E3B6 , 32'hF4B734B0 , 32'hFFFF1459 , 32'h00006BBA , 32'hFFFDB257 , 32'hFB0390A0 , 32'h11ECA6C0 , 32'h000044AA , 32'hFFFFAF66 , 32'h0003A5D4 , 32'hFFFF233C , 32'hF5769600 , 32'h1A429280 , 32'hDD92BC80 , 32'h082EF4A0 , 32'hCAA62EC0 , 32'hFFFC45B2 , 32'hFFFBD266 , 32'hFFFF41F3 , 32'hFC41102C , 32'hFFFC7BDA , 32'hFFFBB27A , 32'hFA8AA810 , 32'h020FD8D0 , 32'hFFFEC764 , 32'h4F526A00 , 32'hFBB58FD0 , 32'h130313C0 , 32'h0B54AC00 , 32'hFFFC9DD8 , 32'h0A22D7F0 , 32'h05F06C28 , 32'hFFA86FB1 , 32'hFFFA57AA , 32'hE4DEDA20 , 32'hF49EEA70 , 32'hF34C1140} , 
{32'h05EFB458 , 32'h0EE42890 , 32'h00035B2D , 32'h10E42660 , 32'h00015CBA , 32'hF883F688 , 32'hFFFC3E00 , 32'hFFFDC132 , 32'hFFFBD9B8 , 32'h0002D8E2 , 32'hE477E6A0 , 32'h04F778C8 , 32'hFB463410 , 32'hFFFB9CF5 , 32'h0001F0D2 , 32'hEC73D1A0 , 32'h00045ACD , 32'h03FFC1A8 , 32'h0CE2DE50 , 32'hFFFF20F7 , 32'h0001F984 , 32'hFC4F5820 , 32'h2EA644C0 , 32'hF7675920 , 32'h00AB0A19 , 32'h0000F317 , 32'h024B7A78 , 32'h0313DF2C , 32'h0004BFFD , 32'hEB03C8A0 , 32'hFFFED7A9 , 32'h04089900 , 32'h0007DAFE , 32'h00019686 , 32'h00042FBF , 32'h9A35B280 , 32'h1EDEEEA0 , 32'hF78FC910 , 32'hFFFE219B , 32'h07602558 , 32'h03FCD770 , 32'hFFFD4536 , 32'h00017630 , 32'h0535DB78 , 32'h4A761180 , 32'h3D3D7540 , 32'hF2273F70 , 32'hFFFBEE40 , 32'h0126EAB8 , 32'h1BAE95C0 , 32'h0081A26A , 32'h0005F13C , 32'h0B836870 , 32'h02636EF0 , 32'h089B0C60 , 32'hFFFD761C , 32'hFBBCF6B8 , 32'hFFF73E68 , 32'h0001E0AC , 32'hFB197230 , 32'h0317338C , 32'hF54CA0A0 , 32'h0B6BBD80 , 32'h000043DD , 32'hB7D07C80 , 32'h0004DC00 , 32'hF2C8C1A0 , 32'h009E0D8B , 32'hFFFDF8B1 , 32'hE27CC180 , 32'h02A14A7C , 32'hD951C240 , 32'h0002A101 , 32'hFFFD1189 , 32'hFFFB61AB , 32'hE33786A0 , 32'h01A53490 , 32'hFFFE3001 , 32'hBC039D00 , 32'h02192778 , 32'h00029744 , 32'hE1B56FE0 , 32'hDC08F900 , 32'hFFFBD80E , 32'h02819C08 , 32'h01FE9524 , 32'hFE1FAEB8 , 32'h00007172 , 32'h0004A70C , 32'h0B9DF510 , 32'hFFFB62CD , 32'h090AD990 , 32'h00010714 , 32'h08B267C0 , 32'h00E1C241 , 32'hFFFAF174 , 32'hFFFD9645 , 32'h0002FA65 , 32'h0004C6B7 , 32'h17AD41A0 , 32'hF89FE140 , 32'hFFFFB39C , 32'hE94B67E0 , 32'h1F4FCD80 , 32'hEE536780 , 32'hFFFC0F3B , 32'hFF2AD11A , 32'hFFFF9A63 , 32'hF7D5CC90 , 32'hDD8C6D00 , 32'hFFFE1196 , 32'hFDB564AC , 32'h0005A574 , 32'h0005D425 , 32'h04DA57E8 , 32'hFAA96E10 , 32'h06141F10 , 32'hFFFF07B0 , 32'hFD0BB4D8 , 32'hFFFC9B45 , 32'hFFFD682C , 32'h0254E25C , 32'hFFFBFE3F , 32'hFFFFB300 , 32'h124BB420 , 32'h06E33B08 , 32'h0001F246 , 32'h0002169D , 32'h0003E1BC , 32'h00005B8F , 32'h00004058 , 32'hF65D6850 , 32'hE947A820 , 32'h00045AC4 , 32'h0002B0F4 , 32'h15DD8560 , 32'hFCD4D200 , 32'hFFFBD313 , 32'h0001340B , 32'h07ED1180 , 32'hFFFA4D6F , 32'h00000414 , 32'hF9811FE8 , 32'hF479A370 , 32'hFC966A8C , 32'h0584A2A0 , 32'hFFFD270B , 32'h000242CA , 32'h03359A0C , 32'hFFF93DC4 , 32'h0000E4DB , 32'hFA359F60 , 32'hFFFBF40E , 32'h0002EF38 , 32'h01A43AD4 , 32'hFFFCA274 , 32'h07EE59D0 , 32'h060865A0 , 32'h0001653F , 32'hFFFE45A7 , 32'hFFFDC53C , 32'h07756B90 , 32'hF70E1DE0 , 32'hFE30ED60 , 32'h02CA3278 , 32'h00024F5A , 32'hF2079500 , 32'hFFFF8AD5 , 32'h00089F46 , 32'h0F3E1210 , 32'hFD567F90 , 32'h01B55150 , 32'h00047826 , 32'hFF60C9BA , 32'h021CA634 , 32'hE04D4080 , 32'hE865E560 , 32'h093741D0 , 32'hFA524DD8 , 32'h028DC620 , 32'hCDCA58C0 , 32'hFFFA243B , 32'h000155ED , 32'h00029EEC , 32'hE8406520 , 32'h2FB90C80 , 32'hFA9578E8 , 32'hF94A3FF0 , 32'h0EA24EB0 , 32'hFCDE4EEC , 32'hFFF7BEBD , 32'h151DD820 , 32'h036F22D8 , 32'h0001A4B6 , 32'hD90A18C0 , 32'hFFFDDEC5 , 32'h02B2C9D4 , 32'hF65CDA20 , 32'h0008C5E9 , 32'hFFF94130 , 32'h00011E85 , 32'hFFFFD53C , 32'h00000031 , 32'h0000EF22 , 32'h0F511780 , 32'hC883D340 , 32'hC1641B00 , 32'hFE8BF5E0 , 32'h15D64800 , 32'hD8FE18C0 , 32'h0001FD85 , 32'h00003F8C , 32'hFFFE976C , 32'h000027FB , 32'h00058D38 , 32'h0A651290 , 32'hEAFB96E0 , 32'hF4BE6450 , 32'hFFFECEBF , 32'h00025EC7 , 32'hFFFFFA5C , 32'h0003D9B9 , 32'h11E157C0 , 32'hE1B3D1C0 , 32'h0000AF56 , 32'h0005D3D5 , 32'hFFFE9351 , 32'h09457200 , 32'hF7C39D40 , 32'hEDB44BA0 , 32'hFFFCA93C , 32'h0006311E , 32'hFFFF388F , 32'h030DFC7C , 32'h02778AD0 , 32'hF7D2E8E0 , 32'hFFFC30A4 , 32'h02BFE11C , 32'h00013ECF , 32'hF89A7AF8 , 32'h00059E92 , 32'h156BB400 , 32'h0001B539 , 32'h0361F568 , 32'hFE5AF568 , 32'hBB5E5180 , 32'hF5B03430 , 32'hFFFEC7B2 , 32'h14D3BE20 , 32'hFECD47C0 , 32'h00010CAE , 32'hF65BB160 , 32'hFFFDC38B , 32'h070E3890 , 32'h276C5600 , 32'h06A569F8 , 32'hFFFA4A8E , 32'hFFFF47F5 , 32'h0EF39E20 , 32'hFFFC9698 , 32'h262F4FC0 , 32'hFFFB0A9C , 32'h03E437E4 , 32'h00010E50 , 32'h160E2A00 , 32'h0006CEAC , 32'h000609F2 , 32'h00011826 , 32'hF8ADBEA8 , 32'hF4D034A0 , 32'h000230CA , 32'h000623A9 , 32'hFFFCFBEB , 32'h0001B772 , 32'h0675C4F0 , 32'h0BD66B60 , 32'h004A8D0E , 32'hF0BA7EC0 , 32'hFBA34028 , 32'hFFF96A38 , 32'hFFF9E684 , 32'h000098A3 , 32'h0052BE77 , 32'h0000F3C9 , 32'hFFF81824 , 32'h03085A00 , 32'h06111D08 , 32'hFFF67507 , 32'hD9C4CCC0 , 32'h04F3AAF8 , 32'hF84CF0D0 , 32'hF5F544B0 , 32'hFFFDE0F6 , 32'h0AA66DB0 , 32'h09667FC0 , 32'hFAA32F48 , 32'hFFFFEFD3 , 32'h0BE63340 , 32'h2ABECBC0 , 32'hF7F422A0} , 
{32'hFD7115F4 , 32'h1683C5A0 , 32'h0001E6A6 , 32'h0A6F9F00 , 32'hFFFB2310 , 32'h06248B40 , 32'hFFFA5A72 , 32'hFFFD7CD1 , 32'hFFFE4E2A , 32'hFFFDFE3D , 32'hEC1CAB40 , 32'hE9E1F400 , 32'h0CB86D80 , 32'h00044700 , 32'h00054C89 , 32'hF90BF8A0 , 32'h0005B777 , 32'hEEA1E640 , 32'h034C73DC , 32'h00037727 , 32'h00013CE9 , 32'hF32FD000 , 32'h01F0DC28 , 32'hFA059AB8 , 32'h033E73F4 , 32'hFFFF12CF , 32'h00C273FC , 32'h0277E678 , 32'hFFFF61F9 , 32'hF6753580 , 32'hFFFF2974 , 32'hF0714F50 , 32'h000504A6 , 32'h00006C66 , 32'hFFFE10C3 , 32'h031C6F68 , 32'h083FDD10 , 32'hF5ED3540 , 32'h0004DC62 , 32'h001D6B4D , 32'h22DBA440 , 32'hFFFEB32C , 32'h0001F8C8 , 32'h0CA546C0 , 32'h04D1AFA0 , 32'hE3AE8DC0 , 32'h2E703D40 , 32'hFFFA82BD , 32'h00C2574F , 32'hFDA2014C , 32'h01593B8C , 32'hFFFA8E41 , 32'h06CC4C70 , 32'h089772F0 , 32'h174CE2E0 , 32'hFFFE4E2B , 32'hFD9141F8 , 32'hFFFCEDF5 , 32'h000167AF , 32'hF3CAF870 , 32'h0BAB4540 , 32'hED07EAE0 , 32'h16E82240 , 32'hFFFFDD37 , 32'hEB6C9680 , 32'hFFF99ADB , 32'hDD4289C0 , 32'hF67B18C0 , 32'hFFFD75E6 , 32'hF3446BE0 , 32'h0F5D21D0 , 32'hFAC83B50 , 32'hFFFFCCF6 , 32'hFFFC5032 , 32'h00011389 , 32'hF4F5C2F0 , 32'hFF784D5B , 32'hFFFD138C , 32'hBCE9CA00 , 32'h010A255C , 32'h000436A4 , 32'hDB56B800 , 32'hFBDF7458 , 32'hFFFFAA26 , 32'h07EEA4B8 , 32'h08CC9F10 , 32'hEFCEE920 , 32'hFFFDC969 , 32'h0000A0BA , 32'hE2CC8120 , 32'h00037802 , 32'h056FF320 , 32'hFFFE2631 , 32'h135976E0 , 32'h012A2390 , 32'h00037319 , 32'hFFFEB367 , 32'h000180A9 , 32'h0002ED62 , 32'h00F19B65 , 32'h04E88C70 , 32'hFFFF75F7 , 32'hFEF7FCB0 , 32'h1DDB5000 , 32'hF0D500E0 , 32'hFFFF266D , 32'hFD386844 , 32'h0003DBB2 , 32'hF1B834E0 , 32'hD7AA5B00 , 32'hFFFE870E , 32'h0D82A770 , 32'hFFFBB6F3 , 32'h0001807E , 32'hF195ABE0 , 32'h099991B0 , 32'h016252C0 , 32'hFFFE71AF , 32'hE9C14C60 , 32'hFFFEE3ED , 32'hFFFD368E , 32'h05AFC9C0 , 32'h0001A93F , 32'h0001D9D3 , 32'h24A62EC0 , 32'h0A430A70 , 32'h0000AE84 , 32'h000654A8 , 32'h00003166 , 32'h000181A0 , 32'hFFFBE4C0 , 32'hFDB3161C , 32'h06B8E960 , 32'h0000B0A0 , 32'hFFFD1A7C , 32'hD06B3B00 , 32'hF8CFA348 , 32'h0003CCB9 , 32'hFFFEF494 , 32'h08E38870 , 32'h0002AE84 , 32'hFFFED64F , 32'hFCD0CE88 , 32'hFC6686A8 , 32'h02D586B4 , 32'hFAD432E8 , 32'hFFFED9B6 , 32'h000092C8 , 32'hFBCE5AE0 , 32'hFFF9B440 , 32'hFFFE547A , 32'hFC50C480 , 32'hFFFC8FEE , 32'hFFFBAD2D , 32'h29789A40 , 32'hFFF823C5 , 32'hE74AE140 , 32'h0026337D , 32'h000252C1 , 32'hFFFED0F0 , 32'hFFFEB0A6 , 32'h097A04A0 , 32'hF278A530 , 32'hF4C84D50 , 32'hEE15D1C0 , 32'hFFFFA15B , 32'hEC3240E0 , 32'h00017174 , 32'hFFFEE19F , 32'h0016B3EC , 32'hFFCDA66C , 32'h00EF1CD6 , 32'hFFFD4414 , 32'hFC4FC920 , 32'h00ABCFE1 , 32'h0AC4B050 , 32'hFC553A0C , 32'h286EB3C0 , 32'h219E9440 , 32'h020B9228 , 32'hF7B3A730 , 32'hFFFB817F , 32'h0003C418 , 32'h000169CF , 32'hFE587C8C , 32'h47C86E00 , 32'hFC216C08 , 32'hFF9534EB , 32'h036C04EC , 32'hF80A6ED8 , 32'hFFFFE840 , 32'h1CE97140 , 32'h0F3C2180 , 32'hFFFBC226 , 32'h357CBC40 , 32'hFFFFCAD5 , 32'h0F715AA0 , 32'h46B16F80 , 32'h0002C1C3 , 32'h00007787 , 32'hFFFF5ADE , 32'h00012C47 , 32'hFFFE56EC , 32'h00006C6D , 32'h03D3488C , 32'h34724780 , 32'h0AD2D2F0 , 32'hFDFE989C , 32'hFA41E470 , 32'h19FB00A0 , 32'hFFFD3C60 , 32'h00002CE6 , 32'hFFFF7CCE , 32'hFFFFBEF6 , 32'h000056AB , 32'hF0215240 , 32'h1A39D500 , 32'hC40D9E00 , 32'h0004D896 , 32'hFFFD5D4F , 32'h000167C8 , 32'hFFFC7ADD , 32'h0F370590 , 32'h0BC414E0 , 32'h0006335E , 32'h0001F825 , 32'hFFF7C4EC , 32'h0327B170 , 32'hF84261F0 , 32'h0A6DBAE0 , 32'hFFFD9B02 , 32'h0007739D , 32'h000001FC , 32'hFED7DEF4 , 32'hFE86A888 , 32'h0182C680 , 32'hFFFFE7F0 , 32'hFE6617D8 , 32'h00018745 , 32'h15C39480 , 32'hFFFE7973 , 32'h115111A0 , 32'hFFFF4243 , 32'hF3601540 , 32'h0B0C4250 , 32'h0ECCE880 , 32'h47957100 , 32'hFFFFFCB1 , 32'h00E9EE7D , 32'h031F62EC , 32'h00041DE6 , 32'hEEE442A0 , 32'hFFFE09AE , 32'h037F5284 , 32'hFC326358 , 32'h191AD540 , 32'hFFFD8FCD , 32'h000300BF , 32'h02642558 , 32'hFFFD344F , 32'h10CBD9A0 , 32'hFFFE1F7F , 32'hFFEF050D , 32'hFFFCB092 , 32'h02C44A34 , 32'h000050A2 , 32'hFFFC5121 , 32'h0000FDAC , 32'h20015540 , 32'h03DD9F80 , 32'hFFFD577C , 32'h0000F0A1 , 32'h0000F833 , 32'h00067889 , 32'h0134EE34 , 32'h10E934C0 , 32'h00303018 , 32'h21B52AC0 , 32'h09091790 , 32'h00032792 , 32'hFFFD3DAB , 32'hFFFD386C , 32'h08B036B0 , 32'h00082486 , 32'h00000087 , 32'h0421D448 , 32'h11142000 , 32'h0005B916 , 32'h3E549F00 , 32'h058CD4C0 , 32'h03BB0018 , 32'hFB139518 , 32'h0004888C , 32'h00BB5ABB , 32'h09E65590 , 32'h03A2D7E8 , 32'hFFFCD5AD , 32'hF1B754D0 , 32'h9228A300 , 32'h223F5CC0} , 
{32'hCBBD1980 , 32'h1B2E3EA0 , 32'hFFFBFCDC , 32'h014811A4 , 32'h000178BA , 32'h01ABC6E0 , 32'hFFFCA00D , 32'h0002E0DB , 32'h000101FB , 32'hFFFF9083 , 32'h02D2337C , 32'h0E331960 , 32'hF5085760 , 32'hFFFE2253 , 32'hFFFC926A , 32'h0F7B6850 , 32'hFFFF5DF2 , 32'hFF14389D , 32'hFA049CE8 , 32'hFFFF2BF3 , 32'h0001CDAC , 32'h0534D858 , 32'hEC935320 , 32'h07E8BC38 , 32'h1BCD4980 , 32'h0000CAB8 , 32'hFEAD35A4 , 32'h03B0AFF8 , 32'hFFFDCD43 , 32'h0956AF10 , 32'h0002734D , 32'hF9DC1890 , 32'hFFFCB8FB , 32'h000440D9 , 32'h0000334C , 32'hE74C2D60 , 32'h0B6FE960 , 32'hE1DDDA40 , 32'h00021FFF , 32'hF766AAA0 , 32'hEE79DF40 , 32'hFFFE6347 , 32'hFFFDB8AF , 32'h06C9BAB8 , 32'h1DF29920 , 32'h715C8F00 , 32'h17ADB8E0 , 32'h000126DB , 32'h05E219B8 , 32'h07E85AA8 , 32'hFE9E46B4 , 32'hFFFA2FBD , 32'hF8BB49D0 , 32'hF756C5F0 , 32'hF0038940 , 32'h0003BFBE , 32'h04953F60 , 32'hFFFDDCEE , 32'h00040CC6 , 32'h0277A3A4 , 32'hFCE8410C , 32'h04A11238 , 32'hEF2F37A0 , 32'hFFFFC1F6 , 32'h193425A0 , 32'h0000106E , 32'h081E7260 , 32'h04FADE88 , 32'hFFFE6D0E , 32'h23BC37C0 , 32'h0C83CE10 , 32'h06EB0608 , 32'h0006225E , 32'hFFFD2B94 , 32'h00074DC6 , 32'h119142A0 , 32'hFEEFB424 , 32'h00019E8B , 32'hEAD87A60 , 32'h00FA18EB , 32'hFFFDE5F7 , 32'hD0354740 , 32'hFE7A90F8 , 32'hFFFC83DC , 32'h05F13CB8 , 32'h02C320B0 , 32'h03FCC7B8 , 32'h00024295 , 32'h00052E90 , 32'hF1DEBE90 , 32'hFFFFE13B , 32'h100A6820 , 32'h000178CA , 32'hF3925420 , 32'h004CA007 , 32'h000318EB , 32'hFFFDAD37 , 32'hFFFD24A7 , 32'hFFFBC3E4 , 32'h075EDD70 , 32'h00ADEFAF , 32'hFFFDB06F , 32'h0345799C , 32'hEC577500 , 32'h03BD0108 , 32'h000330E3 , 32'hFE5DEEDC , 32'hFFFFE5E7 , 32'hFD4F9D10 , 32'h186E21E0 , 32'hFFFCB9DC , 32'h29EE9000 , 32'hFFFB0973 , 32'h0001327D , 32'h0FD3DAD0 , 32'hF0C16660 , 32'hFCE80494 , 32'h0001C1A1 , 32'h0AC20760 , 32'hFFFE52AF , 32'hFFFF85CA , 32'h0BBF6230 , 32'hFFFD4DF7 , 32'h00040EEA , 32'hF8846318 , 32'h00F02C4E , 32'h00039142 , 32'hFFFD86D5 , 32'hFFF61D9C , 32'h00034717 , 32'hFFFD2D4C , 32'h13F650E0 , 32'h0DBA41E0 , 32'hFFFF32C8 , 32'h00057D64 , 32'h1A161760 , 32'hF816A388 , 32'h0002EB46 , 32'hFFFCCA48 , 32'hF894EFC0 , 32'h0000BA59 , 32'hFFFE78A6 , 32'hFB018040 , 32'hF3CF1650 , 32'hFFB80A41 , 32'hFD62006C , 32'hFFFE4BC3 , 32'hFFFFC963 , 32'hFE47F504 , 32'h0004F4F4 , 32'h0000EF20 , 32'h10145980 , 32'h000033DE , 32'h0002BC85 , 32'hEFA12C20 , 32'h00045B9F , 32'hFC258214 , 32'hFB9B9380 , 32'hFFFBAB35 , 32'h00010EF0 , 32'hFFFFD747 , 32'h0F192B10 , 32'hF04E2440 , 32'h049BB3A0 , 32'h05335A98 , 32'hFFFD5671 , 32'h1E2A1FC0 , 32'hFFFE8571 , 32'hFFFDD862 , 32'hFE79051C , 32'h008E60D5 , 32'hF55A3CC0 , 32'h00035D77 , 32'hCF8F3C80 , 32'hF6827760 , 32'hFE643934 , 32'hF595C1B0 , 32'hF97AA6B0 , 32'h23E48C80 , 32'hFFC3FC55 , 32'hFD9A4788 , 32'h0000B1C4 , 32'h00037170 , 32'h00039EF2 , 32'hFFDA837D , 32'hCB096B80 , 32'h0495F678 , 32'h03161EDC , 32'h087007D0 , 32'hF8458C08 , 32'hFFFDFA3E , 32'h010E56C4 , 32'h03057114 , 32'hFFFBB15B , 32'h3D3440C0 , 32'hFFFE84BA , 32'hEF1BEFC0 , 32'h11DACA80 , 32'hFFFCF73D , 32'hFFFDD6DD , 32'hFFFE114C , 32'h0000EC43 , 32'h00011576 , 32'hFFFF417C , 32'h045A2768 , 32'hB53FC080 , 32'h3AFCBEC0 , 32'hFF30AAA7 , 32'h08922910 , 32'hF3112970 , 32'h00025739 , 32'h0000B3FB , 32'h00001B01 , 32'h000144C2 , 32'h0000316A , 32'hF18FF830 , 32'h02895480 , 32'h1C5EF900 , 32'h0000B042 , 32'h00007CFF , 32'h00022012 , 32'hFFFF45CE , 32'h01125494 , 32'h3A8E8A80 , 32'h0003BE09 , 32'hFFFD8675 , 32'h000467F6 , 32'h177AD540 , 32'hFD3E9850 , 32'h13DC0C20 , 32'h0002697F , 32'hFFFE6B4A , 32'hFFFF29F7 , 32'h07FD2920 , 32'hF775F590 , 32'hD77A7680 , 32'h0001F1B6 , 32'h017DBE88 , 32'hFFFB5625 , 32'hFE50ADAC , 32'h00014850 , 32'hEF24BB60 , 32'h00009368 , 32'h16116F20 , 32'h11246DC0 , 32'h24850300 , 32'h3C0E9C40 , 32'hFFFCA674 , 32'h02BFC4C4 , 32'hFFCC3D0A , 32'hFFFF363E , 32'h0F7053A0 , 32'h0001AC38 , 32'h05C87158 , 32'h1F2B1560 , 32'hFA73C550 , 32'h0000BCAF , 32'hFFFA06E0 , 32'h1174B3A0 , 32'hFFFC7870 , 32'h0D6BABB0 , 32'h0002F86A , 32'h00CE8111 , 32'hFFFEBB06 , 32'hF6A423E0 , 32'hFFFC422A , 32'h00011889 , 32'hFFFD785A , 32'h02E6BDAC , 32'hF59477D0 , 32'h00039CAD , 32'hFFFF3944 , 32'h000035CF , 32'hFFF6E73F , 32'hF4F28B20 , 32'h0DBAFE90 , 32'hED27B5A0 , 32'hE66CF1E0 , 32'hF51C6FC0 , 32'h0002F44C , 32'h00012EB8 , 32'h0000910F , 32'hF9B68240 , 32'hFFFCE9CD , 32'hFFFB49B9 , 32'hF8066368 , 32'hF58B63D0 , 32'hFFFF5B66 , 32'hC1B0E7C0 , 32'hFC5500AC , 32'h03C56998 , 32'hF6AC76F0 , 32'hFFFCF319 , 32'hF7E78950 , 32'hF85FDA38 , 32'h03059E44 , 32'h00048A6D , 32'h1E74E9A0 , 32'hB2182C80 , 32'hFE351668}
};

logic signed [31:0] VT_2 [100][100] ='{
{32'h02D91254 , 32'hFBD64850 , 32'h03C8D3DC , 32'h000043AE , 32'hFFFFEA5F , 32'hFD4596B0 , 32'hEEF7B0E0 , 32'hFB97C048 , 32'h0000CC98 , 32'hF46723D0 , 32'hFF183290 , 32'hF115F460 , 32'hE6630380 , 32'h077E4F88 , 32'h0F632A30 , 32'hF5C73340 , 32'hE7D35600 , 32'hF6284A00 , 32'h03CD6CA8 , 32'h0000C932 , 32'hF742A430 , 32'hF0A0E190 , 32'hF9B91038 , 32'h00022A9D , 32'hE3D208E0 , 32'hF2730200 , 32'hF629F6D0 , 32'h012A1F94 , 32'h04AEC388 , 32'h163D5740 , 32'hE8FF6320 , 32'h0B24B100 , 32'hFD87F694 , 32'hE064CEA0 , 32'hFFFFD6A3 , 32'h025FD710 , 32'hFB625E68 , 32'h091937F0 , 32'h00F1B9CB , 32'h0012C9DF , 32'hEEB4AD20 , 32'h00C44AAA , 32'hFE67F504 , 32'hFE352E28 , 32'h043C1628 , 32'hFF35A341 , 32'h0A988530 , 32'h01AEA9A8 , 32'hE5E02FE0 , 32'h0D501650 , 32'hFE806320 , 32'hE8399400 , 32'h0AB87140 , 32'h09656500 , 32'hF7F90ED0 , 32'h0DFFE620 , 32'h0FFECA50 , 32'h1312FD80 , 32'h0A81C700 , 32'h1712A960 , 32'h057B4CD8 , 32'h09315470 , 32'hE83BD900 , 32'h0B247190 , 32'hFBA211A8 , 32'h1B0E4DA0 , 32'hFFFECE3D , 32'hF3D0E960 , 32'h02174A78 , 32'hFF7C969A , 32'hFE9FD280 , 32'hFF319010 , 32'hFDA1EDA0 , 32'hFA2D53F0 , 32'hFBD61018 , 32'hFA1D1400 , 32'hFC269CB4 , 32'h0B24D450 , 32'h1CC00A20 , 32'hFBE433D8 , 32'h14C675A0 , 32'h1916EF80 , 32'h067437D8 , 32'hFFFF8538 , 32'hF5963B20 , 32'hFFAE1455 , 32'hEE27EB00 , 32'hE7D23300 , 32'h0C5935D0 , 32'h0000A828 , 32'hEC22FEE0 , 32'hFADAAD50 , 32'h00095CE5 , 32'hE94EED40 , 32'hFFFFE19B , 32'h11E4B5C0 , 32'h0B6EF620 , 32'h0A0AD9F0 , 32'hF976F888 , 32'hEEB8DCE0} , 
{32'h0DA2FC50 , 32'hEF1641A0 , 32'h01346F88 , 32'hFFFFA1D6 , 32'hFFFFC2BD , 32'h176B31A0 , 32'h016E6AB0 , 32'hF6807B10 , 32'h00006F4B , 32'hD2A325C0 , 32'h1073D220 , 32'h03943834 , 32'hE81F5080 , 32'hF8BB0698 , 32'h0E944B50 , 32'h14700860 , 32'hF3A14EB0 , 32'h023B5A1C , 32'h06B680C0 , 32'hFFFFEAC6 , 32'hFB5C4F48 , 32'h0C3A1D10 , 32'hFC0855D0 , 32'hFFFF5B4D , 32'h07791C68 , 32'hF25BAC80 , 32'h05C87358 , 32'h02D8A110 , 32'h00E441F8 , 32'h0DEBD6A0 , 32'hFA2AE040 , 32'hEDE0E080 , 32'hFC291CA4 , 32'h086CAFA0 , 32'h00009471 , 32'hFFC9C394 , 32'h05AA2148 , 32'hEA3D91E0 , 32'h02DDAA40 , 32'hF227ACF0 , 32'hEF2FF000 , 32'h004E181A , 32'hFCD9E684 , 32'h0DDC82D0 , 32'h19302960 , 32'hFC44F48C , 32'h065328A0 , 32'hF7482C90 , 32'hFCF10610 , 32'hFB51BAF8 , 32'h0710E348 , 32'h0D3A6490 , 32'hE6A801A0 , 32'h05CEF358 , 32'h14201BA0 , 32'h03832D60 , 32'h26C27A80 , 32'hF42193F0 , 32'hEE57DFC0 , 32'h1239A3E0 , 32'hF60F99E0 , 32'h07ED8F18 , 32'h08F8CA70 , 32'h0DE6D110 , 32'h03AC4A2C , 32'hF1AD6840 , 32'h00012485 , 32'hFC42509C , 32'hF9E24778 , 32'hFB039290 , 32'hFE308E30 , 32'hEF330300 , 32'hFC9DD048 , 32'h0A470360 , 32'hEEF70B60 , 32'h09CEED70 , 32'hF28FBEA0 , 32'hEC2EF4A0 , 32'h101189E0 , 32'hF521A110 , 32'h053DB818 , 32'hFEA8EB0C , 32'hFECB7A7C , 32'h00006BA5 , 32'hFDDC574C , 32'h0A086A60 , 32'h09CC85B0 , 32'h108BA840 , 32'h0B815FC0 , 32'hFFFEAEFB , 32'h0B0A5DB0 , 32'hFE5B3BE0 , 32'hFBAE4190 , 32'h16CC10E0 , 32'h000084F4 , 32'h06ED5B90 , 32'hFD38EE48 , 32'hE6CB0980 , 32'h17534760 , 32'hFAB1E138} , 
{32'h0A017320 , 32'h12EDD720 , 32'h0267FD74 , 32'hFFFFCF6F , 32'h00007A37 , 32'hEC9C26A0 , 32'hF1799660 , 32'hE0A834A0 , 32'hFFFFC444 , 32'h00998966 , 32'h02A3E3F4 , 32'hF83D6A28 , 32'h12B4ADE0 , 32'hF1CC1280 , 32'h0C504770 , 32'hFC92D1AC , 32'hF95EE888 , 32'hFA58CA90 , 32'h05B68488 , 32'hFFFF853B , 32'h047C3D10 , 32'h0CB510E0 , 32'h166D8180 , 32'h0001F92B , 32'h0FB29260 , 32'hF484CB00 , 32'hFC979578 , 32'hFA47B510 , 32'hFC3CBF1C , 32'hFFFFD540 , 32'hF45E8F50 , 32'h16BF6A60 , 32'h03150E44 , 32'h0E9F88D0 , 32'h000153C9 , 32'h0C554230 , 32'h02FE233C , 32'h11815EA0 , 32'h09B23EB0 , 32'h09F8CC30 , 32'h00CE53FE , 32'hFFED52D1 , 32'hF595A610 , 32'h21B24E40 , 32'hECC51080 , 32'hFAE5C020 , 32'h11AC6220 , 32'hFA3AF1B8 , 32'hEB3451E0 , 32'h02F155A8 , 32'h150AFFA0 , 32'h0C40F2B0 , 32'hFF6685F0 , 32'hEF7A5FA0 , 32'h01EE9384 , 32'hF5DE69B0 , 32'hF9903D60 , 32'hEF546780 , 32'hF54BD250 , 32'hF576D8F0 , 32'h04EA9658 , 32'h07180F58 , 32'h0E955760 , 32'h03ED8D2C , 32'h0C94D6D0 , 32'h0E237D90 , 32'h00019BBF , 32'hF7EEBEC0 , 32'hFF07492A , 32'hF47B46F0 , 32'h0937EFE0 , 32'hF1495810 , 32'h0168A908 , 32'h0FCBCC50 , 32'h00C0EB6B , 32'h0148BF7C , 32'h0675ADD8 , 32'hEE283100 , 32'h172E7440 , 32'h1F4ECBC0 , 32'hF1A505F0 , 32'h12D76040 , 32'hEFF45D20 , 32'hFFFF47D6 , 32'hF5A5E190 , 32'hFA637558 , 32'h09426230 , 32'h1A0E8960 , 32'h112F39A0 , 32'hFFFF3C77 , 32'h07BCB800 , 32'hFF24FEBE , 32'hEC507840 , 32'hF0486440 , 32'hFFFFA065 , 32'h0814F7A0 , 32'h1900DD80 , 32'h0C60B800 , 32'hEFD870A0 , 32'h038131E0} , 
{32'hE9BD0820 , 32'hF5A52BC0 , 32'h03BF658C , 32'h0000D32B , 32'h000058B9 , 32'hF4034F40 , 32'hFBA69028 , 32'h0B933270 , 32'h00006913 , 32'hFED11738 , 32'hF2380740 , 32'hF8DA4E48 , 32'hF2EE4230 , 32'h0B87D5A0 , 32'hEE42A7E0 , 32'h0AFCBE50 , 32'hF3B35830 , 32'hE7491020 , 32'hEC929260 , 32'hFFFE98CB , 32'hFC7D57A4 , 32'h13126EA0 , 32'h0169E2A4 , 32'hFFFFAD58 , 32'hED4A9700 , 32'hFEC47620 , 32'hFF955C55 , 32'hFE60E28C , 32'h0CEA2250 , 32'h030DC79C , 32'hF18305A0 , 32'h02B5A0E4 , 32'h00D1BA11 , 32'h19C50BC0 , 32'hFFFFCEB2 , 32'hEDE35280 , 32'hFAEFB1C0 , 32'h08BC4660 , 32'h01F46F14 , 32'h0645B0E0 , 32'h14360E20 , 32'hFFA05CF4 , 32'hFDBE0378 , 32'h22B9F800 , 32'hE363BF40 , 32'h017E994C , 32'hE1AC3F00 , 32'hEB0F10C0 , 32'h0421F2A8 , 32'h062DC410 , 32'h1194F0E0 , 32'h0CDC18E0 , 32'hED7C0140 , 32'h00059C6C , 32'h0F8C3270 , 32'h06665608 , 32'hF8A944F0 , 32'hE68BBA60 , 32'h0EC0A7D0 , 32'h03198B48 , 32'hFC8A92C4 , 32'h0F531F90 , 32'hF9B1E428 , 32'hFBCC03D0 , 32'hEC13EC20 , 32'h07647CE8 , 32'h0000E554 , 32'hEE642E60 , 32'hFF90F63B , 32'hEDDB3240 , 32'h0B09FA40 , 32'hF43C28B0 , 32'h13368A60 , 32'hFAF56890 , 32'hFDEDC2CC , 32'h1230E2A0 , 32'h170CD5E0 , 32'h00C94219 , 32'h0683FD68 , 32'hFA6C2410 , 32'h0C958410 , 32'hECEDCA60 , 32'h131287A0 , 32'h00000CCF , 32'h08E06C20 , 32'h16F16180 , 32'hFA807898 , 32'hEE756040 , 32'h03FB46BC , 32'hFFFF9275 , 32'hFBBEDCF0 , 32'h01EDD794 , 32'h007CA165 , 32'hFF22863F , 32'hFFFF9874 , 32'h002721F5 , 32'hE9F13500 , 32'h02D96CC8 , 32'h02B2CD94 , 32'hF59D53B0} , 
{32'h19A2E540 , 32'hEFC818E0 , 32'h0E567420 , 32'h0000FD8A , 32'hFFFF5074 , 32'hFE462D70 , 32'hF70654E0 , 32'hF5CFF170 , 32'h0000E549 , 32'hFD0F6120 , 32'h04438D80 , 32'h0C38A830 , 32'hF6DA8A70 , 32'hF437B5C0 , 32'h03434DAC , 32'hF9D073C0 , 32'hF4C58150 , 32'hF4928DF0 , 32'h042781B8 , 32'h00001420 , 32'hFBB37A28 , 32'hE6EA7000 , 32'h00A647D8 , 32'hFFFDE2BF , 32'h0ED5DD70 , 32'h06D334E8 , 32'hFD6AD524 , 32'hFA829638 , 32'h013E6718 , 32'h1DC1FAC0 , 32'hF2A11FA0 , 32'h0E62C650 , 32'hFA28EAC0 , 32'hF2BBE460 , 32'h000040DE , 32'h073B9C40 , 32'h0508A478 , 32'hFD8905D0 , 32'hFFD574B4 , 32'h0E7DF780 , 32'hFDCB0C94 , 32'h01116800 , 32'h0008B631 , 32'hF90F1600 , 32'hE971D1E0 , 32'h07ABD0D0 , 32'h12953880 , 32'hF9EC9BF8 , 32'h0524FD30 , 32'hF4933D30 , 32'h093682A0 , 32'h12114780 , 32'hFE4C4C38 , 32'h0BBE4790 , 32'h0D7F1630 , 32'hF4C41B50 , 32'hF6DBCCF0 , 32'hFA482780 , 32'hF920BB70 , 32'hF2BBB5A0 , 32'hF06F2870 , 32'h112D0380 , 32'hFB5AD3F8 , 32'h00970615 , 32'h1079FC80 , 32'hF1E5CC70 , 32'hFFFFFF70 , 32'h14D95B40 , 32'hFC4833A8 , 32'h1738BD20 , 32'h053968D0 , 32'h06078E90 , 32'h155D68A0 , 32'hF585B1A0 , 32'h163AB9C0 , 32'h002DD5BC , 32'hFE105380 , 32'h0F7DEE60 , 32'hF0D83760 , 32'hFBFF5630 , 32'hFBC1D750 , 32'hEFE4B780 , 32'hF513F3B0 , 32'h0000ABA5 , 32'h170BF5E0 , 32'h10039FA0 , 32'h1FA61740 , 32'hFECC6054 , 32'hEA53DC60 , 32'hFFFF70A3 , 32'hF3D405D0 , 32'h019F2E54 , 32'hFE8B1FEC , 32'hE2CF6A20 , 32'hFFFFFDE5 , 32'h1967DCC0 , 32'hE8DD9200 , 32'hF462A030 , 32'hFCD44CE0 , 32'hE1E27FE0} , 
{32'hFE765994 , 32'hF0C29C10 , 32'h145166A0 , 32'hFFFEFAF6 , 32'hFFFF7232 , 32'hFF5784BE , 32'hF3077E20 , 32'hFDB8D5A0 , 32'h0000D0F7 , 32'h078F0B60 , 32'h0D7DE120 , 32'h195BF300 , 32'hF854D6B8 , 32'hFBF359C8 , 32'hEEB1B160 , 32'hECD7CCC0 , 32'h03A1229C , 32'hF8788790 , 32'hDEF2A5C0 , 32'hFFFFA810 , 32'h157EE400 , 32'h063A9BD8 , 32'hFA8C74A8 , 32'hFFFFCBFE , 32'hEDE8CBA0 , 32'hFBC92AE8 , 32'hEE34A9A0 , 32'hFBEF7330 , 32'hF1436410 , 32'h1FB52280 , 32'h17952AC0 , 32'hF4039F40 , 32'hF729AFC0 , 32'h0ADE47F0 , 32'hFFFFA8B9 , 32'hF50A6800 , 32'h06966210 , 32'hEE45F5E0 , 32'hF5B437E0 , 32'hF885AC60 , 32'h118175C0 , 32'h01002B14 , 32'hFF2571A6 , 32'hF2157AC0 , 32'hFC71BB50 , 32'h0FB5D090 , 32'hEA0D8940 , 32'hF84CA958 , 32'h14EC0240 , 32'h175D2FC0 , 32'h14913D20 , 32'h0A9CF1E0 , 32'hF6AABEE0 , 32'hF3BC67D0 , 32'hEA850720 , 32'hF51519C0 , 32'h07E7C1D0 , 32'h0C6B0F10 , 32'hFB53F370 , 32'h108DD6A0 , 32'hFA33E9E8 , 32'h09DE1F40 , 32'h0D03E1D0 , 32'h08CE0CC0 , 32'h05C569D8 , 32'h0DC4A280 , 32'hFFFFFC41 , 32'hFE0FF190 , 32'h02D4573C , 32'h073B9AB8 , 32'hF858AD68 , 32'h0465C198 , 32'hFDA19B28 , 32'h04FD5880 , 32'hFABD8238 , 32'hF00FB370 , 32'h05C82030 , 32'hEC0177A0 , 32'h021C8818 , 32'h0389223C , 32'hF82C2068 , 32'h18127180 , 32'h040068C0 , 32'h00009A79 , 32'h0C6FC040 , 32'hE63110A0 , 32'hFC88BEDC , 32'h1EC9E5A0 , 32'hFF5BAECA , 32'h0000E58E , 32'hE9EDAEC0 , 32'h00C190E8 , 32'h09D12FC0 , 32'hF4DA8BB0 , 32'h000318A4 , 32'h00658862 , 32'h0AB2E090 , 32'hFFAF1D8C , 32'hFBEDBF70 , 32'hF42B2E50} , 
{32'h095CFE40 , 32'hF5B1BA70 , 32'hF6A6ADA0 , 32'h0000123A , 32'h00006C88 , 32'hED9AAE40 , 32'h04267FC0 , 32'hE1870FA0 , 32'hFFFFEDE3 , 32'h0DB2D480 , 32'h0B0C0360 , 32'hF93FF990 , 32'h116F1FA0 , 32'h0992B4D0 , 32'hF7CA54C0 , 32'hF374F1B0 , 32'hEC6CC080 , 32'h024EEE5C , 32'h08C3B990 , 32'hFFFEEE46 , 32'h21B00AC0 , 32'h09E53D90 , 32'hE8F74560 , 32'h0000964F , 32'hFE8A794C , 32'h14711320 , 32'h0A8795F0 , 32'h12EFE4E0 , 32'hF1F41B10 , 32'h0B4F5760 , 32'h199D2B80 , 32'h0DAE42D0 , 32'hFAD3AEB8 , 32'h00FF3682 , 32'h000048F2 , 32'h0751E7D0 , 32'hF6E27910 , 32'hE702C260 , 32'hF8B57958 , 32'h0236F2D4 , 32'hFBD1AF10 , 32'h000E6362 , 32'h037E79D8 , 32'h012795B8 , 32'hECB72920 , 32'hD8F8A5C0 , 32'h06BB3E80 , 32'h17E4A3A0 , 32'hF16ED470 , 32'hFD59485C , 32'h07B9F4D0 , 32'hEED257A0 , 32'hF219DC00 , 32'hFA9C59C8 , 32'h05F34678 , 32'h0B62DAB0 , 32'hFEDAA09C , 32'hF184E330 , 32'h04A75118 , 32'h0B10C3B0 , 32'hEB9D66E0 , 32'h062D6FA8 , 32'hF4AC1670 , 32'hF7DE0B20 , 32'hFB4BD180 , 32'hF42AB170 , 32'h00002A77 , 32'h17A25320 , 32'hF6340800 , 32'hEF424700 , 32'hF956A130 , 32'hFB3BA018 , 32'h0675B498 , 32'h02D88614 , 32'hF6B47FC0 , 32'h0B0C29A0 , 32'h092C75C0 , 32'h07AA9D90 , 32'hFF6716F8 , 32'h0D51DC10 , 32'h17490BE0 , 32'h12CD17A0 , 32'h070176D8 , 32'hFFFF7B8E , 32'h0D86AE50 , 32'hF6B96AA0 , 32'hF4EB3720 , 32'hF4B4CF00 , 32'hF98046D8 , 32'h0001AFCF , 32'h0FD80020 , 32'h01DD74BC , 32'h1392A4E0 , 32'h0F8C79B0 , 32'hFFFE8145 , 32'h07F42ED8 , 32'hFDFEDB64 , 32'hF075BBC0 , 32'hFBA14BA0 , 32'hFCA841C8} , 
{32'hFAF09CA8 , 32'hFE18B02C , 32'h0DC0AFB0 , 32'h00004B42 , 32'h0000AFA7 , 32'hFCD3D4CC , 32'hFD52974C , 32'hF6D4E670 , 32'h000038D3 , 32'hEF9F05E0 , 32'hF28F8D20 , 32'hF1B0BCA0 , 32'hEFCF84A0 , 32'hF37D8D60 , 32'h12E9D500 , 32'hFCC33688 , 32'hF8DFE648 , 32'h0223E114 , 32'hF581ECA0 , 32'hFFFFC581 , 32'h04AC2568 , 32'h11F42D20 , 32'hF0717C00 , 32'h0000F97D , 32'h0097258D , 32'h08E22630 , 32'h05EBE660 , 32'hF3447310 , 32'hECB34F40 , 32'hF8F84E48 , 32'h0B4DA4B0 , 32'hEF9C5000 , 32'h1FB7D080 , 32'hFB227A90 , 32'h00015BE1 , 32'h07B54068 , 32'hFB054978 , 32'h03B06E6C , 32'hF4249E20 , 32'hDD4E3600 , 32'h0553B750 , 32'hFFCB4FA0 , 32'hFEDE9A3C , 32'h0EC370C0 , 32'hFB661FE0 , 32'h07213C50 , 32'hF8328E80 , 32'h0D0D4700 , 32'h018D44D8 , 32'h0AD05860 , 32'h0DA0F320 , 32'h0A078910 , 32'h0A3A1990 , 32'hFDAB5BD8 , 32'hECB10AE0 , 32'h0A9CECD0 , 32'hDE8384C0 , 32'h041D9000 , 32'h10118DE0 , 32'h04E8C6F8 , 32'hF9590AD8 , 32'hF5FE73C0 , 32'h0EE8FB50 , 32'hF8854D70 , 32'hF01BA010 , 32'hE5103020 , 32'h000047F3 , 32'hF705A450 , 32'hF4AB92A0 , 32'h0C3D23F0 , 32'h0DD199B0 , 32'h07D8B208 , 32'hEF0A3100 , 32'h001A4A06 , 32'h0C3B9F40 , 32'hF2454E00 , 32'h05121AF8 , 32'h03CF7038 , 32'hF869E130 , 32'h0258EA24 , 32'h1388E940 , 32'hFCB60430 , 32'hEF655800 , 32'h0000B083 , 32'hED28B4E0 , 32'h08102B40 , 32'h03862CE8 , 32'hF2DC1240 , 32'hFB90CAC0 , 32'h00022CB9 , 32'hFBBCD6C0 , 32'h060F6548 , 32'hE630AD00 , 32'hF58A4250 , 32'h000057DF , 32'h1C2295E0 , 32'h102EC580 , 32'hD75134C0 , 32'hFD98483C , 32'h046F9968} , 
{32'h0B8AE530 , 32'h185F14A0 , 32'hF97063F0 , 32'h00019BA7 , 32'hFFFF9F5A , 32'hFC18660C , 32'hFA6118A8 , 32'h1DBCB560 , 32'hFFFE8823 , 32'hEC82C260 , 32'h018F3278 , 32'hF082A810 , 32'hDF377380 , 32'h077900E8 , 32'hF7494B10 , 32'h073F6968 , 32'hFC2EA730 , 32'hDD93BD80 , 32'h0EE436B0 , 32'hFFFF3280 , 32'hFA871468 , 32'hF9226988 , 32'h0376FB10 , 32'h0001136D , 32'h19ECE620 , 32'h0CFEC080 , 32'h039B2950 , 32'h09B5B220 , 32'hF1E08640 , 32'hE8102640 , 32'hF4079210 , 32'h1163F660 , 32'hD9219540 , 32'hF9F9B020 , 32'h00010426 , 32'hF9EBD318 , 32'hFDD5FDEC , 32'hFB0A0670 , 32'h04813F88 , 32'hFCDCB040 , 32'h0B014F50 , 32'hFF58C991 , 32'hF989C090 , 32'h038EFE40 , 32'hFDD792B4 , 32'h09D9B220 , 32'hF40E4EB0 , 32'h099CBC20 , 32'h09DCBA10 , 32'h0B8D57C0 , 32'h11787780 , 32'h08159C60 , 32'hF6F1DD10 , 32'hF4EE38D0 , 32'hF83A1EC8 , 32'h0B297DC0 , 32'hFDCB16E4 , 32'h052F5F68 , 32'hF8C0E880 , 32'hF6CF3F60 , 32'hEFE6D280 , 32'h02C9DD80 , 32'hF0C4A640 , 32'hFA2040A0 , 32'h1069F0E0 , 32'hF80CE4A8 , 32'h00000158 , 32'hEA3A3EC0 , 32'h048B7908 , 32'hFEF86290 , 32'hFE3026FC , 32'h040379D0 , 32'h0CC0BA90 , 32'hFE2B104C , 32'hF49A2920 , 32'hF62BC7A0 , 32'hF928A680 , 32'h193EBEC0 , 32'hEC7A6C40 , 32'h11D8DC60 , 32'h0346B8F8 , 32'h1625DEE0 , 32'h09AA0C90 , 32'h0000FA5A , 32'h06EA5DF0 , 32'hF766A170 , 32'h045E8050 , 32'h07A2FDC0 , 32'hF093E7D0 , 32'hFFFE96AD , 32'hFFA9F6FF , 32'hF6C6BF00 , 32'h0BA83E40 , 32'h0C44E360 , 32'hFFFF1474 , 32'h013F58CC , 32'h2334EE40 , 32'hF52AA320 , 32'h07DB3230 , 32'h09A8AEE0} , 
{32'hF910CE48 , 32'hF901F120 , 32'hE6399460 , 32'hFFFE7555 , 32'hFFFEF61D , 32'h14792600 , 32'h0831DFC0 , 32'hDE957780 , 32'hFFFE6023 , 32'hE4B41AA0 , 32'hF12C4E40 , 32'hF853EB20 , 32'hE7E9C140 , 32'h008E1B1F , 32'hF3A010E0 , 32'hF31F7FF0 , 32'h258507C0 , 32'h01CB7C2C , 32'hFABF5B50 , 32'h0001E2D4 , 32'hF365B0A0 , 32'hF5BE34E0 , 32'h075F57A8 , 32'h00005985 , 32'h03D2D208 , 32'hFA665868 , 32'h03BC69AC , 32'hF911C8D8 , 32'h03D1CE20 , 32'hF3DF59A0 , 32'hF473BC90 , 32'h09441570 , 32'hEC2A2D40 , 32'h016EFB30 , 32'hFFFEF2A0 , 32'hF2DB5D10 , 32'h05285318 , 32'h0230B5BC , 32'hEEFDC2E0 , 32'hF0E10F00 , 32'h00E4BF24 , 32'h0011F376 , 32'h03E154B0 , 32'h0770F8E0 , 32'hF65C7350 , 32'hEE93A360 , 32'hF9D1DA60 , 32'hFAF30B68 , 32'h05FBB528 , 32'hE1ED0B00 , 32'h0C3BC2B0 , 32'hEA06D340 , 32'hF31C14D0 , 32'h0470CB90 , 32'h052A2250 , 32'hF59CE020 , 32'hF4BED3D0 , 32'hF7B6E890 , 32'hF4198300 , 32'hFA79C040 , 32'h0484D0F0 , 32'hFB9D2168 , 32'h00D528DE , 32'h057C4048 , 32'hED03FDA0 , 32'hEF7172C0 , 32'h00017EC4 , 32'h0E1B6190 , 32'h010EE900 , 32'h0B578960 , 32'h081D6780 , 32'hF61C59A0 , 32'h02094050 , 32'h01D89468 , 32'hFAD0C920 , 32'hFAEE8320 , 32'h03487CC4 , 32'hE90C6B00 , 32'h0070CDF5 , 32'hFAA895F8 , 32'hEAE2B0A0 , 32'h07492678 , 32'hFC76A4F0 , 32'hFFFE9C14 , 32'h0338C158 , 32'hE12B11E0 , 32'hE8DBCAE0 , 32'hE88657A0 , 32'hFCFDBBB0 , 32'hFFFF8A3B , 32'hF579D800 , 32'hFCCBA3B0 , 32'h10554CC0 , 32'hE5D1DB00 , 32'h0000F0A5 , 32'hFB1B8350 , 32'h08719DF0 , 32'hF58A1060 , 32'hEA1C03A0 , 32'hF86A39B8} , 
{32'h247B0880 , 32'hF589F720 , 32'hFEC1E96C , 32'h00003946 , 32'hFFFF1193 , 32'h07CB5F10 , 32'hFDDDFC10 , 32'h11F79900 , 32'h0000207E , 32'h07B2E890 , 32'hFF41EC8A , 32'h0AFEA200 , 32'hF481EEC0 , 32'h05C0FF80 , 32'h0362D0CC , 32'h03B3DFA4 , 32'hFFE481F7 , 32'hF9469FF0 , 32'hF7887FD0 , 32'hFFFFF9F7 , 32'h21DE9F80 , 32'h009467E7 , 32'h11530480 , 32'h0000D2B3 , 32'hF3B767C0 , 32'hFD77CB50 , 32'hF7F579B0 , 32'hF67E8260 , 32'h15480400 , 32'hEFE8E1E0 , 32'h27077900 , 32'hDD226000 , 32'hE4D47120 , 32'hDC3CBB00 , 32'h00011A38 , 32'h0AF02D80 , 32'h01B947DC , 32'h04AC3168 , 32'h00DF0EFC , 32'hF8A48DC0 , 32'hF563CC60 , 32'h00005965 , 32'hFB60C258 , 32'h0F3F9860 , 32'h0243DC90 , 32'h0621C670 , 32'h100B6060 , 32'h004AE681 , 32'h011F52AC , 32'hFB9328E0 , 32'h0C5DF680 , 32'hF8EC20D0 , 32'hF86F1348 , 32'hEEB6B260 , 32'h0DB3BE20 , 32'h042A5AD8 , 32'hF3FBED80 , 32'hE4DAAFE0 , 32'hF558F490 , 32'h00F6BC60 , 32'h0097C304 , 32'hF0A40DC0 , 32'h038F76A4 , 32'hFC78AFBC , 32'h00004B2B , 32'h002C0867 , 32'hFFFCE50B , 32'h04822A08 , 32'h00CFD4B6 , 32'hFD232D54 , 32'h07BB2640 , 32'hF27901B0 , 32'h02917C2C , 32'h04599780 , 32'h034452F8 , 32'hFE770880 , 32'h002D88D3 , 32'hFEB90AE4 , 32'h061491D8 , 32'h071B2E90 , 32'h10CF9760 , 32'hE99E50A0 , 32'h1339D8E0 , 32'hFFFD509F , 32'hFCA5EE9C , 32'hF0F8BD00 , 32'h0F161860 , 32'hEA7189A0 , 32'h00471488 , 32'h00021A34 , 32'hF6140660 , 32'h025BDF40 , 32'hF5006F70 , 32'hEF810AE0 , 32'hFFFE7844 , 32'h020E8C50 , 32'h0B1232C0 , 32'h1D5632E0 , 32'h06A90BE8 , 32'h0D939BB0} , 
{32'h156E8F80 , 32'hF754F150 , 32'hF7856BE0 , 32'hFFFE46A0 , 32'h000361B2 , 32'hF6492140 , 32'h07814EF8 , 32'h083FBE70 , 32'h0001B5D9 , 32'h034AE21C , 32'hF44693F0 , 32'hFC6900F4 , 32'h08925FB0 , 32'h09C31CE0 , 32'hF63BCA00 , 32'hF7C33100 , 32'h0A89EB00 , 32'h0AD01C70 , 32'hE209F8A0 , 32'h0001AF82 , 32'hE7983A60 , 32'hFC937C38 , 32'h07EA64C0 , 32'hFFFE1E25 , 32'h136E54C0 , 32'h08DDCCB0 , 32'h0312F214 , 32'hFF0666D4 , 32'hEE66C920 , 32'h05BFF728 , 32'hDE1852C0 , 32'hFCC7BACC , 32'h137D15A0 , 32'hD5EDEE80 , 32'hFFFF14DD , 32'h14B7CE60 , 32'hFCFCBE24 , 32'hF3007660 , 32'hF96C9DE8 , 32'hF9FEC0F0 , 32'h0B54AF90 , 32'hFF170685 , 32'h00652F08 , 32'h0CBFC840 , 32'hFFBC72FE , 32'hF6A6B750 , 32'h1C423F80 , 32'h012354F4 , 32'h1557E860 , 32'h118B4020 , 32'h08AAE130 , 32'h031A357C , 32'hE8C79A00 , 32'hFB296A38 , 32'hEF51C800 , 32'hF9849348 , 32'hEAEC41E0 , 32'h00CAFFDC , 32'h0F959F20 , 32'hFC3EA23C , 32'h0053E999 , 32'h0A098600 , 32'h01A52F38 , 32'h0A03BCF0 , 32'h09B2C110 , 32'h0C8605F0 , 32'hFFFC5053 , 32'h085E56B0 , 32'h03708674 , 32'h00086A1C , 32'h0123C754 , 32'h07EECAA0 , 32'h0BB4CC50 , 32'hFE07C0A0 , 32'hF2257620 , 32'hFF9557BA , 32'h11A5BDC0 , 32'hEC5CE480 , 32'h1707CE20 , 32'hDFB72900 , 32'h08D77B80 , 32'hF4B248C0 , 32'h0C3E5AA0 , 32'h00023F56 , 32'hFCE8CD54 , 32'hFEA86AE0 , 32'h041E0318 , 32'h02FF82D8 , 32'h01B8A4E4 , 32'hFFFD0D22 , 32'h0D769FD0 , 32'h02485B18 , 32'h0E15CA90 , 32'h1D13C4C0 , 32'hFFFE9966 , 32'hFBCBC858 , 32'h0F6AFE70 , 32'h05923D80 , 32'h00C82DDB , 32'hFF266FB9} , 
{32'hF004FA70 , 32'hF300FFB0 , 32'h061BA7C8 , 32'h0002EBC5 , 32'hFFFF8282 , 32'h02B29590 , 32'hFD0DAAD0 , 32'hEDFA2FA0 , 32'h0002C59E , 32'hFC69CA50 , 32'hEF0488A0 , 32'h09B20230 , 32'h0A1AA390 , 32'hF327B1E0 , 32'h023200A0 , 32'hF1243020 , 32'hEFC62E00 , 32'h0690AD90 , 32'h0BA815E0 , 32'h00000D84 , 32'hF4147EF0 , 32'hF7279010 , 32'h0B4F4D70 , 32'hFFFEF504 , 32'h0B3361D0 , 32'hFAC65AE8 , 32'hF6B21100 , 32'h0924DF80 , 32'hF947D870 , 32'hF8F2FDD0 , 32'h07778CF0 , 32'hE56A1140 , 32'hEB939060 , 32'hF6144470 , 32'h00008612 , 32'h124993E0 , 32'h1171EA40 , 32'h3B748D80 , 32'h12B60BC0 , 32'hFA27CE68 , 32'h1DA82400 , 32'hFF5C29B5 , 32'hFC9B9738 , 32'hFAA1F2C0 , 32'h109A0340 , 32'hF4B17740 , 32'hEFEC2820 , 32'h10425800 , 32'hEA323820 , 32'h155F7080 , 32'h050E6BD8 , 32'h0788F968 , 32'hDA637100 , 32'hF84B7D90 , 32'hF5202250 , 32'h002553DF , 32'hFEB7BF5C , 32'h080E4D30 , 32'hF8D57880 , 32'h06851EA8 , 32'hECE458A0 , 32'h03E5ECBC , 32'h0BA5B380 , 32'hFEBA8728 , 32'hFC3F0F4C , 32'h08E2EC50 , 32'hFFFDA323 , 32'h0653FB00 , 32'hF6263820 , 32'hFADD1230 , 32'hEF664AE0 , 32'hF5163BB0 , 32'h09892530 , 32'hFB7D34F0 , 32'hFE6A9068 , 32'hFE52A540 , 32'hFC41B2AC , 32'h054AF3C0 , 32'hEFC88C00 , 32'hF8302EA0 , 32'hF5EBA7E0 , 32'h05526040 , 32'hF09E9E60 , 32'hFFFF30ED , 32'hFBA2AC88 , 32'h024FA454 , 32'h05D8E458 , 32'hE882E760 , 32'h00D60337 , 32'hFFFE0510 , 32'hFEE66694 , 32'hFA6DF9F8 , 32'h0AEC3770 , 32'h0E161550 , 32'h00003D24 , 32'hFD09A27C , 32'hF23C7DF0 , 32'h03E8ED74 , 32'h03129864 , 32'hF60B77D0} , 
{32'h101A7480 , 32'hF2DDF6D0 , 32'hEF734200 , 32'hFFFF8455 , 32'hFFFE905E , 32'hFA161328 , 32'hF0B58F30 , 32'hE7121980 , 32'h0000DCBF , 32'h0E786F10 , 32'h084437C0 , 32'h0FBF7EE0 , 32'h170313A0 , 32'h01487B4C , 32'h003AEB68 , 32'h05098A80 , 32'h0D51D6F0 , 32'hFB16F218 , 32'hF9B73418 , 32'hFFFFD709 , 32'h0E5F4460 , 32'h063E84C0 , 32'h010E1D18 , 32'h000243F4 , 32'h02B6DBC0 , 32'h10CEC660 , 32'h04E4D9D8 , 32'hF9C57E80 , 32'hF41BF230 , 32'hF88D4A50 , 32'hDF073540 , 32'hFADA2CA0 , 32'hE48FA100 , 32'h1A6BA6A0 , 32'h00022E0C , 32'hF1EC47C0 , 32'h0696A770 , 32'h008D53CC , 32'hFDAA1AB4 , 32'hF1836470 , 32'hE7DC5E40 , 32'hFEDA0660 , 32'h04077928 , 32'hF101D0D0 , 32'h067F4C40 , 32'h09E8EF10 , 32'h00133F04 , 32'hED7E9A60 , 32'hE795B460 , 32'h07D5F1E0 , 32'h11E761E0 , 32'h251CE640 , 32'h15EC2240 , 32'h0EBEBDA0 , 32'h068D7120 , 32'h014FAA38 , 32'hF5AF7F40 , 32'hFEAD7D80 , 32'h031D4C1C , 32'h0F2B61F0 , 32'hFC090CE0 , 32'hF7B541A0 , 32'h03EBC058 , 32'h0130A2A8 , 32'h054E3208 , 32'h0D4FF9A0 , 32'hFFFE3BF8 , 32'hF67F4F00 , 32'h030ACA4C , 32'h0DCD9010 , 32'h0314B2B8 , 32'h06E78830 , 32'h04096BC0 , 32'h01C1CF4C , 32'h0BA7DC30 , 32'hF19D9F90 , 32'h072EEE60 , 32'h1786EBE0 , 32'h0AB31B10 , 32'hEBE8F640 , 32'h00AF72D8 , 32'h001F22B0 , 32'h07B42BB0 , 32'h0001D5EE , 32'hF43E6F10 , 32'hE91536A0 , 32'hFEE06EA8 , 32'hDD176380 , 32'h03455E5C , 32'h000193E0 , 32'h0C1CFF10 , 32'hFE43B988 , 32'hFC3F8668 , 32'h0CB95610 , 32'hFFFC0D7F , 32'hF2132C90 , 32'h03A7C520 , 32'hF6D785B0 , 32'h152A7340 , 32'hFF7AC8FD} , 
{32'hE9224200 , 32'hF91B6EE8 , 32'hFB116DE8 , 32'h00005431 , 32'h000182B4 , 32'hF39A6630 , 32'h0C293A00 , 32'hFFED48DA , 32'hFFFECD9E , 32'h115E0500 , 32'h0510C200 , 32'h08AEC070 , 32'h1A75DBA0 , 32'h00F65F92 , 32'h04B0E4A8 , 32'h15E44460 , 32'h086E9C50 , 32'h0106E5A0 , 32'h06ED7408 , 32'hFFFF9319 , 32'hFB30E210 , 32'h09180130 , 32'h173154A0 , 32'h00002E95 , 32'hF2F2F500 , 32'h0659E378 , 32'hFCABCB90 , 32'hF9930048 , 32'h08C43890 , 32'h1AE74540 , 32'h0E305A70 , 32'hFB69E118 , 32'h10613060 , 32'hF07FED60 , 32'h0002E560 , 32'h00444BCF , 32'hEF9CC9E0 , 32'hFE255E68 , 32'h033EA0B8 , 32'h05630CF8 , 32'h06DE0830 , 32'h0202439C , 32'h01499D9C , 32'hFB22B270 , 32'h0CDCB230 , 32'h04959408 , 32'hFA2C9048 , 32'hEAA0FDE0 , 32'hFC072C04 , 32'hFE1D84B4 , 32'hFBAD6E30 , 32'h0415DA90 , 32'hE45EBFC0 , 32'hFC1F1F60 , 32'h06C41698 , 32'h03B812FC , 32'hFDE7F894 , 32'hFAE2E718 , 32'hE750C4C0 , 32'hDF6F67C0 , 32'hFD1601E4 , 32'h0466B290 , 32'hF7274CA0 , 32'h088947A0 , 32'h01C8C9B0 , 32'hE58197E0 , 32'hFFFEECAE , 32'hF82AEAE8 , 32'hFF71201B , 32'h12F138A0 , 32'hFEC7AA64 , 32'h0A45A660 , 32'h0443BF58 , 32'h03537C70 , 32'hF7DBDF00 , 32'h08CF75D0 , 32'hF2498BB0 , 32'h17177940 , 32'h13FA1A00 , 32'h08A3E5B0 , 32'hF57E1670 , 32'h0B2F1EE0 , 32'h0D7EBAE0 , 32'hFFFE0B01 , 32'hF7166120 , 32'h0BD9D5F0 , 32'hF373B680 , 32'hEAFAB520 , 32'hFEEEBC28 , 32'h0000197D , 32'hF0F35D80 , 32'h03DC2A60 , 32'h02E8CAE4 , 32'hFE2A7CA0 , 32'hFFFDB46F , 32'hFA664970 , 32'h31A16680 , 32'hE8E359A0 , 32'h05E95500 , 32'hE7925100} , 
{32'h059CAB08 , 32'h1A525140 , 32'hF41AAFE0 , 32'hFFFE7B5C , 32'h0001339F , 32'h004C5174 , 32'hFF5F7E5C , 32'hFDDDA6B0 , 32'hFFFF6BD4 , 32'h119EBE40 , 32'h0D668070 , 32'hFFAF61ED , 32'hF6C86B90 , 32'hFBEC7AC0 , 32'hF77566B0 , 32'hE422E640 , 32'h150B30C0 , 32'h0D1C8FE0 , 32'hFB8E1DB0 , 32'h0002E6BF , 32'h04068B28 , 32'h1A94C3A0 , 32'h0119BE1C , 32'h0001B8FA , 32'hF318A310 , 32'h011EB560 , 32'hF60D7520 , 32'h021F8860 , 32'h060A8FA8 , 32'h06019C20 , 32'hECEE0860 , 32'h09F1AC10 , 32'hFF0F4C8F , 32'hEAD8A900 , 32'hFFFCC83B , 32'hF5156DE0 , 32'h01252F1C , 32'h14D5EA60 , 32'h094DCF40 , 32'h0DD72810 , 32'hF9E26BF0 , 32'hFFA7F7F7 , 32'h05090C38 , 32'hFE0884FC , 32'h074582D0 , 32'h1F151680 , 32'h05698B30 , 32'h0BCAE490 , 32'hFC044090 , 32'h20D6BF00 , 32'h11869FC0 , 32'hD8491240 , 32'h0175DA90 , 32'hEDDB1620 , 32'h109EFA00 , 32'hFA1C0318 , 32'h0D82B820 , 32'hF39A37A0 , 32'hFCBE5378 , 32'h0CA15B10 , 32'hE9BA6840 , 32'h01CEC8A8 , 32'h046A43A0 , 32'h0ADC4BF0 , 32'h084A31A0 , 32'hF55EB490 , 32'h00028853 , 32'hF98E0328 , 32'hFEECC8B4 , 32'hFB278CB8 , 32'hFC1EC758 , 32'h0163FC04 , 32'h00ACABA2 , 32'h0667AB78 , 32'h0A57E400 , 32'h1243D860 , 32'h03E7ECD0 , 32'h04694C08 , 32'hFF476684 , 32'hFBC91448 , 32'hF728E080 , 32'hE7F68E80 , 32'hF9558068 , 32'h00007D37 , 32'h03CE2D48 , 32'h055F1640 , 32'hFB6BC650 , 32'h03F6475C , 32'hFEDF3A18 , 32'h000074E1 , 32'h0348769C , 32'h02646C7C , 32'h01554144 , 32'hF51980B0 , 32'h0001F83A , 32'hF3046CC0 , 32'hF51800D0 , 32'hCE1EBF80 , 32'h03EEEE58 , 32'h131227C0} , 
{32'hF33FA150 , 32'h1617A540 , 32'h063AF500 , 32'h00011784 , 32'h00000388 , 32'hEE2A1180 , 32'hEBB1BB60 , 32'hFBEF9FA8 , 32'hFFFF576A , 32'hF76E40C0 , 32'hFEA190D0 , 32'h183F7780 , 32'h00C7384F , 32'h1278F820 , 32'h03E2FC7C , 32'h145E0900 , 32'hF074DC40 , 32'h00F6EF1B , 32'h1FCEE0A0 , 32'h0003AF38 , 32'h004BCD63 , 32'hF9793250 , 32'h04B5E640 , 32'hFFFEE1FA , 32'h05F134B0 , 32'hFD6A38B8 , 32'hF4356670 , 32'hFD06E1C0 , 32'hFBDB1B28 , 32'h0F202D00 , 32'h056397A8 , 32'hFB0251B0 , 32'h080DBA60 , 32'h0B5C6610 , 32'h000062E3 , 32'hED79D060 , 32'hF61B6FF0 , 32'h0512B580 , 32'h0BA60220 , 32'hF61EE7B0 , 32'hEB4529C0 , 32'h006ECC8F , 32'h041B7580 , 32'h045C4D60 , 32'hFDD0D9E4 , 32'hE9A6D200 , 32'hF5B2B350 , 32'h053DEFB0 , 32'h0D72E8B0 , 32'h0D709780 , 32'h09856120 , 32'hF6D80A30 , 32'hF7B291A0 , 32'hF00ACDE0 , 32'h03E8A41C , 32'hE98D8080 , 32'h13802B20 , 32'hF18D8490 , 32'h188E79A0 , 32'h055722B0 , 32'hFE10441C , 32'hF8C2D630 , 32'hE2C46040 , 32'hF8CA1E60 , 32'hFC745768 , 32'h055D74C8 , 32'h0004BD25 , 32'h0D9137C0 , 32'hFE2DD15C , 32'h042AA900 , 32'h0ACAD6F0 , 32'h09844A40 , 32'hF1856400 , 32'h04BC97D8 , 32'h06F4E5F0 , 32'hF61EFCA0 , 32'h08B39A40 , 32'hFA92F850 , 32'hF6A9B640 , 32'hD666AD80 , 32'hEEDA9CA0 , 32'hE0246D80 , 32'hF2DADD30 , 32'h000243E4 , 32'h035C9234 , 32'hF1358460 , 32'h09748860 , 32'hFCE106AC , 32'hF5B0BC30 , 32'hFFFD6443 , 32'hFFD993C7 , 32'h00CB2AF6 , 32'h082DCCB0 , 32'hFE1E2B60 , 32'hFFFF5C47 , 32'h0E509030 , 32'h231DD580 , 32'h086B23B0 , 32'hF89380F0 , 32'h0A25E660} , 
{32'h02682648 , 32'hFC961100 , 32'h001BA2CA , 32'hFFFE0946 , 32'h0001DBEC , 32'h06B4D7B8 , 32'h09ABF2A0 , 32'h0713C158 , 32'h000037DC , 32'h24DD5240 , 32'hF9FF27D8 , 32'hE0AEF1C0 , 32'hF76EF3E0 , 32'hE1021CE0 , 32'h192CA180 , 32'h0A1AF220 , 32'h08D9F740 , 32'h08B660B0 , 32'hFBB43F00 , 32'hFFFFAED8 , 32'h1F43C9C0 , 32'hFCAE6174 , 32'hEEACFB60 , 32'h00025279 , 32'h2E41A880 , 32'hF28EEB00 , 32'hF0439750 , 32'hFFA8B037 , 32'h17D1D3A0 , 32'hFCAC547C , 32'hFCE7EBF0 , 32'hFCE0C118 , 32'hFBADC978 , 32'h0E4F1970 , 32'h00000C7D , 32'hED514F00 , 32'hF8D029E8 , 32'hF45F9800 , 32'h03CE182C , 32'hFF0A2AF6 , 32'h28BFBA40 , 32'h0060D4C6 , 32'hFF91841E , 32'h011FA41C , 32'h04E45D78 , 32'hEFA25C80 , 32'h0B113140 , 32'hF3060470 , 32'hF838BE88 , 32'hF17A8BB0 , 32'hF845B0C0 , 32'hFBA8AED8 , 32'hF5177C90 , 32'hFB7A2478 , 32'h081B2110 , 32'hFA086E70 , 32'h0FCCA870 , 32'h1243DA20 , 32'h10461680 , 32'h0B5334F0 , 32'hF545F160 , 32'h03542A7C , 32'h081A11F0 , 32'hFAC13110 , 32'h06916158 , 32'h123E03C0 , 32'hFFFB5D08 , 32'hF5DA4AE0 , 32'hF8579AA8 , 32'hFC3504C4 , 32'hF6094A00 , 32'h09FD19C0 , 32'h0C181EB0 , 32'h0432CB10 , 32'h03217FDC , 32'hF66BA400 , 32'hFD1A4C88 , 32'h01859D10 , 32'h09F68810 , 32'hED998C40 , 32'h06DF6EA0 , 32'hF2A594F0 , 32'h01199BA0 , 32'hFFFD8D55 , 32'h06901448 , 32'h013C2120 , 32'hFC3AB3A8 , 32'hF86A19E8 , 32'h01E6F8EC , 32'h00014EBE , 32'hF52283B0 , 32'hFB0EA990 , 32'h0515D928 , 32'hEF656360 , 32'h00040F15 , 32'h08217310 , 32'h12434480 , 32'hF3406330 , 32'hFBC26C60 , 32'h0562D9A0} , 
{32'hFCBD5A28 , 32'hFA2FF600 , 32'hFDBBFAEC , 32'hFFFE0845 , 32'hFFFEC14D , 32'hF4EBBDD0 , 32'hF580B9F0 , 32'h00D5BE6D , 32'h00022876 , 32'hFC5E12D4 , 32'h03E256D4 , 32'hE4E5FDE0 , 32'hE0C76EC0 , 32'h0AF8E740 , 32'hEF925380 , 32'h09074160 , 32'hFDDD8564 , 32'hE5E31100 , 32'hFA4FD760 , 32'h0000C7AC , 32'h10EC78E0 , 32'h009E88BD , 32'h0D438F10 , 32'h0002934C , 32'hFB269AD0 , 32'hF3564DA0 , 32'hF9F05160 , 32'h06621A88 , 32'h0089C649 , 32'hE7934840 , 32'h16FDB3C0 , 32'h0128BF00 , 32'h1BEC07A0 , 32'hEDEE0420 , 32'hFFFF957D , 32'hFCE58A44 , 32'hF825DDB8 , 32'h0E5EED60 , 32'hFC4AB66C , 32'h05AC86F0 , 32'hEB3DF3C0 , 32'h00CB322D , 32'h068FE7E8 , 32'hE8A1EC40 , 32'h03513208 , 32'hF5CCE270 , 32'h055E5978 , 32'hFD39B13C , 32'hF9B89558 , 32'h0C7F8B30 , 32'hE2F0B440 , 32'h1FDBA020 , 32'hFB1F36C8 , 32'h0F3E6DC0 , 32'h09B37FA0 , 32'hFC723C94 , 32'hFE7FAD10 , 32'hF7C3B5F0 , 32'h0B9E6DF0 , 32'hF19EBFC0 , 32'hF4A2A090 , 32'hFDB2CC0C , 32'h139B0840 , 32'h094FFCC0 , 32'hF5EE1C60 , 32'h19932480 , 32'h00018B8E , 32'h1191E000 , 32'h0460FD50 , 32'h0475ED18 , 32'h0269FEF8 , 32'h09D71990 , 32'h0CB30BD0 , 32'h0477E8A8 , 32'h0BD0F1D0 , 32'h08C319B0 , 32'h0404E870 , 32'hF6D054D0 , 32'h02B14160 , 32'hF667C590 , 32'hEEBA2740 , 32'h16DA3640 , 32'hF58EE930 , 32'h000568F6 , 32'h1C70CEA0 , 32'hFD93E9C4 , 32'h0AF5FAB0 , 32'hFD3CF13C , 32'h149E3A20 , 32'h00029936 , 32'h1130AE40 , 32'h06690D08 , 32'h077CE528 , 32'hF722C680 , 32'hFFFE08F4 , 32'hF1658180 , 32'h07A04638 , 32'hE6F16320 , 32'h01F0D56C , 32'h08A67450} , 
{32'h040A66A0 , 32'hFCA2CCE0 , 32'h096C9E70 , 32'hFFFFDC43 , 32'hFFFDAE50 , 32'h0ED421F0 , 32'h01EBCB10 , 32'hF87C13E8 , 32'h0000B8FA , 32'hFE09E700 , 32'h0A13B970 , 32'hF2002E80 , 32'hF969AAE0 , 32'hFB4FB790 , 32'h04F554A8 , 32'h05362BA8 , 32'h0F0F2BB0 , 32'h0BCABE70 , 32'h07018DD0 , 32'hFFFF69D0 , 32'hF2B50E50 , 32'h1AC9CFA0 , 32'h1CED10A0 , 32'hFFFEFA34 , 32'h1E30A940 , 32'hF9220828 , 32'h004CE08F , 32'hFD6287CC , 32'hEC9CE240 , 32'h107057E0 , 32'h13C4EF40 , 32'h0137B714 , 32'h0B1FD800 , 32'h014EE8E8 , 32'hFFFDF92C , 32'hFFBBEFB2 , 32'hFCB81DE8 , 32'h04D08300 , 32'hF73336D0 , 32'hF64DB290 , 32'hFDEE9C34 , 32'hFED89170 , 32'h0B36C560 , 32'h05289DD8 , 32'hEF7DA8E0 , 32'h09259910 , 32'hF48DC550 , 32'h24BE3600 , 32'h013F56A0 , 32'h145159C0 , 32'h1316EC00 , 32'h010C0EAC , 32'hFEC0CEBC , 32'h1C5EECE0 , 32'h0D6C6270 , 32'h072DC7A0 , 32'h1CE1B560 , 32'h1507CD60 , 32'hFDCC66AC , 32'h068FD2F8 , 32'h170DBA40 , 32'hFEBC8494 , 32'h064B0E58 , 32'h0877DA10 , 32'hF3603900 , 32'hFF965E0F , 32'h0003B461 , 32'hFF3B4B96 , 32'h01C41F24 , 32'h0FCD9B60 , 32'h015A1368 , 32'h0B6CC630 , 32'h132B4340 , 32'h04527010 , 32'h0EAB6360 , 32'hFDAD7000 , 32'h025D8538 , 32'h150DC240 , 32'h0E0229F0 , 32'h12FCF160 , 32'hFCD03B74 , 32'hF1A659E0 , 32'h1A826860 , 32'hFFFE0FDB , 32'h1B83B0A0 , 32'hFE19CB24 , 32'hF809D348 , 32'hF272BB60 , 32'hF98CF878 , 32'h0000FD9E , 32'h0E145360 , 32'h0B00CFE0 , 32'h0091E089 , 32'h04D457C8 , 32'h0000ACEB , 32'h01CA626C , 32'hFDFB80D8 , 32'h1D43A580 , 32'hF2AD9B30 , 32'h07D8DFD0} , 
{32'hEA182220 , 32'h0F3A9900 , 32'h09FADA60 , 32'h000097E7 , 32'hFFFF01CB , 32'h00EE7F26 , 32'hFD7BDA44 , 32'h06474FF0 , 32'hFFFF5857 , 32'h26B226C0 , 32'h05ED6C40 , 32'h06CD23C8 , 32'hDE4182C0 , 32'h05FBF990 , 32'hFC1DF928 , 32'h028BF78C , 32'h13390AC0 , 32'hEE5E31C0 , 32'h08650730 , 32'hFFFC63B9 , 32'hEA8BF9E0 , 32'h18FEEEC0 , 32'hF215B120 , 32'hFFFD89A9 , 32'hF4264E30 , 32'hFADFDCB8 , 32'hF6357690 , 32'hFF8564BE , 32'hFEB577EC , 32'h05D46EF0 , 32'hF5A81E40 , 32'hF8F77998 , 32'hEF940080 , 32'hFA09BF50 , 32'h0000C1C0 , 32'h05848850 , 32'h06828958 , 32'hF86293C0 , 32'h0447E5B0 , 32'hF0961030 , 32'hEE41CCA0 , 32'h0083B9C6 , 32'hF869B108 , 32'h04B10EC8 , 32'hE272BBC0 , 32'hEC911980 , 32'h174CD920 , 32'h15F61FA0 , 32'h027B8CA4 , 32'hF9BE3830 , 32'hED959020 , 32'h27ADE880 , 32'hFDF7E67C , 32'hE9F42C60 , 32'hF9F3F460 , 32'hF47A5660 , 32'h0B9F1920 , 32'h0FF6B920 , 32'hFC6AF5F8 , 32'hF8F812E0 , 32'hF637F290 , 32'h02CBD048 , 32'h09E08410 , 32'hF7AEF4C0 , 32'h0CF4F000 , 32'hF6761620 , 32'hFFFE9281 , 32'h0AA51070 , 32'hF73D4EB0 , 32'h0487DCB0 , 32'hE9B26780 , 32'h01825490 , 32'hFBD53820 , 32'h059B1750 , 32'hFE13BD4C , 32'h0D24E3C0 , 32'hFA548390 , 32'hF4CFA860 , 32'h02FBD604 , 32'h0C6E8EB0 , 32'hF8141B58 , 32'hF264C390 , 32'h04B40F58 , 32'hFFFFDE7B , 32'hE51E4CC0 , 32'hF6889AE0 , 32'hED98DE60 , 32'hEE55DE80 , 32'h059EC6B8 , 32'hFFFE5EDC , 32'h02F3E59C , 32'hFE10DA90 , 32'hFB3DC258 , 32'h0394E540 , 32'hFFFE8AA6 , 32'h0FC2DB10 , 32'hF44FD700 , 32'h04B04F80 , 32'h03988A00 , 32'hF700C020} , 
{32'h06DED9E0 , 32'h049F0FC0 , 32'h16EBB7E0 , 32'h000043F3 , 32'h00028343 , 32'hFC42DB34 , 32'hF9913960 , 32'hF4AF4D70 , 32'h0000920B , 32'h0246D4BC , 32'hF3FCD570 , 32'h0AB9E680 , 32'h0A5CA240 , 32'hF2ADF290 , 32'hE3F34C80 , 32'h0088A2BC , 32'hE4D613C0 , 32'h086B9F20 , 32'hD55DEAC0 , 32'h000414F4 , 32'hE2DB91E0 , 32'h0364AB18 , 32'hF2C72470 , 32'h0000E2F3 , 32'h0209F2F0 , 32'hFD329E1C , 32'hF289B960 , 32'h09A64190 , 32'h14976E80 , 32'hDC794A80 , 32'hF4FE1F30 , 32'hF2EAFEC0 , 32'h17D93F80 , 32'hF3046730 , 32'hFFFEC675 , 32'hE16F1DA0 , 32'h0B1E88A0 , 32'hF68955C0 , 32'h034FE0AC , 32'hFB73C758 , 32'hF8EB8558 , 32'hFFDC8ABC , 32'hFFDA9295 , 32'h0356CD48 , 32'hF83B6040 , 32'hFB728D68 , 32'h03742E44 , 32'h04295A08 , 32'hEEC4BFE0 , 32'hF7E2D3D0 , 32'h07FA0868 , 32'hFE806478 , 32'h05A4E180 , 32'hEFA5A920 , 32'h0B4C9540 , 32'hF841CB10 , 32'h164BC9C0 , 32'h095B69C0 , 32'hEA4C5AC0 , 32'hF92FA0F0 , 32'h14304460 , 32'hF78F9D90 , 32'h040616A0 , 32'hFA402E28 , 32'h01B7A708 , 32'hF9727540 , 32'hFFFDA13A , 32'h08BDB8F0 , 32'hF9BA6B30 , 32'hFAE831A8 , 32'h0BFF4940 , 32'h0462CD90 , 32'h0481BE10 , 32'h0306ADD0 , 32'hEC755D80 , 32'h0751E420 , 32'hFB023618 , 32'h24057EC0 , 32'hF899F108 , 32'h028B166C , 32'h0664B5C8 , 32'h025FD31C , 32'hF1A6B350 , 32'hFFFE945C , 32'h193647A0 , 32'hE9A13F60 , 32'hFF82ADE6 , 32'hFE0DA198 , 32'h03B9339C , 32'h00010F6D , 32'hF803B608 , 32'h0073DAB1 , 32'hFDE0BC9C , 32'h07FB20B8 , 32'hFFFF7D09 , 32'h09C10110 , 32'h0AE016E0 , 32'hFE15E48C , 32'h03729D70 , 32'hFD1C4444} , 
{32'hFDCD42A8 , 32'hFBB4CA10 , 32'h01445234 , 32'hFFFFBCEE , 32'h0001D8DE , 32'hF51DE590 , 32'hF9EBC258 , 32'hF8009898 , 32'hFFFF5B65 , 32'h04914178 , 32'h0EF7C4F0 , 32'h051F7310 , 32'h194FF680 , 32'h03A66294 , 32'h04882408 , 32'h065DF0C0 , 32'hF4D0EAF0 , 32'hEEFB2FC0 , 32'h23BAE980 , 32'hFFFDF62C , 32'h00B387DE , 32'hF3F2B5E0 , 32'hFF721901 , 32'h0004C358 , 32'hFB9DC5A0 , 32'hF3B77A60 , 32'hF4E6AAC0 , 32'hFA5AE5C0 , 32'h13CD1480 , 32'hF3EFF720 , 32'hDC93F500 , 32'hE1674880 , 32'hFD104D2C , 32'hF4B07CF0 , 32'hFFFEECE6 , 32'h18FDD540 , 32'h0B8CCA20 , 32'hF8D87298 , 32'hEFC198E0 , 32'hF77C1CD0 , 32'h02B46394 , 32'h0023A761 , 32'h007E3D3D , 32'h05A71B00 , 32'hDE4DE800 , 32'hF7D727A0 , 32'hEBAA0D00 , 32'h0C7CEE10 , 32'h15659920 , 32'h05638910 , 32'hF62FD210 , 32'hFB9EEE50 , 32'hF282E8D0 , 32'h12BAB5A0 , 32'h08645230 , 32'h164CF9E0 , 32'hF89721B0 , 32'h0FC908B0 , 32'hF9D5C8A8 , 32'h0B96ABE0 , 32'h0916F9B0 , 32'hF60106F0 , 32'h1455D820 , 32'h01E8CF30 , 32'h05DB03D8 , 32'h00546522 , 32'h00004D5A , 32'hFF77D87B , 32'hFF328DBF , 32'hFAE387C0 , 32'h038D1BD4 , 32'h00106533 , 32'hFFE8FF03 , 32'hFAB43360 , 32'h07EE19E8 , 32'h08EA7970 , 32'hFD66C668 , 32'hFC45209C , 32'h03067584 , 32'hFCDF0680 , 32'h0E9B0720 , 32'hF7EAA5B0 , 32'hFB0E6AA0 , 32'hFFF9B79D , 32'h11AC2C40 , 32'hF5D3D5B0 , 32'hE5FB1920 , 32'h1A28CFC0 , 32'hF455D7B0 , 32'h0001B37C , 32'hFD774314 , 32'h03DD8428 , 32'hFA577DB0 , 32'hE6CE3020 , 32'h00054C0A , 32'hE534EE00 , 32'h0B429EF0 , 32'hEF9FAC20 , 32'h11BAAC20 , 32'h06559E68} , 
{32'h108FC920 , 32'h10AA96C0 , 32'h142F6140 , 32'h00032D35 , 32'h000358E2 , 32'hEA5C71C0 , 32'hE7A01620 , 32'hFEC7095C , 32'h0004A6FA , 32'hEDE556E0 , 32'hFF5C7DB2 , 32'h0F2E0330 , 32'hF12591C0 , 32'hF242B080 , 32'hFBEBAB70 , 32'hFF41F788 , 32'h0B073580 , 32'h0476F088 , 32'hFE4D3044 , 32'h0000B06C , 32'h06935F60 , 32'h09475350 , 32'hEC56F180 , 32'hFFFEF21D , 32'h078E4F08 , 32'hF9BE48B0 , 32'hF6EAA9E0 , 32'h0C61F6F0 , 32'h0486FD18 , 32'hEF07D920 , 32'h0DF55710 , 32'hFA86A818 , 32'hF99EA7A0 , 32'h033E9314 , 32'h00015CDF , 32'hF0A0BAA0 , 32'hFFEC6241 , 32'h065D39C8 , 32'hF875B000 , 32'h15305780 , 32'hF9EF14C8 , 32'hFF78D974 , 32'h00E706AC , 32'h02B02DF4 , 32'hF0045FD0 , 32'hE0642300 , 32'hFC1EE104 , 32'hFD909A48 , 32'hE9D55A20 , 32'h0A79FD10 , 32'h0140DE38 , 32'hF1775CE0 , 32'hF98EC820 , 32'h1EEB8000 , 32'hEE053A40 , 32'h00C62D43 , 32'hE79721A0 , 32'hFF1BF010 , 32'hEAB7A980 , 32'hF5A9CD40 , 32'hFDB81060 , 32'hF827F170 , 32'h0351D2B4 , 32'hFF8E446B , 32'h0EE4FD50 , 32'hED34B5A0 , 32'h0000C2A0 , 32'hF7937A40 , 32'hF35E6DB0 , 32'h191ECC00 , 32'hF45E11C0 , 32'h083203D0 , 32'hEF88CDA0 , 32'hFB73F100 , 32'h00A49DB7 , 32'hF951DC60 , 32'hFE8F25DC , 32'h064F6618 , 32'h18A119C0 , 32'hE90168E0 , 32'hF8F57CB0 , 32'hF7CB5A80 , 32'h1E7863E0 , 32'h00035DBB , 32'hF24C5530 , 32'h1DF2B600 , 32'hFA6B37F8 , 32'h12BAFBA0 , 32'h0DF04F50 , 32'h0000E2D0 , 32'hF8296730 , 32'hFE234174 , 32'h103861C0 , 32'h03AEBDC4 , 32'h0000B27F , 32'hF1626CF0 , 32'hF683ADB0 , 32'h066EFF00 , 32'hF9664410 , 32'h0132B030} , 
{32'hF40B6690 , 32'h020229A8 , 32'h0169E640 , 32'hFFFC7AE0 , 32'h00017421 , 32'h11A43620 , 32'hFFFFCF13 , 32'hF1247AC0 , 32'h0000EE7D , 32'h11D6C940 , 32'h0295FEBC , 32'hF5D011E0 , 32'hF1822FC0 , 32'hF618BC60 , 32'hFEBC3D24 , 32'h0EBD6BD0 , 32'h001A2C5C , 32'h0BD889B0 , 32'h091D03C0 , 32'hFFFA95BD , 32'h0F0C1000 , 32'hFBDA0C80 , 32'hEA7ECDC0 , 32'h0002613A , 32'h0EE51390 , 32'h091F98E0 , 32'hEF056CE0 , 32'h02944D28 , 32'h028A26D4 , 32'h05AB5B68 , 32'hF4EA3160 , 32'hF86AC2D8 , 32'h0B4A0B50 , 32'h0081180A , 32'h0000106F , 32'hFFB2E050 , 32'hFF9DD488 , 32'h05C9B280 , 32'h0C977880 , 32'hFD933BB0 , 32'hE962B3A0 , 32'h009E96EC , 32'hF7CE3800 , 32'h0EFC8840 , 32'h09D23640 , 32'hF4135320 , 32'h0AE817C0 , 32'hFCFD2FC8 , 32'h1E3A4E40 , 32'h1A2FF640 , 32'h15307E40 , 32'h03D77B94 , 32'h111AA580 , 32'hF62C7FC0 , 32'hF35F26A0 , 32'h02FB2DC0 , 32'h04FFD208 , 32'hEF524920 , 32'hEF48EEA0 , 32'hDF1B9580 , 32'h0D401570 , 32'h06656A08 , 32'h0B857410 , 32'h0AEDC840 , 32'hFDA3EDE4 , 32'hFCD75868 , 32'h0000AF18 , 32'hFC02AFA0 , 32'hFC751188 , 32'hEE569860 , 32'h0CF783C0 , 32'hF70321D0 , 32'hF7BF1B00 , 32'hFA9F9B78 , 32'h0E3D65C0 , 32'h02A96988 , 32'hF98BCD30 , 32'hFD7EB944 , 32'hFFEAD347 , 32'hED064F20 , 32'h0709AB00 , 32'h2DF1CF00 , 32'h058219C8 , 32'hFFFF3527 , 32'h080912A0 , 32'h0D70D120 , 32'hFDE03A88 , 32'hEECE2F60 , 32'hD8F2F680 , 32'hFFFE6A03 , 32'hECEA7B00 , 32'h06747180 , 32'h05BC2E00 , 32'h01372070 , 32'h00006B7A , 32'hEB6CA3E0 , 32'hEFC97020 , 32'h0F400000 , 32'h04FAA048 , 32'h070C9E70} , 
{32'h0129A380 , 32'hFBDC0698 , 32'h1343BF80 , 32'h0004C03E , 32'hFFFFAE94 , 32'h02B7DFC4 , 32'hF93FCAB0 , 32'hFCC562E4 , 32'hFFFCE3E2 , 32'h0E235460 , 32'h09F95070 , 32'hF00D42D0 , 32'hF31F50D0 , 32'h06181950 , 32'hF788AB00 , 32'h18B52120 , 32'hF9ED8578 , 32'hF86E4598 , 32'h00C501E3 , 32'hFFFED4D1 , 32'h2A75A9C0 , 32'hF944C638 , 32'h01AEFC20 , 32'h0002A442 , 32'h0C97E880 , 32'h02B9F170 , 32'h09ECC100 , 32'hF321B6E0 , 32'hFACB5E48 , 32'h04B7DB18 , 32'hF12F9DE0 , 32'h0B295B60 , 32'h0251EBD0 , 32'hE33FAEE0 , 32'h00003FF2 , 32'hF72F53A0 , 32'h034AB098 , 32'h0B767DE0 , 32'hF18DB710 , 32'hFBB17DF0 , 32'h073E6880 , 32'h03028AF8 , 32'h00E2750A , 32'h100CE000 , 32'h0AB34FB0 , 32'h0CD63780 , 32'hDC748700 , 32'hFFEE4815 , 32'hFBD67960 , 32'hF854AF08 , 32'hF86EE328 , 32'hEBCF5D20 , 32'hFB517048 , 32'hFA2189A8 , 32'hFE2F5528 , 32'hFC231878 , 32'h02B8EA6C , 32'hEF888160 , 32'hF7E0AA00 , 32'hFDB36694 , 32'h1ADA2440 , 32'h10331E00 , 32'h0C538BC0 , 32'h000D6576 , 32'h1B177D80 , 32'h0AC045A0 , 32'hFFFEB049 , 32'h11757860 , 32'hF9E8A3C8 , 32'h1CCBFFC0 , 32'h11A5D160 , 32'h04A524A0 , 32'hF5085820 , 32'h05EC7090 , 32'hFB99D7C8 , 32'h03E60608 , 32'h010BD010 , 32'h07E7E230 , 32'hEFE6C860 , 32'hFF265E0F , 32'hFB8091C0 , 32'hFB2019E8 , 32'hF0A8BF90 , 32'hFFFF1792 , 32'hE494EBC0 , 32'hF7678960 , 32'hE472E8A0 , 32'h047F6C68 , 32'h06586830 , 32'h000238A1 , 32'h1784F7E0 , 32'hFFAB1467 , 32'h01953644 , 32'h1745FF60 , 32'hFFFDD264 , 32'h06B48A58 , 32'hEEEEE5E0 , 32'h05AE26B8 , 32'hFE8535D0 , 32'hE9F5B800} , 
{32'h074715A8 , 32'hF582A420 , 32'hF3DDB120 , 32'hFFFB17F9 , 32'h0002033A , 32'h1735F0A0 , 32'hF71BE290 , 32'h015053C8 , 32'hFFFF1C1F , 32'h135285E0 , 32'h0AA22720 , 32'h069A2A10 , 32'h0233E854 , 32'h12EA05A0 , 32'hF4218A60 , 32'hE5A89140 , 32'hFB9C84B8 , 32'hD02AAD40 , 32'hFE8EA0A8 , 32'hFFFCE5AF , 32'h0A293C00 , 32'h090358E0 , 32'hFEF835A4 , 32'h00018825 , 32'h12E3B760 , 32'hEFA4E7A0 , 32'h0CD6CB70 , 32'h0C44B8B0 , 32'hFEE6E138 , 32'h05AE1540 , 32'hF7BE27C0 , 32'hE9709300 , 32'h13508C80 , 32'hF9029C90 , 32'h0002F0C7 , 32'hF5D00290 , 32'hFD1732A8 , 32'h126AE5C0 , 32'h0FA54890 , 32'hFFEF46E6 , 32'h09ABB1B0 , 32'h005D01AD , 32'hF977F088 , 32'hF2746790 , 32'hEA7F5360 , 32'hFF559BD2 , 32'hFFCF5E95 , 32'hF0926220 , 32'hF0E38920 , 32'hF097A840 , 32'h09D8F5F0 , 32'hED305DE0 , 32'h16E55220 , 32'h114857A0 , 32'hEFD63BE0 , 32'hF927DD98 , 32'h16F4B060 , 32'h023352D4 , 32'h0C817270 , 32'hF9CE8E08 , 32'h08F7C8E0 , 32'h00BF4175 , 32'h0669FD10 , 32'h0D5376A0 , 32'hF4022FF0 , 32'hDD180B00 , 32'h000139BA , 32'hFD3F90D4 , 32'hFC7A5FA0 , 32'hFDEF1344 , 32'hEFB1B140 , 32'hF34790B0 , 32'hF897C658 , 32'hFDFC754C , 32'hF49A4DF0 , 32'hF9330A58 , 32'h0745E230 , 32'hF2157650 , 32'hF93FE6A0 , 32'hFE9A5E50 , 32'h03A5915C , 32'hFE858068 , 32'hF9C46F50 , 32'h00057012 , 32'hF8051218 , 32'h11212CC0 , 32'h10BB6A80 , 32'hFDBF5530 , 32'hF05EF570 , 32'h0002C61A , 32'h13DB7DE0 , 32'hFD69B924 , 32'hFD3316B8 , 32'h0524A1C8 , 32'h0002B20E , 32'hF76286E0 , 32'h1B0B8660 , 32'h09A96900 , 32'h031BDEEC , 32'hF5AFEED0} , 
{32'hD90BBC80 , 32'h006C7879 , 32'h0767CB48 , 32'h0001452F , 32'hFFFBCD85 , 32'hFE3C8448 , 32'h06E58F80 , 32'h04A8A590 , 32'hFFFCBACC , 32'h02D653E8 , 32'hF5C6CCC0 , 32'hF5FCA750 , 32'h08217AE0 , 32'hFEBBF774 , 32'h0F136720 , 32'hE46561A0 , 32'hF0085AE0 , 32'hFAD6BBC8 , 32'h039D59BC , 32'hFFFD092E , 32'h02C41980 , 32'hF5AFA080 , 32'h074808A8 , 32'h0000BA06 , 32'h06F540F0 , 32'h092AA4E0 , 32'h08AC6500 , 32'h07770A08 , 32'h00CA5AE1 , 32'h01D64ECC , 32'hF71C9FA0 , 32'hE39A9D40 , 32'hFE4C567C , 32'hF7010C10 , 32'hFFFE9439 , 32'hEBB7D140 , 32'hFFBC3772 , 32'hE0F8F920 , 32'h0A846D80 , 32'h16BA60A0 , 32'hEB102360 , 32'hFFFAF706 , 32'hFCCE6BB0 , 32'h0D025EF0 , 32'h0DB12490 , 32'h190CB260 , 32'hEFB63880 , 32'h103364C0 , 32'hECDA6420 , 32'hF676E7A0 , 32'h10C77F40 , 32'h04361D90 , 32'h02376500 , 32'hFB1EEDB0 , 32'h0206D2E8 , 32'h08A60240 , 32'hEDD7FFA0 , 32'h087C8120 , 32'hF772C2C0 , 32'hEDC58180 , 32'h009E4439 , 32'h0123EA68 , 32'h0D444CC0 , 32'h0015C7DE , 32'h025D05B8 , 32'hFC6F1BFC , 32'h0001D729 , 32'h04359530 , 32'h0C10D5D0 , 32'hFB6352E0 , 32'hF99D35A8 , 32'hF8A064B0 , 32'h012A67D4 , 32'h08459C70 , 32'h0EA0B140 , 32'hFB1996B0 , 32'hF9C8AF40 , 32'hF1F82CA0 , 32'h05693660 , 32'hED1FC980 , 32'hF73930A0 , 32'h02285398 , 32'h18A07060 , 32'hFFFCF765 , 32'h01EF5740 , 32'hF9616E78 , 32'h02648E10 , 32'h04FD2BA8 , 32'h0865D5F0 , 32'hFFFD6B76 , 32'h230FB740 , 32'hFAE325D8 , 32'h21200440 , 32'hE7A9F0A0 , 32'h0002EF75 , 32'h20B437C0 , 32'hFCE68CA4 , 32'h0387185C , 32'h06308DE8 , 32'h095176D0} , 
{32'h06DD2060 , 32'hFA0EB9E8 , 32'hF5D4AD10 , 32'h00001C44 , 32'h0003507A , 32'h1B2086E0 , 32'h023324C4 , 32'h08993BD0 , 32'h0003C1D3 , 32'h035750B4 , 32'hF215D460 , 32'hFDA34080 , 32'h06492240 , 32'hF7ADF5E0 , 32'h03E75C6C , 32'hEC7ECF40 , 32'h0AF49110 , 32'hEB283880 , 32'h09894280 , 32'hFFFED8E4 , 32'hEC64CEC0 , 32'hFE49E300 , 32'hE54066E0 , 32'hFFFF96FB , 32'h075E06A8 , 32'hF2ACFDA0 , 32'hFDFCDF6C , 32'h01D88EB8 , 32'hF111E9A0 , 32'h0699A3F0 , 32'h1E532BC0 , 32'h0C6CDC80 , 32'h20F2A580 , 32'h0174A79C , 32'h000145F4 , 32'h0B6504A0 , 32'hFC71736C , 32'h03312D08 , 32'hEB5FAB60 , 32'h102E36C0 , 32'hFC6BF34C , 32'hFD720194 , 32'hEC33C5E0 , 32'hFE3BC954 , 32'hE77F5560 , 32'hFFF909D8 , 32'hF98CB0B0 , 32'hED04F160 , 32'hF304D5C0 , 32'h0C274710 , 32'h00CD2ADB , 32'h07D8A480 , 32'hFFCC9051 , 32'hEF8BF3E0 , 32'h07811650 , 32'h1447DC40 , 32'hFB370120 , 32'hEF7DBC80 , 32'hE508B500 , 32'h12230280 , 32'h07235920 , 32'h02D9DC84 , 32'hF3548590 , 32'hFB89ABB0 , 32'h0B509F20 , 32'h18821EA0 , 32'h0000789A , 32'hFEEC4B54 , 32'hFEA308D4 , 32'hF6CDDC30 , 32'h0B946990 , 32'hEFFF8600 , 32'h0B6E2760 , 32'hF56FED90 , 32'h05D571F8 , 32'hFB94C730 , 32'hDDFE3640 , 32'h09149280 , 32'hF4DDDE30 , 32'hE3DD9240 , 32'hEECA51E0 , 32'hF4325D60 , 32'h0BF94E80 , 32'hFFFD4620 , 32'hF04E56D0 , 32'hEB7C14A0 , 32'hF1338570 , 32'h0321CB40 , 32'hF64EEE40 , 32'h0005D437 , 32'h074A6530 , 32'h0507BD50 , 32'hF8748700 , 32'h055C5CA0 , 32'hFFFC897E , 32'h032295F4 , 32'h060CF468 , 32'hF7E13350 , 32'h0576FFD0 , 32'h04B7ED88} , 
{32'h19D9A9C0 , 32'hF64814F0 , 32'h0370E044 , 32'hFFFE265D , 32'hFFFE557F , 32'h0E688690 , 32'hF8DEBA20 , 32'hFF9D2410 , 32'h0001AAB5 , 32'h057330C0 , 32'hFDB92CCC , 32'hFCACC8F8 , 32'hFDE8089C , 32'hE5166CC0 , 32'hDF840C40 , 32'h03F9C5FC , 32'hEE2FCA60 , 32'hFABE0220 , 32'h22FAD140 , 32'hFFFE18F7 , 32'hFD53765C , 32'h01078470 , 32'h00093B3F , 32'hFFFF8E04 , 32'hF33715B0 , 32'h03494F50 , 32'hEE51B780 , 32'h045DF2E8 , 32'hE48B2040 , 32'hF64ECE90 , 32'h07DD9C50 , 32'h0457B558 , 32'hF692E680 , 32'h0D1AF360 , 32'hFFFC94FF , 32'h06D6C6E8 , 32'h08080EC0 , 32'hD9DC4780 , 32'h13830B80 , 32'hF98AE628 , 32'h03BE0A2C , 32'h000904B7 , 32'h05C79D00 , 32'h1367A720 , 32'hF03A3160 , 32'h1DD90F40 , 32'h012E3534 , 32'hF7C47590 , 32'hF62D4F80 , 32'h09E640F0 , 32'hED3C8240 , 32'hE2ED2D00 , 32'h017F6134 , 32'hFA5E9480 , 32'hFF8FBD24 , 32'hF835C880 , 32'hEF9672E0 , 32'h159F88A0 , 32'h00BC2C7E , 32'hED9D3B60 , 32'h08E0BB40 , 32'h027EC378 , 32'h0C7DBD40 , 32'h0019044B , 32'hE2641D00 , 32'h11540AA0 , 32'h0002D85A , 32'h01DE6CC4 , 32'h01C2198C , 32'h00C75549 , 32'h01AAAFF4 , 32'h0221DAFC , 32'hFCAAFB94 , 32'h0BDDB570 , 32'h05A91D38 , 32'h08C500A0 , 32'hF99EC248 , 32'hF5D3A470 , 32'h0DADCB40 , 32'hFD0B3D84 , 32'hEEC0B5C0 , 32'hF30E1C00 , 32'hF18A7F80 , 32'h00009A6A , 32'hFB26BDB0 , 32'h0BBCDA30 , 32'h08F41510 , 32'hE97401A0 , 32'h01D65014 , 32'hFFFF1A5B , 32'hF6B30BB0 , 32'hFB7002D0 , 32'h0EC73DA0 , 32'h1150B040 , 32'h000233A6 , 32'hFB789760 , 32'h084144D0 , 32'hF8CC90E0 , 32'h03BE77F0 , 32'hF75B33A0} , 
{32'hFA52A188 , 32'hF73CAEA0 , 32'h01EEF1D4 , 32'h0001BD8E , 32'h0000B381 , 32'hF2D5B3D0 , 32'h044D85E8 , 32'hFBD85928 , 32'h00008F91 , 32'hF7CF7510 , 32'h01AB4E08 , 32'hF98B1F30 , 32'h0E8C91C0 , 32'h0161EFD4 , 32'hECE65CC0 , 32'hE77DE1A0 , 32'hEAF09F40 , 32'h0008B3E4 , 32'h0619C640 , 32'hFFFF240B , 32'hFEC6DA18 , 32'h1FD86F80 , 32'h0156B994 , 32'hFFFDB2D1 , 32'h173A6D20 , 32'hF7CA4EC0 , 32'hFE6E3EB4 , 32'h07BC6C60 , 32'h0EE36790 , 32'hF1815940 , 32'h12372FC0 , 32'h03D87D80 , 32'hED3A6840 , 32'hF0C240D0 , 32'h00011185 , 32'hF9E64E80 , 32'hFBE29AA0 , 32'h0FE01B40 , 32'hF23EB470 , 32'h0048D025 , 32'hF5FA8EA0 , 32'hFFD4277E , 32'h004182B4 , 32'h10C52460 , 32'h0C7E9BA0 , 32'h08BF1DD0 , 32'hFBDDCD90 , 32'hE4FD0E20 , 32'h187A5940 , 32'hF927AF40 , 32'hEE7DF000 , 32'h0BB83F10 , 32'h08A0C010 , 32'h048ECB68 , 32'hF656EB30 , 32'hF2877E10 , 32'hFBD07A60 , 32'h1B03B780 , 32'hF17F28C0 , 32'h0CF4F5A0 , 32'h00BA1A0B , 32'h0C3425D0 , 32'hD9C32840 , 32'hFBBF69E0 , 32'h1AF71A20 , 32'hFC5EDF98 , 32'hFFFE0431 , 32'hF2A08840 , 32'hFF5393D7 , 32'hFC46FFD8 , 32'h03661650 , 32'h03AF5CE8 , 32'hEBCBBD40 , 32'h0C19B4E0 , 32'h1C0FD1C0 , 32'h068D92B0 , 32'hFA1CFF00 , 32'hE49F7380 , 32'h128E76A0 , 32'h00A17964 , 32'h0A010E90 , 32'hFC67F9BC , 32'hFBF10968 , 32'h00006ED0 , 32'h1354D040 , 32'hFB177578 , 32'hFB44D230 , 32'hEC1017A0 , 32'hEDB582C0 , 32'h0002ED7D , 32'h0AF20550 , 32'h04A3D7A8 , 32'hF76779E0 , 32'h0A176920 , 32'h00048426 , 32'h0330A594 , 32'hFBE637C8 , 32'hF671D850 , 32'hF3A088A0 , 32'hF666AFF0} , 
{32'h0D4B4B90 , 32'hEA539EE0 , 32'h1788D9E0 , 32'hFFFF8A04 , 32'hFFFD20E8 , 32'hFF3E9034 , 32'h0FA58400 , 32'hFAB26AC0 , 32'h0001FEB4 , 32'h17E69280 , 32'hFBE188D0 , 32'hE9E51260 , 32'h034B6CA4 , 32'hF796CB20 , 32'h0C52F070 , 32'h03A42644 , 32'hFC55A7FC , 32'hF09B4C20 , 32'hE95F18A0 , 32'hFFFF3C7D , 32'h01537DBC , 32'hFCE9B74C , 32'h12580520 , 32'h0002454C , 32'h00B18BDE , 32'h19C67560 , 32'h0FE21A00 , 32'h08068D80 , 32'h03501FBC , 32'hF7BCAC00 , 32'hFC575024 , 32'h00E2828C , 32'hF17F17B0 , 32'h17202BA0 , 32'hFFFF7536 , 32'h04A032E0 , 32'hFBE43D98 , 32'h1A5C6C80 , 32'h027769E8 , 32'hEA7BDFA0 , 32'hE37AC940 , 32'hFED0E014 , 32'hFACAA0D0 , 32'hFCA51548 , 32'hFBD2F260 , 32'hFD12C5C0 , 32'hFA123EB0 , 32'h03E81798 , 32'h10844FE0 , 32'h190A8300 , 32'hFE15FA7C , 32'hF34BF660 , 32'h0B91B8F0 , 32'h0342E214 , 32'hFA844768 , 32'h124B02A0 , 32'h087D7FE0 , 32'hF616A980 , 32'hF0EF0170 , 32'hE9ECDD40 , 32'h0412B330 , 32'hF99C3338 , 32'hE0D61EA0 , 32'hF5733870 , 32'hEDE137C0 , 32'hFED77190 , 32'hFFFF08FC , 32'h028191A8 , 32'hFA101518 , 32'hFF01E250 , 32'hEB148140 , 32'h0F1148E0 , 32'h0B9D3310 , 32'hF2853580 , 32'hEE0C8AA0 , 32'hFF9956FF , 32'hE3403420 , 32'hEB8368C0 , 32'h10C8BAA0 , 32'hF9006678 , 32'hFF41757E , 32'hEAE5DDE0 , 32'hF1980D80 , 32'hFFFF1945 , 32'hFF0F0592 , 32'hF9AE8DA0 , 32'hFE38AEF4 , 32'h18857840 , 32'h0A958680 , 32'h00008FC2 , 32'hFD19B398 , 32'hF5DCE2A0 , 32'h0A8A9AF0 , 32'hF97CE3E0 , 32'h00025C85 , 32'h08A9FD50 , 32'hFEAD813C , 32'hF57E8B90 , 32'hFC597C18 , 32'hF817DE30} , 
{32'h11166320 , 32'h065BE588 , 32'h06631340 , 32'hFFFFEF04 , 32'hFFFF1D1E , 32'h0A54A190 , 32'h28822380 , 32'hEB433080 , 32'hFFFB05EA , 32'hF7A53930 , 32'hF83D6118 , 32'hE772C0E0 , 32'h003D8EFB , 32'h01D8DEDC , 32'h20101F80 , 32'h112B9D20 , 32'hFE08C530 , 32'hFB1F4A18 , 32'h0D5522F0 , 32'hFFFC215D , 32'hF4BB27E0 , 32'h042A8C20 , 32'hF7EE6EA0 , 32'hFFFCF1A4 , 32'hEBAA7780 , 32'h03AE4DE8 , 32'hF7F0A8D0 , 32'hF82BBA48 , 32'h044A3BA0 , 32'h14478960 , 32'h01769D70 , 32'hF22DA950 , 32'hF11F7670 , 32'hECE5C720 , 32'h00049BA7 , 32'hDA0FA580 , 32'hEBAC3060 , 32'h0ED85A70 , 32'h170211A0 , 32'h07113B50 , 32'h023D2EA4 , 32'hFEABF12C , 32'hFF516E52 , 32'hF1623120 , 32'hDAECFFC0 , 32'h0EC67DF0 , 32'hF914B948 , 32'hF93AB540 , 32'hF65D6250 , 32'hF3C7F9D0 , 32'h07B4D848 , 32'h02818A64 , 32'h0214D9BC , 32'hF261BA60 , 32'hEB924F60 , 32'hFAFB1368 , 32'hEF8B52A0 , 32'h0A310F10 , 32'hFBFA2B58 , 32'h03CE4D18 , 32'hFC444004 , 32'hFA791C90 , 32'hF9951B20 , 32'hF913AE30 , 32'h02D8A6A4 , 32'hFF072849 , 32'hFFFD23BF , 32'h147AC240 , 32'hFC02452C , 32'hFE6610C8 , 32'h08CD3B20 , 32'h0D05C860 , 32'h037CDD58 , 32'h0BC7D020 , 32'h03B46754 , 32'hFBB763F0 , 32'h0BD716D0 , 32'hF4EB4A10 , 32'h00372E01 , 32'hF9072478 , 32'hFF4B6BB1 , 32'h0A2279E0 , 32'h05E63988 , 32'h00001A09 , 32'h13F0D2A0 , 32'hFB8834D0 , 32'h01B5BB9C , 32'h0CF9D0E0 , 32'h0BE3BC60 , 32'hFFFEC075 , 32'hFBEF4B98 , 32'h059C29F0 , 32'hEFE9F980 , 32'h1EEB7C80 , 32'h00050EA9 , 32'hECE25100 , 32'hFADCC100 , 32'h01C942CC , 32'h080D55F0 , 32'h069E7A38} , 
{32'hFAFD0FD0 , 32'hF69EC590 , 32'h16B54900 , 32'h00000FE4 , 32'hFFFFD290 , 32'h028D1EA8 , 32'h000680CC , 32'h12F658E0 , 32'h0001BABE , 32'hE32AA980 , 32'h18C89CA0 , 32'hEFF180A0 , 32'h2E932480 , 32'h05261968 , 32'h045CD1C0 , 32'hFE79B270 , 32'h13153E80 , 32'h01ABEFD8 , 32'hF1EEC830 , 32'hFFFC1053 , 32'h0E644250 , 32'h05D1DA68 , 32'hEA9DDDC0 , 32'hFFFDBB5B , 32'hEF9C0C60 , 32'hF8754C48 , 32'hEFA5C8E0 , 32'h0D73D290 , 32'hF3B7A5D0 , 32'hF92458C8 , 32'hF710E490 , 32'h23BD1780 , 32'hF8861B20 , 32'hE9633E40 , 32'hFFFDD300 , 32'hEA7896A0 , 32'h0CBC1370 , 32'h0D521100 , 32'h0D53F6D0 , 32'hED559440 , 32'h07813360 , 32'h01104AA8 , 32'h0063D031 , 32'h059A6FC0 , 32'hF8123310 , 32'hF2B7E6E0 , 32'h00DED66D , 32'h171B38A0 , 32'h01EB1894 , 32'hF00EB530 , 32'hF796E400 , 32'h08B492D0 , 32'hF7C08B90 , 32'hFE6724F4 , 32'hF9284390 , 32'h04B647A0 , 32'h1355BDE0 , 32'hF9D949C0 , 32'hF659B050 , 32'hF7D11D30 , 32'h0C2A85A0 , 32'hFDC2BC4C , 32'h00B78E02 , 32'hF77CB4D0 , 32'hEB843F80 , 32'h0EBC68C0 , 32'hFFFD2451 , 32'hFDE70330 , 32'h07806FE8 , 32'h06E70CF0 , 32'hFE558C80 , 32'hF8AF0C88 , 32'h040CE3E0 , 32'h084E6190 , 32'h12FD6400 , 32'hFB8A6340 , 32'h0098A02E , 32'hF614F830 , 32'h01F3A2C0 , 32'hFD8ADF14 , 32'hFB4EC630 , 32'hFB72D4B8 , 32'h1065C560 , 32'h0002B69F , 32'hED0CFD40 , 32'h02AFA064 , 32'h1B396320 , 32'hFD0F7424 , 32'hE9907840 , 32'hFFFAE636 , 32'hFDE15400 , 32'hFF89247D , 32'h05CD61F8 , 32'hF477E710 , 32'hFFFE8797 , 32'h014935EC , 32'h056238C0 , 32'hF45975D0 , 32'h13DFAC00 , 32'hFEC6BB1C} , 
{32'hEC307960 , 32'hF5043260 , 32'h06E59040 , 32'h000481FD , 32'h0001D1F7 , 32'h0EB37340 , 32'h0A7448A0 , 32'hF7C05320 , 32'h0000BEE4 , 32'h10A44F40 , 32'hE5EADF80 , 32'h09328320 , 32'hF5C326D0 , 32'h18B5C1A0 , 32'h06BFD218 , 32'h0E628050 , 32'hEAD4AE40 , 32'h14C8BB80 , 32'h081938E0 , 32'h0000D439 , 32'h0F510110 , 32'h128A2CE0 , 32'hF7869F80 , 32'hFFFED74C , 32'h0498A5D8 , 32'h02637C0C , 32'hF46E43C0 , 32'hFF9F1CAA , 32'hEE165B00 , 32'hDA8828C0 , 32'hF154D250 , 32'h19B4BCA0 , 32'h092CE140 , 32'hF05A3950 , 32'hFFFE594D , 32'h01DE7A14 , 32'h074D2048 , 32'hED218DA0 , 32'h02523DB4 , 32'h191F6FA0 , 32'hFE393700 , 32'hFEA1F710 , 32'h02955798 , 32'hF16B58C0 , 32'hFF5A19EB , 32'h10E83F20 , 32'h04459908 , 32'h0185D6C4 , 32'hF470B930 , 32'h06C77B00 , 32'h0D39AFB0 , 32'h026CFEC4 , 32'hEC993660 , 32'h1A64C0E0 , 32'hF13E4760 , 32'hFD021F58 , 32'h0A717720 , 32'hF4DAEFC0 , 32'hF8101060 , 32'h00E00724 , 32'hDAA2A500 , 32'hF7380630 , 32'hFAF6A8B8 , 32'hFE8BECC0 , 32'hEED3E920 , 32'hFC4772BC , 32'h00012D28 , 32'hF5932870 , 32'hFDCC25C0 , 32'h0671CB30 , 32'h05CF6990 , 32'h01CF2224 , 32'h003D4A28 , 32'hFECCFC58 , 32'hFF4FD1B0 , 32'hF9AC50B0 , 32'hF47B90C0 , 32'hED7556A0 , 32'h00B25494 , 32'h049A5D98 , 32'h01FBE1E4 , 32'hF0455BD0 , 32'h034EB358 , 32'h0005BDEF , 32'hFFAFED52 , 32'hECB60D40 , 32'hFFC19DAB , 32'h0B4063E0 , 32'hF53275B0 , 32'hFFFF27FD , 32'hFCB32518 , 32'hF804CB38 , 32'hE41507A0 , 32'hF7E0D360 , 32'h0003DC0F , 32'hF1ACA3C0 , 32'h03EE04A0 , 32'h11FD59C0 , 32'hFC49719C , 32'hE8407E60} , 
{32'h03B796DC , 32'h04BD5C50 , 32'h180EE340 , 32'hFFFD231E , 32'hFFFAD83B , 32'h06E7E228 , 32'h11A85F20 , 32'hEEF7E8E0 , 32'h00002DCA , 32'h02492C04 , 32'h110A39C0 , 32'h04948070 , 32'hF79493F0 , 32'h09B5E110 , 32'h0DDB7960 , 32'hED0BEB00 , 32'hFFC516EC , 32'hFE318D9C , 32'h07C46780 , 32'h000005B8 , 32'h029CB068 , 32'hE66E4300 , 32'hFF23AAC9 , 32'h0001A2FD , 32'hF1C6CBA0 , 32'hF1A6F580 , 32'hFE5CFB9C , 32'hFD6C563C , 32'h00E74A40 , 32'hED2DC440 , 32'hF6BA9C60 , 32'h10405300 , 32'h12122580 , 32'h0C361480 , 32'hFFFE7040 , 32'hF7232EA0 , 32'hF5236CF0 , 32'hF9557610 , 32'hF7680D60 , 32'hEBDEC420 , 32'h08FF6090 , 32'hFE8BE8C0 , 32'h0AE31A30 , 32'hEBA7D900 , 32'h00F5B667 , 32'hFA74CF48 , 32'hF7171950 , 32'hF35FCC20 , 32'hFE36DD04 , 32'h191A38E0 , 32'h0B6318C0 , 32'h0083FCA4 , 32'hF0379930 , 32'hF47663E0 , 32'h1D461B80 , 32'hF8AD4508 , 32'hFE441684 , 32'h132B48C0 , 32'hF9367F20 , 32'hED18C220 , 32'h04FC2EB8 , 32'hF8ED26E0 , 32'hFFF745E7 , 32'h072BB7A8 , 32'h1C6D6140 , 32'hFBC48070 , 32'h0004FA56 , 32'hFC0124CC , 32'hF684B890 , 32'hF02CD7A0 , 32'h0DD21120 , 32'h0204BC98 , 32'hF34AF9B0 , 32'hDD504180 , 32'h0E211790 , 32'h001ABDED , 32'hFF1220CE , 32'hE8F14540 , 32'hF6DF5380 , 32'h17BDE800 , 32'h15851040 , 32'hF35715D0 , 32'h13D47760 , 32'hFFFF884A , 32'hF36469B0 , 32'hFFD78BDC , 32'h19D51AE0 , 32'hEA433A60 , 32'h123A4560 , 32'hFFFFCA30 , 32'h08D60820 , 32'h017C9B5C , 32'h10E90200 , 32'h098F2F90 , 32'hFFFF0A67 , 32'hF6E74360 , 32'h04ED6080 , 32'h02F4D180 , 32'hF5653090 , 32'hFC98A454} , 
{32'h0E254D20 , 32'h07319EB0 , 32'hF6635DA0 , 32'hFFFED0E3 , 32'hFFFF1081 , 32'h058F51E0 , 32'h04485478 , 32'hFC9F7570 , 32'h0002DB5D , 32'h05C6BA10 , 32'hF6A29E40 , 32'h15CE6F60 , 32'hFDA19988 , 32'hFAE6C968 , 32'h12B851A0 , 32'h0BD4D7B0 , 32'hF566DB10 , 32'h0744CBB0 , 32'hF7615860 , 32'hFFFC8ADA , 32'h11832B80 , 32'h1DA90780 , 32'h0BFE8820 , 32'h0001309A , 32'hE19C5B00 , 32'hEBCCC5C0 , 32'h07DADBF8 , 32'h07086AC8 , 32'hE0D05C20 , 32'hF21E1C30 , 32'hEEFC0280 , 32'hF994F888 , 32'hF285FE40 , 32'hED474720 , 32'hFFFE0D87 , 32'hF4E76830 , 32'hFF642C31 , 32'hF6C01D90 , 32'hF9BD8D60 , 32'h08F911F0 , 32'h1F919920 , 32'hFDAD8CD4 , 32'hF1A59380 , 32'h04EB66D8 , 32'hFB8E6468 , 32'hF166B9E0 , 32'h0369F410 , 32'hEE489760 , 32'h171D93C0 , 32'h05E2CFF8 , 32'h0CFECCC0 , 32'h09F64DE0 , 32'hFEBF8A50 , 32'h09DFA990 , 32'h13577640 , 32'h0B851250 , 32'h01F4FF8C , 32'h0D3CE4D0 , 32'h00D4AC2C , 32'hF74D3E50 , 32'h12F10640 , 32'hEDCFC0E0 , 32'hE73324E0 , 32'h081A79A0 , 32'hFE2AD0D8 , 32'h0A204E40 , 32'hFFFE6BEF , 32'h1729E120 , 32'hFD1C58C0 , 32'hF6B2F790 , 32'hEE0107C0 , 32'h0359F398 , 32'hF4ABB150 , 32'hFB2BD5E8 , 32'hFDFCC264 , 32'hF77BC3D0 , 32'hEF15ECA0 , 32'h0A122250 , 32'hF6764110 , 32'hFB616790 , 32'hE82A5020 , 32'h11109320 , 32'hF4EFA360 , 32'hFFFE42E6 , 32'h01716AEC , 32'h18588900 , 32'hF9B3C5C0 , 32'hFA31C0C0 , 32'hFB9C31C8 , 32'hFFFCABB6 , 32'h173656E0 , 32'h01945014 , 32'hFF66872E , 32'hF2895570 , 32'hFFFF9423 , 32'h10DFB400 , 32'hF82C8218 , 32'hF9FC2DC0 , 32'hF4E3F7A0 , 32'h0E1C2DE0} , 
{32'hF85BAEE0 , 32'hFC87B668 , 32'hFBC38768 , 32'hFFFDC77D , 32'h00042508 , 32'h08BF1140 , 32'hF539E990 , 32'h00EF0D5B , 32'hFFFE6166 , 32'hF3E4DD50 , 32'h10228F40 , 32'hFD095E94 , 32'hF6DDF2D0 , 32'h1A50D400 , 32'h02671580 , 32'h023DFD24 , 32'hF8C3CA30 , 32'h0132D3FC , 32'h021B7E60 , 32'h00065D31 , 32'h017E6D14 , 32'hF25C8460 , 32'h1E53E9A0 , 32'h0001038F , 32'hEE5072E0 , 32'h1D84AE00 , 32'hFB0F7660 , 32'h03654E80 , 32'h12B2F7E0 , 32'hF0D25E70 , 32'h0E282D00 , 32'h07F52930 , 32'h11A655C0 , 32'h098CE3F0 , 32'hFFFD5B0A , 32'h0A3960F0 , 32'h04639870 , 32'hF2DD7C70 , 32'hF3734110 , 32'hE53D75A0 , 32'h2582AB00 , 32'h00037A86 , 32'hF8ECFA68 , 32'h006083FE , 32'hF49B5BD0 , 32'h02DFD460 , 32'h11FEE920 , 32'h10A47840 , 32'hEA2EBD20 , 32'hF2B2E460 , 32'h197C2720 , 32'h04665040 , 32'h0E521130 , 32'hE4156340 , 32'hF18F4CB0 , 32'hF2F7F450 , 32'h08492960 , 32'h00D82380 , 32'hF2F34110 , 32'hFA43E218 , 32'hFDC7AC5C , 32'h02D0C200 , 32'hF3BA6EE0 , 32'h01B5FCA4 , 32'h0E078950 , 32'h057F2E98 , 32'hFFFE7E38 , 32'hF9E0A4E0 , 32'hFA026B30 , 32'h0047A083 , 32'hF1A9CD00 , 32'h02BDD82C , 32'hFCA32170 , 32'h0DE27400 , 32'h107C37A0 , 32'hEB5896C0 , 32'hF2256610 , 32'h05275E88 , 32'h12868880 , 32'hE6821BE0 , 32'hFF5879B0 , 32'hFA7F3CB0 , 32'hF57CEDD0 , 32'hFFFDFED1 , 32'h0E879510 , 32'h14FD1940 , 32'hECCDB440 , 32'h0100D078 , 32'hFD3B2924 , 32'h00006FE0 , 32'h113F86C0 , 32'hFAC2D9A0 , 32'hFD481388 , 32'hFA884EF0 , 32'hFFFCB173 , 32'hE7CB6FE0 , 32'hF12814F0 , 32'hFD162FC8 , 32'h03F28F50 , 32'hF8BBAA80} , 
{32'hFD00726C , 32'h0E987220 , 32'h119C2D40 , 32'hFFFEAB64 , 32'h0000194C , 32'h000285DA , 32'hFFA64FCD , 32'h0AC5B580 , 32'h000291DD , 32'hF5BFCE50 , 32'hF80C21F8 , 32'hF4ABC910 , 32'h1238FD60 , 32'h10F5F8A0 , 32'hFDD9EC84 , 32'h05D04B20 , 32'h12AC4380 , 32'hF37BC2F0 , 32'h035E2DD0 , 32'hFFFFE297 , 32'h13BB7C60 , 32'hF35B3290 , 32'hFF7B29DD , 32'hFFFF9425 , 32'hEDF129E0 , 32'h072D39E8 , 32'h06328D60 , 32'hFCDF5BA4 , 32'hEF117340 , 32'hF7A429A0 , 32'h010D4FCC , 32'hF142A980 , 32'h011CCAE0 , 32'h0B397C30 , 32'hFFFF1831 , 32'h001BD42C , 32'h07C07FE8 , 32'h151134C0 , 32'hF021D9B0 , 32'h08A48B80 , 32'hF2999F30 , 32'hFF095C7A , 32'hFE88311C , 32'hF62175A0 , 32'hFF356FB5 , 32'h041CAD88 , 32'h26373400 , 32'hE55DBF80 , 32'h06F9AD20 , 32'hFC73593C , 32'h10062BE0 , 32'hF1EC6D80 , 32'hF349DB80 , 32'h0568F4C8 , 32'h0346E3B4 , 32'hEFCF8C20 , 32'h0C89AC60 , 32'h1C3BC6E0 , 32'hF5EABB80 , 32'hFF64D07C , 32'hEC1B4E20 , 32'hEBCEDA60 , 32'h164285E0 , 32'hF8E5C9F8 , 32'hFA889750 , 32'h0235AD60 , 32'h00022343 , 32'hF421A100 , 32'hF810B6A0 , 32'hFD3FDA78 , 32'h13B45400 , 32'hF2FE3700 , 32'h1497A3C0 , 32'h002544C8 , 32'h0C05A4D0 , 32'h02F23230 , 32'h049F02C0 , 32'h0052F335 , 32'h051891F8 , 32'h01926B18 , 32'h0322289C , 32'hFD9C6C54 , 32'hF3254B60 , 32'h0001A2ED , 32'h09DE8320 , 32'h0E9B9EF0 , 32'hDAAE9C80 , 32'h06251E30 , 32'hF2CE9350 , 32'h00019015 , 32'hFDEBFE30 , 32'h075BDDA8 , 32'h0EC70E50 , 32'h1793F140 , 32'h0002F2FD , 32'h29F49440 , 32'h01E5FA40 , 32'h05FD4580 , 32'hFFD06EA3 , 32'hFCEF244C} , 
{32'hE50E8040 , 32'hF9DE8BA0 , 32'h0600BF68 , 32'h00003014 , 32'hFFFBF94B , 32'h0E3C7BB0 , 32'hF8E13608 , 32'h0BC1A3A0 , 32'h00069063 , 32'hF7C01720 , 32'h01818E18 , 32'h03B9B500 , 32'h045D9038 , 32'hF4B30970 , 32'h037ED070 , 32'hE6AC97C0 , 32'h06B81C10 , 32'h010964B8 , 32'hF7CFAD20 , 32'hFFFEA673 , 32'h0C7EE8B0 , 32'hE6E7F180 , 32'h107CBB20 , 32'h00002840 , 32'h0D281E20 , 32'h024A1688 , 32'hFCEFFC48 , 32'hEC08F160 , 32'hF3390260 , 32'hF94545E0 , 32'h01DCEEDC , 32'hFDD05474 , 32'hF93C7EC0 , 32'hED67D0C0 , 32'h00032E89 , 32'h01771018 , 32'h008C777F , 32'hE7868600 , 32'h24774240 , 32'h0540F538 , 32'hEAD9FF00 , 32'h0099FE8C , 32'hF5073880 , 32'hF636D790 , 32'hF7A2E400 , 32'hDA710C40 , 32'hF2442430 , 32'hF8CF5C70 , 32'h0B01D190 , 32'h04986330 , 32'h0F6B7480 , 32'hFA350040 , 32'h095797F0 , 32'h0A24ACA0 , 32'hF00D0790 , 32'hF2D50C70 , 32'hFE0314D0 , 32'hF295F9C0 , 32'h07953880 , 32'h0B363DD0 , 32'h0A0CBA80 , 32'hFD7B6708 , 32'hFC0BF9F0 , 32'hF7BEAFB0 , 32'h0D98D980 , 32'h0DBFD570 , 32'hFFFC2A32 , 32'hFDBCEADC , 32'hF4E667A0 , 32'hF07E5B70 , 32'h0C036DB0 , 32'h07E05A40 , 32'h0542A350 , 32'h027082A0 , 32'hF5D94BF0 , 32'hF6C3BA30 , 32'hF9583C20 , 32'h0243123C , 32'h09BFFE80 , 32'h22888300 , 32'hEB39F8A0 , 32'hEDB0FC20 , 32'hFF049AE9 , 32'hFFFD74E0 , 32'h0FED8D10 , 32'h171C6980 , 32'hEF85BDE0 , 32'hEFB6DEE0 , 32'h0ECE6380 , 32'hFFFDCDC2 , 32'hFAD6EC70 , 32'h0232F498 , 32'hE9B53E40 , 32'h0C53C930 , 32'h00025A17 , 32'hFBD1E660 , 32'hFC5A9638 , 32'hEA05B540 , 32'h0FED8700 , 32'hFD44F00C} , 
{32'h124F8860 , 32'hFE569B8C , 32'hFA442E28 , 32'h000655E1 , 32'hFFFF575C , 32'h14AAB100 , 32'h02359E44 , 32'h05E1D0D8 , 32'h00049F14 , 32'h097B0970 , 32'hFE4188E8 , 32'hE88B52E0 , 32'h10440E40 , 32'h0ECD5FC0 , 32'hF840E750 , 32'hECF14EE0 , 32'hE345D3A0 , 32'h14128620 , 32'h12642200 , 32'h000218AB , 32'hF6FFE870 , 32'h1B3C7DE0 , 32'hFB9AF388 , 32'hFFFB07FE , 32'hF1FC72F0 , 32'hD9EF4780 , 32'hEEC57CE0 , 32'hED2ECDC0 , 32'h166DE120 , 32'hFD3D6CFC , 32'h01E8D938 , 32'h070F2B00 , 32'hF493F110 , 32'h07C61298 , 32'h0000811B , 32'h03DEC5F0 , 32'h032EB5F8 , 32'h00812DF4 , 32'h01619E54 , 32'hF32897F0 , 32'hFD2369A4 , 32'h01AD5A9C , 32'hFF449589 , 32'hEF29F1C0 , 32'h0A5495D0 , 32'hEDAA4200 , 32'h04C10D00 , 32'h09BF5DB0 , 32'h14BD21C0 , 32'hF8EA16F8 , 32'h14D005C0 , 32'h0600EF88 , 32'h135B2EC0 , 32'hFE2BB6C4 , 32'h017C7064 , 32'h02F2F240 , 32'hEF03E8A0 , 32'hED27EFA0 , 32'hFCACE270 , 32'hF47E7080 , 32'hF425E8D0 , 32'h19B23840 , 32'h0A44CFA0 , 32'h05499F60 , 32'hF7F54940 , 32'h01F3B5A8 , 32'hFFFEF2A5 , 32'hEA6E5CE0 , 32'hFBD64FD0 , 32'h1AED42A0 , 32'h0721D9B8 , 32'h0CEC8500 , 32'h02BD9770 , 32'hF16D3260 , 32'hF81678E0 , 32'hF347AD80 , 32'h07381B48 , 32'h04858280 , 32'hEDDD9560 , 32'hFC2225EC , 32'hF4D02560 , 32'hFDE63058 , 32'h0077DA62 , 32'h00035D9F , 32'h06A19408 , 32'h0A1EA930 , 32'hEF7C7080 , 32'h08B0A0C0 , 32'h1605DEA0 , 32'hFFFF7813 , 32'h09E49EA0 , 32'h0379203C , 32'h1427A200 , 32'h05618EE0 , 32'h000830A3 , 32'h11EE4300 , 32'h0924BFC0 , 32'h06484C28 , 32'h0D072490 , 32'hF78EFAB0} , 
{32'h01218458 , 32'hFE806A30 , 32'h13540600 , 32'hFFF9D1B8 , 32'hFFFC9B4C , 32'h0527B530 , 32'h15995380 , 32'hD80D2E80 , 32'hFFFF6D2A , 32'h0724F568 , 32'h0A0ACEE0 , 32'h0F2A0B50 , 32'h01060D10 , 32'h068735D8 , 32'hDE7AE440 , 32'h0FDC0F00 , 32'h06DD1AF8 , 32'hDFE03080 , 32'hF5773420 , 32'h0001F72E , 32'h0896C600 , 32'hF6C8DA90 , 32'h117F4BA0 , 32'hFFFDC7BF , 32'h0AB93000 , 32'hEF574A80 , 32'hFF3C53F3 , 32'hF409D280 , 32'h0FF78EC0 , 32'h0331F12C , 32'hF38711A0 , 32'h09FAADD0 , 32'h030BCF28 , 32'hFD1F4EB4 , 32'hFFFB838B , 32'h00977D48 , 32'h00B81F22 , 32'hFC1F1340 , 32'hEB579DE0 , 32'h11ABECC0 , 32'hFFCDB88C , 32'hFFFF7BC1 , 32'hF5AC6820 , 32'h047F4C78 , 32'h19ABDEC0 , 32'hF2FF2910 , 32'h016E2F78 , 32'h1CDA1B40 , 32'h01A03B80 , 32'hFBC133D8 , 32'h030A2140 , 32'hFA11AE08 , 32'h0BAAF6F0 , 32'hED302240 , 32'h0070142F , 32'h0BB27470 , 32'hEDBA1AA0 , 32'h19407240 , 32'h03519D1C , 32'h162AE7E0 , 32'hEC04D3E0 , 32'hFDBC280C , 32'hF5B04E50 , 32'hF93BC118 , 32'hE6C561E0 , 32'h009C5C05 , 32'h00000D8F , 32'hFA8C9538 , 32'hFF1B98D8 , 32'hF958C9A0 , 32'h0ACC47C0 , 32'h07819DB8 , 32'h02607B4C , 32'h0EDA8E20 , 32'h04296D08 , 32'h00230FB5 , 32'hEA5EE300 , 32'hFC7D31C4 , 32'hF5E61E50 , 32'hF8A518C8 , 32'hEC871460 , 32'h024364CC , 32'h1753BCE0 , 32'hFFFEB982 , 32'hF7C62C10 , 32'h1BC7FD40 , 32'h0B624EF0 , 32'h029C0924 , 32'h031AF06C , 32'hFFFFC6D9 , 32'hF5B95C60 , 32'h06C79868 , 32'hF09F91C0 , 32'h09C81450 , 32'h0000D421 , 32'h069C7250 , 32'h03F0D6A0 , 32'h03999B28 , 32'h07319970 , 32'h0A07DE80} , 
{32'hFB198DE8 , 32'hED662F40 , 32'hF8BABA10 , 32'h00037820 , 32'hFFFF9F33 , 32'hFC79B5CC , 32'hE5DB0660 , 32'hF6EF14F0 , 32'hFFFEA7C0 , 32'hFCCE0B70 , 32'hF54D0500 , 32'h07639720 , 32'hFBCAD9F8 , 32'hEBA9F040 , 32'hF2FC1E60 , 32'h1DB5A540 , 32'h03DC31E8 , 32'h133767C0 , 32'hF27D0D00 , 32'hFFFB1296 , 32'h0A116D20 , 32'hF14DB080 , 32'hF0822EA0 , 32'h000407E6 , 32'hF32A6640 , 32'hF357F670 , 32'h0E6A78D0 , 32'h133ABBC0 , 32'h1FAF34C0 , 32'h001E1282 , 32'h04DF3C80 , 32'h14EFEA00 , 32'hF71A8380 , 32'hF96D2100 , 32'h0004397C , 32'h1FFAA880 , 32'hE2F45F20 , 32'h07C2C3A0 , 32'h16BA53C0 , 32'h10CA9E60 , 32'hFC6BB428 , 32'hFFAE3B56 , 32'hF9D25968 , 32'hF4823170 , 32'hEC4ABD00 , 32'h11C11660 , 32'h013947D4 , 32'h0AB2A340 , 32'h07B813A0 , 32'hF558FA60 , 32'h1BAF9E40 , 32'h0C17F150 , 32'hFDB04E40 , 32'hFF057435 , 32'hF2AC5C50 , 32'h14A4A6A0 , 32'h08CC7530 , 32'h0ECC0D90 , 32'h11E9AA00 , 32'hFBEBE390 , 32'h1299AC60 , 32'hF126C990 , 32'hFF682EB9 , 32'h1364B7E0 , 32'h07221FD0 , 32'hF4FBEEA0 , 32'hFFFFEEAA , 32'hED09F960 , 32'hF9759628 , 32'hFD6ADE98 , 32'hFFF0BC56 , 32'hFCFDDCA8 , 32'h0224F3BC , 32'h092C7B60 , 32'h12A282E0 , 32'h02363E6C , 32'hF96B8428 , 32'hEE539DC0 , 32'hF0196D10 , 32'h006E9550 , 32'hF96A4650 , 32'hF3215860 , 32'h0069D2F3 , 32'hFFFB4B05 , 32'hFEE8C45C , 32'hF63EA7E0 , 32'hF92525B8 , 32'hFBEA2EB8 , 32'h0AF591D0 , 32'h00043616 , 32'h0946E700 , 32'h0586D7E0 , 32'h10AFF360 , 32'h12E1A0A0 , 32'h0005B390 , 32'h07C23CB0 , 32'h0A7064D0 , 32'hF5E3CC70 , 32'hFC340AC0 , 32'h01F93288} , 
{32'hED947580 , 32'hF52449B0 , 32'hF2083F80 , 32'h00029723 , 32'hFFFD3438 , 32'hF709A230 , 32'hFCD58640 , 32'hE4A72B40 , 32'h00033D8D , 32'h05F2D1B8 , 32'h03DAC7A8 , 32'h00F84F01 , 32'hFEB3BE54 , 32'hF8BF9D58 , 32'h0A279530 , 32'h0269F3A0 , 32'h08F99920 , 32'hF96AEBC0 , 32'h0594B028 , 32'h0003369F , 32'hF806F9F8 , 32'h089BF8E0 , 32'hF0A2EE40 , 32'h0000BAD3 , 32'h003304EE , 32'hFDBEBC68 , 32'h03CCCC1C , 32'h079DED80 , 32'hF95D9C38 , 32'hE3944080 , 32'h0CC95070 , 32'h19F35AC0 , 32'hF8D5B600 , 32'hE8345240 , 32'hFFFF78B1 , 32'h102E3980 , 32'h09CD12C0 , 32'hFD170F0C , 32'h0C63A880 , 32'hE1B9BF40 , 32'hE6938E60 , 32'hFF981D5B , 32'hFDA8EDA8 , 32'hFF0583C3 , 32'h07375BD0 , 32'h12A8BF80 , 32'hF0A8F220 , 32'hE0757D00 , 32'h0211AF50 , 32'hF9BA09C0 , 32'h04C61070 , 32'hFAA62A30 , 32'hF97A5C20 , 32'hE03E95E0 , 32'h0D3CE8F0 , 32'hF233FF80 , 32'h00199BE5 , 32'h00FD72F3 , 32'h0F1B2230 , 32'h1A7A0A00 , 32'h0D647920 , 32'hFD1305C0 , 32'h10BA4980 , 32'hECFBD320 , 32'hFF20238D , 32'hF509B510 , 32'h0002DF66 , 32'h075CFFB0 , 32'hFF000A20 , 32'h04EA5440 , 32'hE9F41F60 , 32'h0F48C650 , 32'h1339C560 , 32'hEEAF99E0 , 32'hFEC0F3E8 , 32'hFCF33A1C , 32'h04F80060 , 32'h0A7CEFF0 , 32'h029F36DC , 32'hF3329470 , 32'h027493D0 , 32'h0625C4D0 , 32'h0EDA1560 , 32'hFFFAF796 , 32'h09ECA560 , 32'h2502B8C0 , 32'hFF4E6CF4 , 32'h1A4278A0 , 32'hFE4E3B40 , 32'hFFFED865 , 32'h007C0CC7 , 32'h07E04688 , 32'h0392B088 , 32'hF74CE570 , 32'hFFFFD8E8 , 32'h01E85AC4 , 32'h06F5D098 , 32'h159451C0 , 32'hFD3DD7AC , 32'hFA340150} , 
{32'h035DB1C0 , 32'h0753CA68 , 32'hE3C82EC0 , 32'h00010C5A , 32'h0008E123 , 32'hF630CEE0 , 32'h06999AA8 , 32'hF5A93D70 , 32'h0000CB96 , 32'hE7B34BC0 , 32'hFFE6F2A9 , 32'hF56638D0 , 32'hFA9739C0 , 32'hEADA11E0 , 32'h00785819 , 32'hF692DE40 , 32'h060E7100 , 32'hF670E6B0 , 32'hFF7622EA , 32'h00044759 , 32'h1B4C7440 , 32'hFED7B88C , 32'h17120F40 , 32'hFFFCF826 , 32'hF01B6760 , 32'hFB51C158 , 32'hECA7B3A0 , 32'hF448A550 , 32'hF8A6ED28 , 32'hF8BBBBC8 , 32'hFFDB4855 , 32'h03110544 , 32'h08E6F310 , 32'h01696A24 , 32'hFFFF3F54 , 32'h011161AC , 32'hFD237C14 , 32'h0262EEF0 , 32'h1465BEE0 , 32'h0AC94B10 , 32'h05DB0C48 , 32'hFFBA66BD , 32'hFDDA012C , 32'hFDBD3A70 , 32'h0A1E1F10 , 32'hE90829A0 , 32'h0B643270 , 32'hF7049ED0 , 32'hF8BA5BB0 , 32'h17EC9AA0 , 32'hF48EF4D0 , 32'h06A847D8 , 32'h00DF1C6A , 32'hF2ADEDC0 , 32'h0556A8C0 , 32'h021AEC30 , 32'hFDB0A91C , 32'h17377F40 , 32'h10D42E00 , 32'hEE360A40 , 32'h14045060 , 32'h1670E1E0 , 32'h0042D57E , 32'hFB2D5830 , 32'hF2D5E720 , 32'hE1881420 , 32'hFFFD782A , 32'hF2EEADC0 , 32'h072EC048 , 32'hF98F0AB0 , 32'hF9442200 , 32'h048703E8 , 32'hF759A8B0 , 32'h063102F8 , 32'hFDDE4E70 , 32'h00F5BE3D , 32'hFC976630 , 32'h0C351930 , 32'hF65B8E00 , 32'hF3982CA0 , 32'h094CFEF0 , 32'hEB1C3980 , 32'h129F09A0 , 32'h0001A452 , 32'h05460C68 , 32'hD91D6980 , 32'hF6320930 , 32'h16F53660 , 32'hF058C1F0 , 32'hFFFFCE74 , 32'h0581E348 , 32'h020F7AEC , 32'hF28DEDA0 , 32'h032B40C0 , 32'h00002B37 , 32'h09CEFBC0 , 32'hED1EEBA0 , 32'h08387600 , 32'h116C53E0 , 32'hDF179380} , 
{32'h00DE8C8B , 32'hF2E36880 , 32'h0DF82140 , 32'hFFFEE8B8 , 32'hFFFE336D , 32'hE293BC40 , 32'h1CF67660 , 32'h04ECC2D8 , 32'h00049F3A , 32'h0697F8C8 , 32'hF3E52510 , 32'h03A14F54 , 32'hF30CA500 , 32'hF2EE6640 , 32'hF46C4170 , 32'hFEF97344 , 32'h01229360 , 32'h03FBB2A4 , 32'h05549DC8 , 32'hFFFE33C9 , 32'hE3953C20 , 32'hF9484078 , 32'h0051A169 , 32'h0001F58F , 32'h0102168C , 32'h0B6D2CF0 , 32'h114D9F80 , 32'hF9242CF0 , 32'h04C7CA70 , 32'h090DF690 , 32'h18D7BAA0 , 32'h06278490 , 32'hE32223C0 , 32'hF27362D0 , 32'h000437B4 , 32'hED934280 , 32'h07F363B8 , 32'hF3EF38E0 , 32'hF65C6A30 , 32'h06DF8D78 , 32'hF98D7520 , 32'hFF3C3141 , 32'hEE846B60 , 32'hFC312C14 , 32'h024FFC1C , 32'hE18A2F40 , 32'h044A2FD8 , 32'hF0FFF2D0 , 32'h00ADC678 , 32'h0A4C27D0 , 32'h13960900 , 32'hF7B2DC20 , 32'h02422348 , 32'hFE9D51E4 , 32'h0237529C , 32'h04460188 , 32'h153F0900 , 32'h0A141410 , 32'h00173576 , 32'hF93A32F0 , 32'h01DA87E8 , 32'h055F6918 , 32'h12336380 , 32'h10E2F320 , 32'hE99B8340 , 32'h0CD6C880 , 32'hFFFE1821 , 32'hF5A640D0 , 32'h08B0B850 , 32'hFFCA8A1B , 32'h07A4B770 , 32'hFCB51558 , 32'hFE887248 , 32'h04CBC8C0 , 32'h1EADFE60 , 32'hFBD79310 , 32'h0DFA7BA0 , 32'h08BA78B0 , 32'hF19E7C60 , 32'hFE4922B8 , 32'h12220760 , 32'hFB38ADD0 , 32'hE95C8F20 , 32'hFFFE2703 , 32'hE478D160 , 32'h06EAB2D8 , 32'hFD55BD30 , 32'h0BE15CC0 , 32'hFFE442FC , 32'h0000C2D3 , 32'h2217B1C0 , 32'h012C41C8 , 32'hF35D4BA0 , 32'hF1836770 , 32'h00007FE6 , 32'hE656E3C0 , 32'h0A977290 , 32'hFECA2054 , 32'h06421908 , 32'hF55E8180} , 
{32'h02C3BCC8 , 32'hF9B1D250 , 32'h0CD28890 , 32'hFFFDABA1 , 32'hFFFCFA84 , 32'hFBB783E8 , 32'h04A87BA8 , 32'hFFB7638E , 32'h00018CD1 , 32'h13B94540 , 32'hFD547770 , 32'hFA8E2FB8 , 32'hED239080 , 32'hFE90A224 , 32'h09C04A60 , 32'hE0D375A0 , 32'h1892CE80 , 32'hFE24AE38 , 32'h049D3950 , 32'h000025A6 , 32'h0970B690 , 32'hF46260F0 , 32'hEF8FEF60 , 32'h000173DB , 32'hE47DC6A0 , 32'hF7DB5610 , 32'h09004D50 , 32'h10F11A00 , 32'hF13941E0 , 32'hFF43B69E , 32'hEFE97A40 , 32'hEE784400 , 32'h015EB6E8 , 32'h09D8F960 , 32'h00006B7C , 32'h0DA95740 , 32'hF5F37B20 , 32'hF9F30440 , 32'h0C5029F0 , 32'hFB18C140 , 32'h027708E8 , 32'h0174C4C0 , 32'h0B2A9C40 , 32'h0A57D440 , 32'h0C360150 , 32'hF60879A0 , 32'hF9871BF0 , 32'h0EC868B0 , 32'h0FA6E7A0 , 32'hEC1372A0 , 32'hFB61B700 , 32'hFD64EB04 , 32'hEF7D01E0 , 32'hFF09357B , 32'hFE472648 , 32'hF9C2DEB0 , 32'hFA647150 , 32'hF6FA3E70 , 32'hF24D9E10 , 32'h098FCFA0 , 32'h063827C0 , 32'hFA4C0AF8 , 32'hED292320 , 32'hFA039780 , 32'hFB3493A0 , 32'hFDCAA36C , 32'hFFFDFE00 , 32'hD7D5A540 , 32'hF600FA20 , 32'h0D78B9C0 , 32'h0C695640 , 32'hFC154FB0 , 32'h0316DEB0 , 32'h0FC4CCB0 , 32'h0FC52B20 , 32'h17E8CA40 , 32'hFD17BA0C , 32'h1F241900 , 32'h09142C50 , 32'hF0488010 , 32'hF2F55550 , 32'h0A309CA0 , 32'hEECE51C0 , 32'hFFFF03DB , 32'h1606C1C0 , 32'hF98F7DC8 , 32'h1AA88FC0 , 32'h07F98F90 , 32'h0B49CF30 , 32'hFFFF2C9B , 32'h15BA3320 , 32'h07DD1640 , 32'hEEA16EA0 , 32'h092986D0 , 32'hFFFA7831 , 32'hF68D6CA0 , 32'h09686590 , 32'h0FECCD30 , 32'hF0F5A1E0 , 32'hF19412F0} , 
{32'h015447B4 , 32'hFE9733F8 , 32'hFFD0C41F , 32'hFFFF8BDD , 32'hFFF7EF18 , 32'hEE9E9B80 , 32'hE47ECF20 , 32'hFED62448 , 32'h0003524A , 32'hF57A6240 , 32'hE48071A0 , 32'hC773A740 , 32'h0B5C4A80 , 32'h09424170 , 32'h0B2C5A70 , 32'hEFEB71A0 , 32'hFE54823C , 32'hFFE9D20D , 32'hF34BBCC0 , 32'h000007C8 , 32'h0D46E670 , 32'hFC499BE8 , 32'hFB9EB170 , 32'hFFFC476C , 32'hFD38EA1C , 32'hEF4B8660 , 32'hF9C34CE8 , 32'hF69D3B20 , 32'h07BFD0C8 , 32'h11597D20 , 32'hF4BB4A70 , 32'hF8FCEC18 , 32'hF5CCE7F0 , 32'h077C2230 , 32'hFFFBC3A0 , 32'h0CC10FA0 , 32'h09B284C0 , 32'hE7E73C20 , 32'hE5671300 , 32'h0A97E2B0 , 32'hEDBB8C80 , 32'h00D0CAB5 , 32'h021FE2F4 , 32'hFF0B835D , 32'h06940528 , 32'h0541E530 , 32'hF71168F0 , 32'hFD6C0F24 , 32'hFA593630 , 32'h0BCDC930 , 32'h0430B2D8 , 32'h0FBDC9A0 , 32'hFB825508 , 32'hEBE3AEA0 , 32'h000327B5 , 32'hF6E0E260 , 32'h09F25250 , 32'h0A6AC170 , 32'hF1595C40 , 32'hFAA92378 , 32'h009CA2AD , 32'hED16EB60 , 32'hF6782790 , 32'h0F2C2BB0 , 32'hF5BD7370 , 32'hF900F590 , 32'hFFFC1608 , 32'h161B77C0 , 32'h002DA72A , 32'h03E499E4 , 32'hE7DD1440 , 32'hF6AC2120 , 32'hF8E7E4A8 , 32'h09167880 , 32'hF75D1240 , 32'h008A0531 , 32'h03670070 , 32'h06F0AC78 , 32'hE6AF3280 , 32'h066EA020 , 32'hF8246CB8 , 32'hEB116900 , 32'hFF84E479 , 32'hFFFE7E4E , 32'hFD28D810 , 32'h1482BA60 , 32'h056A5A18 , 32'hF8FB1A20 , 32'hF46BAAD0 , 32'h00018D99 , 32'hF552E500 , 32'hFD478CD8 , 32'hF4E26AA0 , 32'h0E155220 , 32'hFFFEF364 , 32'hE16F84A0 , 32'h07C42F20 , 32'h05BBF9A8 , 32'hEE19DF20 , 32'h005806E2} , 
{32'h0445C680 , 32'h16D91B00 , 32'hF111E580 , 32'h00000A54 , 32'hFFFC53CF , 32'h1037C840 , 32'h22FD6580 , 32'h042E1B48 , 32'hFFFC7F00 , 32'hF1862560 , 32'h035208F4 , 32'h08716CE0 , 32'hFE4A7A10 , 32'hFCB95AD8 , 32'hF875AB70 , 32'hFDD6BA0C , 32'hF9EF18A8 , 32'h06C81790 , 32'hE59EF680 , 32'h0008AE5D , 32'h17E831A0 , 32'h0E64D0E0 , 32'h072BC938 , 32'h00073D72 , 32'h0D7D9140 , 32'h094B2D50 , 32'h0CA1EC20 , 32'hF3DC6190 , 32'h172B12E0 , 32'h0DB797C0 , 32'hFB2107B0 , 32'h028B3954 , 32'h0B249AC0 , 32'h0087D8DE , 32'hFFFF8FF3 , 32'h0F3DBC60 , 32'h03360864 , 32'hF70CD920 , 32'h13629EE0 , 32'hED612BA0 , 32'hE46CBD40 , 32'hFDD12494 , 32'h0E0F8F00 , 32'h0002CE45 , 32'hE3BD2580 , 32'h00675A18 , 32'hFEB7E2BC , 32'hF6690B70 , 32'hECF2A3C0 , 32'h0B6D3E40 , 32'hF6A28530 , 32'h0849C070 , 32'hE4CC2F40 , 32'hFE728180 , 32'hF460C950 , 32'h09962550 , 32'hFCE7E8AC , 32'h17049720 , 32'hF72AC020 , 32'h07A708B8 , 32'hF8169068 , 32'hF97DC600 , 32'hF1659930 , 32'hF1CAF030 , 32'hFF8A9D4C , 32'h17386E40 , 32'h0001F26A , 32'hED8E9200 , 32'hF24E56B0 , 32'h11493E60 , 32'h06E54DD8 , 32'hF527B7F0 , 32'hEC151CC0 , 32'hFD82DB3C , 32'hF7EA5950 , 32'h0A2F59E0 , 32'h0949B020 , 32'h0601BCB8 , 32'hEB042FE0 , 32'hFFB11D9E , 32'hF48A4980 , 32'h04DDCAE8 , 32'hEEF76680 , 32'h00010F2B , 32'hFDDCB468 , 32'h0FEA6CE0 , 32'h00DB50E9 , 32'hFE97CDF4 , 32'hF4ABA210 , 32'h0001D8EE , 32'h0B429AC0 , 32'h06826F48 , 32'h19528500 , 32'hE7BEF920 , 32'h0000B118 , 32'hF7D9E860 , 32'h012D6984 , 32'h0EEDC970 , 32'h066A5B28 , 32'hFDE7012C} , 
{32'hF9343858 , 32'h02814640 , 32'hFCEE6690 , 32'hFFFA3F38 , 32'h0003B6BF , 32'hFFC8B234 , 32'hF3D6E5C0 , 32'hF8EC8520 , 32'hFFFB1B09 , 32'hF1931F50 , 32'hF79C0230 , 32'hFC70F524 , 32'h071C67D8 , 32'hFB428798 , 32'hE8E60EE0 , 32'h0DC3BE00 , 32'h13F95A20 , 32'h22842000 , 32'h16EF6AC0 , 32'h00030DE8 , 32'h09A622C0 , 32'hFBDBDA58 , 32'h08BEB780 , 32'h00005801 , 32'hFA6CEB70 , 32'hF8178388 , 32'h15CC3D00 , 32'hF0D40880 , 32'h05591C50 , 32'h0198CE5C , 32'hFC0FC258 , 32'hEC72B700 , 32'h04A994D0 , 32'hEB1D71C0 , 32'hFFFE9B17 , 32'hE99C2140 , 32'h00F50A36 , 32'hF716C550 , 32'hF7CECB90 , 32'h00F360C9 , 32'h080BEC00 , 32'h01B98924 , 32'hFFFEC1DE , 32'hFD5F2008 , 32'hE7952180 , 32'hF6CAC310 , 32'hEEFF2480 , 32'hFC13F8BC , 32'h00CC1524 , 32'h15DA1EE0 , 32'hEC4FD1E0 , 32'h006A07D1 , 32'h266A4040 , 32'hE793B1E0 , 32'h02EABA08 , 32'h061F4028 , 32'h041BA038 , 32'hFB5467C8 , 32'hFF436B16 , 32'h02F79BE4 , 32'hE9F28240 , 32'hF21F9850 , 32'h01035FC8 , 32'hFCB16D3C , 32'h088BBB10 , 32'h05007028 , 32'h00029D8C , 32'hE580E2C0 , 32'hF4DCF730 , 32'h0DF97B90 , 32'hF0674C40 , 32'hF4A062A0 , 32'h263AC5C0 , 32'hF7D62000 , 32'hEC7A2480 , 32'h0216F80C , 32'hF38CE4F0 , 32'hF2444FC0 , 32'h0A891140 , 32'h00FB9984 , 32'h0C0498D0 , 32'h09DFDBD0 , 32'hFC4DA8E0 , 32'hFFFE0ACC , 32'hFFF20B98 , 32'hFE73D8D8 , 32'h1C7E1A00 , 32'hFDB34CAC , 32'hF507B810 , 32'h0000C410 , 32'h0F126110 , 32'hFB887450 , 32'hFF8EF843 , 32'h0098125A , 32'hFFFFCAA6 , 32'h0B5036B0 , 32'hFBF7F058 , 32'h033DD788 , 32'hF2F5AEE0 , 32'hF025BD80} , 
{32'hFFA0A14C , 32'hFB329DF8 , 32'h130512C0 , 32'h00043A16 , 32'hFFFB6934 , 32'h05F3B538 , 32'hEAB333C0 , 32'hF3C36AD0 , 32'h00044365 , 32'h06723E20 , 32'hF96C6328 , 32'hF0176AA0 , 32'hE8143EE0 , 32'h0DAB3C50 , 32'hF7139310 , 32'hE205DCC0 , 32'h031FCA9C , 32'h1A260B00 , 32'h0B818B00 , 32'hFFFFC6A5 , 32'h0684F688 , 32'h20072740 , 32'h1E740E80 , 32'hFFFEB966 , 32'h00048AB1 , 32'h218F0EC0 , 32'h00024C7E , 32'hF5B9B2C0 , 32'h0C8AD3F0 , 32'hFD8FA2E0 , 32'h0134F264 , 32'hFD77F2D0 , 32'h013E2BE0 , 32'h070ADD68 , 32'hFFFCBFBF , 32'h0B3CA0F0 , 32'h0F598D20 , 32'h06486800 , 32'h1025F220 , 32'h15E5C460 , 32'h0199AC64 , 32'h03586974 , 32'h00B69762 , 32'hFA58FB30 , 32'hF33015C0 , 32'hFB9D43F8 , 32'hF8CB5958 , 32'hFC87DD1C , 32'h0D56E490 , 32'hDF713A40 , 32'hFA47C868 , 32'h02C02644 , 32'hF887FAF0 , 32'hFD9AB000 , 32'h0DA147B0 , 32'h08415750 , 32'h0990B4C0 , 32'h14C54A20 , 32'h0C170030 , 32'h022012B4 , 32'h0AB54D50 , 32'hF267DA40 , 32'hF8298650 , 32'hFF7FEA76 , 32'h02B37764 , 32'h08551940 , 32'h000408AF , 32'h0F64E3B0 , 32'h02DE0F7C , 32'hF8B25170 , 32'h17226F60 , 32'hF59C6340 , 32'h01DA4580 , 32'hE6CB9280 , 32'hFFCFB221 , 32'hF5A86440 , 32'h000C9327 , 32'h0BE7B2D0 , 32'h072FD220 , 32'hF0E9DEF0 , 32'h032EFFC0 , 32'h0E7C3520 , 32'h0BED4D50 , 32'h0000B43A , 32'hE2812AE0 , 32'hFE26468C , 32'h12162560 , 32'h138D6CE0 , 32'hFB419E30 , 32'hFFFF0B2F , 32'hF10CB350 , 32'h088769A0 , 32'h03641A1C , 32'h0C769B20 , 32'hFFFAB374 , 32'hFFD9C43E , 32'h09AE4150 , 32'hF0C87360 , 32'h10348600 , 32'hFD436B8C} , 
{32'hF249F8A0 , 32'hE4BFBFC0 , 32'hFC1DF6E0 , 32'h00088F08 , 32'hFFFE2D05 , 32'h05FEA760 , 32'h110D7AA0 , 32'h0B0FB000 , 32'hFFFED778 , 32'hEEA7E260 , 32'h14712100 , 32'h0BEBE890 , 32'hEDF9F680 , 32'hE8634DE0 , 32'hF3000ED0 , 32'hFD8C1194 , 32'hF784F790 , 32'h08E85C90 , 32'h080EDC30 , 32'h00027485 , 32'h0BBAEBD0 , 32'h1039E360 , 32'hF4B25320 , 32'h000218E1 , 32'hF18A1E40 , 32'h01882600 , 32'hFD9B06D0 , 32'hE751A3A0 , 32'hFA8C9488 , 32'h01B1C5F4 , 32'hEDF4F1C0 , 32'hFDAD6970 , 32'hF76F01D0 , 32'h0A60E670 , 32'h000073A0 , 32'hFB9AB058 , 32'hF3F00670 , 32'h13BA04A0 , 32'hEBB29B60 , 32'h06699920 , 32'hF293BF80 , 32'hFF661787 , 32'hE60E6120 , 32'hED047180 , 32'h0A9198C0 , 32'h06557508 , 32'h066A7390 , 32'h163C20E0 , 32'hEFEFA5E0 , 32'hF0653A70 , 32'hFDF40310 , 32'h05E40008 , 32'h00B24433 , 32'hFBDF5390 , 32'hF6F10E20 , 32'h05969440 , 32'hF4EAE090 , 32'hFDC9911C , 32'hFE5830C0 , 32'hF1186970 , 32'h07D10A80 , 32'h02F118D4 , 32'h0D8EC770 , 32'hF3F39C50 , 32'h0DB38630 , 32'h12B5C720 , 32'h000025D2 , 32'h0813F230 , 32'hFC995010 , 32'hE136C920 , 32'hFE3E81FC , 32'h028F71C0 , 32'hFEEEBE7C , 32'hF5D38360 , 32'hEEA75360 , 32'h021EABD4 , 32'h0EA2A9E0 , 32'h0DFD8CD0 , 32'h0EEC4FF0 , 32'hFD94CAD8 , 32'hFF01F3DF , 32'hE6826340 , 32'hFF7920B4 , 32'h0002163A , 32'h0B002AB0 , 32'h09FA94F0 , 32'h0331D868 , 32'h079397A8 , 32'hE4974060 , 32'hFFFA3CC7 , 32'h084C3EB0 , 32'h03283500 , 32'h023646DC , 32'h038B538C , 32'h0002193B , 32'hF9A8AC60 , 32'h1D6D2860 , 32'h00010765 , 32'hD88C7100 , 32'hFB952560} , 
{32'h194AF2C0 , 32'hDCA5C980 , 32'h0A73C150 , 32'hFFFD1C99 , 32'hFFFC79C7 , 32'hEC599DE0 , 32'h07415EA8 , 32'h0A902490 , 32'hFFFDC697 , 32'hFCEE004C , 32'h1A63B420 , 32'hE6C4C320 , 32'hF9619F98 , 32'hFF1D9D33 , 32'hE1905960 , 32'h06C8F8B0 , 32'h027FC708 , 32'h12BA1B80 , 32'h13B67FA0 , 32'h0002DE04 , 32'hFA995AD0 , 32'hFE614F38 , 32'hF6374650 , 32'h00033609 , 32'h00448FA9 , 32'h08687890 , 32'hFB2C4030 , 32'hFFED5D3A , 32'h0090795A , 32'h027428F0 , 32'hEC56F140 , 32'hF00CB620 , 32'h1B754680 , 32'hFB36BAF0 , 32'h0003A7EF , 32'hFCE583D0 , 32'hF7EE2B60 , 32'h0209DA3C , 32'h05E0F870 , 32'hFC1608A4 , 32'h01177828 , 32'h00669AE3 , 32'h01D5DD24 , 32'h0B2E8C40 , 32'h06EB6258 , 32'hFCE45334 , 32'hFD21F394 , 32'hE919C7A0 , 32'hF74C44E0 , 32'h00A7FCC6 , 32'h03E2BF40 , 32'h044E1F80 , 32'hF510EB80 , 32'hFCF444DC , 32'hF1B00050 , 32'hFDE0D344 , 32'h0443AC98 , 32'hFB06D2B0 , 32'h00E990D6 , 32'h0CDE5BE0 , 32'hEFE13FA0 , 32'hEFC95560 , 32'hF0ABEF30 , 32'hF9486860 , 32'h011CBAD4 , 32'hE7555620 , 32'hFFFF37D3 , 32'hFCC0DA14 , 32'h0A7939F0 , 32'hE4439EA0 , 32'hF03E3DB0 , 32'h063DB2B0 , 32'h016FEA80 , 32'hF48AA510 , 32'h0E5A5040 , 32'hE6A51360 , 32'h05D72740 , 32'h075D55A8 , 32'hFA04CDA0 , 32'h17575DE0 , 32'hD4CF1C00 , 32'h010D5BA0 , 32'hFFCCA4A4 , 32'hFFFA65C8 , 32'hF4A9F340 , 32'hF413F510 , 32'hF22B8420 , 32'hFFC25857 , 32'h07DD7F78 , 32'hFFFAA60E , 32'h0378632C , 32'h0C0FBE90 , 32'h046DDDB0 , 32'hECE376A0 , 32'h0004D18D , 32'h062645E8 , 32'hF46D4F90 , 32'h1161B6C0 , 32'h077E1390 , 32'h0BD7C220} , 
{32'h01947478 , 32'h0B0A0D90 , 32'h08C45D30 , 32'hFFFC364F , 32'hFFFEBA64 , 32'h0949A670 , 32'h1024D320 , 32'h11FBFD00 , 32'h0000668A , 32'hFBF8F258 , 32'hEED23880 , 32'hFBDA0970 , 32'hFF85D431 , 32'h0CC4EE50 , 32'hE6B78FE0 , 32'h08134BC0 , 32'h01C280C0 , 32'h17B9B320 , 32'h02847F54 , 32'h000014EB , 32'h13708600 , 32'hF4100690 , 32'h017CE5D8 , 32'h0000429C , 32'h05E9E568 , 32'hE4B06960 , 32'h10C65AE0 , 32'h05655E60 , 32'hEB64BDE0 , 32'hF8A31050 , 32'hFF9D9701 , 32'hFC1AE070 , 32'hFC7C6298 , 32'h1669CD60 , 32'hFFFE2B57 , 32'hFD085E4C , 32'h0755BB10 , 32'h0B2447D0 , 32'h02C185B8 , 32'h0F3C56B0 , 32'hF6314E20 , 32'hFF258300 , 32'h127D3360 , 32'hF24ABFE0 , 32'hF21A3920 , 32'h09C86330 , 32'h08E4B550 , 32'h0FBE2050 , 32'h059313F0 , 32'h094A6BA0 , 32'h03DBFCBC , 32'h0C41A230 , 32'hFAA99288 , 32'hF3F7AE40 , 32'h014CDD24 , 32'hFE59D700 , 32'hF5F5C860 , 32'h00125AD5 , 32'hF1E71F10 , 32'h1D1232C0 , 32'h1D86DF20 , 32'h1C67FCE0 , 32'hF9172788 , 32'hFA7CD7D0 , 32'h09AAE8E0 , 32'hE20254A0 , 32'hFFFF102C , 32'h16F0EA20 , 32'h07462540 , 32'hE8DAF940 , 32'hFB670E60 , 32'h0DD7C0D0 , 32'h0FD48440 , 32'h0EB13100 , 32'h05B1B240 , 32'hFA25C800 , 32'h008DA9A1 , 32'h00DD0840 , 32'h0CB6F010 , 32'hF3936CB0 , 32'h11F7FF40 , 32'h07976E80 , 32'hF1573210 , 32'h0001F80E , 32'hF0C760A0 , 32'h0FE28660 , 32'hFD8BF0A4 , 32'hF7462FA0 , 32'h11AA1DA0 , 32'hFFFD85E0 , 32'hFC4BEA84 , 32'h01207C80 , 32'hFF715B1F , 32'hE554E380 , 32'h0001103B , 32'hF682DBA0 , 32'h117FD7E0 , 32'hFEEC9660 , 32'h105C59A0 , 32'hEE1E3040} , 
{32'h021CE8F0 , 32'h09C874F0 , 32'hF9A1A270 , 32'h0002E49F , 32'h0005100A , 32'hFEF059F0 , 32'h0C077810 , 32'hDF5CC900 , 32'hFFFB8145 , 32'hFF7328AC , 32'h08CB4640 , 32'hFE90B558 , 32'hF8B8B160 , 32'h15EED060 , 32'hEF109000 , 32'hF2BD1D50 , 32'hFDE36CA8 , 32'h0E9AD900 , 32'hF6AD50C0 , 32'hFFFC1FB2 , 32'hFD20DF28 , 32'hF2711810 , 32'h04DA2C80 , 32'h000324A5 , 32'h17DA4260 , 32'hF1A6E1A0 , 32'hEFF6CAA0 , 32'h07387470 , 32'hE020EAE0 , 32'h063FF8B0 , 32'h015EF43C , 32'hF1C40BA0 , 32'hF0C36DC0 , 32'hF3A881A0 , 32'hFFFC3E53 , 32'hF8693560 , 32'hE47FC560 , 32'hFF958941 , 32'hFD49AD44 , 32'hFDA3417C , 32'h045D67C8 , 32'h012B5468 , 32'h0234BFF0 , 32'hF744C3F0 , 32'hF8066DB8 , 32'h09F2EB30 , 32'hF78E9DB0 , 32'hFEC3056C , 32'hF68BF360 , 32'hEF7D7C40 , 32'hEF6D3E80 , 32'h19D8AE20 , 32'hFE61D50C , 32'hF7D0FCD0 , 32'h01B31274 , 32'hFC1A33C4 , 32'hFEE5B200 , 32'hE2008420 , 32'h0934AC40 , 32'hF153D0B0 , 32'h06B6A470 , 32'hEA4AA380 , 32'hFB175608 , 32'h14A63600 , 32'hF2885A50 , 32'h0EDA1080 , 32'hFFF81FC8 , 32'hE8427360 , 32'h07518D00 , 32'hF736E430 , 32'hF74D8E90 , 32'hFB75E190 , 32'hF18009D0 , 32'h006DF1A9 , 32'h0EE7D350 , 32'h0544A560 , 32'hEC09B800 , 32'h0F19BE30 , 32'h071D8EA0 , 32'h085383B0 , 32'h1B5F2CC0 , 32'hEADFBF60 , 32'hF0485160 , 32'hFFFBB338 , 32'hF90CB548 , 32'h0ED15990 , 32'hECB00340 , 32'h16FC50E0 , 32'hFD67ECA4 , 32'hFFFF6C5D , 32'hE8935D00 , 32'h07DF1E20 , 32'h1443E520 , 32'h00D31D57 , 32'h00030EA3 , 32'h0AADA780 , 32'hFBCCDBF0 , 32'h01100FB8 , 32'h07EAD0F8 , 32'h03AA868C} , 
{32'hEE7A3860 , 32'hF0357A80 , 32'h012EA360 , 32'h00023B34 , 32'hFFFDB2DB , 32'h00326FF0 , 32'hFB139F48 , 32'hE8F62AE0 , 32'hFFFD5C80 , 32'hFFA20AF2 , 32'h04E75C70 , 32'hE6D6D620 , 32'hFC7F2F44 , 32'h07609B80 , 32'hEF035AC0 , 32'h018E33A0 , 32'h06D26580 , 32'hFFA08BB6 , 32'hF26DBC00 , 32'hFFFFB5DB , 32'hEB19F3A0 , 32'hFFCB0226 , 32'hF7D30410 , 32'hFFFEAF0C , 32'hEB1F74A0 , 32'h00889B90 , 32'h004A9A1E , 32'hEB8C3E60 , 32'hF5F17350 , 32'hF79B5CB0 , 32'h096E1CA0 , 32'hE78EC8C0 , 32'hF140F100 , 32'h12DF5DA0 , 32'hFFFF917E , 32'h01967A08 , 32'hFE833CB0 , 32'hFD4A36AC , 32'h142BE980 , 32'h064D2D68 , 32'h11A24540 , 32'hFE63B014 , 32'h0FD44210 , 32'h0E8C4C00 , 32'h05F07DD0 , 32'hFD7DE43C , 32'h1D953E80 , 32'hFD2AA1D8 , 32'hE9440700 , 32'h0C54D470 , 32'hFF0530BF , 32'hF3FF8700 , 32'hFE4083C8 , 32'h130B8840 , 32'h019BEF28 , 32'h0A194720 , 32'h031F7364 , 32'hF0339910 , 32'h06C54DB0 , 32'h08826F60 , 32'h0ACCDA70 , 32'hFEBAB3B4 , 32'hF4BE12E0 , 32'hFDF45E38 , 32'h266AA300 , 32'h0B503560 , 32'hFFFFB9CF , 32'h05620460 , 32'h00615F1D , 32'h139ED480 , 32'h0A0299E0 , 32'h23495780 , 32'h01FE8220 , 32'h05696A90 , 32'hFF6ADACE , 32'h1344A680 , 32'hF1D85DD0 , 32'hEC047600 , 32'hE2EF0A80 , 32'h0650B308 , 32'h0414ADD8 , 32'h015A7B38 , 32'h0852C0E0 , 32'h00020DFE , 32'hFCD3A988 , 32'h0B69DB50 , 32'h01A95128 , 32'h07A893F0 , 32'hDF3BAB80 , 32'h00009AB1 , 32'h085251B0 , 32'hFC70E8C4 , 32'hFE24A000 , 32'hF4B49080 , 32'hFFFEC3A9 , 32'h04186B20 , 32'h117A3A80 , 32'h06EC8508 , 32'h0B7EFF30 , 32'h09FE00A0} , 
{32'hF844EB48 , 32'hF28EE060 , 32'hF502F680 , 32'hFFFB08F8 , 32'h000069B2 , 32'h15B97AC0 , 32'hEEB86B80 , 32'h0E9EA5E0 , 32'h00067797 , 32'h0B6B38B0 , 32'h094BFBA0 , 32'hFD54E020 , 32'h0F423460 , 32'hFD2C97C8 , 32'h00E5BD4E , 32'h08521060 , 32'hFB3B6C40 , 32'hEE0C9720 , 32'h00D13484 , 32'h00045EE9 , 32'hF8E63FB0 , 32'h20EEBE00 , 32'h0CAFA720 , 32'h000060BB , 32'h015AA38C , 32'hF1647B80 , 32'h21457D80 , 32'hF2E471A0 , 32'h035D43A8 , 32'hFDF02008 , 32'hF9C00CF8 , 32'h0807D780 , 32'hF0D35E30 , 32'hFF1750B5 , 32'h0001632E , 32'hF9CF65E8 , 32'hF37BC940 , 32'hEB426AE0 , 32'h05A1BFA8 , 32'hF35E6AF0 , 32'h00B6C647 , 32'h014161EC , 32'hFE6B9D5C , 32'hF7B04D20 , 32'h089AFEE0 , 32'hEBE4DAC0 , 32'h016235C4 , 32'h0A876890 , 32'hE72CF3E0 , 32'h16121D40 , 32'hF10CEFB0 , 32'hF6621F50 , 32'hEC1BAA20 , 32'hF94F3FD0 , 32'hE79800A0 , 32'hEF5B7840 , 32'hF86AB5B0 , 32'h00191D1B , 32'hF867B548 , 32'hFB5178A0 , 32'h07DEEBE8 , 32'hE5B413E0 , 32'hFAD7C7C8 , 32'h10DA1460 , 32'h0C5B8840 , 32'hF00CB500 , 32'h00005A56 , 32'h00D1CD7D , 32'h1646C220 , 32'hF4B7F8A0 , 32'h1CD38460 , 32'hF90DF108 , 32'h151A4100 , 32'hFEF3C0A0 , 32'h19E26EA0 , 32'hFAA420D0 , 32'h023E197C , 32'h04F5F658 , 32'hF7B08970 , 32'hEE24FA80 , 32'h0D5648B0 , 32'h06473470 , 32'hF45443C0 , 32'h000B138E , 32'h014582C0 , 32'hFDA424C0 , 32'h04D1ED60 , 32'h0E5777E0 , 32'h0BBFFB60 , 32'hFFFF9BDB , 32'hE48A9F40 , 32'h0A0D7350 , 32'h015CDF08 , 32'hFDA1FF08 , 32'hFFFE2D80 , 32'h08631F30 , 32'hEC68E440 , 32'hFE5FCC30 , 32'hED5616C0 , 32'hFF959F2D} , 
{32'hF5AA4560 , 32'h0D505450 , 32'h018066AC , 32'h0006812C , 32'hFFFEA415 , 32'hE7BA3960 , 32'hFA8C7248 , 32'hFE2029E0 , 32'h00031D15 , 32'hFACC6698 , 32'h0AEA1930 , 32'hF6AB47E0 , 32'hFDFFBC80 , 32'h0CE64140 , 32'h018FDFA4 , 32'h109B4900 , 32'hED59FEC0 , 32'hFF8A3A94 , 32'hE2BE25E0 , 32'h00027405 , 32'hFE9CFBEC , 32'h05E52758 , 32'hF8193F98 , 32'hFFFABEFA , 32'h057E2E00 , 32'hE90C0840 , 32'h14A1A8A0 , 32'hF7B67720 , 32'hE7446D40 , 32'h08B72B40 , 32'hFE7E2C80 , 32'hED8AEBE0 , 32'hEE75AD60 , 32'hFDB624F0 , 32'hFFFFDBB8 , 32'h1BE2C360 , 32'h041DB060 , 32'hFB14BC58 , 32'h07BC4CC8 , 32'h03B8B288 , 32'h03A03418 , 32'hFF427921 , 32'h0826D670 , 32'hEC30E2E0 , 32'hF3D9E1C0 , 32'hFCCDB2F4 , 32'hFE16C86C , 32'hF56FAF70 , 32'hF7C10D70 , 32'hEC31C2E0 , 32'hFF454F95 , 32'hEA6F36A0 , 32'h0097BEFF , 32'hE9E0D420 , 32'h061F62D8 , 32'h0CC649B0 , 32'h0E01AA90 , 32'h0653D3C8 , 32'hF93F0448 , 32'hF0AC28A0 , 32'hF5A65960 , 32'h22745C00 , 32'h0D64B020 , 32'hED8BA000 , 32'hF86FD748 , 32'hF830F850 , 32'h0006BB1B , 32'hF155E960 , 32'h08DE8980 , 32'h025FE270 , 32'h14E57900 , 32'h0C272D90 , 32'hFCC11FF0 , 32'hE317BA60 , 32'h05EAC708 , 32'hEB2997E0 , 32'hEC4B6840 , 32'hFD0186CC , 32'h17BA3160 , 32'hF9EB0A50 , 32'hEF128B40 , 32'hF9F41578 , 32'hFD0DB4BC , 32'hFFFFA2EB , 32'h0296FF58 , 32'hF0D1CBC0 , 32'h0AAC6FE0 , 32'hF1C2D330 , 32'hF7B9E620 , 32'h0008920F , 32'h01A3B5DC , 32'h0CEF3170 , 32'hFA774818 , 32'h00FD6D0C , 32'h0001FC04 , 32'hEF015B40 , 32'hEF3BFDA0 , 32'hFC81F488 , 32'hF4ED3780 , 32'h18823AC0} , 
{32'h14979EA0 , 32'hF9EA5F08 , 32'hECF314E0 , 32'hFFFE9996 , 32'h0002C7D0 , 32'hD4EA2480 , 32'h0450F760 , 32'hFCCD55B0 , 32'h0001CB77 , 32'h05421D50 , 32'hF8CAE588 , 32'hFDA2EC54 , 32'hF44492C0 , 32'h02A9ED08 , 32'h0AD0B920 , 32'h0C70C2C0 , 32'h130798E0 , 32'hFB229B18 , 32'hFFC355D1 , 32'hFFFDA07C , 32'hF6190970 , 32'h08E0B450 , 32'h0241A368 , 32'h00000E6C , 32'h05709F70 , 32'hE5ADF6C0 , 32'h12A49640 , 32'hFE427E40 , 32'hF3C95870 , 32'hF78559C0 , 32'h03DFEF18 , 32'hFC3FF100 , 32'h10888A40 , 32'h083B9620 , 32'h00091965 , 32'h0CF81AC0 , 32'h03317D20 , 32'hFD6B6120 , 32'h1CD6AF00 , 32'hFE685270 , 32'h0BFF95A0 , 32'h001C8D2D , 32'hF681EC50 , 32'hF89DF768 , 32'h0B6D5610 , 32'h05880950 , 32'hEC8F6AE0 , 32'h13474220 , 32'h057BDB30 , 32'hF8298D28 , 32'h057BF178 , 32'hFA24BCE0 , 32'h1DB23C60 , 32'hFFF506BD , 32'hF829E6A0 , 32'hF9ECD4F0 , 32'h0B74E150 , 32'h0359FDD8 , 32'hDA290D40 , 32'hFFA6CA89 , 32'hEEA39100 , 32'hEBD86040 , 32'hFFB3A8DB , 32'hF8AA3150 , 32'h07DADB10 , 32'h1936EEA0 , 32'hFFFC3EC3 , 32'h0EFFDBD0 , 32'h016CD590 , 32'hF03CF8E0 , 32'h12893020 , 32'hFAA119B8 , 32'hEBBC8E20 , 32'h039D7BDC , 32'hFBB9ECC0 , 32'h0336F528 , 32'h13A0BCA0 , 32'hF8EF1B48 , 32'hFD42FD90 , 32'hFE8EAF10 , 32'h05BA8A30 , 32'hF8010CE8 , 32'h0F6F8C90 , 32'hFFFD7F98 , 32'h07BB4A58 , 32'h07841488 , 32'hFB4B1648 , 32'hFAD982C0 , 32'hF7CBD0C0 , 32'hFFFAA72B , 32'hF74BF620 , 32'h029C5A38 , 32'h11BBC9C0 , 32'hF4C38EC0 , 32'h00017289 , 32'h09273860 , 32'hFF0858EF , 32'hFA6F4538 , 32'h13513120 , 32'hD958C0C0} , 
{32'h031DC240 , 32'hF3211D50 , 32'h0553A538 , 32'h0001F8BD , 32'hFFFF160F , 32'hE9950620 , 32'h0A9A4840 , 32'hFB4E69B8 , 32'h00056BF2 , 32'hF9D53498 , 32'h00D26F71 , 32'hFC1DCB50 , 32'hFB29D3D0 , 32'h046F2760 , 32'h086D9510 , 32'hFD1D2698 , 32'hE2B11D60 , 32'hFF9F4F43 , 32'hFDAFE480 , 32'hFFFACF9B , 32'h041550F0 , 32'h00FFC48C , 32'h0F1E28A0 , 32'h00012C02 , 32'h0112B150 , 32'h1333DD40 , 32'hE80EACE0 , 32'h10E7D300 , 32'hF113A260 , 32'h0BE9E5E0 , 32'h0023F858 , 32'h0DFAF180 , 32'hFCCAAF3C , 32'h007B75F0 , 32'h0001DE8F , 32'hFC91C324 , 32'h09679F90 , 32'h00ACC5F0 , 32'h103B1DA0 , 32'hF4441220 , 32'h0748D8D8 , 32'hFFEB490F , 32'h02D2CC68 , 32'hE9E43BE0 , 32'hF8A9E718 , 32'hFDC48008 , 32'h05E29030 , 32'hFBBD7818 , 32'h12292340 , 32'hFD6316C8 , 32'hEDC71180 , 32'h02A35F28 , 32'h11CB1640 , 32'h07EB1208 , 32'h00AA3077 , 32'hF8961388 , 32'hFCE68C68 , 32'h01147BBC , 32'hEFD94580 , 32'h1060A740 , 32'h0533B468 , 32'hF25173C0 , 32'h1750FA00 , 32'h0B3E06D0 , 32'h10397960 , 32'hED90C680 , 32'h000BA1FD , 32'hE73CD320 , 32'h02ECD368 , 32'hF6EE14D0 , 32'h158CDA00 , 32'hF5CFCAC0 , 32'h1708F7E0 , 32'h1CE53A60 , 32'hDCCB8C00 , 32'h0D724840 , 32'hF34ED240 , 32'hFC76C5F8 , 32'hE79C6F20 , 32'hE9860440 , 32'hFA4AFC30 , 32'hF711E430 , 32'h0EFFF980 , 32'hFFFAF17F , 32'hEC4B70A0 , 32'h05C34228 , 32'hF597FEB0 , 32'hF1370410 , 32'h05D52B30 , 32'hFFFD7971 , 32'h05485A18 , 32'h13D78020 , 32'h028B3618 , 32'hEEA22B40 , 32'hFFFF9381 , 32'hFB1B0ED8 , 32'hFEE90460 , 32'h03D08530 , 32'hE299A0E0 , 32'h1256C140} , 
{32'h18333820 , 32'h0D5A0820 , 32'hFE42E430 , 32'h00050A65 , 32'hFFFD7895 , 32'h0149D424 , 32'hFB17DBC0 , 32'hFE6AB290 , 32'h0007DA38 , 32'h036AADFC , 32'hD504D9C0 , 32'hFD5DEBA0 , 32'h0735A380 , 32'h050A2B60 , 32'h034F2C80 , 32'hFB80FA90 , 32'h0365F3BC , 32'hF4B79CF0 , 32'hF7FC2A90 , 32'h000445EB , 32'hFE135760 , 32'hFD650C24 , 32'h03891270 , 32'h00012764 , 32'hEE899CE0 , 32'h020519C8 , 32'hFB5867F8 , 32'hF52E4F90 , 32'h0DC92AB0 , 32'h0A0777C0 , 32'h0ABD1A40 , 32'h174C7140 , 32'hF7F1CA80 , 32'hFC35E3F0 , 32'h0003CC1C , 32'hEFA1FBE0 , 32'hF6E20DA0 , 32'hF8B82400 , 32'hFCEB5830 , 32'hEF420EA0 , 32'h023E7994 , 32'hFEB82090 , 32'h107C1060 , 32'h05A6ED08 , 32'h0E43BCC0 , 32'hFC28B130 , 32'hEA4960A0 , 32'h0C1C1250 , 32'hFC509BC8 , 32'hFD0961C4 , 32'hFB8DDDB8 , 32'h0B2E02B0 , 32'hFF1DC9F3 , 32'h0E6AE640 , 32'hF2149560 , 32'h0982A000 , 32'h065E11D0 , 32'hFE92CA34 , 32'h1302D680 , 32'h0AE6C730 , 32'hF32EDE20 , 32'hFF3F2084 , 32'h1F803260 , 32'h0753B710 , 32'h14AD5D80 , 32'hEBF0E7A0 , 32'hFFF8926A , 32'h052CAEE0 , 32'hF8141E08 , 32'hDC9FE480 , 32'h0CBD11C0 , 32'h0A533510 , 32'hFBDDAEC0 , 32'hEF9005C0 , 32'h0311BA60 , 32'h0F198A50 , 32'hE3B21320 , 32'h055E34B0 , 32'h23003FC0 , 32'h01FA8058 , 32'hE7BEAB00 , 32'hFC33F230 , 32'hEA73F460 , 32'h00015C80 , 32'hFC7C5FAC , 32'h030E3C14 , 32'h041DDC10 , 32'h004CCFDE , 32'hE00B6580 , 32'h0004E8CD , 32'h0A71FEE0 , 32'h04F61248 , 32'h0CF3E690 , 32'hFCD1B92C , 32'h000429E7 , 32'hFF02C6DF , 32'h01E34984 , 32'h111ABC40 , 32'h0CBE32B0 , 32'hFB46F868} , 
{32'hF4B5CAC0 , 32'h0516F6E8 , 32'h03A4D9C8 , 32'hFFFA891C , 32'hFFFDC706 , 32'hEE085C40 , 32'h095BA170 , 32'h0F0AA0F0 , 32'hFFF95982 , 32'h101D4460 , 32'hE08EB020 , 32'hF11FE570 , 32'h0EB0E7E0 , 32'hE35B4D00 , 32'hE2BF0BA0 , 32'h0A3A4650 , 32'h0470BE88 , 32'hF61E5E30 , 32'h13841B00 , 32'h00068A90 , 32'h0A498950 , 32'hFFD7965B , 32'h128F38E0 , 32'hFFFF5C5A , 32'hF7B8BCD0 , 32'hFE317F58 , 32'hFA8AF658 , 32'hF3C24600 , 32'hEA625BC0 , 32'h05E4F718 , 32'h01041D98 , 32'hFC73778C , 32'h08873E20 , 32'hF0A5CF70 , 32'h00048018 , 32'hFBFA1510 , 32'hF38B7100 , 32'h04294950 , 32'hF9B7E268 , 32'hE1F2A3A0 , 32'hF610C930 , 32'h0022F2CD , 32'hF2F2D970 , 32'h015608F4 , 32'hFA0ACCA0 , 32'h01FAFB58 , 32'h12EC7DE0 , 32'h0B71E540 , 32'hF20CF810 , 32'hE829C3A0 , 32'h2089DB80 , 32'h0586DD58 , 32'hFCFB0884 , 32'h15FB9D20 , 32'h1113DAE0 , 32'hF3080670 , 32'h07D22EC8 , 32'hFE9B7DC8 , 32'h04E97488 , 32'h15252B00 , 32'h045079C0 , 32'h06DB0000 , 32'hF7FCAE10 , 32'hF9BD9830 , 32'h0BC06CA0 , 32'hFED067AC , 32'h0005606F , 32'hF1606B10 , 32'h10289A20 , 32'h06C985F0 , 32'hFBE35BC0 , 32'hF1BD78F0 , 32'hE328B840 , 32'hEE1533E0 , 32'hF2C27630 , 32'h001A43A6 , 32'hED5B6860 , 32'hF7712310 , 32'hF2ABB950 , 32'hF8E6CE28 , 32'h0644C5E0 , 32'h09718340 , 32'h07D95140 , 32'h000729B2 , 32'h07657C48 , 32'hFF0A2474 , 32'h11379620 , 32'h09A11CF0 , 32'h0AEE4F80 , 32'h000163A0 , 32'hED7A7160 , 32'hFB1669E8 , 32'h0C6F8DA0 , 32'h02A3EE48 , 32'hFFF88116 , 32'hEF0008E0 , 32'hEEDC84E0 , 32'hF5035DF0 , 32'hF790A050 , 32'h0172646C} , 
{32'hF5733E10 , 32'hE8AFF7E0 , 32'hF6CBDC50 , 32'hFFF90CA9 , 32'hFFFC78E1 , 32'hFFF090D8 , 32'h1718A8A0 , 32'hF785D8C0 , 32'h00039134 , 32'hE0AC21E0 , 32'hCF91C900 , 32'h040952E0 , 32'h07E28A38 , 32'h08CE0310 , 32'hF113B670 , 32'h059388A8 , 32'hFE67DCB8 , 32'hE5003B40 , 32'h0A1BC530 , 32'hFFFEE96D , 32'h0C613DC0 , 32'h13850D20 , 32'hEDA3DA80 , 32'hFFF98B7A , 32'h0A534110 , 32'h11761080 , 32'hFA4E44D8 , 32'h030B8370 , 32'h0C7C58E0 , 32'h02BE9CB0 , 32'hF0DCD8D0 , 32'hF682B5D0 , 32'hFAB0F160 , 32'h065C3630 , 32'h00036BCC , 32'h1350BD20 , 32'hF6F05780 , 32'hFC2406B8 , 32'hFA3B1000 , 32'h008C5E06 , 32'h0F76C150 , 32'hFE523998 , 32'h048325F0 , 32'hE6F7C160 , 32'hFA7140B0 , 32'h01A8FA78 , 32'h073EA988 , 32'h07B82510 , 32'h0E245910 , 32'h10C26CC0 , 32'hFA0FC850 , 32'hEDCEAEA0 , 32'h079199D8 , 32'hF64B5300 , 32'hFF1C9054 , 32'hDF8B5700 , 32'h130885E0 , 32'hF32E0D00 , 32'hFCE28490 , 32'hF743AF70 , 32'h0F429B70 , 32'h009F97C7 , 32'h03EFAED4 , 32'h0556E880 , 32'h0B184130 , 32'h0CB63800 , 32'h00109E46 , 32'h01009384 , 32'hEC967F60 , 32'h097C8700 , 32'hF66B4430 , 32'h04EEB8E0 , 32'hF43ED8C0 , 32'hFC70578C , 32'h11112E60 , 32'h05A83570 , 32'h02C84480 , 32'h163B3BE0 , 32'h12B2E5A0 , 32'h0E305050 , 32'hF84E7868 , 32'h04CA42F0 , 32'h101972E0 , 32'h000530CA , 32'hF3CA7530 , 32'hFA2C8A80 , 32'h0EBEAEA0 , 32'h03A562D8 , 32'h12AE8A40 , 32'h0001B418 , 32'h0114D354 , 32'h05C82500 , 32'hFCDD40B0 , 32'hF496BEC0 , 32'h00032011 , 32'h1081F020 , 32'hFA9AAEF8 , 32'hFE5579B4 , 32'h0ABDDCC0 , 32'h10D3FB00} , 
{32'hFCB47F40 , 32'hF99C0E68 , 32'hD1904400 , 32'hFFFCC302 , 32'hFFF68D2D , 32'hEFB07B60 , 32'h0654F3B0 , 32'hF6692150 , 32'h000049C6 , 32'h15B228C0 , 32'hFB1B52E0 , 32'h09BF15D0 , 32'hF503A870 , 32'h1ED8B0A0 , 32'h01BBF1B8 , 32'h00BE7FC0 , 32'hFC5DD850 , 32'h05B8EDE8 , 32'h0F5050B0 , 32'h00003F4C , 32'h090E07E0 , 32'hEFA2B9C0 , 32'hF118EB40 , 32'hFFF887F8 , 32'hF9E50B88 , 32'hFD763334 , 32'hF782B7D0 , 32'hF603E350 , 32'h05E5DFC8 , 32'hF669B4D0 , 32'h0A59E670 , 32'hF7B21070 , 32'h093937C0 , 32'hFC69D740 , 32'h00016117 , 32'hEFCB11A0 , 32'h09980E90 , 32'h061ED9A0 , 32'hFBFD5B98 , 32'hF2E408E0 , 32'hF8F95BB0 , 32'hFC827F88 , 32'h0FA87250 , 32'h0FE46100 , 32'h04AF4798 , 32'hFB2B4900 , 32'h03232400 , 32'hF9A84838 , 32'hFF5C70CB , 32'h00AA02B3 , 32'h0DB13EE0 , 32'h09D52000 , 32'hF9DBAB50 , 32'h09BD5710 , 32'hE19E2A60 , 32'h0D742470 , 32'h08A4F100 , 32'h1A2D8440 , 32'hEB5E4A60 , 32'hFFE2DF8B , 32'h19246F80 , 32'h17254DC0 , 32'hF99C4358 , 32'h061EB158 , 32'hFA1ADCA0 , 32'h083913E0 , 32'hFFFEB2C1 , 32'h0139B7C0 , 32'h00F5A604 , 32'h036D5810 , 32'h0E8B0380 , 32'hFB6E0018 , 32'h1ABEDC00 , 32'h09C8BBE0 , 32'hF83B6588 , 32'hF98AD180 , 32'h01C74C60 , 32'h098373F0 , 32'h07F6E7B0 , 32'h1498AF20 , 32'hF5B21570 , 32'hEC2F2440 , 32'h005A8186 , 32'hFFFDDB6F , 32'hF2B47960 , 32'h079CB620 , 32'h1D92F6E0 , 32'h13B85A00 , 32'hFFAD24E6 , 32'h000572F4 , 32'hF4844660 , 32'hF3613300 , 32'h09A5CF80 , 32'h06B0A898 , 32'h0003C446 , 32'h0B7E9090 , 32'hF02A4E90 , 32'hE91215C0 , 32'hF2079660 , 32'h12A531C0} , 
{32'h1BF9FF20 , 32'h0ECBD980 , 32'h015DAC9C , 32'hFFFD8D04 , 32'h0005888F , 32'h062D88B8 , 32'hF86FB768 , 32'h02BAEA38 , 32'hFFFE184C , 32'h002ED4EB , 32'hF2292750 , 32'h00F069A5 , 32'hFF3F0F93 , 32'hFF4E7799 , 32'hFD8CCEF4 , 32'h1833FDA0 , 32'h0CF8F030 , 32'hF8CEECE8 , 32'hFC2137A8 , 32'hFFFFA3E6 , 32'hF7DA28C0 , 32'h10537C40 , 32'h01E5EE90 , 32'h0004D533 , 32'hFA799498 , 32'h10E8FEE0 , 32'hEB307600 , 32'h1AB26440 , 32'h0B8ACD00 , 32'h09138670 , 32'hF4DF4480 , 32'hE7D9A640 , 32'h0D3C9280 , 32'hFC30B770 , 32'hFFFAB84B , 32'h050BB140 , 32'h1384B140 , 32'hF53CFB20 , 32'h142C83E0 , 32'h00276F25 , 32'hF84EF908 , 32'h01E099D4 , 32'h0A0F8B30 , 32'hDFBF5840 , 32'h1612DCC0 , 32'hEFF0B340 , 32'hE8A5D8C0 , 32'h066E6188 , 32'hEFE7EF40 , 32'hF792C0A0 , 32'h079F3DF8 , 32'h04535EA8 , 32'hFBFC16F0 , 32'h0016B44C , 32'h0B98A830 , 32'hF01688A0 , 32'hEA62B080 , 32'hF839D900 , 32'h00EDB9A1 , 32'h07F117D0 , 32'h11436AE0 , 32'h17BA6800 , 32'hF3E87890 , 32'hF54621B0 , 32'hF90723E8 , 32'h0DA24300 , 32'hFFFFBDCA , 32'hF7A4BF80 , 32'h022B2FE8 , 32'hFB6A88D0 , 32'hFCA99ED0 , 32'hF8776C28 , 32'h11ACAEE0 , 32'hFCDE9A60 , 32'h1AAFF8A0 , 32'hF86E8248 , 32'hF58B7AB0 , 32'hE83D7480 , 32'hFA3B4808 , 32'h16DE8820 , 32'h0E249800 , 32'hFFB5A03C , 32'h023FE07C , 32'h0001059A , 32'hF7E2EA20 , 32'h08878FA0 , 32'hEEE575E0 , 32'h08B7E9F0 , 32'hE7F1DBC0 , 32'hFFFBE71C , 32'h0AB7BD20 , 32'hFB23C6F8 , 32'hFE61BA64 , 32'h01EAF1FC , 32'h00070936 , 32'h02D15FAC , 32'h05811268 , 32'hF4010310 , 32'hDC823F40 , 32'hFB0A0B98} , 
{32'h05F6BCB8 , 32'h04C6C778 , 32'h106599A0 , 32'hFFF7948C , 32'hFFF56C4C , 32'h06416D48 , 32'hF1209590 , 32'hF5C1C860 , 32'hFFFB955D , 32'hEFD85080 , 32'h0067F002 , 32'h05E01918 , 32'h035CF1DC , 32'h1B1D5CA0 , 32'hFDD64168 , 32'hFB9CA140 , 32'h0F378B00 , 32'hFB95B048 , 32'h0C925190 , 32'hFFFF429A , 32'h0781D5F8 , 32'h149C8A80 , 32'hDBB5D200 , 32'h000278F0 , 32'h0631D048 , 32'h0CDDF960 , 32'h0EA06300 , 32'hF8ED1B00 , 32'h00E62F32 , 32'h0D65E350 , 32'h0912A9F0 , 32'h02BAB8EC , 32'h0268FB9C , 32'hF363CE90 , 32'hFFFD32DB , 32'h079DE3C0 , 32'hE1F32A60 , 32'h0164B2C4 , 32'h0BA434F0 , 32'h047BE5B8 , 32'h08936F80 , 32'hFF46F090 , 32'hF5D8D200 , 32'h0F802D00 , 32'h19137A40 , 32'hFC9CD648 , 32'hFA8B15E0 , 32'h01CE748C , 32'hFB2BD660 , 32'hFF69EFA4 , 32'h1664AC20 , 32'h088BD2A0 , 32'h06F81AF8 , 32'h0DE74890 , 32'h103A08C0 , 32'hE985F5E0 , 32'hF2070F10 , 32'h21C87B00 , 32'hFDB44A7C , 32'hE797DCE0 , 32'h07C26B28 , 32'h04A30098 , 32'hFEE3E4A0 , 32'hEDFA2A20 , 32'hFE02A050 , 32'h0CD8D280 , 32'hFFF5DFF4 , 32'hFB4FEC28 , 32'h0C0608B0 , 32'hF9244670 , 32'hF6E35920 , 32'h0573DCC8 , 32'h19CCE0E0 , 32'h011EEA84 , 32'hDF17DAC0 , 32'h0A0AA4D0 , 32'hF11825C0 , 32'hFB1ED138 , 32'hF9585238 , 32'hFC988554 , 32'h0A142C20 , 32'hF22E5DB0 , 32'hE62229E0 , 32'h0000576A , 32'h00DDF04B , 32'hF754BAE0 , 32'hFB7410D8 , 32'hFB49B958 , 32'h0F2F38A0 , 32'hFFFF93A5 , 32'hF8DD6F28 , 32'h0F2C35B0 , 32'h00A19593 , 32'hE7E2A7E0 , 32'h00098EF9 , 32'hEA03D4A0 , 32'hFAE18140 , 32'h05750418 , 32'h0F37ECB0 , 32'h04FADF38} , 
{32'h255A6680 , 32'hEC83F260 , 32'h01E0D514 , 32'h0004EA9D , 32'h000642FA , 32'hFC2DCE84 , 32'h03714F64 , 32'hFFAD0514 , 32'h0005FC1C , 32'hFC273CA8 , 32'hFB6FAC70 , 32'h126682A0 , 32'h0DAC2BD0 , 32'h022F3A38 , 32'h14E28640 , 32'hF83BC550 , 32'h09743A80 , 32'hFEBE0CCC , 32'h0181D974 , 32'hFFFCFFC4 , 32'hFA33F2B0 , 32'h077951A8 , 32'h0145D238 , 32'hFFFF1F9E , 32'hFE6376D4 , 32'h096D1420 , 32'h0197F45C , 32'hDEA9A4C0 , 32'hF254EE30 , 32'hE3840B00 , 32'hFF36F5AF , 32'hF5E82BA0 , 32'h081A4150 , 32'h05BE38E0 , 32'hFFFA24EF , 32'hFF383FA6 , 32'hF8E3DE18 , 32'h054F6D10 , 32'hF2423890 , 32'h16ED3FA0 , 32'hE8B12380 , 32'hFF14E6B7 , 32'h16B26460 , 32'h0BE18850 , 32'hF3F41580 , 32'h00897F62 , 32'hEEA0A6C0 , 32'h0BCDD410 , 32'h039EA1F4 , 32'hF21783D0 , 32'hFB14AA40 , 32'hFDA9BB6C , 32'hF38CB400 , 32'hEC2B0DA0 , 32'hED0C6400 , 32'hFAA5E518 , 32'h24DC8EC0 , 32'h007888BA , 32'h1FA57240 , 32'hEB479E60 , 32'hFB2C9EE0 , 32'h16594720 , 32'h077C1FE0 , 32'hFC6545C0 , 32'h0E850250 , 32'h04B979B0 , 32'hFFF6F11A , 32'hEBDA0FC0 , 32'h0A8C55D0 , 32'hFC3D3A68 , 32'hF86EABA8 , 32'hFFAF4388 , 32'h004EFBC8 , 32'h0F775F00 , 32'h02921510 , 32'h0402B3A0 , 32'hEE9AA500 , 32'hFB589028 , 32'hE6036FC0 , 32'hF6C6BF00 , 32'h03E33984 , 32'h115F0540 , 32'h0C98FAA0 , 32'hFFFB00A9 , 32'h03DC5294 , 32'h10E9F640 , 32'hF38DB210 , 32'hF0EB6D70 , 32'h0D81A3D0 , 32'hFFF581DF , 32'hF71C7780 , 32'hF56AFB60 , 32'h01E62230 , 32'hF63A3930 , 32'h0008BF84 , 32'hFD06052C , 32'hFDC45EFC , 32'hF7CD6180 , 32'hF33D5C50 , 32'hFC31C1F8} , 
{32'hF104D820 , 32'hFE987E04 , 32'hDC34DE40 , 32'h00018DCE , 32'h00013D85 , 32'h02319C9C , 32'hF044DDC0 , 32'h04FB2D18 , 32'hFFF98933 , 32'h03443A44 , 32'hFA2E73C8 , 32'hFEFA190C , 32'hF4EB4DD0 , 32'hE9E3B500 , 32'hF8167D88 , 32'h032A58BC , 32'hF61C3370 , 32'h03AEA438 , 32'hF1C8A050 , 32'hFFFEED63 , 32'hFDA5AE44 , 32'h0E183FC0 , 32'h0233B578 , 32'h0006F6C8 , 32'hF5B8A270 , 32'h09597860 , 32'hF17C3E30 , 32'h0B577980 , 32'hED480200 , 32'h14384A80 , 32'hF2149C30 , 32'h064222A8 , 32'h0B1E88A0 , 32'h0439AF70 , 32'hFFFC6E9C , 32'hFA099B58 , 32'hFC9384C8 , 32'h118D8CC0 , 32'hE961B7E0 , 32'hF6D7C290 , 32'hF01E7380 , 32'hFF3D829C , 32'h15995160 , 32'hFFD6EBDF , 32'hFD6609EC , 32'hEE514E00 , 32'hF1A4B160 , 32'hFCEB1A30 , 32'h0AD467D0 , 32'hEAA7DFE0 , 32'h00A094F5 , 32'hE35BF6C0 , 32'hFA28DD90 , 32'h02423338 , 32'h090E3310 , 32'h0764FC40 , 32'hF5B8F480 , 32'h0BDCB9E0 , 32'hF313EBE0 , 32'hEE8613C0 , 32'hEAD1C540 , 32'hF9B75A58 , 32'h054159F8 , 32'hFD1EA8F8 , 32'h15A3ECE0 , 32'h0B364D80 , 32'hFFFBF705 , 32'h03E3F880 , 32'hF9842C20 , 32'hF71A54B0 , 32'hF7D52140 , 32'h04648A10 , 32'h0C5AE0A0 , 32'h1C1868A0 , 32'h1110E020 , 32'hE2E618C0 , 32'hEB6CFC60 , 32'hF82E0538 , 32'hF2D8BDE0 , 32'h09D98870 , 32'h1523D0C0 , 32'hF73B7AE0 , 32'hF9BD9210 , 32'h00017C11 , 32'h044C5F48 , 32'h063BA890 , 32'h11010960 , 32'h022B882C , 32'h107C7320 , 32'hFFFBF039 , 32'h00755BA2 , 32'h08016C60 , 32'hF827B288 , 32'h01D18D08 , 32'h00088498 , 32'hFE387248 , 32'h08790200 , 32'h188C98E0 , 32'h23D82940 , 32'hFF5707B3} , 
{32'hFE1E166C , 32'hFD9A8DE4 , 32'hF32C7730 , 32'hFFFC95FA , 32'hFFFAFA79 , 32'hEE85EB00 , 32'hFBD9E0B0 , 32'h15487480 , 32'hFFFD11B0 , 32'hFD1A7A08 , 32'h091C46C0 , 32'h02D8FD18 , 32'h005D36FE , 32'h1367AE20 , 32'h086B5D80 , 32'h05300290 , 32'hFCFC4F54 , 32'h10AFEA20 , 32'hF24751F0 , 32'h00027113 , 32'hFEF1F278 , 32'h01B4DF70 , 32'hF670F100 , 32'hFFFAC458 , 32'h1E50A940 , 32'hFF976444 , 32'hE03096E0 , 32'hF60C8440 , 32'hF8915748 , 32'hFD6A742C , 32'h07162BA8 , 32'hF2465C70 , 32'hF215E000 , 32'h036CCEA4 , 32'h00060403 , 32'hFA769348 , 32'hFE6FB06C , 32'hFD533D14 , 32'hED9F4E60 , 32'hE72CE320 , 32'hFD75248C , 32'h05388D78 , 32'hF5477770 , 32'hEE8B21E0 , 32'hFAAD4EF8 , 32'h0904E100 , 32'h01DF59C8 , 32'h0879A620 , 32'hEFDEFCE0 , 32'h00F14C3D , 32'h0F3C8590 , 32'hEB4FF1A0 , 32'h06844928 , 32'h01E08A48 , 32'h0F624700 , 32'h0D9754C0 , 32'hF43FB610 , 32'h0C58F760 , 32'h15B63CA0 , 32'hF1C05FC0 , 32'h0A47A280 , 32'hF8EE7968 , 32'hEDE3C160 , 32'hFEBC9520 , 32'h0377A7D8 , 32'hFAB93170 , 32'h0001801A , 32'h01051350 , 32'hEF41B180 , 32'hF2FB0530 , 32'h03AE99EC , 32'hF0399190 , 32'h111EB020 , 32'hF844D5D8 , 32'h1005AC80 , 32'h2FF36F00 , 32'h005F4E45 , 32'hF18EFC90 , 32'hFB3A1380 , 32'hF9260240 , 32'hDD319900 , 32'h165EDBA0 , 32'h00AD1A2E , 32'hFFF926D0 , 32'hF7E6C140 , 32'h0179BA18 , 32'h02BA2A7C , 32'h090B3B70 , 32'h0C0757A0 , 32'h000720CB , 32'hFDE31464 , 32'h0525EE50 , 32'hEBB98340 , 32'h021765D0 , 32'h0003CF75 , 32'h027EA4BC , 32'hFE116EF8 , 32'h010BC714 , 32'h0A104B30 , 32'hDFD7A8C0} , 
{32'hF82F2390 , 32'hEF245380 , 32'hFD0D81AC , 32'h000CBBBC , 32'hFFFD22D1 , 32'hF4528390 , 32'h0095D573 , 32'hF9A663C8 , 32'hFFFEED22 , 32'hF072BB80 , 32'hFDFF12C8 , 32'h08CF6D90 , 32'hF7AC2620 , 32'hF06B5350 , 32'h0B1CBB00 , 32'hF1669D90 , 32'h0E9DCFC0 , 32'hFC022F90 , 32'h0E860900 , 32'hFFFD1853 , 32'h128AC1C0 , 32'h0CF4E580 , 32'h13F23D20 , 32'h00020A31 , 32'h01E0C188 , 32'h015D8E68 , 32'h09DEC940 , 32'h23BE7E40 , 32'h0605CBB8 , 32'h044A34C0 , 32'hFA664EB0 , 32'h014E00E8 , 32'h06B31C70 , 32'hF22CA090 , 32'hFFFCB01A , 32'hF03D45E0 , 32'h12204060 , 32'hEFD2FFA0 , 32'hF3749FC0 , 32'h01BD651C , 32'h0B1AF340 , 32'hFDD15AEC , 32'h1ACA3D40 , 32'hF8337760 , 32'hFDFA6228 , 32'hFDF4A330 , 32'h08ECC720 , 32'h001FD601 , 32'hF97B0ED0 , 32'hFF8953EF , 32'h0C46AAB0 , 32'h0A5ADB20 , 32'h0F876130 , 32'hFC2D2DB0 , 32'hF10B79E0 , 32'h19ED5240 , 32'h07FC3C50 , 32'hF77329F0 , 32'hF3639770 , 32'hF9B30610 , 32'h00755281 , 32'h129FDEA0 , 32'h010E5DA8 , 32'hEB0A0A60 , 32'h0380A624 , 32'h048B96F0 , 32'h000271B9 , 32'hFD3BAE84 , 32'h1819A0C0 , 32'hFF09DD10 , 32'hFF5DC2E6 , 32'h0C9F1EC0 , 32'hFF1B5D78 , 32'hE10B8D80 , 32'h08E6AEC0 , 32'h24E02280 , 32'h09397A80 , 32'hF3FD1FB0 , 32'hF124BA40 , 32'hF8C78318 , 32'hFB1569D0 , 32'hF4F411A0 , 32'hE5E02580 , 32'hFFFB0184 , 32'h00DD3FEB , 32'h05EA4750 , 32'hF28C6F70 , 32'hF96ECBF8 , 32'h0DA5B960 , 32'h0000FF16 , 32'hE0597F40 , 32'hFECB789C , 32'hF7D2C8F0 , 32'h11348F60 , 32'hFFF734F8 , 32'h07BA5CF0 , 32'h106A1E40 , 32'h1434D200 , 32'h09462DE0 , 32'h1365FC00} , 
{32'hF4758E80 , 32'hFE3587C0 , 32'h1E609420 , 32'hFFFB12E8 , 32'h0004B12F , 32'h04775BB8 , 32'hFDEB60E4 , 32'h006C7BF3 , 32'h0002DA88 , 32'h0001CE22 , 32'hF851A248 , 32'h0B33B950 , 32'hF6A7AD20 , 32'hEFD5C880 , 32'h14421C40 , 32'h0F5B1F70 , 32'hFE5E1ED4 , 32'hFE286604 , 32'h0427CFE8 , 32'hFFF872BE , 32'h038FE0D8 , 32'h118075C0 , 32'hFBFC0F98 , 32'h00064E00 , 32'h01AA8380 , 32'hF880C938 , 32'h03048988 , 32'hF8226120 , 32'hEE48AE80 , 32'h08A201A0 , 32'hFE9F62FC , 32'h001E1483 , 32'h015F0208 , 32'hF7A0A100 , 32'hFFFC160F , 32'h0F4F2F20 , 32'h1BD09780 , 32'h0BDE0820 , 32'hEBFCDD20 , 32'hFED0FBC8 , 32'h03FF1D14 , 32'hFEE2DF4C , 32'h17ABB380 , 32'h03F7C628 , 32'h0873DD70 , 32'hF7D306C0 , 32'h0C3E1690 , 32'hEE4A4500 , 32'hF3351DC0 , 32'hF22D0CB0 , 32'hFBD0C448 , 32'h012B9014 , 32'h1B5911C0 , 32'hED1F8640 , 32'hEB429C20 , 32'hF3E318B0 , 32'hF30B9910 , 32'hFE833DA4 , 32'h100221A0 , 32'h038D92D0 , 32'h05271FD0 , 32'hFD384260 , 32'hE4DC9A60 , 32'h1B82AD40 , 32'hF73EC2C0 , 32'hF6EF7780 , 32'hFFFC4001 , 32'hFCF522F0 , 32'hF4090930 , 32'hF554DF40 , 32'h12886020 , 32'hF71723C0 , 32'h0EFAC2B0 , 32'h007B6991 , 32'hFF0F4981 , 32'h0FD45E20 , 32'hFF991313 , 32'h0795B840 , 32'hFBB54700 , 32'h12B46920 , 32'hFD2B1AC4 , 32'hF30A6750 , 32'h0CAD88A0 , 32'h0008D092 , 32'h126B2520 , 32'hF4755320 , 32'hFF5670D9 , 32'h0897B530 , 32'h0122FF70 , 32'h0005A73F , 32'h0B9B6A20 , 32'hE87B4DE0 , 32'h2BDBCFC0 , 32'hF5E86DA0 , 32'h00042B9E , 32'hE6E42960 , 32'h048FFE08 , 32'hFAFAE570 , 32'h191D6F20 , 32'h03AB898C} , 
{32'h002B1439 , 32'hF09C43D0 , 32'hFB8613B8 , 32'h0006483B , 32'hFFFA7C87 , 32'hEE9EFA20 , 32'hEB962B60 , 32'hFC1B500C , 32'h000BB05D , 32'hFA6FFF78 , 32'h01EE52F0 , 32'hFF7845CF , 32'h025F48EC , 32'hEA6180E0 , 32'h0E3262B0 , 32'hF3DBCF20 , 32'hF6EE2EA0 , 32'hF06C8750 , 32'h0A676A40 , 32'h0003A5E0 , 32'hFDB9A13C , 32'h05235F20 , 32'hFEAE82C0 , 32'hFFFDC952 , 32'h07AD6858 , 32'hF5B512F0 , 32'h1E650960 , 32'h06F9E998 , 32'h05BF1E20 , 32'hF25F0BC0 , 32'h048B0C50 , 32'hF62625F0 , 32'h1372C320 , 32'h02A0ACD8 , 32'h0000C07A , 32'hD8472EC0 , 32'hFB944DD0 , 32'hFD5F28D8 , 32'h02669F54 , 32'hFE49710C , 32'hF98699B8 , 32'h00094331 , 32'hFEC7A328 , 32'hE3B9A5A0 , 32'hFE4A8FC4 , 32'h118D1A00 , 32'h18B25520 , 32'h168C41C0 , 32'h17ED1940 , 32'hFA029B50 , 32'h054B4BF8 , 32'hFDC87320 , 32'hE2B1CFA0 , 32'hED562BA0 , 32'h11BDCDC0 , 32'h00223453 , 32'hEDC8E9C0 , 32'hFECD4314 , 32'h0FCEB670 , 32'h0180B15C , 32'hFEDEAF0C , 32'h06468D10 , 32'hF07E9930 , 32'h1028D7A0 , 32'hFB136188 , 32'h0CAC6F70 , 32'hFFF7F695 , 32'hF531F430 , 32'hED5ABBE0 , 32'h0BA5C790 , 32'h0BB4D850 , 32'h08B0ED70 , 32'h05022478 , 32'h0D40B100 , 32'hEDD30F60 , 32'hF9599890 , 32'hFBCA49B8 , 32'hFDFF5378 , 32'h0D60A720 , 32'h12D2B7A0 , 32'hF638FA70 , 32'h01EF6750 , 32'hF76EE9D0 , 32'hFFFD8989 , 32'hE53E1260 , 32'h01506418 , 32'hF20DAE10 , 32'h00206DF9 , 32'hE5265D20 , 32'h000F1C85 , 32'hF9047E40 , 32'h01684298 , 32'h04E72F68 , 32'hFC551EC0 , 32'h00051A37 , 32'hEC8AED40 , 32'hE9BBF0A0 , 32'h0EFEA270 , 32'h0D5544B0 , 32'hFECEF714} , 
{32'h01DFB7F4 , 32'h0CB577C0 , 32'h0C4D1120 , 32'h00041D2E , 32'hFFFE3844 , 32'hFB4D3130 , 32'hFED788BC , 32'h010A1204 , 32'hFFF8F25C , 32'hFACE2300 , 32'hF374AF50 , 32'h1044F700 , 32'hFDED4490 , 32'hF10E90B0 , 32'hF6AAD860 , 32'hECC8CF60 , 32'hFBC6D2D0 , 32'h13609FC0 , 32'h0267B324 , 32'h00084CA3 , 32'h0F0103E0 , 32'hF84124F8 , 32'h03D61C20 , 32'hFFFE36C8 , 32'hFC8D365C , 32'hEF7FF220 , 32'h0E549030 , 32'h19F40620 , 32'h0B098DF0 , 32'hFC17DF2C , 32'hF4B34AE0 , 32'hF61EC7C0 , 32'hFA5098E0 , 32'h0B3E19C0 , 32'h00032370 , 32'h03F95F04 , 32'hDBAD7D40 , 32'h03756EC8 , 32'h0423B0C0 , 32'hD5BD16C0 , 32'hFE8905D0 , 32'h01B7A2B0 , 32'h04C471A8 , 32'h0B235D10 , 32'hFDC81CD4 , 32'h0A6F5600 , 32'h03D8E864 , 32'hF83CED70 , 32'hFAB52DB8 , 32'hFF05B620 , 32'hF50674A0 , 32'hFE661694 , 32'h05639040 , 32'h0615E420 , 32'hEEE65BE0 , 32'hF0E43EB0 , 32'h09B0F9A0 , 32'h020070E0 , 32'h049D0C38 , 32'hF09E1D10 , 32'hE5913520 , 32'h15058960 , 32'hFACB0A78 , 32'h0A6E51A0 , 32'hF6A3BF30 , 32'h0D05FF90 , 32'hFFF783CE , 32'h242DF740 , 32'h129B84E0 , 32'h054500F0 , 32'h13331F80 , 32'hF48936A0 , 32'h17F57320 , 32'hF9DD36E0 , 32'h00BEC43F , 32'h012D2860 , 32'hEFE523C0 , 32'h08AC2F20 , 32'hF52D1C10 , 32'h042E5760 , 32'hFE22EC34 , 32'h016F4450 , 32'h25B04840 , 32'h0007324D , 32'hF850C928 , 32'h071419D8 , 32'hEA2EB7C0 , 32'h0CEA3810 , 32'hF7476AD0 , 32'hFFFF96DB , 32'h0D331020 , 32'h06AF72A8 , 32'hE3B2AAA0 , 32'hFE178764 , 32'hFFFD07FB , 32'hF94E8088 , 32'h075756E8 , 32'hFB2DF878 , 32'h0145AC18 , 32'h027E6F8C} , 
{32'h0B755750 , 32'h0DF02730 , 32'h0B46E5A0 , 32'hFFF9B6BC , 32'hFFF14493 , 32'hFAFE7068 , 32'h0F20A8C0 , 32'hF85EC4D0 , 32'h000A2C87 , 32'hFFC62E63 , 32'hDC93B780 , 32'h149AACE0 , 32'hF9AB0DC8 , 32'h04EA2F08 , 32'hF83D7B10 , 32'hF2085A00 , 32'hF1B7F0A0 , 32'hF96FCD40 , 32'h02E291EC , 32'h000648B1 , 32'h0E40E380 , 32'hFF939D4C , 32'hFFDD3BB5 , 32'hFFFF5E86 , 32'hFF1AAB8D , 32'hF5DBA6F0 , 32'hFADCE788 , 32'hFF5DEB6A , 32'hF3F826E0 , 32'h0E5B5510 , 32'h0123E56C , 32'h06F87C50 , 32'h0ACD8270 , 32'h0A5F1750 , 32'h0005C9E2 , 32'h027FB1FC , 32'h06ADE3B8 , 32'hFDAB6B4C , 32'h04ECBBE8 , 32'hF5A13760 , 32'hF8280968 , 32'h03711294 , 32'hE3B68B60 , 32'h0CC36E00 , 32'h11AC9F40 , 32'h010E2540 , 32'h02E34B3C , 32'h094D3C90 , 32'hF3DA1C20 , 32'hEF753C80 , 32'hEA8E6640 , 32'hFAF18E68 , 32'hF7E696C0 , 32'hF672D730 , 32'h04D5D980 , 32'h1C362880 , 32'h0E58F360 , 32'hFB2DDF00 , 32'hFF37CB09 , 32'hF1732160 , 32'h117215C0 , 32'hE548DE60 , 32'hF9F07BD0 , 32'h058AEBE8 , 32'h17413540 , 32'hF9298030 , 32'hFFF81E6B , 32'hEB4152C0 , 32'h059A9370 , 32'h107553E0 , 32'hF26372B0 , 32'h11DE04C0 , 32'h27657340 , 32'hF59E6D70 , 32'h08600CC0 , 32'hE9FC7720 , 32'h29DD72C0 , 32'hE8B8FFA0 , 32'h013D3A48 , 32'h014C1D68 , 32'hF8ECB3E0 , 32'h02DEDE60 , 32'h0096E640 , 32'h0001207D , 32'h0ABF3F40 , 32'h00D00B8D , 32'hF1A7A480 , 32'hF789F5F0 , 32'hF690B940 , 32'hFFF924F2 , 32'hFA140740 , 32'hFAAB9600 , 32'hF57102A0 , 32'h03314B54 , 32'hFFFC024E , 32'hF4415860 , 32'hF6E4A7D0 , 32'hF48E14B0 , 32'h0D0E8260 , 32'h069266C0} , 
{32'h01DF83CC , 32'hEAE4EFA0 , 32'hFD27E758 , 32'hFFFFE29A , 32'h0000FAE5 , 32'h19088000 , 32'hF0E1EAF0 , 32'hFCC692BC , 32'h0000AAD1 , 32'h0B1D7240 , 32'hF8571278 , 32'hF85B99A8 , 32'h0A239680 , 32'hFF10F78F , 32'h02B1D9A8 , 32'h17690B80 , 32'h069FF658 , 32'h02A5D910 , 32'hF67F1E00 , 32'hFFF26EA8 , 32'hFBFF1D98 , 32'hF3520870 , 32'h07686110 , 32'h00024AC3 , 32'hFBB254A8 , 32'h10E95B00 , 32'hEF692760 , 32'h14C05840 , 32'hE651A060 , 32'hEFCC02C0 , 32'h084032E0 , 32'hFD6A7C88 , 32'hF7F411C0 , 32'h01288CF4 , 32'hFFF16D8B , 32'hFB491ED0 , 32'hE1897EE0 , 32'h03705CF4 , 32'hFD0BF764 , 32'h0B671840 , 32'hF4E4E9B0 , 32'h021D7604 , 32'h0187B2B0 , 32'h043E5BA8 , 32'hFFD07D0D , 32'hF1F45C60 , 32'hF302D300 , 32'h0DFCD850 , 32'hFA57E6B0 , 32'hFC4CD138 , 32'hF4A1CC10 , 32'h00F9C4BF , 32'h054E4930 , 32'hEB86ADA0 , 32'h08911180 , 32'hFA0DD2A0 , 32'hFBC00148 , 32'h1C886540 , 32'hEEF7AFC0 , 32'h083E7EB0 , 32'hF251E330 , 32'h19C37980 , 32'hF51B82B0 , 32'h227897C0 , 32'h0B5E95E0 , 32'hFB1A13F8 , 32'h0004ADA9 , 32'hF4523510 , 32'h02F8C6B8 , 32'h0B581610 , 32'h094BE850 , 32'hEF43CBE0 , 32'hF07F7200 , 32'hE0D06BE0 , 32'hEDC1DF80 , 32'h06EAB858 , 32'h2BF93A40 , 32'hFBF1B3E0 , 32'h03D843E4 , 32'h00CC69B0 , 32'hF7EC5F40 , 32'hF7ADA9E0 , 32'hF8C05F20 , 32'hFFF5C60A , 32'h02977884 , 32'h0B4E5D60 , 32'hFD512264 , 32'h07394F40 , 32'hF7A79700 , 32'hFFFE4AB2 , 32'h06E00E38 , 32'h06AFEFF8 , 32'hF008AB20 , 32'hEAF9B080 , 32'hFFF32B0A , 32'h072B07F0 , 32'h01F75064 , 32'h00C022D5 , 32'h0E27B670 , 32'h0F8D79D0} , 
{32'hFE915DCC , 32'h1965A340 , 32'hFC911A7C , 32'h0002450B , 32'hFFFE7D0D , 32'hF55D2260 , 32'h01A4F594 , 32'h08800910 , 32'hFFFEBD7C , 32'h02D59158 , 32'h0C9A6A40 , 32'h03F01EB0 , 32'hFBF54718 , 32'hE17CA640 , 32'h09770050 , 32'hF5A04880 , 32'hFABB54D8 , 32'hFE017E4C , 32'h0230481C , 32'h0005D4ED , 32'h02E7EA1C , 32'hFC0109BC , 32'h05321AB0 , 32'h0007434B , 32'hF938C8D0 , 32'h084E5710 , 32'hF55A8610 , 32'hE87CBE60 , 32'h0830D6C0 , 32'hED750780 , 32'hFCB22EE4 , 32'hFDF71328 , 32'hFF05D386 , 32'hFBF2CB98 , 32'hFFF8FCFF , 32'h18CA9280 , 32'hEDC8C700 , 32'hFA97A1C8 , 32'hE77274E0 , 32'h07823D10 , 32'h0383FA94 , 32'hFFF6623C , 32'hFE152738 , 32'hF61C2750 , 32'hF78EC690 , 32'h0177903C , 32'hEB0D4D40 , 32'h0024D865 , 32'hF268FC10 , 32'hF2CAA0E0 , 32'h07A1C590 , 32'h040E41D8 , 32'hFEFBF3FC , 32'h0D7FBA00 , 32'hF91643A0 , 32'hE15AAC40 , 32'h0F2283C0 , 32'hF3AF1360 , 32'hE4878B00 , 32'h0B7B0960 , 32'h077CF498 , 32'h057CE9F8 , 32'hF0D99C60 , 32'h15443AE0 , 32'hE3613C80 , 32'hFE6D3330 , 32'h00005672 , 32'hFAEDA5C8 , 32'hFA7DB078 , 32'hF569E440 , 32'hFA667378 , 32'h2BF3E540 , 32'h17D31A40 , 32'h015C81B0 , 32'hF8A9C778 , 32'h0B618D50 , 32'h0D3FCE90 , 32'hEB6D2540 , 32'hFCBCAB88 , 32'hF69E8BE0 , 32'h05D448A0 , 32'h0EB24750 , 32'hF8FF32E8 , 32'h0008B28C , 32'hEA832CC0 , 32'hFC74BADC , 32'h0BCCA8B0 , 32'hF6AD4C10 , 32'hEF81A6C0 , 32'hFFF6E973 , 32'h02967448 , 32'h196A8BC0 , 32'h06C0B5F0 , 32'h09272B20 , 32'hFFF930F7 , 32'h1195B160 , 32'hF9372D70 , 32'h059C6938 , 32'h112884A0 , 32'h0B2D4D80} , 
{32'hFC47CF08 , 32'h129F1C00 , 32'h01349A40 , 32'h0005A887 , 32'h00057E8D , 32'hEE9CBEA0 , 32'h184E8FC0 , 32'h0E480B90 , 32'h000E9F52 , 32'hFAE53D88 , 32'h0A01EEC0 , 32'hFF4B00CE , 32'h0311E828 , 32'h032ECDA8 , 32'hFEA8DCC8 , 32'hF3848100 , 32'h0816D670 , 32'hFEDD9A74 , 32'h08F16A30 , 32'hFFFF2314 , 32'h04798780 , 32'h137EE840 , 32'hEA8C7500 , 32'h00043095 , 32'hFF83D94C , 32'h242BF540 , 32'h07DC2688 , 32'h10FAB2A0 , 32'h03DD9528 , 32'hF06E4F90 , 32'hF3B35730 , 32'hF4EE01C0 , 32'hFA84EE30 , 32'hFF21C180 , 32'h000F8E2C , 32'h0BE5F8F0 , 32'hEEDFBDE0 , 32'h038A4390 , 32'hFB6DE578 , 32'h032D69E0 , 32'h05E8E158 , 32'hFD799A3C , 32'hFB0F12F0 , 32'h00C8BD59 , 32'h02ABF4F4 , 32'hF49AF240 , 32'hFC180904 , 32'hFD4BC97C , 32'hF20EDCD0 , 32'h08299790 , 32'hFD24B8A4 , 32'h08B69F30 , 32'h09D90300 , 32'hF1344830 , 32'h11921920 , 32'h19C12C40 , 32'h04DB1298 , 32'hFAFE3B58 , 32'h08E70300 , 32'h14118340 , 32'h0CB7B800 , 32'h06609138 , 32'h0FD24C20 , 32'h2EDFE940 , 32'hFE2DE698 , 32'hFF8A87C5 , 32'hFFFECAD1 , 32'h0D511CF0 , 32'h028FE12C , 32'h11013E20 , 32'h18BC85A0 , 32'hFFBF650C , 32'hFD078BB4 , 32'h0A357C00 , 32'hFAA8A4B8 , 32'hE48B97A0 , 32'hED3DA200 , 32'hED2253A0 , 32'hFE3B64B0 , 32'h04DF2B80 , 32'hEBBED520 , 32'hF4AC3700 , 32'hF8184500 , 32'hFFFBFCEC , 32'h1976C440 , 32'h0B6DE960 , 32'h07F760A0 , 32'hF7DFBC00 , 32'h04FD32F0 , 32'hFFF71BDC , 32'hE505E2A0 , 32'hF874C468 , 32'h029CA4EC , 32'h029D4550 , 32'hFFFD9D12 , 32'h05D85FB8 , 32'h0407E980 , 32'h105A7640 , 32'hFD6CC13C , 32'hE457AD80} , 
{32'hFA0BFDB8 , 32'h01C814C4 , 32'h0F84BF40 , 32'h00037142 , 32'hFFF8C8E8 , 32'hFE9B4568 , 32'hEFFF43E0 , 32'hF0117B60 , 32'hFFFE047A , 32'h0427DE20 , 32'hF3711560 , 32'h036FC118 , 32'h0373B028 , 32'hF3E8B930 , 32'hFF878BC1 , 32'hFD5A8778 , 32'h216D5AC0 , 32'hF7B11A20 , 32'h082682B0 , 32'hFFFFD764 , 32'hFAA505F0 , 32'h03EC4EF4 , 32'hF9C3EE40 , 32'hFFFAECAB , 32'h04C659E8 , 32'hFEFB8A8C , 32'hDBF54580 , 32'hF44D2B60 , 32'h06DEE108 , 32'hF7E5FAF0 , 32'hFD232348 , 32'hFD46B994 , 32'hF7F570E0 , 32'hFBBD3B00 , 32'hFFF4BECC , 32'h075B2878 , 32'hFDF4C15C , 32'hF43B5260 , 32'hF61FE3D0 , 32'hF5EBA550 , 32'h09A76DB0 , 32'hFC56F118 , 32'hF63EBD20 , 32'hE3DDE620 , 32'h0205CE5C , 32'h113EB340 , 32'h037CE3C4 , 32'hF861A400 , 32'hFD0A8C2C , 32'h0C01FBD0 , 32'hF52F6EA0 , 32'hFFC1ED8A , 32'hF8860208 , 32'h03CD82F0 , 32'hF8C71BA8 , 32'h23F97C00 , 32'h1046FE60 , 32'hF421B030 , 32'h05FD39F8 , 32'hF1FC31F0 , 32'hFC4E9E20 , 32'h0EABA420 , 32'hE2B2A220 , 32'hE7C6C160 , 32'h01A6F1FC , 32'hF10828B0 , 32'h00043535 , 32'h0A366E10 , 32'h1364DC00 , 32'hFC83FCEC , 32'h1CF83300 , 32'hEA710C40 , 32'hFB000C00 , 32'h1D072DC0 , 32'hED64AD40 , 32'hE9051140 , 32'h0EE3A7B0 , 32'hFECF6098 , 32'h078857A0 , 32'h043D55E8 , 32'h0C5787F0 , 32'h005BFBE8 , 32'hEE388A00 , 32'h0007D6FE , 32'h05D19810 , 32'h1154ED60 , 32'h04C27E90 , 32'hFD8ECC1C , 32'h0C125F40 , 32'hFFFCB825 , 32'h17DFBF80 , 32'h1A08FF80 , 32'h0EBB0520 , 32'hFAFF5D50 , 32'h00050B63 , 32'h04F30CB8 , 32'hF77D92C0 , 32'h08E3A040 , 32'h034663DC , 32'h04C240B0} , 
{32'hF9DDE888 , 32'hDD613480 , 32'hFCCF08D0 , 32'h0009E5DE , 32'hFFF76282 , 32'hFD5DEFBC , 32'hFBC342F8 , 32'h0E6E7BF0 , 32'hFFFC8667 , 32'h0213C9E0 , 32'hEE271DA0 , 32'h1213AB60 , 32'hFB612678 , 32'h150CD460 , 32'h158740C0 , 32'hFC989CB8 , 32'h12AF4300 , 32'h0ACC3CD0 , 32'hFEE47408 , 32'h000B090A , 32'h05362718 , 32'hFEF23780 , 32'h08EE4C60 , 32'h000E1CEC , 32'h05DC1E20 , 32'hF3E42D70 , 32'hF78C47E0 , 32'h1A8E5740 , 32'h0D72D410 , 32'h0DC9C270 , 32'hFC6D92E8 , 32'hFDCD1AF4 , 32'hF25964B0 , 32'hF9704950 , 32'h00002E4A , 32'hFF0E5ECA , 32'h011BE8EC , 32'h03EC252C , 32'hF33E8AB0 , 32'h00315E40 , 32'hF694B190 , 32'h02368F9C , 32'hFFB2D4AB , 32'h1EADD700 , 32'hECDB8300 , 32'h06C8E3C0 , 32'h0CB538B0 , 32'h09732B20 , 32'hE86F13C0 , 32'h0FD818C0 , 32'hEBD7D6E0 , 32'hFE12A614 , 32'h084603B0 , 32'h00EA9451 , 32'h1C063DC0 , 32'hEA7574A0 , 32'hFAE5D400 , 32'hFFA2478C , 32'hFD174A64 , 32'hFDE03604 , 32'h035B982C , 32'h029CC298 , 32'h06036390 , 32'hF18C9DE0 , 32'hF311A840 , 32'hFDFBF810 , 32'h00187834 , 32'hEC0EB0A0 , 32'hF96CC770 , 32'hE96F63C0 , 32'h1702BA60 , 32'h26F26800 , 32'hF1687D70 , 32'hFFC366A5 , 32'hF425A950 , 32'hDD63B880 , 32'hFC616738 , 32'hFCD6C1F8 , 32'hEBD62620 , 32'h07FB78E0 , 32'hFA691C58 , 32'h105737A0 , 32'hFC3840B0 , 32'h0003B857 , 32'h02B00AC0 , 32'h041C6B58 , 32'h013F4674 , 32'h0BE15450 , 32'hF7A96010 , 32'h0009B826 , 32'h047DE468 , 32'h0DAC1A20 , 32'h0DA74400 , 32'h0FC66730 , 32'h0007C387 , 32'hFC12F9D0 , 32'hFF0C071B , 32'hF31E5360 , 32'hFEE7D7B4 , 32'hF4B8CBF0} , 
{32'h056AB6A0 , 32'hFFFA77D6 , 32'h169B6C80 , 32'hFFF56933 , 32'h0009748D , 32'h0A3CD610 , 32'hF4CCA250 , 32'hFFCF569F , 32'h00088BAA , 32'h029EAB88 , 32'hF19AE560 , 32'hFCF3AC58 , 32'h0053DFDD , 32'h195A62C0 , 32'h03173740 , 32'h0529E240 , 32'h0E5DDA20 , 32'h121FB3C0 , 32'h0AA3D010 , 32'h00094672 , 32'hFF03A4BB , 32'h02FD1010 , 32'h0EA7EBA0 , 32'hFFFFD231 , 32'h00F4C040 , 32'hFD774EAC , 32'h16A40E40 , 32'h0B505070 , 32'hFEF4F2D4 , 32'hFB938B40 , 32'hF9AA4030 , 32'h02CD387C , 32'h080F9360 , 32'h050F2AF8 , 32'hFFFF168B , 32'h009FB858 , 32'h0DC0CC10 , 32'hFF738BDD , 32'hFE05F818 , 32'hE96E58A0 , 32'hF5B7A3F0 , 32'hFE4102DC , 32'hD32D9E00 , 32'hEE2E3240 , 32'hF923C128 , 32'hF6FA3740 , 32'hF702AA10 , 32'hE471A300 , 32'hF4AEE6B0 , 32'hF76B3E00 , 32'h00BD57E9 , 32'hEFD986A0 , 32'hF4D4B170 , 32'hFFDA75AA , 32'hF75EE410 , 32'h12DA0C40 , 32'hF262B0A0 , 32'h01BFD83C , 32'h01F286A0 , 32'hFCDFB618 , 32'hFA27E2D8 , 32'h1D825DE0 , 32'h09DD2CE0 , 32'h179C89C0 , 32'h06D31FC0 , 32'h0B03F760 , 32'h00081685 , 32'hF9DECFE0 , 32'hFFB91339 , 32'hF0D818E0 , 32'hEA560E20 , 32'h1AD4B360 , 32'hEBBB2AE0 , 32'h276D8840 , 32'h00947164 , 32'h1AC9B840 , 32'h0441B3E0 , 32'h0B1F4E40 , 32'hF6746070 , 32'h04183090 , 32'h0047FEE1 , 32'hFADACEB8 , 32'h0BC62E50 , 32'h000B370E , 32'h0BDF8CD0 , 32'hF2B754D0 , 32'h12CF3080 , 32'hFE2D95F8 , 32'hF5358F30 , 32'hFFFB9CCD , 32'hEFC989A0 , 32'h0E7C6DE0 , 32'h0184245C , 32'hFA1BDAC8 , 32'h0007A7D8 , 32'h0E70CB90 , 32'hF9C602F0 , 32'hFFCA8A4C , 32'h00BE7932 , 32'h0BC42FE0} , 
{32'h02492754 , 32'h0F064F90 , 32'h0670EF98 , 32'hFFF89918 , 32'hFFEB3F03 , 32'h0132DACC , 32'h08D26350 , 32'hF0E8B0A0 , 32'hFFFE1389 , 32'h07F17590 , 32'h0CC453A0 , 32'hEFEE0CC0 , 32'hFFA43FB2 , 32'hFD7B2AD8 , 32'hF759A380 , 32'h05A30480 , 32'h02F4E030 , 32'h048B3CB0 , 32'h089CA970 , 32'hFFF79EAA , 32'hF91DE640 , 32'h069ED850 , 32'h00EE901C , 32'hFFFF830C , 32'hFE31D55C , 32'hF6E86140 , 32'h028B5578 , 32'h22B186C0 , 32'h0B6BB2A0 , 32'h0A165990 , 32'h0C1577B0 , 32'hFD101BF0 , 32'hF6DAE2F0 , 32'hFE3EB21C , 32'h00025543 , 32'h0D8520D0 , 32'h0018160C , 32'hFEE76AB0 , 32'hE11549E0 , 32'h0148DA34 , 32'hF8A3C250 , 32'h03BEFB54 , 32'h11D46B00 , 32'hEC40EC20 , 32'hFB37D160 , 32'h01661EC0 , 32'hFB07F5B0 , 32'hFC110A24 , 32'h00625C6E , 32'h0224AB08 , 32'h0E3D9A90 , 32'hF97668F8 , 32'hEAEC7100 , 32'h0273A7D8 , 32'hEF4BAE40 , 32'hEFF84E60 , 32'hFADA3960 , 32'hFBC92100 , 32'h0D9B6620 , 32'hF0C38AB0 , 32'h14EA5020 , 32'hEAB52A80 , 32'h08DC8F10 , 32'hF836B460 , 32'h0AD5DEB0 , 32'h0BB05AD0 , 32'hFFE5B735 , 32'hEC025BA0 , 32'h1A07F660 , 32'hEE27D520 , 32'h0C351360 , 32'h04B43838 , 32'hFA972A90 , 32'h01FB5280 , 32'hDCADA440 , 32'hF7085270 , 32'h086E1FF0 , 32'h03682EC4 , 32'h016E3E34 , 32'hF56E0050 , 32'hF2CA9CD0 , 32'hFEF0D3E0 , 32'h068313C0 , 32'h000A96B0 , 32'h040AA8E8 , 32'h04BB4038 , 32'h0D271440 , 32'hF3A35AF0 , 32'hF2C40B80 , 32'hFFFBFD8C , 32'h0B9F2D60 , 32'hD1705640 , 32'hE2904D60 , 32'hF3051E70 , 32'hFFFFBEC3 , 32'h146D51A0 , 32'hF087E970 , 32'hF5F4FDE0 , 32'h142A2E60 , 32'hF3693340} , 
{32'h07B21948 , 32'h09099350 , 32'hFD9B8D3C , 32'hFFFB5AA2 , 32'hFFFCBD79 , 32'hFD2A6A34 , 32'hE2AD3DE0 , 32'hF1117A60 , 32'hFFFFF9F4 , 32'h0DA4B940 , 32'hF569B060 , 32'h01DBF484 , 32'hF7567740 , 32'hFDB585B8 , 32'hFE0A6398 , 32'hFBB1F920 , 32'hF4596B80 , 32'h0C0C6C60 , 32'hFE09A094 , 32'h00152ABD , 32'h0136DB44 , 32'hF7128440 , 32'hEC0118E0 , 32'h00000676 , 32'h00BD005C , 32'h1E444F20 , 32'h25268B00 , 32'hDC90ED80 , 32'h0086EF91 , 32'h09D1E650 , 32'hFE60C930 , 32'h06168B18 , 32'hFA5EE0D0 , 32'hEFE201C0 , 32'hFFF98CDE , 32'hF1F335C0 , 32'h03E13F08 , 32'h092D3DF0 , 32'hFCC0B7C8 , 32'hEF8881C0 , 32'h11ACFD20 , 32'hFF4674DD , 32'h04C55BA8 , 32'hED881620 , 32'hFC3C33C8 , 32'h05227570 , 32'h0A1BCFF0 , 32'h094AA070 , 32'hFF9C5411 , 32'h09B72EB0 , 32'hE16357C0 , 32'h079D5638 , 32'hF5C16A30 , 32'h09E7FC70 , 32'h108DA9C0 , 32'hF7091F40 , 32'hFFF84ADA , 32'hFA8734F0 , 32'hE54F7200 , 32'h006ED4AF , 32'h114CA8E0 , 32'h0F446380 , 32'hFEF2D2E8 , 32'hF7F4B290 , 32'hEC415B20 , 32'hFB3A30B0 , 32'hFFFA0BFE , 32'hEBF66AA0 , 32'h02F886B4 , 32'hE782B8A0 , 32'hFB3910F8 , 32'hEFFAED40 , 32'hF0D9CE30 , 32'h022B1CF4 , 32'h0B49B3C0 , 32'hFA032CA0 , 32'h05E72B98 , 32'hEF6A0580 , 32'hF5B46E20 , 32'hFD28AA24 , 32'hEC00DBE0 , 32'hFCB4D22C , 32'h17D20B00 , 32'h000C7D24 , 32'h1843D8C0 , 32'h0E49B850 , 32'hF4957970 , 32'h03E492C8 , 32'h07FD8BA0 , 32'h000242E8 , 32'h0152258C , 32'hEE922140 , 32'hF4089E60 , 32'h02F13708 , 32'h0003B5F5 , 32'h0AB15810 , 32'h13B0C180 , 32'h05928E70 , 32'h0FD50420 , 32'h06AB7240} , 
{32'hF6EF6D00 , 32'h0BE409D0 , 32'h0507AFC8 , 32'h0009C051 , 32'hFFFA6FB8 , 32'h19DCBD40 , 32'hFD152B50 , 32'hFF17C7FF , 32'hFFF9B9F2 , 32'hFBE48880 , 32'hF80BAE40 , 32'h04000158 , 32'h07AAAE58 , 32'hF7B62D70 , 32'hFD3E65C0 , 32'h0486AE00 , 32'hF6FE0000 , 32'hEFB31000 , 32'h028119A0 , 32'hFFF35584 , 32'h03CF9430 , 32'hF6707180 , 32'hEBD37600 , 32'h00008251 , 32'h08B6AFD0 , 32'h0865CF10 , 32'h06FE6558 , 32'hF745D9E0 , 32'h0241B6A0 , 32'hFBA92768 , 32'h0AEB9320 , 32'hF5B6AF00 , 32'hFF255916 , 32'hF504D660 , 32'hFFEF972B , 32'h04B50F00 , 32'h10459500 , 32'h08956680 , 32'h07DC5E58 , 32'hF4347100 , 32'h02FBC248 , 32'hFF06A1C3 , 32'h3275A600 , 32'h05CF23F8 , 32'hFBA1D710 , 32'hF9BD4F50 , 32'h0857A750 , 32'hFF63B981 , 32'h07544EC8 , 32'hF8E47E18 , 32'h0D533B40 , 32'h0274ADA4 , 32'h0CA23B30 , 32'hFD15C600 , 32'h16337520 , 32'h15B8FC00 , 32'h00DCEFDF , 32'hFEAD4734 , 32'hFD17E68C , 32'hF6616E80 , 32'hECA03C60 , 32'hF18F6470 , 32'hF653E7C0 , 32'h16028220 , 32'h061E7BA0 , 32'h0E02AF40 , 32'hFFFD24C2 , 32'hF9462A48 , 32'h2901BB80 , 32'hEAA408C0 , 32'hF0DA9AA0 , 32'h19569AA0 , 32'hF645D980 , 32'h0DB4E990 , 32'hFABBD770 , 32'hFFB01964 , 32'h17517180 , 32'h082721B0 , 32'h07C64C18 , 32'hFE9AA874 , 32'hF0DFCB90 , 32'hFD525F70 , 32'h0B82E6A0 , 32'h0006A414 , 32'hF116B530 , 32'hFDFFE718 , 32'hFDE46D64 , 32'h0D3D5490 , 32'h03079794 , 32'hFFFFDD08 , 32'h0049832D , 32'h1ECDC700 , 32'hFA8DF288 , 32'h05C4B988 , 32'h0004E3CB , 32'hFD8C29CC , 32'hF9DB4350 , 32'hF5C6A4D0 , 32'hE385DF00 , 32'hE0D5E360} , 
{32'hF6F23F60 , 32'hFAFE5268 , 32'h171E6FA0 , 32'h0015622D , 32'hFFFB5516 , 32'hF85DC628 , 32'h1AA6E220 , 32'hF819C278 , 32'h00000489 , 32'h060F3670 , 32'h03D504A0 , 32'hFDACB470 , 32'hF6C3B7A0 , 32'h026FA03C , 32'h0B9B2700 , 32'h02027A38 , 32'hFB73ED08 , 32'hFFD6A121 , 32'hF8275420 , 32'h0006285D , 32'hF79E68A0 , 32'h043521C0 , 32'h0A5172E0 , 32'h00039420 , 32'hF349D450 , 32'hF0485E00 , 32'h0D3D8F30 , 32'hFF37F455 , 32'h0606AD10 , 32'hEE481DA0 , 32'h04B23D10 , 32'h04766710 , 32'hFDD0F4E8 , 32'hF8A34458 , 32'hFFFD7DA0 , 32'h0D4433A0 , 32'hF09F2880 , 32'hF2D77440 , 32'hFAC3B3C8 , 32'hFDC13B64 , 32'hFCD276D4 , 32'h01D0B57C , 32'h19A0EF20 , 32'h00C1513C , 32'hFDB7A73C , 32'hFE065698 , 32'hFAF5A720 , 32'h01AC9AAC , 32'hF92ED3C8 , 32'h0ACD57D0 , 32'h00572C6F , 32'hF85433E0 , 32'h13734DC0 , 32'h1A31A100 , 32'h13CB73C0 , 32'hF766FBF0 , 32'hF7919DD0 , 32'hFA6430A0 , 32'h09D73E40 , 32'hFA4D2810 , 32'h038C9798 , 32'h168DA1E0 , 32'hFFF7A85E , 32'hF7A9A430 , 32'h16CC99E0 , 32'h01BCF2B4 , 32'h00025F28 , 32'hFA99E808 , 32'hF333CC00 , 32'hFA9A39E8 , 32'hE15FB320 , 32'hCCF60640 , 32'h0DD30970 , 32'h19473BC0 , 32'h04E29930 , 32'hE6B88920 , 32'h14C11EE0 , 32'h08124920 , 32'hFE2D8A54 , 32'hF5CB8940 , 32'hEB109B60 , 32'hFF261580 , 32'hF3CB4390 , 32'hFFFD0E0F , 32'hF572DD90 , 32'hF6B111B0 , 32'h004811EE , 32'h04AA3038 , 32'hE494D500 , 32'h000A682B , 32'hE0F34FA0 , 32'h0B26F4A0 , 32'h07096D98 , 32'h122D5280 , 32'h0005D22E , 32'h0266A60C , 32'h075E9700 , 32'hFD3B8E30 , 32'h0C071DA0 , 32'h07356E30} , 
{32'h0820EE30 , 32'h10035EC0 , 32'hED488140 , 32'hFFFA0ADD , 32'h000D2C5C , 32'h1E8EC360 , 32'hFBE928E8 , 32'hF74BB7F0 , 32'h0006BC00 , 32'h06455748 , 32'hFF85FD70 , 32'hF217D890 , 32'h03BDBB1C , 32'hF48161D0 , 32'h02956FB0 , 32'hFE841F10 , 32'hE3BAD220 , 32'h06E368D0 , 32'hFCC78438 , 32'hFFEBE06E , 32'hF9296A18 , 32'hF4E98C90 , 32'h0220AAE0 , 32'hFFF92866 , 32'hF29DB690 , 32'h0CBE4B00 , 32'h149252E0 , 32'h1D73B9E0 , 32'hF5665530 , 32'hFCE91DF0 , 32'hFDC6FF40 , 32'hEE1E1200 , 32'hFD1E9E38 , 32'hF643C170 , 32'hFFF972EF , 32'h02E4B018 , 32'hFC41AA78 , 32'h03526940 , 32'hE27DDE20 , 32'h0878A160 , 32'h06C81D50 , 32'h0572D0A0 , 32'hE49C0BC0 , 32'h01FDE5D4 , 32'h08EA77D0 , 32'hF66717B0 , 32'hFA827698 , 32'hFE5A4830 , 32'h016D083C , 32'h09461EF0 , 32'h01C75270 , 32'h1030B780 , 32'h0AD0A190 , 32'h0172FBA0 , 32'hFFC27101 , 32'hF7E17EF0 , 32'h1A4AE5C0 , 32'hFF242D04 , 32'h1239ACE0 , 32'h00584D9E , 32'hFED8D030 , 32'hFF1982EE , 32'h01BFF47C , 32'hD024C240 , 32'h06296840 , 32'hF8D48B00 , 32'h0012D045 , 32'hFAC311B0 , 32'hFB790C10 , 32'h0B47A6D0 , 32'h181482A0 , 32'h07A1B978 , 32'h025481AC , 32'h14A32FE0 , 32'h0C3889B0 , 32'h0DF908C0 , 32'h119830C0 , 32'hF9CD9760 , 32'h0634FE20 , 32'h0C92B500 , 32'hEE1C32E0 , 32'hF667FFD0 , 32'h113E2B60 , 32'h00044B83 , 32'hF026EBB0 , 32'h021D7F30 , 32'h059B0EE0 , 32'h07E03000 , 32'h05095DE0 , 32'h000835AB , 32'hEB1409E0 , 32'h1192DEE0 , 32'h177F0B40 , 32'hF2BDF740 , 32'h00053B0D , 32'hEB72BDA0 , 32'h045CBCD8 , 32'hFD204B4C , 32'h000AD4EF , 32'hF0323E30} , 
{32'h055916D0 , 32'hF78C3CD0 , 32'h0CF62EA0 , 32'h00082E24 , 32'h000D4689 , 32'hFF1AEE4E , 32'hF12326D0 , 32'h135A26E0 , 32'hFFFD1CE0 , 32'h09BB4200 , 32'hF3E8F9D0 , 32'h0E6E5040 , 32'hF40BDFE0 , 32'h0A200330 , 32'h06C9B498 , 32'hFB799CB8 , 32'hF0ED8E40 , 32'h03BB0B2C , 32'h0AF88050 , 32'hFFF1A6FF , 32'hF4496720 , 32'h004E8FF7 , 32'h0EFB9D70 , 32'hFFFBC717 , 32'h0C697FC0 , 32'hFF9507D1 , 32'hFCC97088 , 32'hF9FF99A0 , 32'hFF407A45 , 32'h00C2EF02 , 32'hEF95DDC0 , 32'h0D26F200 , 32'hFC9E6144 , 32'h0934DE10 , 32'h0009E857 , 32'hFB0A46C0 , 32'hD21D4200 , 32'h079392F8 , 32'hF8763A90 , 32'h064B9170 , 32'h041FD950 , 32'h05A497D0 , 32'h21C13940 , 32'hF4EB5D90 , 32'h0B400F60 , 32'hEE368E60 , 32'h0D4CC0B0 , 32'hEEAF3700 , 32'hF8B36CD8 , 32'h00503D41 , 32'h0C01A8B0 , 32'hFACBDCF8 , 32'hFE42BF18 , 32'hE304B600 , 32'hF50F7EE0 , 32'h1290F960 , 32'hF9218058 , 32'hFD210564 , 32'hF1FA3150 , 32'h14B2D040 , 32'h19D9AEA0 , 32'hEB8EA7A0 , 32'h18A77D20 , 32'hE1914F60 , 32'hEDB8CD40 , 32'h067C9348 , 32'h0003602E , 32'h05109760 , 32'h0AE6EE00 , 32'h182303A0 , 32'hEEF23E40 , 32'hF562ADB0 , 32'hF4CC3970 , 32'h08FE8B90 , 32'hFA72B688 , 32'h0C542B60 , 32'hFD7D1ADC , 32'hF233DB20 , 32'h03F8D8F8 , 32'h0E0E2AB0 , 32'hFFE91565 , 32'h0534BF28 , 32'h087D0B40 , 32'h0001C8A6 , 32'h0C993850 , 32'hFE7A0EB8 , 32'h042BFAF0 , 32'hFEF0DD40 , 32'hEB421D20 , 32'h000F9F2D , 32'h083EDB70 , 32'h1858C380 , 32'h02FC8508 , 32'hFDFF03C8 , 32'hFFEEA20E , 32'hFF5B85A7 , 32'hF566D150 , 32'hEED3AD60 , 32'h08EC5EC0 , 32'hF9E2DD98} , 
{32'hF6A5C820 , 32'h071AF588 , 32'h04A741C8 , 32'hFFF6BEC0 , 32'hFFFEE6BD , 32'h03228BDC , 32'hF6E98C40 , 32'hEB243AA0 , 32'h0006FA4E , 32'hF3C0A670 , 32'hFF15257A , 32'h029AC250 , 32'hFCBAEA34 , 32'h0593B300 , 32'h176F4560 , 32'h08422680 , 32'hFB1978A8 , 32'hFEE7D0D4 , 32'hEDB42140 , 32'hFFF6CA7D , 32'h05509C18 , 32'h0CBA2630 , 32'h0369E264 , 32'h00013666 , 32'h02C3F46C , 32'h04820AC0 , 32'hEE041740 , 32'hF9CF0300 , 32'h06F24A18 , 32'hF70A38B0 , 32'h00FF6595 , 32'hF1DF32F0 , 32'h0A2EEBA0 , 32'h04CE1440 , 32'hFFF7B52B , 32'hFE628704 , 32'hDF4C79C0 , 32'hFADB6A00 , 32'hFE9F44BC , 32'hFF3C7924 , 32'hFB7E7C68 , 32'h00432D5E , 32'hE3AFC1C0 , 32'h030F5560 , 32'hF2FDC6E0 , 32'hFFA3D3F6 , 32'h107D7CA0 , 32'h01CFFFAC , 32'h1A585900 , 32'h003FA1E3 , 32'hF21DBEA0 , 32'hEB20D780 , 32'h02D859B8 , 32'h06136CD8 , 32'hFD151CE8 , 32'hFE76C0AC , 32'hF75EFA90 , 32'hFCDE0B18 , 32'hF06400A0 , 32'h1E0A1EC0 , 32'hFB6B8860 , 32'h095E2790 , 32'h0A905AE0 , 32'hFBDC03A0 , 32'h02B4498C , 32'h00E476EB , 32'hFFFD108F , 32'hFA2A1770 , 32'h39A20900 , 32'hF9BBB9B8 , 32'hF2A84510 , 32'h029238FC , 32'h0D867CA0 , 32'hF7A58290 , 32'h1388AC00 , 32'h02FDE92C , 32'h0102D5BC , 32'h10BC3500 , 32'hF5A82740 , 32'h0EF6BAD0 , 32'hF3AB05D0 , 32'hFC3E6EF4 , 32'hF3B75BF0 , 32'h0010089E , 32'hF152C230 , 32'hFF530BBF , 32'h0D2C1BB0 , 32'hF7824C90 , 32'h005C6CB4 , 32'hFFF5AE85 , 32'h08A5B770 , 32'hDC664440 , 32'h1ACBD640 , 32'h0C6BB060 , 32'hFFE3510E , 32'hF42B1810 , 32'h02F6D88C , 32'h03A38770 , 32'h01568480 , 32'hE94E18C0} , 
{32'hFB64C7F0 , 32'h18CBA8E0 , 32'h08053D70 , 32'h000DA7B3 , 32'h00121080 , 32'h02DB2D34 , 32'hF0B754F0 , 32'hF24720E0 , 32'hFFF95352 , 32'hFA1C3248 , 32'h05663860 , 32'hFA7070C8 , 32'h0F4D74F0 , 32'h026EBD78 , 32'hFA923188 , 32'h06BCEA90 , 32'h09E16E70 , 32'hF3DB0680 , 32'h059212C0 , 32'h000FA070 , 32'hF8847440 , 32'h0B7497A0 , 32'h11827C80 , 32'hFFE8E562 , 32'h03118014 , 32'h05787BB8 , 32'hFD9D719C , 32'h0ACA3FE0 , 32'hF9A8BD10 , 32'h000A293E , 32'h04F29978 , 32'hF564A1C0 , 32'hF80E5E00 , 32'hF94C6250 , 32'h000C1BA0 , 32'hF7C76020 , 32'hE754F980 , 32'hEFA69A40 , 32'hFD579B24 , 32'h009B187B , 32'hFC92E028 , 32'hFDBA9080 , 32'h0DF8E7B0 , 32'h09834A20 , 32'h0F452700 , 32'h0FA499A0 , 32'h18CE2260 , 32'hF9760740 , 32'h0C097170 , 32'hF45DA8A0 , 32'hF79B2090 , 32'hFC78C848 , 32'hFBE95DB0 , 32'h0732EC40 , 32'hE6B71AE0 , 32'h18EB9740 , 32'h07A3AF28 , 32'hF6CF2760 , 32'hF4200BA0 , 32'h0693BF58 , 32'h08C4A630 , 32'h0CA49A10 , 32'h0AC4EF80 , 32'h0043915D , 32'hFA1C37A8 , 32'h0E78C1C0 , 32'h00057F5D , 32'hFCA43A08 , 32'hC054FB00 , 32'hE1C38AC0 , 32'hF7639E80 , 32'h0547AB58 , 32'h06FD2728 , 32'hEADFF720 , 32'h02929390 , 32'hEE585880 , 32'h0E8EBDD0 , 32'h06242070 , 32'hE2992F80 , 32'hF7B8F540 , 32'hFF137C06 , 32'hF79EE540 , 32'h07B205E0 , 32'hFFF08704 , 32'hFD112F14 , 32'hF7788670 , 32'h079B5EA0 , 32'hFD018B6C , 32'h11769EE0 , 32'hFFF5F54F , 32'hFFC161F2 , 32'h06000128 , 32'hFC7B2E1C , 32'hF12AD740 , 32'hFFEDBF22 , 32'hF65BC3C0 , 32'hFA66F338 , 32'hF932F278 , 32'hF200DCC0 , 32'hE7AD4140} , 
{32'h00EADD63 , 32'h0CE76980 , 32'hF9A81A98 , 32'hFFEF77B2 , 32'hFFF414C5 , 32'hF80961B0 , 32'h071F01E8 , 32'hF33FABD0 , 32'hFFF302FB , 32'h056131B0 , 32'h03B11778 , 32'hFBCE5098 , 32'hFA6BE300 , 32'h005B891D , 32'h0B7FEC80 , 32'h0CBA0E60 , 32'hFCD112DC , 32'h01823E80 , 32'hFE4FADC4 , 32'hFFFF1530 , 32'h00DABF70 , 32'hFD710F48 , 32'hFA2C9720 , 32'h0004EE8D , 32'hFABF8F18 , 32'h04D0E548 , 32'h0674A488 , 32'h08563840 , 32'h07632EE8 , 32'hFD2324B8 , 32'h0443F3F8 , 32'hFD20426C , 32'hFD3B5594 , 32'h0D390D10 , 32'hFFFAD5F6 , 32'hEF181F80 , 32'h223518C0 , 32'h00B88389 , 32'hF3874820 , 32'h0AC5F4E0 , 32'hFDD2F67C , 32'hFFB15C75 , 32'hF3D4A220 , 32'h0AC50110 , 32'hFF870FAC , 32'h07E46FC8 , 32'h0B09D3A0 , 32'h0DF91380 , 32'h02BCC0FC , 32'h03646060 , 32'hF8FA34E0 , 32'hF4F37BB0 , 32'hF3E69880 , 32'h03A413C4 , 32'hE1DE3140 , 32'hED215800 , 32'hF7E41610 , 32'hF7A82C30 , 32'h0DA9A6E0 , 32'h04497FA0 , 32'h0FBAAC30 , 32'h0274BC18 , 32'hFD938EE4 , 32'h0DC4CE60 , 32'h0649EB18 , 32'h09284280 , 32'hFFFA35D5 , 32'hF765BB10 , 32'h174FFAA0 , 32'h07566E50 , 32'hEE66FCC0 , 32'hE9232DA0 , 32'h00E4A937 , 32'hE0D1FE20 , 32'hF77224E0 , 32'hF7A1AAA0 , 32'hEBD95880 , 32'hFCF50390 , 32'hFA19C450 , 32'h0A888120 , 32'hFC9FD364 , 32'hF6840370 , 32'h02F75800 , 32'h000BD1BC , 32'h10E7A6E0 , 32'hFF249260 , 32'h08CB31E0 , 32'hF2054230 , 32'h04C44750 , 32'hFFF97875 , 32'h08625B60 , 32'h4AE61700 , 32'hFE24D2C8 , 32'h0103DCB4 , 32'h0001EF96 , 32'h028748F0 , 32'h0B4BC700 , 32'hF6949360 , 32'h1150DFA0 , 32'hEE845DE0} , 
{32'hFF598037 , 32'h00BBC3D4 , 32'hFE560388 , 32'h001042CC , 32'hFFE64E1A , 32'hFF172674 , 32'h02F29D44 , 32'hFDF7A4E8 , 32'h00047E74 , 32'hFDECE5A0 , 32'hFE9FE60C , 32'h01702F58 , 32'h011EDE6C , 32'hFEE65718 , 32'h00A249D8 , 32'h003CFA49 , 32'h0335C1E8 , 32'hFD0E4AB0 , 32'h00159C9D , 32'h0010762B , 32'hFFB219AE , 32'h0149A784 , 32'hFD37E2CC , 32'h001605B4 , 32'hFF2AC528 , 32'h016C649C , 32'h012D7E38 , 32'hFD9A6700 , 32'hFF4CEAA3 , 32'hFD573AF0 , 32'h0083A3EB , 32'h00CD1156 , 32'h00CF3D8C , 32'h0060091C , 32'h007C9517 , 32'hFFAE7490 , 32'h02DB7AA4 , 32'h001D2951 , 32'h019B17C0 , 32'h00208899 , 32'h00B6640B , 32'h7FFFF800 , 32'h00CF14ED , 32'h001EA268 , 32'hFE325CF4 , 32'h01CE50F4 , 32'h0212FF60 , 32'hFE48E6C8 , 32'h0095D118 , 32'h025005A8 , 32'h01542874 , 32'h0109C89C , 32'hFF1CC4AB , 32'h0216B864 , 32'hFDFCF340 , 32'h038E4800 , 32'h00818015 , 32'h00FCCC55 , 32'hFDE462E8 , 32'h01056D04 , 32'hFE4B2F0C , 32'h0329CCE8 , 32'hFEC9BACC , 32'h031800CC , 32'hFFC76C20 , 32'h00D249CA , 32'hFFC845BA , 32'h01A00D94 , 32'hFEEB45C0 , 32'hFCD0AFD4 , 32'hFFCCD710 , 32'h01A5E9FC , 32'hFE984E98 , 32'h00639712 , 32'hFF86C012 , 32'hFE246F14 , 32'hFD0313F0 , 32'h01524888 , 32'hFF56C95D , 32'hFFB0D9DD , 32'h022B91E4 , 32'hFC7882C4 , 32'hFE81835C , 32'hFFEC2720 , 32'h019F6CEC , 32'h00291A2B , 32'h00BADBA3 , 32'hFEC661A4 , 32'h0259DA60 , 32'hFFB248EA , 32'h01622EDC , 32'hFFA2E0E0 , 32'h01CC5A10 , 32'hFFD44118 , 32'h001296AB , 32'h0050E867 , 32'h003FB5C3 , 32'h032D9C1C , 32'hFE43FC24 , 32'h0464ED88} , 
{32'hFFFA487F , 32'hFFF235DB , 32'hFFFA91CD , 32'h04BBAA28 , 32'h0B4CBDA0 , 32'h000036C0 , 32'hFFFE1910 , 32'h000598B6 , 32'h184A8760 , 32'h0000DE04 , 32'hFFF9BDEA , 32'h0000ACEE , 32'hFFFDE938 , 32'h0008BD50 , 32'hFFFD55CF , 32'h0001C445 , 32'hFFFB978F , 32'h00030E60 , 32'h0002DA89 , 32'hE35A7AE0 , 32'h00009D20 , 32'hFFFB5DC2 , 32'h000214B7 , 32'h07B9A560 , 32'h00045D3F , 32'hFFFA5CC7 , 32'h00039964 , 32'h00032437 , 32'h0005B2DB , 32'h00072B15 , 32'h00000118 , 32'hFFFFEC37 , 32'hFFFD6D6F , 32'hFFFDA152 , 32'hFDEBB17C , 32'hFFFFD856 , 32'h0006E500 , 32'h00000C37 , 32'hFFFDC68C , 32'hFFFB6C05 , 32'h000007B0 , 32'hFFC2416E , 32'h0001A3F3 , 32'hFFFE4677 , 32'hFFFA00E4 , 32'h000628BF , 32'h0000BA1B , 32'hFFFED393 , 32'hFFF7D495 , 32'h00089CD8 , 32'h000099B2 , 32'hFFFBCDC6 , 32'h00085BF0 , 32'h0001D982 , 32'h001121AC , 32'hFFFB944C , 32'h000018E9 , 32'h00056CA7 , 32'h00047998 , 32'hFFFC865B , 32'hFFFEBA35 , 32'h0004A511 , 32'h00000C9C , 32'hFFF0F5C3 , 32'hFFFD4A9C , 32'hFFF8FF14 , 32'hAC471F80 , 32'hFFFB30D4 , 32'hFFE84BF7 , 32'h0002FF45 , 32'h0007DAC4 , 32'hFFFF5BF8 , 32'hFFF991C6 , 32'h00054E13 , 32'h0002EFE2 , 32'hFFFF507B , 32'hFFFE8226 , 32'hFFFC3D8C , 32'h00023F26 , 32'h0003A7E0 , 32'hFFFA6683 , 32'h00053973 , 32'h0002930F , 32'h13D51F60 , 32'hFFFD4844 , 32'hFFFAC159 , 32'hFFFF93A2 , 32'h000BA884 , 32'hFFFFDEB3 , 32'hBA50BF80 , 32'hFFFBA6C3 , 32'h0012EE68 , 32'h00063C3C , 32'h00013414 , 32'hCB68C5C0 , 32'hFFFDFD6F , 32'hFFFFDC20 , 32'hFFFC31DC , 32'hFFF93FC8 , 32'h00092DA6} , 
{32'hFFF89248 , 32'hFFF8E55E , 32'h00041447 , 32'hCE0CFD00 , 32'h473DF080 , 32'hFFFE271B , 32'h0001C850 , 32'hFFFD8DCF , 32'hDD842D00 , 32'hFFFCD0B4 , 32'hFFFD017D , 32'hFFFDA66F , 32'h0000C272 , 32'h00026849 , 32'h0004F16E , 32'hFFFABA28 , 32'hFFFC63C3 , 32'hFFFAE177 , 32'h0002E3D8 , 32'h2AC60B00 , 32'hFFFE7BEA , 32'h0002435D , 32'h000211E3 , 32'h3986F900 , 32'hFFFF7F69 , 32'h00000360 , 32'hFFF87317 , 32'h0005AB08 , 32'hFFFC3928 , 32'hFFFCDCFE , 32'h000403E5 , 32'h00003646 , 32'hFFF79498 , 32'h00020F94 , 32'hFF84830F , 32'h00030755 , 32'hFFFAE146 , 32'hFFFB11AA , 32'h00002F1F , 32'h00052BC6 , 32'hFFFCE9EC , 32'hFFFD809B , 32'h00052025 , 32'hFFFF0279 , 32'h0000C80B , 32'h0001A161 , 32'h0002B234 , 32'h000276D3 , 32'h0007EC35 , 32'hFFFFC552 , 32'h00022AB5 , 32'h0001B2A2 , 32'h0001B5B3 , 32'hFFFE4412 , 32'h0003F740 , 32'h000A26F5 , 32'h0006C871 , 32'h00004E38 , 32'hFFFCDF7D , 32'h00010C48 , 32'h0002EE57 , 32'hFFFF75B4 , 32'h00038709 , 32'hFFFAF56A , 32'h00049C22 , 32'hFFFF44C5 , 32'hD8AEC480 , 32'h0003691B , 32'h00016D7E , 32'h00051BB1 , 32'h0006CD52 , 32'h00015BAF , 32'h000227CB , 32'hFFFA0693 , 32'hFFFC29E4 , 32'hFFFE6F4E , 32'h000C768F , 32'h0002338D , 32'h00017104 , 32'hFFFFF7D4 , 32'hFFF438C8 , 32'hFFFE9816 , 32'hFFFF5F8F , 32'h0DF41EB0 , 32'hFFF4E4DF , 32'h00043C42 , 32'h00050907 , 32'hFFFD1007 , 32'h0001182A , 32'h0F043AD0 , 32'hFFFD0333 , 32'h0000D048 , 32'hFFFF8D60 , 32'h0003FD6D , 32'h1C02BA60 , 32'h00000930 , 32'hFFFBE7ED , 32'h000003E3 , 32'hFFF9DD13 , 32'h0001711A} , 
{32'hFFF84426 , 32'h0002BEE3 , 32'h0002CDDE , 32'hC20B9FC0 , 32'hC1A1D200 , 32'h00099B15 , 32'hFFF24196 , 32'h000342F0 , 32'h288F2BC0 , 32'hFFFFD816 , 32'h0002BAB4 , 32'h0001855E , 32'hFFFF6B06 , 32'hFFFC1813 , 32'h00033BAB , 32'h00031EDB , 32'hFFF97266 , 32'h00014009 , 32'hFFFCDAD0 , 32'h09D01450 , 32'hFFFC9835 , 32'hFFFF93CA , 32'h000F0247 , 32'h1329AD80 , 32'h00002BA0 , 32'h0001BCEE , 32'hFFFB0779 , 32'h0003E4C3 , 32'hFFFBC1B1 , 32'hFFFB8DEC , 32'hFFFDA79F , 32'hFFFFDD1E , 32'hFFFE581F , 32'hFFFC91D9 , 32'h29CA4880 , 32'h0000189C , 32'hFFEF14AD , 32'h00004439 , 32'hFFF9E047 , 32'h00048C3F , 32'h0004B87D , 32'hFFA7B9A0 , 32'h000EB17B , 32'h00009528 , 32'hFFFE9065 , 32'hFFFE8DF0 , 32'h0007BCFF , 32'hFFFD05FC , 32'hFFFE6B66 , 32'hFFFCAC18 , 32'hFFFAD54C , 32'h0000C3FC , 32'h00083967 , 32'hFFFC5A92 , 32'h0001D042 , 32'h0004D921 , 32'h000165DE , 32'hFFF73C81 , 32'hFFFA6991 , 32'h000704C9 , 32'hFFFB6801 , 32'h000869F6 , 32'h0003EAE8 , 32'hFFF37551 , 32'hFFFA29CA , 32'hFFFFC8F2 , 32'hEDE8EC40 , 32'h00027509 , 32'hFFFDFC6D , 32'h00074A4A , 32'hFFFDCAB0 , 32'hFFFC4860 , 32'hFFF79E7C , 32'hFFFD7669 , 32'h00047E36 , 32'h0006F354 , 32'h0008240E , 32'h00038EB0 , 32'hFFFCF9A1 , 32'hFFFD5785 , 32'h0003B213 , 32'h0001E023 , 32'h0004BEB2 , 32'hDE95A680 , 32'hFFF861CC , 32'hFFF94649 , 32'h00004AEC , 32'h000745E3 , 32'hFFF97AD3 , 32'hE1A8A940 , 32'hFFFEDFF9 , 32'h00076A99 , 32'h00052D5E , 32'h000696B3 , 32'h33FA32C0 , 32'hFFFD1176 , 32'h0000EAC9 , 32'hFFFC265C , 32'hFFF92987 , 32'hFFF97554} , 
{32'hFFFBC7A4 , 32'hFFFFA589 , 32'hFFFFA5A9 , 32'h12A27D40 , 32'hE2A43CE0 , 32'hFFFDE8C4 , 32'h0001DEC1 , 32'h00076731 , 32'hE386BBC0 , 32'hFFFBA693 , 32'hFFFCCDE9 , 32'h0005159E , 32'hFFFF080E , 32'h0001ADF6 , 32'h00017229 , 32'h0002B7DB , 32'h00021C08 , 32'hFFFDC08E , 32'h00026E97 , 32'hF82C4018 , 32'h0000ED49 , 32'h000556AB , 32'h000B7118 , 32'hD673E8C0 , 32'hFFFF25AB , 32'h00098ED2 , 32'hFFFE76E4 , 32'h00061BFD , 32'hFFFB7B05 , 32'hFFFDDC7E , 32'hFFF836EF , 32'h00020D26 , 32'h00045BC2 , 32'h0004C0EA , 32'hCCA77D80 , 32'h000423A3 , 32'hFFF90923 , 32'hFFFEF0D7 , 32'h00039660 , 32'hFFFFBD26 , 32'h0000A737 , 32'h001CF96A , 32'hFFEE6CF6 , 32'h0001948F , 32'hFFFC5043 , 32'hFFFA56D7 , 32'h000552E4 , 32'hFFFA1F7E , 32'hFFFCABA9 , 32'h000583ED , 32'hFFF91D01 , 32'hFFFC444E , 32'h0005ABAD , 32'hFFFF5118 , 32'h0000C2D4 , 32'h00009397 , 32'h0004B4F7 , 32'hFFF8E3AC , 32'hFFF65726 , 32'h0010D1A1 , 32'h00021DB8 , 32'h0000CF2C , 32'h000A0FA0 , 32'h0002AE02 , 32'hFFFDA3EC , 32'hFFFB4575 , 32'hB27C9900 , 32'h00019315 , 32'hFFF8BEE2 , 32'h00038D1B , 32'h00047A6A , 32'h0006969F , 32'hFFFADB16 , 32'hFFFB2C9B , 32'h00082496 , 32'h00014516 , 32'h00021B31 , 32'h0000B149 , 32'hFFFA136E , 32'hFFFE8275 , 32'h0001248F , 32'h0005182B , 32'h0002B81B , 32'hED6E8A20 , 32'h00013E25 , 32'hFFFC9B7E , 32'h0009C3FD , 32'hFFFD66BF , 32'h00048EDE , 32'h24E6CE80 , 32'hFFFE0F48 , 32'h0001BF4A , 32'h000A75EF , 32'h00004760 , 32'h31E83DC0 , 32'hFFFF093A , 32'h0002E30C , 32'h00004B65 , 32'hFFF83B62 , 32'hFFFF2EA0} , 
{32'hFFF9508F , 32'h00068E71 , 32'h00010609 , 32'hEDF82B80 , 32'h37337E40 , 32'hFFFAFD7D , 32'h00052D4F , 32'hFFFB3AF2 , 32'h4F442500 , 32'hFFFCF30E , 32'h00016755 , 32'h0002A5B7 , 32'hFFFC5178 , 32'hFFFF10E3 , 32'hFFF9C941 , 32'h0000D45C , 32'h0008FBA4 , 32'h0003BA0B , 32'h00019AFB , 32'hC8915140 , 32'h0005C2B8 , 32'hFFFFC036 , 32'h00003B26 , 32'hF0EDD380 , 32'hFFFD08C6 , 32'h00016D9B , 32'hFFFD2FD1 , 32'hFFF8C376 , 32'h0007A1E5 , 32'h0004990D , 32'hFFFCE993 , 32'h00017987 , 32'hFFFEBF45 , 32'h0000766B , 32'h07E283D0 , 32'hFFFF88CE , 32'h000554D3 , 32'hFFFD9D0A , 32'h0000AA92 , 32'hFFF5E870 , 32'hFFFC9A5A , 32'h00240343 , 32'h00036A61 , 32'h0005A18D , 32'hFFFD579B , 32'h000C951A , 32'h0001CD84 , 32'h00069843 , 32'hFFF8CAAB , 32'hFFFE4109 , 32'hFFFC302E , 32'hFFFCE11E , 32'hFFF8C70D , 32'h000C2F98 , 32'hFFFFE030 , 32'hFFF80A8D , 32'hFFFD9402 , 32'hFFFD7C6B , 32'hFFF990A5 , 32'hFFFABB5C , 32'hFFFDE8C9 , 32'h00036847 , 32'hFFF711E7 , 32'h0000D1E0 , 32'h00001095 , 32'h00046327 , 32'hF6B3FF70 , 32'hFFFFE8EC , 32'h0007A59D , 32'hFFF43CD1 , 32'hFFF8533F , 32'h00032351 , 32'h0001AF73 , 32'hFFF6AACA , 32'hFFF94FA2 , 32'hFFF4055E , 32'h0000A5D2 , 32'hFFFF4144 , 32'hFFF4F014 , 32'hFFFBA797 , 32'h0002A839 , 32'h00026CBD , 32'hFFFD4D35 , 32'hEB6B3CC0 , 32'h0003FDFE , 32'h0001D7E1 , 32'h00047DE3 , 32'hFFFF18FA , 32'h0004B40F , 32'h373EB180 , 32'h000818DD , 32'h00068C8C , 32'hFFF97C10 , 32'h00034788 , 32'h085B1300 , 32'h0006B5C7 , 32'h0004D56D , 32'h0002B322 , 32'h00007763 , 32'h00036E55} , 
{32'hFFFC5AD7 , 32'h0000EFE5 , 32'hFFFF8D34 , 32'h0BCAE460 , 32'h26A56E40 , 32'hFFF67798 , 32'h000236F5 , 32'h00023071 , 32'h1F03AEA0 , 32'h0004AEF0 , 32'hFFFEA00E , 32'h00001C5D , 32'hFFFB4904 , 32'h00012F21 , 32'hFFFFA4FC , 32'hFFFEF6E9 , 32'hFFFE9AC7 , 32'hFFFB7B99 , 32'h00000EC1 , 32'h0C21A470 , 32'h0002AEDD , 32'hFFFE13C3 , 32'hFFFE722B , 32'hF6CBC8B0 , 32'h0003414F , 32'hFFF9D9BB , 32'h00066424 , 32'h0001E83A , 32'h00059A4F , 32'h000711AF , 32'h00059019 , 32'h00024E47 , 32'hFFFEABDA , 32'h000278A6 , 32'hB9DF2F00 , 32'hFFFCB1BA , 32'hFFF66AB4 , 32'h0001788D , 32'hFFFE8706 , 32'hFFFA2756 , 32'h00007004 , 32'h0023C43E , 32'h000439B3 , 32'h0000CB3B , 32'h0000427F , 32'h00025389 , 32'h000940AC , 32'hFFFE1366 , 32'hFFFCB807 , 32'h00005AAD , 32'h0005DE22 , 32'h00005E2D , 32'hFFFDDD46 , 32'h0001B10B , 32'hFFFB6114 , 32'h0000DAB0 , 32'hFFF9D70A , 32'hFFFF9FC8 , 32'hFFFDE1D4 , 32'h00052347 , 32'h0008C63D , 32'hFFF4721B , 32'h00016D0B , 32'hFFFE36DB , 32'h00004D42 , 32'h000294A0 , 32'h20124C40 , 32'h0002F7CF , 32'h0005BEC9 , 32'h0006D7A2 , 32'h0001966A , 32'hFFFA03D2 , 32'h0000C079 , 32'hFFF6AD84 , 32'hFFFAE618 , 32'h00021807 , 32'hFFFC154B , 32'h0001B4B3 , 32'h00029345 , 32'h0002FD79 , 32'hFFFCA642 , 32'h0002CF61 , 32'hFFFD9ACB , 32'hEC913B60 , 32'h000069A0 , 32'hFFFB5FB5 , 32'h0003E9C3 , 32'hFFFBC942 , 32'hFFFBD431 , 32'hBAB4D080 , 32'h00053B8C , 32'hFFF8C6A6 , 32'hFFF90D0B , 32'h000472AC , 32'h33EF1800 , 32'hFFFC92C9 , 32'hFFFCE09B , 32'hFFFC5E08 , 32'h0008FDFA , 32'hFFFE46AA} , 
{32'hFFFF33ED , 32'hFFF63023 , 32'h000039CB , 32'hBECD5580 , 32'h02D029B0 , 32'hFFF4C43E , 32'h0003A88E , 32'h000408F9 , 32'hEFA9EB60 , 32'hFFFEE2E6 , 32'h00067193 , 32'h0004727A , 32'hFFFD8BD3 , 32'hFFFB49C3 , 32'h00059494 , 32'hFFF9CD5F , 32'h0002B134 , 32'h00020132 , 32'hFFFD19E9 , 32'hE74A9660 , 32'hFFFFD76E , 32'hFFFD7A19 , 32'h0005652D , 32'hBDA7BE00 , 32'h00004622 , 32'h00000158 , 32'hFFFEFB89 , 32'h00024024 , 32'h0002926B , 32'hFFFACF63 , 32'h000167E2 , 32'h0003F6A2 , 32'hFFFE4023 , 32'hFFFBBC82 , 32'hFE459878 , 32'h00019841 , 32'hFFF98FBE , 32'hFFFD647D , 32'h00056DC0 , 32'h00025165 , 32'hFFFC3DDF , 32'h00208A78 , 32'h000EA8D6 , 32'h000719DC , 32'hFFFE516F , 32'h0002DC67 , 32'hFFFA2239 , 32'h0001890C , 32'hFFFC23B3 , 32'hFFFCAF96 , 32'h00011405 , 32'h0005014B , 32'h00025BD2 , 32'hFFFC81FA , 32'h000B5460 , 32'h000CF8BE , 32'hFFFEDC23 , 32'h00003053 , 32'hFFFD7AA5 , 32'h00022BA0 , 32'hFFFE6B53 , 32'h0001F209 , 32'h0004246E , 32'h0003F239 , 32'h00025A33 , 32'h00028DE4 , 32'h0DDDCB30 , 32'hFFFFC8D2 , 32'hFFEEA9FB , 32'hFFFD9730 , 32'hFFFFC12F , 32'hFFFEF04A , 32'hFFFFF681 , 32'hFFFB1A8E , 32'hFFFE4728 , 32'hFFF8F68D , 32'hFFFE67BD , 32'h0001C005 , 32'hFFFD457A , 32'hFFFB4CDC , 32'hFFFE9F03 , 32'hFFFF2FD4 , 32'hFFF480D0 , 32'h502EB880 , 32'hFFFDED25 , 32'h0000E672 , 32'hFFF15DA4 , 32'h0000D849 , 32'hFFF9DADE , 32'hF24B03C0 , 32'hFFFB36C4 , 32'hFFFDC948 , 32'hFFFE311B , 32'h000305A0 , 32'h114C3600 , 32'hFFFF4608 , 32'h0003621E , 32'h000679FA , 32'hFFFC9389 , 32'h00049103} , 
{32'hFFFD24DB , 32'hFFFA520E , 32'hFFFD48A5 , 32'h20C40100 , 32'h07D3A360 , 32'h000C4E48 , 32'h0002B8A0 , 32'hFFFD88CD , 32'h35557580 , 32'h0004150D , 32'h00073F7E , 32'hFFFC91D2 , 32'hFFFE4DAB , 32'hFFFD79EB , 32'h000319A7 , 32'h000B22B5 , 32'hFFFF9840 , 32'hFFFFD70A , 32'hFFFF3EC5 , 32'h5AD71800 , 32'h00009E61 , 32'hFFF78881 , 32'hFFFDDB81 , 32'hD49AC3C0 , 32'h00009419 , 32'h0004C511 , 32'hFFF4AE4B , 32'h000D1DE5 , 32'hFFF9D86A , 32'h00036DB9 , 32'hFFFE11BE , 32'hFFFA3881 , 32'hFFFFD856 , 32'h0000200D , 32'h1C8D7A80 , 32'h000297E1 , 32'h00019376 , 32'h0003E8F7 , 32'hFFFC366D , 32'h000B9C9A , 32'h00004DC0 , 32'hFFDF805E , 32'h00031CEE , 32'h000752C7 , 32'hFFFBFD13 , 32'hFFFCDDC7 , 32'hFFF71BF0 , 32'h00014D99 , 32'h0004DB16 , 32'hFFFE6762 , 32'h00067FDC , 32'h000151C0 , 32'h000987C4 , 32'hFFFA2139 , 32'h0002CC8D , 32'hFFFAF34C , 32'hFFFED965 , 32'h000607B7 , 32'h0000D77B , 32'hFFFFC222 , 32'hFFFFAE77 , 32'hFFF543B6 , 32'hFFFCF87B , 32'hFFFD33C9 , 32'h0002D435 , 32'h00003129 , 32'hEBAC3A80 , 32'hFFFE9C7F , 32'h0011C8F1 , 32'h000589A7 , 32'hFFFE28B7 , 32'hFFFB4682 , 32'hFFFE0C94 , 32'hFFFF4C72 , 32'hFFFE1558 , 32'h000B6C82 , 32'h000303F5 , 32'hFFFCB5D8 , 32'h000255E7 , 32'h0007B175 , 32'h0005F716 , 32'h0001FDB3 , 32'hFFFDD1A7 , 32'h2266FFC0 , 32'hFFFAC839 , 32'h00019F8E , 32'h000136CD , 32'hFFFE7133 , 32'h00033704 , 32'h0A667B90 , 32'h00061A60 , 32'h0008A905 , 32'h0004DA00 , 32'hFFFA6DC3 , 32'h03D55DB4 , 32'hFFFEDC51 , 32'h0003378B , 32'hFFFBE045 , 32'h0000DE5A , 32'h0000D0C6} , 
{32'hFFFE9716 , 32'hFFF98736 , 32'h000545A0 , 32'hDDC9BD00 , 32'h20588F00 , 32'h0005C693 , 32'hFFFFA323 , 32'h00016807 , 32'hDEAF4C00 , 32'h00036B4B , 32'hFFF95FC1 , 32'h00023300 , 32'hFFF8CBFF , 32'hFFFC2BFB , 32'h0006729C , 32'hFFFD01FB , 32'hFFFA0B16 , 32'h00004813 , 32'hFFFD8FDB , 32'h16E5C1C0 , 32'h00064D7B , 32'h0004873E , 32'hFFF7E390 , 32'hBD070780 , 32'hFFFD7A14 , 32'hFFFC60A0 , 32'h00059AA9 , 32'hFFFFE2DB , 32'h00059DFD , 32'hFFFFE746 , 32'hFFFE8E3C , 32'h0003C739 , 32'hFFFE0A32 , 32'hFFFF01C5 , 32'h166C94A0 , 32'h0004E090 , 32'h000AF424 , 32'h000622D5 , 32'hFFFA1ED8 , 32'hFFFEDE4B , 32'hFFFBFBA8 , 32'hFFEC1BEC , 32'h0003BBBA , 32'hFFF958BF , 32'hFFF9F76C , 32'hFFFC437E , 32'hFFFAC74A , 32'h00027A63 , 32'hFFF9E423 , 32'h00054A3E , 32'hFFFF327B , 32'hFFFF0992 , 32'hFFFF968B , 32'h0006A519 , 32'h00082137 , 32'hFFF3D8BD , 32'hFFFB76EC , 32'hFFFF5346 , 32'h00068BE7 , 32'hFFF8E000 , 32'hFFFDC44F , 32'hFFFE49CF , 32'hFFFC5D58 , 32'h0001DA08 , 32'h0001BD1E , 32'hFFFEEF07 , 32'hFD752D3C , 32'hFFF962C0 , 32'h00177EB0 , 32'hFFFE1787 , 32'h0006D6AC , 32'h0005D5FF , 32'hFFFEFFF0 , 32'h000B0024 , 32'hFFFCA915 , 32'hFFFBC60E , 32'hFFFFB4B9 , 32'hFFFD8127 , 32'h00059FEF , 32'h0005339C , 32'hFFFC53A4 , 32'h000107AF , 32'hFFFA7E4A , 32'hB1656780 , 32'hFFFED99A , 32'h0003D010 , 32'hFFFF82CF , 32'h00034893 , 32'hFFF6A810 , 32'hED872480 , 32'h0001475E , 32'h00044F3E , 32'h0009360F , 32'h0005EDD0 , 32'hDC2AEAC0 , 32'h00001092 , 32'h00036BED , 32'hFFFFF8DD , 32'h0007AAD6 , 32'h0003691A} , 
{32'hFFFE6179 , 32'h0001E8F8 , 32'h000386B6 , 32'h36A82100 , 32'h20395B00 , 32'h00063E77 , 32'hFFF5CA4C , 32'hFFF9C617 , 32'hE135BE60 , 32'h0003977F , 32'hFFFCCE53 , 32'hFFFDC950 , 32'hFFFD8975 , 32'h00021078 , 32'hFFFFEDDC , 32'hFFFF6D72 , 32'hFFFFEB20 , 32'h00008F2E , 32'hFFFA9706 , 32'hDCDC0680 , 32'h0005D891 , 32'hFFFACA8F , 32'h00058D74 , 32'hF5C204D0 , 32'hFFFEF93A , 32'h00028FBA , 32'h000047FD , 32'hFFFD94DC , 32'h0000C763 , 32'h0000CDC7 , 32'h00021840 , 32'h00007D98 , 32'h0004F1FE , 32'h000206BD , 32'h4D344A80 , 32'hFFFFEED4 , 32'h0002DA06 , 32'hFFFB6B15 , 32'hFFF814D3 , 32'hFFFB7FEE , 32'hFFFE832C , 32'hFFA1B331 , 32'hFFF694DA , 32'hFFFF9893 , 32'hFFFF9E02 , 32'hFFFE2CC2 , 32'h00036F10 , 32'h0005ADE8 , 32'h000002EC , 32'h0003062A , 32'hFFF7B094 , 32'hFFFB551E , 32'hFFFB5D60 , 32'hFFFCF45A , 32'h0007AABA , 32'hFFF55429 , 32'hFFFE09EF , 32'h00036664 , 32'hFFFAE0D4 , 32'h0005CAD8 , 32'h0003DD50 , 32'hFFFED0B8 , 32'hFFF88239 , 32'h00004A01 , 32'hFFFCFFCF , 32'hFFFE2158 , 32'hFA63BE48 , 32'hFFF973F6 , 32'h0010CA66 , 32'h0003553A , 32'hFFFE33B7 , 32'hFFFEDBFF , 32'h000513D6 , 32'hFFF7D254 , 32'h00000AFE , 32'h0005FB82 , 32'h00076BD2 , 32'h00032ECF , 32'h0001E8DB , 32'hFFFFE4ED , 32'hFFFB59B3 , 32'h0004FD71 , 32'hFFFDF017 , 32'h02B69148 , 32'hFFFC7A7C , 32'h0002EEE4 , 32'h0006B2F1 , 32'hFFFDF78E , 32'hFFFE14F1 , 32'hE3CFC400 , 32'h00034104 , 32'hFFFDBC9F , 32'hFFFF50FD , 32'h00004A21 , 32'h3B8327C0 , 32'hFFFCFF49 , 32'hFFFEC284 , 32'hFFFD3F76 , 32'h00051819 , 32'h00040862}
};

logic signed [31:0] VT_3 [10][10] ='{
{32'hB2067880 , 32'hBD469900 , 32'h1452A4A0 , 32'h36BD7880 , 32'h06931100 , 32'hFABEFA78 , 32'hA4B4E200 , 32'h2FB52B00 , 32'hFEC60BE8 , 32'h302908C0} , 
{32'h34628EC0 , 32'hA7DC8D00 , 32'h0B5F7AA0 , 32'h36A12040 , 32'hD221D9C0 , 32'h17886B00 , 32'h094EBB20 , 32'hC06C47C0 , 32'h4FCFC500 , 32'hF34B58C0} , 
{32'hB99F6C00 , 32'h27F40800 , 32'h028C4248 , 32'h419D3000 , 32'hCA85AAC0 , 32'h20F81000 , 32'h1D2A9EC0 , 32'h20E708C0 , 32'h0B6A8440 , 32'h9BA33B80} , 
{32'h4EBBB180 , 32'h05AABB70 , 32'h05C769A8 , 32'h2FD13500 , 32'h074D6628 , 32'h955A3680 , 32'hE6351760 , 32'h40396A80 , 32'h036EA5A8 , 32'hD17AA700} , 
{32'h2A435600 , 32'hD6E785C0 , 32'hB89D7280 , 32'h0E0C0A70 , 32'hC624B5C0 , 32'h2DF93280 , 32'h2ACFFE80 , 32'h4F7D3B00 , 32'hC941D900 , 32'h2794AD40} , 
{32'h0E37A0F0 , 32'hD5C74280 , 32'h7FFFF880 , 32'hCDC13600 , 32'hD5D46680 , 32'h0A3A5CD0 , 32'h0F073060 , 32'h199C2280 , 32'hCBD09040 , 32'hE847CA40} , 
{32'h1C1D0E80 , 32'h28068640 , 32'h09BA2650 , 32'h482A7380 , 32'hE0D64980 , 32'h07ECC888 , 32'hD5008640 , 32'hB1D84280 , 32'h9B98F080 , 32'h0D5102C0} , 
{32'h05E8A340 , 32'h434AAC00 , 32'h07F6B4E0 , 32'hDD88E4C0 , 32'h8F8C2800 , 32'hEF660420 , 32'hD0126C80 , 32'h0BBDB2D0 , 32'h383C3BC0 , 32'h33193000} , 
{32'h32DF21C0 , 32'h0530E2E8 , 32'hEC13B5C0 , 32'hDA9ACB80 , 32'h16159A20 , 32'h56314880 , 32'h9B8D1580 , 32'h1491AC80 , 32'h060059C0 , 32'hC03887C0} , 
{32'h2793A8C0 , 32'h3AE03C40 , 32'h41C78A80 , 32'h3E175C40 , 32'h33832580 , 32'h3E943C40 , 32'h1AB000E0 , 32'h2A216140 , 32'h25D4F840 , 32'h38EDC080}
};

logic signed [31:0] US_0 [784][37] ='{
{32'hFFFB507D , 32'h0000A155 , 32'hFFFE30CD , 32'hFFF56C3D , 32'hFFFE0623 , 32'h0000D612 , 32'hFFFF5106 , 32'hFFFFC67E , 32'h0001CE1E , 32'h000078CA , 32'h0000F761 , 32'h000181DF , 32'hFFFF48AF , 32'hFFFD87E0 , 32'hFFFDEC83 , 32'h00022293 , 32'hFFFE97FA , 32'hFFFCF205 , 32'h00094A29 , 32'hFFF9D5E6 , 32'h0002D1A9 , 32'hFFFA2B6A , 32'hFFFDE897 , 32'hFFFD6421 , 32'h00008EBE , 32'hFFFE8AE0 , 32'hFFFB8102 , 32'h00085AB9 , 32'hFFFD7A29 , 32'hFFFF4A4C , 32'hFFFEA6E2 , 32'hFFFBFA0B , 32'hFFFFF117 , 32'h0000BF1F , 32'h0001FC0D , 32'h000209B3 , 32'hFFF8EF0B} , 
{32'h00013FF1 , 32'h0002A0E4 , 32'hFFFB2A7A , 32'h000A4441 , 32'h0003D5C4 , 32'hFFFD4D41 , 32'h0002033E , 32'hFFFE0ED8 , 32'h0004002F , 32'h0000532E , 32'h0003A93A , 32'h0002F9FA , 32'hFFFEF6E3 , 32'h00034430 , 32'hFFFD9CD0 , 32'hFFF8CCF9 , 32'hFFFBB974 , 32'hFFFD7DED , 32'h00015799 , 32'h00023B1F , 32'hFFFFBA4D , 32'h000156CF , 32'h00029107 , 32'hFFFB22BA , 32'h00059B24 , 32'h000061FF , 32'h0004FFA6 , 32'h0000B9EB , 32'hFFFFF9D5 , 32'hFFFE947E , 32'hFFFDDC61 , 32'h00011800 , 32'h000339B5 , 32'hFFFB5CA5 , 32'hFFFF9736 , 32'hFFFCAB67 , 32'hFFF9F0CA} , 
{32'hFFFAD66D , 32'hFFFE3CEE , 32'hFFFE3EF0 , 32'h00067DD7 , 32'hFFFECE85 , 32'h00061A9E , 32'hFFF9D4FB , 32'hFFFE6DB7 , 32'hFFFEB58D , 32'hFFFD5473 , 32'hFFFFEC81 , 32'hFFFC8BE4 , 32'h0001BE6B , 32'h0000058C , 32'h0007720F , 32'hFFFEA0D2 , 32'h0000191E , 32'h00046089 , 32'h000039C1 , 32'hFFFE3212 , 32'h0000E1E1 , 32'hFFFEC4C9 , 32'hFFF7DE62 , 32'hFFFD21E3 , 32'hFFFDFA2C , 32'hFFFD42F4 , 32'h0002F8BB , 32'h000123C2 , 32'hFFFE8155 , 32'h0002EED9 , 32'h0005BB52 , 32'hFFFDBA76 , 32'hFFFC1D7E , 32'hFFFF0C3A , 32'hFFFA7667 , 32'hFFFD03D1 , 32'h0005F5AD} , 
{32'hFFFC8778 , 32'h0004D755 , 32'hFFF857E6 , 32'hFFFDB807 , 32'h00012615 , 32'h00004C65 , 32'hFFFA3BF9 , 32'hFFFEA7AE , 32'h0005CE05 , 32'hFFFD8FC7 , 32'hFFFF8CF3 , 32'h00007273 , 32'h00006474 , 32'hFFFFA839 , 32'hFFFA2DC8 , 32'h000C04A3 , 32'h00005208 , 32'h00023C9D , 32'hFFFE6DAB , 32'hFFF9D810 , 32'h0000B88F , 32'h0005E6FF , 32'h000588A3 , 32'hFFFEE786 , 32'hFFFE983A , 32'hFFFEA1F1 , 32'h000249F5 , 32'h0003859D , 32'hFFFCF0E7 , 32'h00019635 , 32'hFFFF8D5C , 32'h000052B4 , 32'h0002BC0B , 32'hFFFD7377 , 32'h000043A8 , 32'hFFFFA2D5 , 32'h0001E88A} , 
{32'hFFFF9600 , 32'h000112F5 , 32'hFFFDDF07 , 32'hFFFE8C33 , 32'hFFFFA1EB , 32'h00068716 , 32'h0004E48C , 32'h0000764B , 32'h000210D1 , 32'hFFFC154B , 32'hFFFD28DE , 32'h0001732A , 32'h00054128 , 32'hFFF81E86 , 32'hFFFF02F2 , 32'hFFFC08A6 , 32'hFFFBED58 , 32'h0000E5FD , 32'h0004EA15 , 32'hFFFE2A69 , 32'hFFFDDC50 , 32'h0006AB83 , 32'h000227B6 , 32'h00018229 , 32'hFFFB2AD3 , 32'h000268A6 , 32'h00025529 , 32'hFFFDE47A , 32'hFFFC6DF7 , 32'hFFFA4A88 , 32'h00043196 , 32'hFFFC96A0 , 32'h00052372 , 32'h000140C4 , 32'hFFFE213A , 32'hFFFE9BC4 , 32'hFFFC395C} , 
{32'h00063B5A , 32'h00088932 , 32'hFFFD2C01 , 32'h0002685C , 32'h000582AF , 32'hFFFCB4FF , 32'hFFFC11AF , 32'h0001CA63 , 32'hFFFF66A6 , 32'h0000A074 , 32'h00051098 , 32'h00017BBF , 32'h00024BCE , 32'hFFFA5902 , 32'h00037242 , 32'h0004C3BF , 32'hFFFFF6CD , 32'h0000A363 , 32'hFFFCC66B , 32'h00073F75 , 32'hFFFD64A5 , 32'h00005D97 , 32'h000154C9 , 32'h0002F2C1 , 32'hFFFD3090 , 32'h00026564 , 32'h00004052 , 32'h00013D88 , 32'hFFFE38F6 , 32'hFFF9513A , 32'h000168C8 , 32'h000051D4 , 32'h0005AF9D , 32'h0000EB7B , 32'h00021FBA , 32'h0002E4F5 , 32'hFFF82B12} , 
{32'h00010C15 , 32'h000182F3 , 32'hFFFF0E90 , 32'hFFFC8B19 , 32'hFFFC6410 , 32'hFFF90F22 , 32'hFFFC62D9 , 32'h00017F95 , 32'h00042669 , 32'hFFFFE287 , 32'h00018351 , 32'hFFFECC5E , 32'h0003D656 , 32'h0002F90F , 32'hFFFAE708 , 32'hFFF81BDB , 32'h00011BA7 , 32'h00003873 , 32'hFFF7FA74 , 32'h0002BCB7 , 32'h0001B612 , 32'h0007E69D , 32'h00012484 , 32'hFFFA3B8B , 32'hFFFCD329 , 32'hFFF8349E , 32'hFFFE7670 , 32'hFFFA1759 , 32'hFFFECA90 , 32'hFFFD7362 , 32'h0000E339 , 32'hFFFF68F2 , 32'h00068C8A , 32'hFFFE18F6 , 32'h000015B2 , 32'h00038DA9 , 32'hFFFF3886} , 
{32'h00016E76 , 32'hFFF9CEED , 32'hFFFB895B , 32'hFFF93AFA , 32'hFFFF5786 , 32'hFFFE09D5 , 32'h00041912 , 32'hFFFC7A62 , 32'h000115BC , 32'h000317AD , 32'hFFF82191 , 32'hFFFED961 , 32'h0002D5A1 , 32'hFFFBD2B8 , 32'hFFFD8DCA , 32'h0001F3AA , 32'h00057DAC , 32'h0000A493 , 32'hFFFC58F8 , 32'hFFFC1D53 , 32'hFFFE4B8B , 32'hFFFEB219 , 32'hFFFEE149 , 32'h000280AA , 32'hFFFC116E , 32'h00008797 , 32'h00048F62 , 32'hFFFC623F , 32'hFFFFDDD2 , 32'hFFFC78BA , 32'h00067DF2 , 32'h0003D494 , 32'hFFFB17E2 , 32'hFFFFFD6D , 32'hFFF749BA , 32'hFFFF4091 , 32'hFFFDF5EA} , 
{32'hFFFB4DE8 , 32'hFFFA9023 , 32'hFFFDC73F , 32'hFFFFACCE , 32'hFFFE3E25 , 32'h0001E205 , 32'hFFFE2BA9 , 32'hFFFB5070 , 32'h00055FAB , 32'hFFFD670A , 32'h0000F952 , 32'hFFFDC978 , 32'h0000F294 , 32'h000248A3 , 32'hFFFA6371 , 32'hFFFE9340 , 32'hFFFBE11B , 32'hFFFF1A1E , 32'hFFFEBC25 , 32'h00013606 , 32'h00031578 , 32'h000046F6 , 32'hFFFFC2AC , 32'h0000F7BF , 32'h00033047 , 32'h00037072 , 32'hFFFB6126 , 32'hFFF9E417 , 32'h00018608 , 32'h0001AA30 , 32'h00007DCE , 32'hFFFCD4F9 , 32'hFFFAC234 , 32'h00007D00 , 32'h00056339 , 32'h00067CC3 , 32'hFFFD4579} , 
{32'h0004C34D , 32'hFFFBE4ED , 32'h00007BD5 , 32'hFFFEEB5B , 32'h000384CE , 32'h00031A98 , 32'h0004D172 , 32'hFFFDD877 , 32'h0004293A , 32'h0002C3D6 , 32'h0000D3D1 , 32'hFFFF9CB4 , 32'hFFFE0A22 , 32'hFFFAA98C , 32'h00032C4B , 32'h000387CB , 32'h0003CD6C , 32'hFFFE442E , 32'h00009450 , 32'h0002213D , 32'hFFFDF27F , 32'h0005BE19 , 32'hFFFD26C1 , 32'h0003780C , 32'hFFFFF08D , 32'h0005BBCE , 32'hFFFDC2F8 , 32'hFFFF2FE6 , 32'h0002A0AB , 32'hFFFFF28E , 32'h0004FE9B , 32'h00024552 , 32'h00002338 , 32'h000404AE , 32'h00030759 , 32'h00051A75 , 32'h0004C44B} , 
{32'hFFFEDF2C , 32'hFFFAD090 , 32'h0000395D , 32'h0002E107 , 32'hFFFFD948 , 32'hFFFBDA87 , 32'h00029074 , 32'h000587EE , 32'hFFFDED70 , 32'hFFFFDE25 , 32'hFFFFB781 , 32'hFFFC603B , 32'hFFFE7DA2 , 32'hFFFDE1D3 , 32'h00038F5F , 32'h00020F6C , 32'hFFFE5A3E , 32'hFFFB4D77 , 32'h0001EACB , 32'hFFFD27A1 , 32'h00010A1F , 32'hFFFEF810 , 32'h0002C696 , 32'hFFFF52EC , 32'hFFFE5A50 , 32'hFFFB56C2 , 32'h00039D3E , 32'h00004EA1 , 32'hFFF74F97 , 32'hFFFF09E4 , 32'hFFFF32FE , 32'hFFFF68DC , 32'h000216F9 , 32'hFFFF8F5E , 32'h0003D146 , 32'hFFFFF0F8 , 32'h00043A8A} , 
{32'hFFFDBBCE , 32'h0003F985 , 32'h0001F75D , 32'hFFFF5E7F , 32'h0001B7C2 , 32'hFFFFCA12 , 32'hFFFB3440 , 32'h0000E567 , 32'hFFFFA0F9 , 32'hFFFE58C3 , 32'h0005428A , 32'hFFFC4EC4 , 32'hFFF9E946 , 32'hFFFC5B1F , 32'h0000C5F9 , 32'hFFFCD2C7 , 32'hFFFDC7DC , 32'h000481D2 , 32'h0002A6CB , 32'h00051DF8 , 32'h000592A5 , 32'hFFFF8978 , 32'h00062CFC , 32'h0000F0BE , 32'hFFFFA161 , 32'h00029F2A , 32'hFFFFF441 , 32'h00021CCF , 32'hFFFC9BB7 , 32'h0003AFB3 , 32'h0002FB0F , 32'h0001565D , 32'h00007AF7 , 32'h0002CDAA , 32'hFFFE1457 , 32'hFFFE2D3E , 32'hFFFFD00D} , 
{32'h000274D5 , 32'h0001DE63 , 32'h00062507 , 32'hFFFDCDE5 , 32'hFFFBCE0B , 32'h0006A547 , 32'h000207AD , 32'hFFFCA7A4 , 32'hFFFDB453 , 32'h0003438C , 32'h00023735 , 32'hFFFFA250 , 32'hFFFA8000 , 32'hFFFCE4BF , 32'h00016A26 , 32'h0000E4CE , 32'h00001BA9 , 32'h0002C149 , 32'hFFFEE97E , 32'h0006DF55 , 32'hFFFDE2DC , 32'h00004330 , 32'hFFFFC8B5 , 32'hFFFD6F8B , 32'h00034A55 , 32'hFFF9C34F , 32'hFFFD83F3 , 32'hFFFD1ACE , 32'h00011F68 , 32'h00040AC2 , 32'h000599DB , 32'h00017A9B , 32'h00049042 , 32'h000285FC , 32'hFFFCC13E , 32'hFFFE908E , 32'hFFFCECF9} , 
{32'hFFFDDF92 , 32'hFFFC71E3 , 32'h00005F89 , 32'hFFFE1BA7 , 32'hFFFECFA7 , 32'h000721F6 , 32'hFFFE872A , 32'hFFF7B21B , 32'hFFFC2D7E , 32'hFFFBD451 , 32'hFFFCD5DC , 32'hFFFE993E , 32'hFFFE7063 , 32'hFFFEC019 , 32'hFFFC6124 , 32'h000212B9 , 32'h00030055 , 32'hFFFF4400 , 32'h0004BE5B , 32'h000261E4 , 32'hFFFF3B7D , 32'hFFFF993D , 32'hFFF9D73C , 32'h0001FA0C , 32'h0000BFE0 , 32'h000499D5 , 32'hFFFCE88D , 32'h0000215B , 32'h00060B4F , 32'h0002F4D0 , 32'hFFFF4C73 , 32'hFFFE3B79 , 32'hFFF70C79 , 32'hFFFFFE7F , 32'h000163C5 , 32'hFFFB860B , 32'hFFFF17BF} , 
{32'h00027D94 , 32'hFFFED277 , 32'h00058308 , 32'h0000D1E7 , 32'h00005846 , 32'h0000E332 , 32'h00004BF7 , 32'hFFFBA9D8 , 32'h0004694C , 32'h0004BB68 , 32'hFFFEE3F8 , 32'hFFFED452 , 32'hFFFC9E6B , 32'hFFFF9C30 , 32'hFFFC8B0F , 32'h000095A1 , 32'hFFFFD9B6 , 32'h000024BE , 32'hFFFAE3DD , 32'h0005BC3F , 32'hFFFDECF1 , 32'h000341B3 , 32'h00021319 , 32'h0000A8D1 , 32'hFFFB67F3 , 32'hFFFFC5C8 , 32'h0001D878 , 32'hFFFD3332 , 32'hFFFD1293 , 32'hFFF9C01D , 32'h0008837D , 32'h0001E243 , 32'hFFFD8ADB , 32'hFFFF421C , 32'h0001765B , 32'hFFFD9BD0 , 32'hFFFCE678} , 
{32'h00020D52 , 32'h0003499E , 32'h00004F2B , 32'h00001B51 , 32'hFFFF003F , 32'h00033A01 , 32'hFFFD7812 , 32'hFFFAE2AA , 32'h000ADA83 , 32'h0002DC38 , 32'hFFFCE6DE , 32'h0004BCAF , 32'hFFFDB7FD , 32'hFFFF7E11 , 32'h00026847 , 32'hFFFF16F3 , 32'h0001116D , 32'hFFFD2CA1 , 32'h0001E26D , 32'h0005E18A , 32'h0005A861 , 32'hFFFFEE80 , 32'h0005458C , 32'h00001FA1 , 32'hFFFF50F9 , 32'hFFFDE5B0 , 32'h0003CAD2 , 32'hFFFED10E , 32'h0003675E , 32'hFFFE06E2 , 32'hFFFF7E4C , 32'hFFFFE4C0 , 32'h000308A4 , 32'hFFFD3F44 , 32'hFFF9FD05 , 32'hFFFC5BC2 , 32'h00050249} , 
{32'h00043FBA , 32'h00061756 , 32'h0006BABD , 32'hFFFFE275 , 32'h000535B6 , 32'hFFFD9267 , 32'h0007478A , 32'h00061C61 , 32'hFFFF6B3F , 32'h000558CC , 32'hFFFFBBA4 , 32'hFFF7A35B , 32'hFFFFB19B , 32'hFFFF26B1 , 32'hFFFC9FC9 , 32'h0000353A , 32'h0004DA82 , 32'hFFFF492D , 32'h00032403 , 32'h0007CB38 , 32'h000432C2 , 32'h00060C08 , 32'hFFFB8844 , 32'h00002700 , 32'h00008017 , 32'hFFF9AB11 , 32'hFFFE3A97 , 32'h0003203A , 32'hFFFF0F72 , 32'h0001750F , 32'hFFFAEE44 , 32'h0001AB92 , 32'h0003F426 , 32'h0000996A , 32'h0001930C , 32'hFFFBE287 , 32'hFFFEE0F1} , 
{32'hFFFD5654 , 32'hFFFFF354 , 32'hFFFFB39A , 32'h00022650 , 32'h00010ECB , 32'h000288F7 , 32'hFFF720BA , 32'hFFFB2C32 , 32'hFFFB762D , 32'hFFFE218E , 32'h000085A9 , 32'h00006881 , 32'hFFFC2A44 , 32'hFFFFF242 , 32'h00002E69 , 32'h00002C52 , 32'h0005506F , 32'hFFFDA822 , 32'h000391EE , 32'h000595F5 , 32'h00015FF0 , 32'h00019CED , 32'hFFFEE744 , 32'hFFFCE16B , 32'h0002A7E0 , 32'hFFFDE4C5 , 32'h0003C934 , 32'h0000894B , 32'h00016633 , 32'hFFFEA56C , 32'h00031D4A , 32'hFFFC8490 , 32'h00026088 , 32'hFFFF047C , 32'hFFFDBB5D , 32'hFFFE874F , 32'h000116DD} , 
{32'hFFFC233E , 32'h0004F769 , 32'h00005A4F , 32'hFFFDC612 , 32'h00022ADD , 32'hFFFC32E1 , 32'hFFFA49EA , 32'h00035B8A , 32'h0005C35B , 32'hFFFEA48A , 32'hFFFDFD87 , 32'h0000A9A2 , 32'h00040C77 , 32'h0001B3C4 , 32'hFFFD8734 , 32'hFFFC47EF , 32'hFFFABFAA , 32'hFFFAEB82 , 32'hFFFF3E01 , 32'h00031E2B , 32'hFFFF3D67 , 32'hFFF984FA , 32'h0001E05D , 32'hFFFC58DF , 32'h000368EA , 32'h00030146 , 32'h00007798 , 32'h00017955 , 32'h0003D2BC , 32'h000024CC , 32'hFFFDEF35 , 32'h0000E609 , 32'hFFFD78EE , 32'h0003565C , 32'h00024FF5 , 32'h00023F28 , 32'hFFFDBA89} , 
{32'hFFFE8838 , 32'h000767BE , 32'hFFFD4276 , 32'h0001BC11 , 32'h000159C6 , 32'h0005A03D , 32'h0003280E , 32'h0000B39E , 32'hFFF6CED3 , 32'hFFFD87CE , 32'hFFFE5951 , 32'h0000FCC1 , 32'h00024588 , 32'hFFFB4DE3 , 32'h000A313D , 32'hFFFEF422 , 32'hFFFF0691 , 32'hFFFCB0A2 , 32'h0002DF07 , 32'h0002EF26 , 32'h00023887 , 32'h0000C179 , 32'hFFFF4F9B , 32'hFFF9C974 , 32'hFFFDD210 , 32'h0001367C , 32'h00028051 , 32'h00038F99 , 32'hFFFF19DC , 32'hFFFE1296 , 32'h00002501 , 32'hFFFD6E20 , 32'h000428CF , 32'hFFF8C22F , 32'h00023D98 , 32'h0004D9D2 , 32'hFFFDE4C8} , 
{32'hFFFFA043 , 32'hFFFB5E89 , 32'h0002290D , 32'h0000AB9D , 32'hFFFE2F5E , 32'hFFFE62E2 , 32'h0000DD76 , 32'h0001AB42 , 32'h00010FB0 , 32'h000508E7 , 32'h00033A82 , 32'h0003FF17 , 32'h0003DEDA , 32'h0000CF76 , 32'h000113E1 , 32'h0008895E , 32'hFFFBB0D5 , 32'h0000F026 , 32'hFFFD8989 , 32'h00017D67 , 32'h000176DE , 32'h00009AC8 , 32'h00062146 , 32'h00003F21 , 32'hFFFF453E , 32'h000148BB , 32'hFFFD0AAA , 32'hFFFE1E93 , 32'hFFFA5B26 , 32'hFFFC63E4 , 32'hFFFF85B6 , 32'hFFFD30C7 , 32'h000493D6 , 32'hFFFEE9BD , 32'h00042FD2 , 32'hFFFD95EE , 32'hFFFFDFF3} , 
{32'h00007D90 , 32'hFFFF1BDD , 32'hFFFFD040 , 32'h000278E4 , 32'hFFFD9389 , 32'hFFF7CE4E , 32'hFFFB0D0F , 32'h0002EA77 , 32'h00033D2D , 32'hFFF653CD , 32'hFFFC7F7C , 32'h0002BF2A , 32'hFFFEDDE1 , 32'h0002371F , 32'hFFFFADD3 , 32'h0000B99D , 32'hFFFB710A , 32'h00003895 , 32'hFFF9FA52 , 32'h0000883A , 32'h0001A2B5 , 32'h0005A1EE , 32'hFFFAC3F4 , 32'h0003509E , 32'h00012BD3 , 32'h0003728A , 32'hFFFF9C00 , 32'h0008356D , 32'hFFFDE015 , 32'h0001DCC8 , 32'h0001EFD2 , 32'hFFF8A12F , 32'hFFFE1C1C , 32'hFFFC3040 , 32'hFFFA654C , 32'hFFFA8B29 , 32'hFFFD6639} , 
{32'h0007A17E , 32'hFFFBAC58 , 32'hFFFC2330 , 32'hFFFFB44F , 32'h000135F3 , 32'h000132E0 , 32'hFFFF937B , 32'hFFFB899B , 32'hFFFA725A , 32'h0003DA20 , 32'hFFFF2CB5 , 32'hFFFFA564 , 32'hFFF9E1DD , 32'h0003AC00 , 32'hFFF92B57 , 32'hFFF965A2 , 32'h00007BBB , 32'h00015E2B , 32'h0005874D , 32'hFFFBC93F , 32'h0002B387 , 32'h00016DBD , 32'h00017B76 , 32'hFFFF62E1 , 32'h000596FE , 32'h00049305 , 32'hFFFD3A2E , 32'h0007BE7C , 32'h0002F91C , 32'hFFFFC321 , 32'h000028BC , 32'h0000874D , 32'h00018A63 , 32'hFFFC9B1B , 32'hFFFA541D , 32'hFFFF86D1 , 32'h000239DE} , 
{32'hFFFDD483 , 32'hFFFD24C9 , 32'hFFFE6CCE , 32'hFFF8FE85 , 32'h0000F977 , 32'h00000BA8 , 32'hFFFF3E0D , 32'h00086FAE , 32'hFFFFB963 , 32'h0002CEAC , 32'hFFFBC863 , 32'hFFFE2B95 , 32'hFFFC309A , 32'hFFFE987D , 32'hFFFBD5C5 , 32'h00016B3E , 32'h0000EDA0 , 32'h0000658A , 32'h00041208 , 32'hFFFEEA0D , 32'h00013120 , 32'hFFFF5FA4 , 32'hFFFFA3D2 , 32'hFFFF5663 , 32'h00015DEB , 32'h0005BAC6 , 32'hFFFFF6E3 , 32'h00003A52 , 32'h00035490 , 32'hFFFF7B2E , 32'h000250EE , 32'h0000CA76 , 32'hFFFD239E , 32'h0005C4E0 , 32'h00033C43 , 32'hFFFF3BB3 , 32'h00003BCD} , 
{32'hFFFC7D6E , 32'h0005F978 , 32'hFFFC1DD7 , 32'h000038FC , 32'hFFFB06BE , 32'h0006F9BA , 32'hFFFF7948 , 32'hFFFB9B52 , 32'hFFFE7A2D , 32'hFFFA11CD , 32'h0000AEB3 , 32'hFFFC3D60 , 32'hFFFE21F0 , 32'hFFFE408E , 32'hFFFFD008 , 32'h00036422 , 32'h0002249A , 32'h00069C9E , 32'hFFFEDC96 , 32'hFFFDD6B6 , 32'h0003A1EC , 32'h00029384 , 32'h0004A5D4 , 32'h000018EB , 32'hFFFBEE26 , 32'hFFFE9229 , 32'h0006C573 , 32'h00030A2E , 32'hFFFB5FD8 , 32'h0005D78D , 32'hFFFE9027 , 32'h0004B047 , 32'hFFFB82FA , 32'h00000E62 , 32'hFFFA7550 , 32'hFFFD3707 , 32'h0001194F} , 
{32'hFFFE7F15 , 32'h00057657 , 32'hFFFB279C , 32'h000183CC , 32'h000177B5 , 32'hFFFD97DC , 32'hFFFFFA4B , 32'hFFFC4884 , 32'h0000FD42 , 32'hFFFE4DF1 , 32'hFFFEAB60 , 32'h00022AAB , 32'hFFFEC6FA , 32'h0001EBCE , 32'h0003EDFD , 32'hFFF8D5A0 , 32'h0000F9BB , 32'hFFFEE15D , 32'hFFFE256D , 32'h0002B25C , 32'h0003134C , 32'h000690CB , 32'h00003CDF , 32'h00015E33 , 32'hFFFEB701 , 32'hFFFDEABC , 32'hFFFC958C , 32'hFFFC374A , 32'hFFFBAEAF , 32'hFFFEC751 , 32'h00041983 , 32'hFFFCB378 , 32'h0000E162 , 32'h00012ADD , 32'h0000D902 , 32'h0000B322 , 32'hFFF92952} , 
{32'hFFFD85E6 , 32'hFFFF945B , 32'hFFFB0109 , 32'h0001B1F9 , 32'h0000946E , 32'hFFFBCCCD , 32'h0002494D , 32'hFFFE1B9B , 32'h00007D4B , 32'hFFFDE5A1 , 32'hFFFE364F , 32'hFFFBDBFF , 32'h0002F5EC , 32'h0004FBAC , 32'h000106E5 , 32'h00044F9C , 32'hFFFFC38D , 32'h00054785 , 32'hFFFEB366 , 32'hFFFA9029 , 32'h000441ED , 32'h00053AF3 , 32'h00012FF9 , 32'hFFFD757B , 32'h000359DB , 32'h0004601A , 32'hFFFB9269 , 32'hFFFCC12D , 32'hFFFB01F4 , 32'h000255C8 , 32'h0000E8B3 , 32'h0001CAD6 , 32'h00045CF7 , 32'h0001BD81 , 32'h00007AB7 , 32'h0002D12C , 32'hFFF80CE7} , 
{32'hFFF81C96 , 32'h0002C022 , 32'hFFFE6F64 , 32'hFFFB5467 , 32'h0002C8F9 , 32'h00012B8B , 32'hFFFF3CDC , 32'h0004B2C1 , 32'hFFFE1AE4 , 32'hFFFA01C8 , 32'h0005440C , 32'hFFFCFDBF , 32'hFFF806BE , 32'hFFFC63EF , 32'h0008A5AB , 32'h00013F19 , 32'h0005F7C5 , 32'h00008CA0 , 32'h0001413F , 32'hFFFB5F84 , 32'h0003F643 , 32'hFFFD0919 , 32'h0000A3BC , 32'h00004EBB , 32'hFFFF976C , 32'hFFF9BFC2 , 32'hFFFB9413 , 32'h000196F1 , 32'hFFFDAF47 , 32'h000192B3 , 32'hFFFFAA67 , 32'h0002FDE8 , 32'h00029C7B , 32'hFFFD718F , 32'hFFFE0E03 , 32'h00013E01 , 32'hFFFA6994} , 
{32'h0001FCF5 , 32'hFFF931E5 , 32'hFFFCA03C , 32'hFFFF8C93 , 32'hFFFE806C , 32'h00016101 , 32'hFFFDD59F , 32'hFFFF7F79 , 32'hFFFB417F , 32'h000460CA , 32'h0005FAE4 , 32'h0000D71C , 32'hFFFDCBB1 , 32'h0001A1D3 , 32'hFFF87CB2 , 32'hFFFEA3B4 , 32'h00017DA0 , 32'hFFFD4E6B , 32'h0001168A , 32'hFFF8D5F5 , 32'hFFF574CF , 32'h0002D8A3 , 32'hFFFF49EE , 32'hFFFD1B34 , 32'hFFFC5687 , 32'h00006889 , 32'hFFFC5517 , 32'h0003820D , 32'h00031A38 , 32'hFFFCC1FB , 32'hFFFCA0A4 , 32'hFFF74A53 , 32'h0002AD6A , 32'h0000AA45 , 32'hFFFEDFE8 , 32'h00014729 , 32'h000546ED} , 
{32'h00028496 , 32'hFFF78974 , 32'hFFFE7798 , 32'h00027172 , 32'h000376FD , 32'h0003B310 , 32'hFFFEDFDA , 32'hFFF98BE6 , 32'hFFFF6A13 , 32'h000267FD , 32'hFFFFFFBB , 32'h0004CFAF , 32'hFFFCA0D2 , 32'h00021D15 , 32'h00063D01 , 32'h00015F7F , 32'h0001FA16 , 32'h00004098 , 32'h000194C5 , 32'hFFFBEA7E , 32'h00049815 , 32'hFFFF0570 , 32'hFFFF06CC , 32'hFFFDFEF6 , 32'hFFFF97E8 , 32'hFFFDF6AD , 32'h0002ECD6 , 32'h0002F7ED , 32'h00057AC2 , 32'hFFFF3BE0 , 32'h00021D0D , 32'h0002BCBA , 32'hFFFE1077 , 32'hFFFC2FCF , 32'h0000C950 , 32'hFFFE5D50 , 32'hFFFEE92C} , 
{32'hFFFE84A7 , 32'h00009899 , 32'hFFFF7EF1 , 32'hFFFE5A12 , 32'hFFFC2A91 , 32'h000331CE , 32'h000317A4 , 32'hFFF96BE1 , 32'h0002ACFC , 32'h00024256 , 32'h00028D18 , 32'h00027F68 , 32'hFFFC9ACE , 32'hFFFF96FA , 32'hFFFE6805 , 32'h0004A7B4 , 32'hFFFE860B , 32'h0000DDBB , 32'hFFFFC65F , 32'h0001DF4E , 32'hFFFE07E5 , 32'hFFFFAA79 , 32'hFFF6466D , 32'h0001C483 , 32'hFFFF40F9 , 32'h0002106B , 32'hFFF8352A , 32'h0006D7DC , 32'hFFFDF14C , 32'h0002BD82 , 32'hFFFDF6F1 , 32'hFFFF5F73 , 32'h0000FB87 , 32'h00052877 , 32'hFFFFA9E9 , 32'h0001BB21 , 32'h0000155E} , 
{32'hFFFD514E , 32'hFFFD8FEF , 32'hFFFACFEB , 32'h000450F9 , 32'h0008F9B9 , 32'hFFF9D0E4 , 32'hFFFE2F33 , 32'h000158D3 , 32'h000652A6 , 32'h0002BB53 , 32'h00035DFB , 32'hFFFF09CC , 32'h00020B9C , 32'h000198A3 , 32'h00009FAA , 32'h00029C56 , 32'h0004A4F6 , 32'h00000018 , 32'hFFFD9E2F , 32'h0002889B , 32'hFFF9C2B3 , 32'h00003F83 , 32'h0001E511 , 32'h000250C2 , 32'hFFFEA396 , 32'hFFFA5EA7 , 32'hFFFC5C89 , 32'h0001BEDB , 32'hFFFADC54 , 32'h0005486A , 32'hFFFC8682 , 32'h00007EB0 , 32'h0007E07C , 32'h0004CA42 , 32'h000154A7 , 32'hFFFB3994 , 32'h00028E22} , 
{32'h00003038 , 32'hFFFFED0F , 32'hFFFF27DC , 32'hFFFE2EB1 , 32'hFFFF64B6 , 32'hFFFE0181 , 32'h000378C6 , 32'h00038BDF , 32'hFFFC5D99 , 32'h0001F962 , 32'h00004F89 , 32'hFFF6FAA9 , 32'hFFFFE659 , 32'hFFFE7A48 , 32'h00071342 , 32'hFFFEA1AF , 32'h00002F98 , 32'h00051980 , 32'hFFFDB0B2 , 32'h0005DFAE , 32'h00024E71 , 32'hFFFEE800 , 32'hFFFE8D88 , 32'h00009CC3 , 32'h00020D5A , 32'hFFFD8B2E , 32'h00012470 , 32'hFFFE5938 , 32'h0001265F , 32'h0001B682 , 32'h0004BCEB , 32'h00062F73 , 32'h00026D45 , 32'h0004CDE0 , 32'hFFFC5DFC , 32'h000297F3 , 32'hFFFF1DC2} , 
{32'h0000CAF9 , 32'h00006457 , 32'hFFFCA4EC , 32'h00022391 , 32'hFFF83EF6 , 32'hFFFABA78 , 32'hFFFF466B , 32'h0002815C , 32'hFFFF1CD7 , 32'hFFFD3B54 , 32'h000060D1 , 32'hFFFE81C3 , 32'h0002706A , 32'hFFFE43B9 , 32'hFFFFB578 , 32'h0002F185 , 32'hFFFE5F96 , 32'h000621A1 , 32'h0002841E , 32'h0001F58E , 32'hFFFFC372 , 32'hFFFD1F23 , 32'h0000BC12 , 32'h00041047 , 32'h000929C8 , 32'h00022C1A , 32'h0002F1ED , 32'h00007E7B , 32'h0001EB25 , 32'h00039CB8 , 32'h00010983 , 32'hFFFE5E70 , 32'h00007D9A , 32'h0000E1AB , 32'hFFFFE104 , 32'h00013243 , 32'hFFFF7543} , 
{32'h00061A0D , 32'h000170AC , 32'hFFFD7536 , 32'h00009139 , 32'hFFFB635E , 32'hFFFCEF6B , 32'hFFFC7A6A , 32'hFFFBD396 , 32'hFFFFC953 , 32'h000296E2 , 32'hFFFE6CFC , 32'h0002B220 , 32'hFFFA9500 , 32'hFFF8E1C9 , 32'h000A262B , 32'h0001760E , 32'h0004882A , 32'h0007C33C , 32'hFFFB3D41 , 32'h0002D822 , 32'h00010E98 , 32'hFFFF620C , 32'h0001B9AE , 32'hFFFAF58A , 32'h0009D757 , 32'hFFF7F0B3 , 32'hFFFD39C3 , 32'hFFFD513E , 32'hFFFFB8B2 , 32'hFFFD3185 , 32'hFFFE3510 , 32'h00044208 , 32'h0003216E , 32'hFFFD39E6 , 32'h0000C660 , 32'hFFFE6A02 , 32'hFFFBFC5B} , 
{32'hFFFC07F7 , 32'h0005035F , 32'h00022BD3 , 32'hFFFD1D6E , 32'h0001793F , 32'hFFF9A673 , 32'hFFFB6655 , 32'h00043745 , 32'hFFFEC94A , 32'h0004B11A , 32'hFFF95E58 , 32'hFFFE6B05 , 32'hFFFFA0EC , 32'hFFFC8592 , 32'h00005352 , 32'h0005EFC5 , 32'hFFFE95B2 , 32'hFFFDA21E , 32'h0002E5C3 , 32'hFFF71F2E , 32'hFFFEBF4E , 32'h00062F72 , 32'hFFF9E5BE , 32'hFFFEDCAA , 32'hFFFDECB3 , 32'h0004FD47 , 32'h00000AA7 , 32'h0004D3CF , 32'h00028B5A , 32'hFFFEDCD0 , 32'h0000C21D , 32'hFFFED6AD , 32'hFFFFFE70 , 32'hFFFCE21B , 32'h000148C9 , 32'hFFF926D0 , 32'h00018A12} , 
{32'h00012025 , 32'h00002D8C , 32'hFFFEA44A , 32'h0000D790 , 32'h0001A9D3 , 32'h0000A533 , 32'hFFFFB328 , 32'hFFFD2AFE , 32'h0000DABD , 32'h0001950F , 32'hFFFCFD70 , 32'h00035460 , 32'hFFFC6961 , 32'h0001FF6D , 32'hFFFFE85E , 32'hFFFC2FE1 , 32'hFFFECDA3 , 32'h000456B3 , 32'hFFFEE10D , 32'h0004CDCB , 32'h00034628 , 32'hFFFFF3D2 , 32'hFFF73CEB , 32'hFFFEE7D8 , 32'hFFFD6DDA , 32'h00062E1F , 32'hFFFC1A3A , 32'h0000FD4E , 32'hFFFA3C8A , 32'hFFFB81B6 , 32'h000259AD , 32'h0002233C , 32'hFFFF4AA8 , 32'hFFFD01D4 , 32'h0001D7CE , 32'h00009C03 , 32'h000137C6} , 
{32'h00011BA7 , 32'hFFFF7333 , 32'h0000618F , 32'h00062148 , 32'h00031BFF , 32'hFFFE3057 , 32'h000055CD , 32'h00046196 , 32'hFFFD2C53 , 32'h0002A858 , 32'hFFFF77F3 , 32'h0002FF92 , 32'hFFFC560C , 32'h000019C7 , 32'h0005E8E5 , 32'h00063832 , 32'hFFFD755F , 32'hFFFF49EB , 32'h00037475 , 32'hFFFCE654 , 32'h0002414A , 32'hFFFEAF03 , 32'h0001F134 , 32'h00030B1A , 32'h00022CD2 , 32'h0001C6DD , 32'h00007FA5 , 32'h0000472B , 32'hFFFB9CB5 , 32'h000677C8 , 32'h0003025B , 32'h00015AE0 , 32'hFFFCF329 , 32'hFFFF910E , 32'h000097A1 , 32'h000497CB , 32'h0007EBA5} , 
{32'hFFFF6459 , 32'h0006E71E , 32'h0001A441 , 32'h0001A09B , 32'h000073D2 , 32'h0004792E , 32'h0000F15D , 32'hFFFADCB2 , 32'h000220D4 , 32'h0001EA98 , 32'hFFF940D3 , 32'h0001CED0 , 32'hFFFF7DC3 , 32'h000456D9 , 32'h000396DC , 32'hFFF87D47 , 32'hFFFBE2FA , 32'h00000271 , 32'h0003A70E , 32'h00050BAB , 32'h0002B0F6 , 32'hFFFBD77B , 32'h000332D6 , 32'hFFFDE5E2 , 32'h00066BDC , 32'h00002F38 , 32'hFFFD5F90 , 32'h00025415 , 32'hFFFF53E5 , 32'h00004005 , 32'h000028B6 , 32'h00042799 , 32'hFFFFABE3 , 32'hFFFC8389 , 32'hFFFEF4F3 , 32'h00014CC1 , 32'h0001E656} , 
{32'hFFFD49E2 , 32'h00013013 , 32'hFFFF8D13 , 32'h0004B0D8 , 32'hFFFFB13D , 32'hFFF850C1 , 32'h00015808 , 32'h0004C596 , 32'hFFFF022C , 32'hFFFFDE15 , 32'hFFFB51C0 , 32'hFFFAE68B , 32'h0002E98C , 32'h000397E9 , 32'hFFFE6761 , 32'hFFFEB4CF , 32'h0002B437 , 32'h0000F333 , 32'h000002AF , 32'hFFFF49CA , 32'h0002C867 , 32'hFFFE42AB , 32'hFFFE4B98 , 32'h00008DC6 , 32'hFFFCD6A4 , 32'hFFFD9066 , 32'h0000BA0D , 32'h00018246 , 32'hFFFCCCCC , 32'h0000CF03 , 32'h0006CC26 , 32'hFFFF7CB0 , 32'h0004243F , 32'h00049B3B , 32'h0004E1C7 , 32'hFFFDA1E5 , 32'hFFFF63D2} , 
{32'hFFFB6E1C , 32'h0003F58B , 32'hFFFD3E08 , 32'h0004BAAA , 32'h0002BEFE , 32'h00044EE7 , 32'hFFFDAC8C , 32'h0001BE10 , 32'h00021D6F , 32'h0000FDC6 , 32'h00047ADF , 32'hFFFDC1BD , 32'hFFFCE5BB , 32'h0001F014 , 32'h00000003 , 32'h0002EA0E , 32'hFFFF8E9E , 32'hFFFF3592 , 32'hFFFFA890 , 32'hFFFFD5E3 , 32'hFFFCEC6E , 32'hFFFD3B6B , 32'hFFFC89E8 , 32'hFFFEC057 , 32'h0001F0C9 , 32'h000226AF , 32'hFFFED734 , 32'hFFFF0DA3 , 32'h00020424 , 32'hFFFE0CDF , 32'h0004AC66 , 32'hFFFA0E3C , 32'h0000D92F , 32'h0009EE1C , 32'hFFFEB6EC , 32'h00004353 , 32'hFFFEE74A} , 
{32'hFFFE62B1 , 32'h00020655 , 32'h0004F1E4 , 32'h0004AB37 , 32'h00018C96 , 32'h000044B1 , 32'hFFF85D51 , 32'h00027389 , 32'hFFFF786C , 32'h00036B4B , 32'hFFFA4ECE , 32'hFFFF79BE , 32'hFFFF2B3F , 32'h0001AE68 , 32'hFFFE1B61 , 32'h00040E95 , 32'h0002D2A4 , 32'hFFFE3A6D , 32'hFFFC7135 , 32'h000064F5 , 32'hFFFC3231 , 32'hFFFD0BBC , 32'hFFFD63B2 , 32'h0002D608 , 32'hFFFB68E9 , 32'h00021298 , 32'hFFFBB05F , 32'hFFFFC937 , 32'hFFFBCFFF , 32'h000528ED , 32'h00054A05 , 32'h0004273C , 32'hFFFF4098 , 32'hFFFE3381 , 32'hFFF9E49C , 32'h0000BDA2 , 32'h0002A088} , 
{32'h0001CA7D , 32'hFFFEC84A , 32'h0005A266 , 32'h0003F3B8 , 32'h000129C8 , 32'hFFFD24B1 , 32'h00028A69 , 32'h00011DC3 , 32'hFFFDAAEC , 32'h0006AA18 , 32'hFFFF4660 , 32'hFFFE4082 , 32'h00013917 , 32'h0003368A , 32'hFFFD58FD , 32'h00003EBB , 32'h00009D2D , 32'h0000F2AA , 32'hFFF9E8FC , 32'hFFFD1919 , 32'hFFFEB5D9 , 32'hFFFD06F7 , 32'h0004F93F , 32'h00029608 , 32'hFFFEE2DE , 32'hFFFD3C53 , 32'hFFFD0B77 , 32'h000088FE , 32'hFFFB509C , 32'hFFFD38BB , 32'h000511D8 , 32'h00045BB1 , 32'hFFFFD7D8 , 32'hFFFC9D4D , 32'h00046522 , 32'hFFF9247D , 32'h00021135} , 
{32'hFFFC3E49 , 32'hFFFEA30B , 32'h0004C010 , 32'h00028D94 , 32'hFFFDD75B , 32'hFFFB4C69 , 32'hFFFD80CA , 32'hFFFFF70F , 32'h0003A2AF , 32'hFFFE6850 , 32'hFFFF1909 , 32'hFFFE216F , 32'h00041C70 , 32'h000141AF , 32'hFFFC0AB5 , 32'hFFFD7A82 , 32'h00057A37 , 32'hFFFE8595 , 32'hFFFE05C9 , 32'hFFFC84A0 , 32'hFFFC6042 , 32'h000340FD , 32'h0001F58E , 32'hFFFD2FDA , 32'h0003C4A9 , 32'hFFFF06EC , 32'h00017DD8 , 32'h00064232 , 32'hFFF965CB , 32'h00014488 , 32'hFFFF5262 , 32'hFFFA6F10 , 32'hFFFDA2D5 , 32'hFFFA08A3 , 32'hFFFD1A0B , 32'hFFFD0F1D , 32'hFFF80164} , 
{32'hFFF6FCBC , 32'hFFFE92AE , 32'hFFFF4047 , 32'h000311DF , 32'hFFFC68BC , 32'hFFF755AD , 32'h00005314 , 32'h000008A6 , 32'h000498FA , 32'h00057A39 , 32'hFFFC9249 , 32'h0000C9A3 , 32'hFFFF6139 , 32'h0005A4DF , 32'h00093590 , 32'h00051ACD , 32'hFFFE9B64 , 32'hFFFD60FB , 32'hFFFE5744 , 32'hFFFD525B , 32'h00042434 , 32'h00025A07 , 32'hFFFEDA37 , 32'hFFFDCF3C , 32'hFFFDE5F4 , 32'hFFFE2FC9 , 32'h000422E9 , 32'hFFF8787D , 32'h00050257 , 32'hFFFF42B4 , 32'hFFFC09A0 , 32'h0007D551 , 32'h000052FD , 32'h0001D718 , 32'hFFFE73D2 , 32'hFFFFD5FD , 32'hFFFCB7D3} , 
{32'h0003FC16 , 32'h0001AB2E , 32'h0000BD3F , 32'hFFFDB09A , 32'h0004A3A2 , 32'hFFFF9E1C , 32'hFFF9C8AD , 32'h00063A14 , 32'h00016B7E , 32'h00013885 , 32'hFFFFFBE5 , 32'hFFFFEC40 , 32'h00028182 , 32'hFFFFA9ED , 32'hFFFFC493 , 32'h00030360 , 32'h00016925 , 32'hFFFE6359 , 32'hFFFEF5D1 , 32'h0001C595 , 32'h0000A23F , 32'hFFFEFFE4 , 32'hFFF77DA1 , 32'h0000D8FE , 32'hFFFBC779 , 32'h00004F14 , 32'h0001527F , 32'h000373F9 , 32'h0001BED4 , 32'h00020638 , 32'h00004283 , 32'h00042266 , 32'hFFF7723B , 32'h0003347F , 32'hFFFEBDF2 , 32'h0000CE32 , 32'h00028E8D} , 
{32'hFFFB0185 , 32'h000266BB , 32'hFFFEC8AB , 32'h00001BCB , 32'h0001AAD3 , 32'hFFFA0842 , 32'h00082F87 , 32'h0001BC86 , 32'h00084B68 , 32'hFFFFCAA0 , 32'h00042567 , 32'h0000BD17 , 32'hFFFC5AC6 , 32'h00004A57 , 32'hFFFC552B , 32'hFFFC0ABB , 32'h00025C5E , 32'h000148DA , 32'hFFFDE442 , 32'hFFFE7F65 , 32'h000341FB , 32'h0003D73F , 32'h0000252B , 32'h0001E753 , 32'hFFFBB820 , 32'hFFFCD962 , 32'h0000C019 , 32'hFFFE276F , 32'h0000F135 , 32'h0000F409 , 32'hFFFEE45F , 32'h0001F7F0 , 32'h0003424F , 32'h000183B6 , 32'hFFFC00B4 , 32'h00016F62 , 32'hFFFC6D60} , 
{32'h00024EF6 , 32'h000129B6 , 32'hFFFF68A5 , 32'hFFF7B73E , 32'hFFFEF0FF , 32'h0001169D , 32'hFFFDC9A9 , 32'hFFFCE255 , 32'hFFFD18D9 , 32'h00007DEE , 32'h00052FE3 , 32'hFFFE7E22 , 32'h0008EF28 , 32'hFFFF0612 , 32'h0003ACFC , 32'hFFFFEEB5 , 32'hFFF9A18A , 32'h00032BC9 , 32'h0001B40D , 32'h000103DD , 32'hFFFC4612 , 32'h0003DC8B , 32'h0000AA6E , 32'hFFFE9017 , 32'h0005AD80 , 32'h00057F07 , 32'hFFFB8C20 , 32'hFFFD88D6 , 32'hFFFFF430 , 32'hFFFF4213 , 32'h0000DDBE , 32'h000279EA , 32'hFFFC23F6 , 32'h00043F0E , 32'h00047DCA , 32'hFFFD1985 , 32'hFFF85C4F} , 
{32'h0006D128 , 32'h000363A8 , 32'h0001B6C8 , 32'h000C0666 , 32'hFFFA9D83 , 32'h0003AE10 , 32'hFFFFC0E8 , 32'h0002288D , 32'h0003123F , 32'hFFFE71D9 , 32'h00096BF1 , 32'h00081A7A , 32'h00023BDC , 32'h000783A1 , 32'hFFFF214C , 32'hFFF9964C , 32'hFFFD38DE , 32'h000398F3 , 32'hFFFB7173 , 32'h000442DB , 32'hFFFB3417 , 32'hFFFEB63D , 32'hFFFD9767 , 32'hFFFF2AF8 , 32'hFFF8AA2B , 32'h0000C29F , 32'h0004B649 , 32'h0000DBE6 , 32'hFFFBBEDF , 32'hFFFDB396 , 32'hFFFD6F39 , 32'hFFFC4066 , 32'h0000E4C9 , 32'h00050E6A , 32'h0000C9BE , 32'hFFFCC9D1 , 32'h0002F1B1} , 
{32'hFFFC7C03 , 32'h00005567 , 32'h0001792B , 32'h00050ED3 , 32'hFFFE3F8F , 32'h000567B9 , 32'hFFFFE632 , 32'h0001D445 , 32'h000325C4 , 32'h00010177 , 32'h00075B8B , 32'h0000E942 , 32'h00007088 , 32'hFFFF5DF8 , 32'hFFFE0318 , 32'hFFFBCF44 , 32'h00032F6B , 32'hFFFF1E84 , 32'hFFFCBE13 , 32'hFFFA8648 , 32'hFFFDE9B5 , 32'hFFFDC2C9 , 32'hFFFE7E97 , 32'hFFFC3C04 , 32'h0001B530 , 32'h000019D9 , 32'h0001540A , 32'hFFFF6CB4 , 32'h0000815F , 32'hFFFCAF62 , 32'h0007BB00 , 32'hFFFB3379 , 32'hFFF7F0A9 , 32'h000036C1 , 32'hFFFDD457 , 32'h0000F388 , 32'h000188BD} , 
{32'hFFFFD82F , 32'h0001F6C2 , 32'h000069E3 , 32'hFFFF4F14 , 32'hFFFE2A88 , 32'hFFFEC049 , 32'hFFFFBBDB , 32'hFFFC29E8 , 32'hFFF9E3E5 , 32'hFFFFBEC4 , 32'h0000A9EA , 32'hFFFEB409 , 32'hFFFAE562 , 32'hFFFD355E , 32'h0003BEFA , 32'hFFF89917 , 32'hFFFE0E94 , 32'hFFFF13E3 , 32'h00015C1E , 32'hFFFC0F99 , 32'hFFF9254E , 32'hFFFAF652 , 32'h0002EEA6 , 32'hFFF8C40C , 32'hFFFD9FF6 , 32'h0007434F , 32'h000467AC , 32'hFFFD99C0 , 32'hFFFF232A , 32'hFFFBE0EE , 32'hFFFCFCAA , 32'hFFFECFD3 , 32'h000237A0 , 32'h0004E27F , 32'hFFFF30BA , 32'h0001950B , 32'hFFFE3CCE} , 
{32'h00067C08 , 32'hFFF99D18 , 32'hFFFC61E1 , 32'hFFFB4A07 , 32'h00043FBA , 32'h0001069A , 32'hFFFE5D6C , 32'hFFFBFBAA , 32'hFFFEE3C8 , 32'h0002AACF , 32'h000006AA , 32'hFFFFF622 , 32'hFFFE85F5 , 32'h0001A28B , 32'h0000F527 , 32'hFFFBEBDF , 32'h0001A1C3 , 32'hFFFE81EF , 32'h000423D5 , 32'h0003920F , 32'hFFFCAA7D , 32'hFFF92D70 , 32'hFFFF780A , 32'hFFFC8374 , 32'h000027F5 , 32'h00000A7C , 32'hFFFFE7FB , 32'h0000DC49 , 32'hFFF842D2 , 32'h000292E3 , 32'h00071FCF , 32'h000243EE , 32'hFFFF9B7F , 32'hFFFFDEFE , 32'hFFFFE7FC , 32'h00030C6A , 32'hFFFBFCA4} , 
{32'hFFFC7535 , 32'hFFFFD6AF , 32'hFFFC7F78 , 32'h00043BEC , 32'hFFFA9F3A , 32'hFFFDDC14 , 32'hFFFB179E , 32'hFFFD5D7E , 32'hFFF8147C , 32'h000078F0 , 32'h000272A5 , 32'hFFFDE9CF , 32'h000BCD57 , 32'hFFF9DED8 , 32'hFFFCCA57 , 32'hFFFDDF8E , 32'hFFFDBB62 , 32'hFFFE2111 , 32'h00009ECF , 32'h0004DFF6 , 32'hFFFE9ED6 , 32'h000628DC , 32'h0001C346 , 32'hFFFDE6A5 , 32'h00078BD5 , 32'hFFFEA563 , 32'hFFFF1951 , 32'hFFFCBBC6 , 32'h0002A84E , 32'h00040678 , 32'hFFFE31DB , 32'hFFFB9ECF , 32'hFFFF57FB , 32'h000B3A9F , 32'hFFFC13EA , 32'h00006A53 , 32'h00002D1C} , 
{32'h0003BA3F , 32'hFFFCE342 , 32'hFFFA2535 , 32'hFFFF819A , 32'h000441B1 , 32'hFFFEBA93 , 32'hFFF8AB87 , 32'h00005DCF , 32'hFFFC9234 , 32'h0002252A , 32'hFFFDDF8C , 32'hFFFDA000 , 32'h0003706F , 32'h000059C1 , 32'hFFFF06D7 , 32'h000532A9 , 32'hFFFC9A4C , 32'hFFFD3F32 , 32'h000072A7 , 32'hFFFF23BB , 32'h0006D262 , 32'hFFFC80F0 , 32'hFFFF51A0 , 32'hFFFD37D9 , 32'hFFFE30EA , 32'h00001F44 , 32'h00070698 , 32'h0001C1B0 , 32'h000098B1 , 32'hFFFAEB9E , 32'h0002D4DB , 32'h0001D752 , 32'hFFFF60F8 , 32'hFFFA6A88 , 32'h0001D68A , 32'h0004779C , 32'h0000EFFF} , 
{32'h0000E786 , 32'h0002568C , 32'h00017C94 , 32'hFFFF8CEF , 32'h00014A4A , 32'h00037535 , 32'h0002E3C1 , 32'hFFFEB9A5 , 32'hFFFD9A6A , 32'hFFFD236E , 32'h0000B300 , 32'h00021054 , 32'h000240E0 , 32'hFFFDEF66 , 32'h0002E483 , 32'h0000F916 , 32'hFFFE107F , 32'hFFFBC053 , 32'hFFF91F56 , 32'h00012D5B , 32'hFFFFBECD , 32'hFFFE7AEB , 32'hFFFE4670 , 32'hFFFECD66 , 32'h0001DF51 , 32'h0000F217 , 32'hFFFF3119 , 32'hFFFCBB92 , 32'hFFFE7265 , 32'hFFFF9F61 , 32'hFFFC2BE8 , 32'h000397FC , 32'h0003863C , 32'hFFFEBE72 , 32'hFFFD1C95 , 32'h00031C7E , 32'hFFFDBAFC} , 
{32'h0004B9EA , 32'hFFFD455E , 32'h0000C85E , 32'hFFF97528 , 32'hFFFE74BB , 32'h0006FF17 , 32'h000692DF , 32'h000326D3 , 32'h00013212 , 32'hFFFD380C , 32'h000408B5 , 32'hFFFD6EB7 , 32'hFFF7B934 , 32'h0001010C , 32'hFFFAA5E1 , 32'hFFFAC7D8 , 32'h0004B718 , 32'h0000E914 , 32'h00018538 , 32'hFFFE7EB3 , 32'h00015CD2 , 32'h000193AF , 32'hFFFBF80A , 32'h0001C3CE , 32'hFFFC33B3 , 32'hFFFD6FF3 , 32'h00067009 , 32'hFFFECCAC , 32'h0000A64E , 32'h0003DF7C , 32'h000092E3 , 32'h0001361D , 32'h00002F8F , 32'h00045CB8 , 32'hFFFF4CB2 , 32'hFFFE83B7 , 32'hFFFE3B1E} , 
{32'hFFFB4573 , 32'h0003D24A , 32'h00048C6D , 32'hFFF82911 , 32'hFFFDF27A , 32'h0004B4FE , 32'hFFFC5A3D , 32'hFFFC92AD , 32'hFFFE50B5 , 32'hFFF8E72D , 32'hFFFD5BB1 , 32'hFFFC9FDA , 32'h00010C65 , 32'hFFFEC8E2 , 32'h00004EDF , 32'h0001BD47 , 32'h0000C83E , 32'hFFFC6A9C , 32'hFFFF75D3 , 32'h0001BA1D , 32'h000487F7 , 32'hFFFAFD77 , 32'hFFFD3B03 , 32'hFFFFBAC3 , 32'h0001503F , 32'hFFFFB69C , 32'h00023FFE , 32'hFFF8D7B7 , 32'hFFFFA8E4 , 32'h00053F6E , 32'hFFFB6A1A , 32'h0002B279 , 32'h00023DC0 , 32'h0000005B , 32'hFFFD287F , 32'h00016478 , 32'h00023945} , 
{32'hFFFF44AB , 32'hFFFD9A42 , 32'h00013665 , 32'h00028F3E , 32'hFFFEDF3D , 32'hFFFFC34B , 32'hFFFC9E45 , 32'h000142C8 , 32'h00010248 , 32'h00030054 , 32'h00031082 , 32'hFFFF2999 , 32'h0001195F , 32'h0000F57E , 32'hFFFAA662 , 32'hFFFF760C , 32'h00001356 , 32'h00098098 , 32'h0001B452 , 32'h0008A117 , 32'hFFFB3F26 , 32'h0001B16B , 32'hFFFF2E6B , 32'h0003E0B3 , 32'h00020244 , 32'h00007B7C , 32'h00000FCF , 32'hFFFFB90B , 32'hFFFC3D4B , 32'h000062D4 , 32'hFFFB8529 , 32'hFFFEB78B , 32'h00076644 , 32'hFFFDC143 , 32'hFFFEB4F5 , 32'hFFF58E9A , 32'hFFF899EE} , 
{32'h000168E5 , 32'h000891F8 , 32'hFFFF1013 , 32'hFFFD6CAE , 32'hFFFE40C2 , 32'hFFFD6BE0 , 32'hFFFE9E4F , 32'hFFFEB2D1 , 32'h0001C748 , 32'hFFFC41B9 , 32'hFFFBA4EE , 32'h0004D879 , 32'hFFFE842E , 32'hFFFB40ED , 32'h0000CEBB , 32'h0001B8C3 , 32'h00003944 , 32'hFFFE3053 , 32'hFFFF3222 , 32'h0003146C , 32'h000306A8 , 32'h0000300B , 32'h0003A913 , 32'hFFFD1F4C , 32'hFFFD140F , 32'h000233B0 , 32'hFFFEAE62 , 32'h00000C4F , 32'hFFFF6563 , 32'hFFFD221D , 32'hFFFF130C , 32'h0003650D , 32'hFFFE53E7 , 32'h00044ED6 , 32'hFFFBEDCA , 32'hFFFD6289 , 32'h000182F2} , 
{32'h0001C2CB , 32'h000010AE , 32'h0001140F , 32'h0000B19F , 32'h00040157 , 32'h00004000 , 32'hFFFBD58F , 32'h0001B119 , 32'h0002432D , 32'hFFFF8FF1 , 32'hFFFC38B1 , 32'h00049CDF , 32'h00021245 , 32'h000414D8 , 32'hFFFEB415 , 32'h00004223 , 32'hFFFEB7F5 , 32'h00028A19 , 32'hFFFAD9CC , 32'hFFFEB2F1 , 32'h0000A8D6 , 32'hFFFEE5D0 , 32'h00009346 , 32'h00039890 , 32'h000151E1 , 32'hFFFE0137 , 32'h0000516A , 32'h0006637E , 32'hFFFF8B03 , 32'h000252C8 , 32'h000202A7 , 32'h00040C41 , 32'hFFFDB196 , 32'h0002214C , 32'hFFFB5C98 , 32'h000066B5 , 32'hFFFBA1E3} , 
{32'hFFFC4A88 , 32'hFFFCD2CF , 32'hFFFE18FA , 32'hFFFF325A , 32'hFFFFB6DA , 32'h000103A7 , 32'h00039C05 , 32'h000057D1 , 32'hFFFD1C4D , 32'h0001B79B , 32'h0001391F , 32'hFFFBFC9A , 32'hFFFD6E29 , 32'hFFFE2774 , 32'hFFFE5D75 , 32'h000784D4 , 32'h00002060 , 32'hFFFEDA5B , 32'h00082464 , 32'h000047CE , 32'hFFF71CF4 , 32'h0008BF7D , 32'h00076065 , 32'hFFF986EA , 32'hFFFCB09A , 32'hFFFF0CF6 , 32'h00013DA3 , 32'hFFFFCAA6 , 32'hFFFB3EFA , 32'h0001EA04 , 32'hFFFC8046 , 32'hFFFF5160 , 32'h000792AF , 32'h0001544D , 32'hFFFEC85E , 32'h000105B2 , 32'hFFFD5C53} , 
{32'hFFF9F66B , 32'h0005DF02 , 32'hFFFC06DB , 32'h0000FF44 , 32'h0000F570 , 32'hFFFDC01E , 32'h0000C526 , 32'h00057721 , 32'hFFFC7A36 , 32'h00033F44 , 32'hFFFF8BA7 , 32'h0000A778 , 32'h00033C09 , 32'h00073C5B , 32'h00021244 , 32'h00004224 , 32'h00021F8D , 32'hFFFA9696 , 32'h0005443C , 32'h0000FB4A , 32'hFFFDCB99 , 32'h0002F819 , 32'h000485C4 , 32'hFFFF8442 , 32'hFFFB972E , 32'hFFF9799D , 32'h00035B5D , 32'h0005D2C3 , 32'hFFFF75DB , 32'h0002C82C , 32'h00045F97 , 32'h00031059 , 32'hFFFED2B7 , 32'h000579C3 , 32'h0000C354 , 32'hFFFFEA57 , 32'h000120AC} , 
{32'h00021628 , 32'h0001B556 , 32'hFFFF3659 , 32'hFFFC47BC , 32'h0003F01A , 32'hFFFDAC1E , 32'h00003342 , 32'hFFFEDCB5 , 32'hFFFF2D22 , 32'hFFFA2002 , 32'hFFFFFA34 , 32'h0000DC8D , 32'hFFFF53FF , 32'hFFFE401D , 32'h000089EA , 32'h000357A9 , 32'hFFFE7662 , 32'hFFFAD5E3 , 32'h00056317 , 32'h0002388F , 32'h00047D49 , 32'h00013920 , 32'h0003D2F9 , 32'hFFFF4220 , 32'hFFFBB80E , 32'h00026364 , 32'hFFFEC87F , 32'h0004DBD4 , 32'hFFFEAF3C , 32'hFFFEF474 , 32'hFFFC9CD6 , 32'hFFF8776D , 32'h00001EB3 , 32'h0002D4CC , 32'hFFFC6830 , 32'h0004D428 , 32'hFFFDAB41} , 
{32'hFFFE886F , 32'hFFFE91BB , 32'h0003A34C , 32'h0005DC9A , 32'h00078D5A , 32'h0002A079 , 32'h000473E1 , 32'h00046BED , 32'h00001B8A , 32'h0001599B , 32'h0005E43B , 32'hFFFD6A9E , 32'h00022FA6 , 32'hFFF8627F , 32'hFFFE8651 , 32'h0000B1F8 , 32'h00000E6A , 32'h00038DE1 , 32'h00014C1E , 32'hFFFA8822 , 32'h0000E865 , 32'hFFFFDD79 , 32'h0006697A , 32'h000091F1 , 32'h0000F98E , 32'h00007BF7 , 32'h0001C9A1 , 32'hFFFF3185 , 32'h00019D15 , 32'h0002BA76 , 32'hFFFA2AF6 , 32'h0002F787 , 32'h000296FA , 32'h0001C086 , 32'h0000AC6D , 32'h0002F249 , 32'hFFFC64FB} , 
{32'h00001743 , 32'hFFFD6814 , 32'hFFFECA24 , 32'hFFFEECE3 , 32'hFFFC9181 , 32'h000293EF , 32'h00036B4E , 32'hFFFDF3E0 , 32'hFFFD935D , 32'hFFFFD544 , 32'hFFFD4446 , 32'h00000CF9 , 32'hFFF95724 , 32'hFFFC6624 , 32'h00019994 , 32'hFFF60190 , 32'h000462EA , 32'h0001004F , 32'hFFFA66FF , 32'hFFFA3231 , 32'h000141F9 , 32'h00019DDA , 32'hFFFCAE78 , 32'hFFFF7689 , 32'hFFFFA5A5 , 32'hFFFF48AC , 32'h00036CE7 , 32'h00014D96 , 32'h0004E9EF , 32'h0004684A , 32'hFFFC7B5B , 32'h00005336 , 32'hFFFFBC81 , 32'hFFFCDDE8 , 32'hFFFF166C , 32'hFFFC04EB , 32'h0000EEF4} , 
{32'hFFFF5C08 , 32'hFFFCBF37 , 32'hFFFEA259 , 32'hFFFFBA7D , 32'hFFFEAFD4 , 32'h0001FB09 , 32'h0000B3E4 , 32'h0000F5B5 , 32'h00077DC8 , 32'hFFFDDDE5 , 32'h00061E0E , 32'hFFFC44BD , 32'h00039BF6 , 32'hFFF7C9BD , 32'hFFF9D7D9 , 32'h000550BA , 32'hFFFC3A41 , 32'hFFFE6D23 , 32'hFFFEDD65 , 32'hFFFFEF71 , 32'hFFFCB38E , 32'h0004BACD , 32'hFFFD721F , 32'hFFFE45B6 , 32'h00013F2A , 32'h00018535 , 32'h000173FB , 32'h00040E60 , 32'h000167F9 , 32'h00007BDE , 32'hFFFD4E30 , 32'hFFFB0333 , 32'h000190C5 , 32'h0007BB0C , 32'h00009FCE , 32'hFFFEA9FE , 32'h0004180C} , 
{32'hFFFFFE65 , 32'h0002CC36 , 32'h0002D6FD , 32'hFFFE91E4 , 32'h00024061 , 32'hFFFE55C9 , 32'hFFFF0F67 , 32'h00045C67 , 32'h0002B033 , 32'h00014EE7 , 32'hFFFECE99 , 32'h0001C472 , 32'h00005809 , 32'h0001B0B5 , 32'hFFFF6217 , 32'h0003CF29 , 32'h000183C0 , 32'hFFFFCE03 , 32'h0001B870 , 32'h000121BD , 32'h0004DFE1 , 32'hFFFDF1AA , 32'h0001EDF7 , 32'hFFFFDFAD , 32'h0003793E , 32'h00029381 , 32'hFFFCAB30 , 32'h0000241A , 32'h00018DEE , 32'hFFFE85CD , 32'h00000BE2 , 32'hFFFFBDEB , 32'hFFFCC3DA , 32'h0003276A , 32'hFFFA93B9 , 32'h00005499 , 32'hFFFBF792} , 
{32'h0003A98B , 32'h0000DCAE , 32'h00008C36 , 32'hFFFF9594 , 32'hFFF882AD , 32'hFFFE5E22 , 32'hFFFEA3EE , 32'h00000FF5 , 32'h00046969 , 32'h0004AE43 , 32'hFFFFD1F0 , 32'h000160FA , 32'hFFFC7CF6 , 32'h0000D30A , 32'hFFFF7991 , 32'h00039A92 , 32'h0000FDEA , 32'hFFFC0741 , 32'h0004ED4E , 32'h0000F97D , 32'hFFFD15DF , 32'hFFFDB1F3 , 32'h00015C18 , 32'h0006586D , 32'h0002CD9D , 32'h0003D51B , 32'h00026DA1 , 32'hFFFF3860 , 32'h0000CF15 , 32'hFFFF0EA9 , 32'h000179E4 , 32'h000072F0 , 32'hFFFD96D1 , 32'h000350F6 , 32'h0002EDCE , 32'h0000011A , 32'h000349FF} , 
{32'hFFFD6EBE , 32'h0001E835 , 32'hFFFCF058 , 32'hFFFDF8BC , 32'h0001F700 , 32'hFFFE0D28 , 32'h000167AD , 32'h0000D317 , 32'hFFFF0530 , 32'h000040C0 , 32'h00016492 , 32'h0001AAA9 , 32'h00046A7E , 32'h00033DD8 , 32'h00001E38 , 32'h0004F596 , 32'hFFFFD2BC , 32'h0001D402 , 32'hFFFB680A , 32'h0001C56C , 32'h0001B277 , 32'hFFFF5BB1 , 32'hFFFCBFCA , 32'h000092CD , 32'h000034C8 , 32'h00006FFE , 32'h00042543 , 32'h0000AF2C , 32'hFFFECFEF , 32'hFFFEF193 , 32'h00052691 , 32'h00045F69 , 32'h00003541 , 32'hFFFCE0BA , 32'hFFFDE882 , 32'h0002A55D , 32'hFFFD0626} , 
{32'hFE2DD0F4 , 32'hFFEF4A4A , 32'hFEC76540 , 32'h03EE4F70 , 32'h0044B795 , 32'h0046A147 , 32'hFF6D4159 , 32'h042329B0 , 32'hFF082E29 , 32'h001D4DA8 , 32'h006620A7 , 32'h01C8A06C , 32'h0120343C , 32'hFFF94F93 , 32'hFF09D0A8 , 32'hFF9C5DF8 , 32'h0090AA49 , 32'h00FD3AE9 , 32'hFD34A244 , 32'h00C0943F , 32'hFF647F19 , 32'h016D9B84 , 32'hFDD5C350 , 32'h00347E1B , 32'h00783056 , 32'hFEF71828 , 32'hFEB28D70 , 32'h0074E00E , 32'h0005C5BD , 32'hFF8095B7 , 32'hFF2E9B79 , 32'h00C6E35E , 32'hFEA4CAE0 , 32'hFDAC8370 , 32'h028619F0 , 32'hFCDF1D74 , 32'hFE9BAACC} , 
{32'hFFFD0FC5 , 32'h00040A35 , 32'hFFFF0C77 , 32'hFFFF1A79 , 32'h0000FC18 , 32'h0003E02C , 32'h00012895 , 32'hFFFEEF53 , 32'hFFFF4EDF , 32'hFFFD0A6F , 32'hFFFA5D05 , 32'hFFFF440B , 32'h000046A1 , 32'hFFFF6D38 , 32'hFFFE7438 , 32'hFFFFCB81 , 32'hFFFF513F , 32'hFFFD7C1A , 32'h0002BF27 , 32'hFFFCB580 , 32'h00024573 , 32'h00015D6B , 32'h000014B6 , 32'h00015221 , 32'h000068CC , 32'h00025BB2 , 32'hFFFFD65C , 32'hFFFB901A , 32'h0002C8E5 , 32'hFFFD338E , 32'h00011B8B , 32'h0004AEF7 , 32'hFFFD7DC3 , 32'hFFFC93E8 , 32'hFFFE9EBD , 32'h0003180F , 32'hFFFF9468} , 
{32'hFFFFE4B5 , 32'hFFF9EBF8 , 32'h000182BD , 32'h000039DC , 32'h000537B7 , 32'h00029FA0 , 32'h000512E8 , 32'hFFFF0764 , 32'hFFFC57AE , 32'hFFFFAB86 , 32'hFFFF1E47 , 32'h0002FB3B , 32'h000432F0 , 32'h0000BFEB , 32'h0001D33D , 32'h00011192 , 32'hFFFEDE6E , 32'hFFFF5276 , 32'hFFFEF9EE , 32'hFFFF5FC6 , 32'h0002585C , 32'hFFFEDAF8 , 32'hFFFCDCD9 , 32'hFFFC9F86 , 32'h000258A4 , 32'h000236E0 , 32'h00036671 , 32'h0005193B , 32'hFFFF3B5C , 32'hFFFF8AB2 , 32'hFFFB582A , 32'h0001ECE2 , 32'hFFFD1485 , 32'hFFFB2675 , 32'hFFFD548B , 32'h0007CCC7 , 32'hFFFE4491} , 
{32'hFFFFECDA , 32'h000169EB , 32'h00009D52 , 32'h0000DF75 , 32'h0001AA0F , 32'hFFFF0978 , 32'h000051F9 , 32'h00007003 , 32'hFFFECBB0 , 32'hFFFE749F , 32'hFFFF08B0 , 32'hFFFE5BB2 , 32'hFFFF2F8B , 32'hFFFD7ED1 , 32'h00022A00 , 32'h0004D234 , 32'hFFFD6893 , 32'h0002C8F7 , 32'h00032FF1 , 32'hFFFCFAF3 , 32'hFFFF6997 , 32'h00059B53 , 32'h00049FF6 , 32'h00067C36 , 32'hFFFBE9D7 , 32'h0004A22A , 32'h000503DB , 32'hFFFF4DE5 , 32'hFFFD548F , 32'h0000263E , 32'h0003AED4 , 32'h00001AC7 , 32'h00033D3B , 32'h0001BD89 , 32'hFFFFCAA8 , 32'hFFFF1859 , 32'h00034057} , 
{32'h00035824 , 32'h00016773 , 32'h0000DBE1 , 32'hFFFEFC0F , 32'h0000E14C , 32'hFFFD8163 , 32'h0001D722 , 32'hFFFDE2FF , 32'h0000C21D , 32'hFFFC1E26 , 32'h0000C15A , 32'h0001CC0F , 32'hFFFF9C5C , 32'h0000D91E , 32'hFFFC50BE , 32'hFFFE91E7 , 32'h00009426 , 32'hFFFF97F3 , 32'h0004466B , 32'hFFFCB569 , 32'hFFFB5B28 , 32'hFFFFBC92 , 32'h00028447 , 32'h00010C44 , 32'hFFFA5C45 , 32'hFFFDF25D , 32'h0003250B , 32'h0004819C , 32'hFFFFD577 , 32'h00048415 , 32'h0000539F , 32'h0001FCC7 , 32'h000186CC , 32'hFFFDB972 , 32'hFFFD1BC8 , 32'hFFFCCD81 , 32'h0001F24C} , 
{32'h0001AAEF , 32'h0001A1CD , 32'hFFFF316D , 32'hFFFA2657 , 32'hFFFDEF52 , 32'h0003603C , 32'hFFFCC971 , 32'hFFFBE735 , 32'hFFFEBF64 , 32'hFFFF4296 , 32'hFFFE04E7 , 32'h0001CB97 , 32'h00009942 , 32'hFFFFBBEC , 32'h00039688 , 32'h00045DF8 , 32'hFFFCBA98 , 32'hFFFB7153 , 32'hFFFEB35A , 32'h0000C645 , 32'hFFFE4DE7 , 32'hFFFF0B0D , 32'hFFFD4B74 , 32'h00008B03 , 32'h0001DE93 , 32'h0000D36C , 32'h00018AF1 , 32'h0001D16E , 32'h0000173A , 32'h00006F32 , 32'h00049857 , 32'hFFFE06D7 , 32'hFFFED5F3 , 32'hFFFC7294 , 32'hFFFE9707 , 32'h0001EE08 , 32'h00048743} , 
{32'h00018629 , 32'hFFFD019D , 32'h00038048 , 32'hFFFD9BE0 , 32'hFFFC0D49 , 32'hFFFF4D38 , 32'hFFFA3C6C , 32'hFFFDB37D , 32'h00000B61 , 32'hFFFFDB3D , 32'h0000C850 , 32'hFFFB2CB8 , 32'h000171B1 , 32'hFFFCB5CE , 32'h00012B97 , 32'h0003E912 , 32'h0001A374 , 32'hFFFFDAEE , 32'hFFFE1987 , 32'h0001D193 , 32'hFFFB8C50 , 32'hFFF93E0D , 32'hFFFA983C , 32'h0001AED0 , 32'hFFF89755 , 32'hFFFDE863 , 32'h0000E3F1 , 32'h0001564E , 32'hFFFB5C4E , 32'hFFFCA07F , 32'hFFFDFA8B , 32'h00003BC0 , 32'h0004FD90 , 32'h00014A75 , 32'hFFFE094C , 32'hFFFD8EC4 , 32'h0000E043} , 
{32'hFFFC43C0 , 32'h0006133D , 32'h00023E37 , 32'h0002DF3F , 32'h00011FF6 , 32'hFFFCCA1A , 32'h0000E74F , 32'hFFFEC514 , 32'hFFFB5DA6 , 32'hFFFBDED7 , 32'h00028326 , 32'h00009473 , 32'h00032817 , 32'h00031C4F , 32'h00040D28 , 32'h00025563 , 32'hFFFBACA7 , 32'h0001C830 , 32'h0001746F , 32'h00057F6A , 32'hFFFF2349 , 32'hFFFE7CBB , 32'h00052AE9 , 32'hFFF9A2A2 , 32'hFFFBD7D9 , 32'hFFFDA8D5 , 32'hFFF74437 , 32'h000000DC , 32'hFFFFA40E , 32'h0003746F , 32'h0000A716 , 32'hFFFBB395 , 32'hFFFC5B54 , 32'hFFFFAA8C , 32'hFFFBE382 , 32'h000452EE , 32'hFFFD661A} , 
{32'hFFFF54EA , 32'h00029E10 , 32'h0000B78F , 32'h00021333 , 32'hFFFFBF30 , 32'hFFFEA40D , 32'h0004F0D8 , 32'hFFFA01D3 , 32'h00010853 , 32'hFFFE6BFD , 32'h0000E70B , 32'hFFFDAEAD , 32'h0001636E , 32'h00012271 , 32'h0006BB3F , 32'h00008856 , 32'hFFFB7889 , 32'h00053520 , 32'hFFFF37E5 , 32'hFFFDAC3D , 32'h000526DE , 32'hFFFA15CB , 32'hFFFE18FC , 32'h0003517D , 32'h0004F245 , 32'h00031CBE , 32'h0003EB8D , 32'h0002982E , 32'h00030D3D , 32'hFFFC6A95 , 32'h00030E5E , 32'hFFFF12D8 , 32'h00015FF4 , 32'h0000F376 , 32'hFFFE64DF , 32'h000061F3 , 32'hFFFF031E} , 
{32'h000145CA , 32'hFFFA2BDC , 32'hFFFE9311 , 32'h0000ECA2 , 32'hFFFFC1E4 , 32'h00014A68 , 32'h0005FCAA , 32'hFFFDA693 , 32'hFFFFAD42 , 32'h0002BF58 , 32'hFFFFCBFB , 32'hFFFC19A4 , 32'h00054434 , 32'hFFFB3374 , 32'h00005620 , 32'hFFFFF7E0 , 32'hFFFD2481 , 32'hFFFC961E , 32'h00016BE0 , 32'h000301C4 , 32'hFFFF382D , 32'hFFFE440B , 32'hFFFF0513 , 32'h0003A59D , 32'hFFFDFE7D , 32'h000327EC , 32'hFFFDCD28 , 32'h00004487 , 32'h0001409D , 32'hFFFEB959 , 32'h0002E69C , 32'h0003B764 , 32'hFFFE4782 , 32'hFFFCBBB3 , 32'h00011D5C , 32'h0002257C , 32'hFFFAFBE2} , 
{32'hFFFFF45B , 32'hFFF507FA , 32'h0008E278 , 32'hFFFD42D5 , 32'hFFFA7A3D , 32'hFFFC4EB7 , 32'h0007137F , 32'h0003A7FF , 32'hFFFEBF10 , 32'hFFFE1426 , 32'hFFFFEE24 , 32'h0003A36F , 32'h0005821E , 32'h0003E777 , 32'hFFF9DE93 , 32'h00006CD9 , 32'hFFFC0D69 , 32'h00063B85 , 32'h00021D63 , 32'h000229EC , 32'hFFFEE856 , 32'hFFFBF803 , 32'h00018419 , 32'hFFFD67AD , 32'h0003B1E0 , 32'h00076EC3 , 32'hFFFF15A8 , 32'hFFFDC2CD , 32'h000208D2 , 32'hFFFB5D19 , 32'hFFF897F4 , 32'hFFFEB8B8 , 32'h0007EF9E , 32'hFFFD5E57 , 32'hFFF5174B , 32'h0002D177 , 32'h000049C4} , 
{32'h00021086 , 32'hFFFB98BD , 32'hFFFFC35B , 32'hFFFEF704 , 32'h0004EFB9 , 32'h000346E3 , 32'hFFFD065F , 32'h0001077A , 32'hFFFF317B , 32'hFFFC6691 , 32'h0007413A , 32'hFFFF8EA3 , 32'h0003249F , 32'hFFFBDA24 , 32'h0001FC03 , 32'hFFFA08A6 , 32'h0006285E , 32'h00040E5C , 32'hFFFF3D57 , 32'hFFFB32C0 , 32'h00018FF9 , 32'hFFFCA383 , 32'h0005D182 , 32'hFFF588AD , 32'h0000B85F , 32'hFFFE211F , 32'h00007B98 , 32'h0006DC7E , 32'hFFF9B665 , 32'h00034B43 , 32'h0003608E , 32'h00000965 , 32'h0001CBA2 , 32'h0003A7EB , 32'hFFFBDA1C , 32'hFFF61166 , 32'hFFFD94D4} , 
{32'h000227D5 , 32'h00015532 , 32'h0006A875 , 32'h0001AD39 , 32'h000159D9 , 32'h0004A139 , 32'h00021773 , 32'hFFFEB035 , 32'hFFFF553A , 32'hFFFF8F36 , 32'hFFFF8ED1 , 32'h0003D598 , 32'hFFFCB22C , 32'hFFFF2936 , 32'hFFFA8EDC , 32'h0000047B , 32'h00006A54 , 32'h0001FB83 , 32'h00054C6C , 32'hFFFD5AC6 , 32'h0001F36A , 32'h0000BD26 , 32'hFFFFC51D , 32'hFFFD5B16 , 32'h0002387F , 32'hFFFFA124 , 32'hFFF83F25 , 32'hFFFE148C , 32'h0004EA8D , 32'h000582EF , 32'h00006BC1 , 32'hFFFDF02E , 32'hFFFF7A3D , 32'h00003294 , 32'hFFFC801F , 32'hFFF91F05 , 32'hFFFF71A4} , 
{32'h0001E4D7 , 32'hFFFF732B , 32'h00011812 , 32'h0000A4EC , 32'hFFFC7199 , 32'h0004FF99 , 32'h00011CE5 , 32'hFFFBA432 , 32'h00015250 , 32'hFFFEEAC1 , 32'h0001C65D , 32'h000061A7 , 32'h000015E3 , 32'hFFFE9B19 , 32'hFFFFFEDC , 32'h0000499A , 32'h000046EB , 32'hFFFB934E , 32'h0004328A , 32'h00004F12 , 32'hFFFDB639 , 32'hFFFEF961 , 32'h0000DDED , 32'h000107A4 , 32'hFFFF8FE1 , 32'hFFFBC31E , 32'h00008EFE , 32'hFFFFB3D9 , 32'h0000D44F , 32'hFFFFFB3C , 32'hFFFDCF14 , 32'h00018BE2 , 32'hFFF8CBD6 , 32'h00031EF1 , 32'hFFFEE75D , 32'hFFFFACFF , 32'h0000B177} , 
{32'h00012FB8 , 32'h00017838 , 32'h00047A99 , 32'h00024C4C , 32'h0000ADD2 , 32'hFFFCEB5C , 32'hFFFA431B , 32'h0000BD06 , 32'h0004768E , 32'hFFFF3224 , 32'h0002E11D , 32'h00027F36 , 32'h0001196B , 32'hFFFD1DAE , 32'hFFFE6190 , 32'hFFFFA500 , 32'h000647BD , 32'h00013F1C , 32'hFFFD90AC , 32'h00006FE9 , 32'hFFFEE6C5 , 32'h00015708 , 32'h0000DA97 , 32'h0005654F , 32'hFFFD5D84 , 32'h0003A741 , 32'h0003459A , 32'h00023F33 , 32'hFFFF8318 , 32'hFFFE91CD , 32'hFFFEC0DF , 32'h0003585D , 32'hFFFCC4C3 , 32'hFFFF4B74 , 32'h00014725 , 32'h00017BCA , 32'h00001505} , 
{32'h0002EEA1 , 32'hFFFE13BC , 32'hFFFB5679 , 32'hFFFF1713 , 32'hFFFE908A , 32'h00007FFF , 32'h00008B1E , 32'hFFFEB61B , 32'h0004CD93 , 32'hFFFCF258 , 32'h00049F80 , 32'hFFFDD5A9 , 32'h0001FEA1 , 32'hFFFDCCE6 , 32'h00017FC6 , 32'h000542EA , 32'hFFFDA9EA , 32'hFFFBBF8E , 32'hFFFFA2C1 , 32'h0003B24C , 32'h000107C9 , 32'h00043358 , 32'hFFFECC1D , 32'hFFFF8520 , 32'hFFFFB43C , 32'hFFFD18C4 , 32'h00056C20 , 32'h000251A2 , 32'h0001D33D , 32'hFFFB30F8 , 32'hFFFFB1D3 , 32'h0003CF0E , 32'h00009C87 , 32'h00008A0B , 32'h00004312 , 32'h00021A9B , 32'h0002F3A7} , 
{32'h000204E9 , 32'h00039523 , 32'h00056B52 , 32'hFFFF53BB , 32'hFFFDBEA5 , 32'h000749A6 , 32'hFFFCC443 , 32'h000492C6 , 32'hFFFE9DC4 , 32'hFFFFEFC7 , 32'hFFFCC07E , 32'h00064320 , 32'h000577D3 , 32'h0002AF5B , 32'hFFF86093 , 32'hFFFE3584 , 32'h0004B1DD , 32'hFFF9FD24 , 32'hFFFE71FA , 32'h0001984D , 32'hFFFB469B , 32'h0001748D , 32'hFFFF96B5 , 32'h00011041 , 32'h00002DF1 , 32'hFFFD35F0 , 32'hFFFB35CE , 32'h0003761B , 32'h0001A432 , 32'h0006968F , 32'hFFFA4FB5 , 32'hFFFF0675 , 32'hFFFF9F8A , 32'h0000D4A1 , 32'hFFFDC147 , 32'h00052A34 , 32'hFFFA84FB} , 
{32'h00032163 , 32'hFFF9FF7A , 32'h0001D9FF , 32'hFFFF4CA6 , 32'hFFF91DE7 , 32'h0002D49F , 32'h00027D11 , 32'hFFFCFBED , 32'h0003D3D8 , 32'hFFFD5CE0 , 32'h0002CCE4 , 32'hFFFF60B8 , 32'h00023AC8 , 32'h00001082 , 32'hFFF97E85 , 32'h0000DFFA , 32'hFFFD9BDC , 32'hFFF92BAE , 32'h00081169 , 32'h000051B4 , 32'h000059F8 , 32'hFFFDBD77 , 32'h0004BD72 , 32'hFFFEE524 , 32'h0003626B , 32'hFFFF01D2 , 32'h00037140 , 32'h000109C8 , 32'hFFFDFF21 , 32'h00001FFD , 32'h0001EC2A , 32'h0000EFA7 , 32'h00016F8F , 32'h00026BF3 , 32'h000101C5 , 32'h0002CBD5 , 32'h0002E43B} , 
{32'hFFFFC271 , 32'h00039265 , 32'h00037947 , 32'h0007E0BF , 32'hFFFF3728 , 32'h00023AEC , 32'h0001E5EA , 32'h0000EA1C , 32'hFFFA1439 , 32'hFFF97493 , 32'h000087C3 , 32'hFFFCFA27 , 32'h000056FF , 32'hFFFA79FD , 32'hFFFFA133 , 32'h000224AB , 32'h00002667 , 32'h000319FC , 32'hFFFFD83E , 32'hFFFA1047 , 32'hFFFE03AB , 32'h00027825 , 32'h0000593D , 32'h0001711A , 32'h0004CE3C , 32'hFFFC59EA , 32'hFFFF05C1 , 32'hFFFF2477 , 32'hFFFDC785 , 32'h00002A34 , 32'h00056351 , 32'h0000ED8A , 32'hFFFE8597 , 32'hFFFB4FAC , 32'h00035793 , 32'h00059E1A , 32'h000451EA} , 
{32'hFFFF378F , 32'h00015BDE , 32'h0004EE76 , 32'hFFFFF11C , 32'hFFFEB1B5 , 32'hFFFE959F , 32'hFFFBFF9C , 32'h00026D16 , 32'hFFFE0628 , 32'h00047439 , 32'h0000837A , 32'hFFFC539F , 32'h00024696 , 32'hFFFE5E7B , 32'h00012741 , 32'hFFFCB2F7 , 32'hFFFE273C , 32'h00015134 , 32'hFFFC6EAD , 32'hFFFD663C , 32'hFFFE55FB , 32'hFFFF46D7 , 32'h0001555E , 32'h00025F97 , 32'hFFFD61BF , 32'h000198B1 , 32'hFFFB2E28 , 32'hFFFE47D6 , 32'h000245F4 , 32'h00070111 , 32'h00002A52 , 32'h000507B8 , 32'h0005E0A2 , 32'hFFFF390E , 32'hFFFB63FC , 32'h00037E56 , 32'h0001F1EC} , 
{32'h0005374D , 32'h0000D17F , 32'hFFFFF132 , 32'h0002B04A , 32'hFFFD1A2F , 32'hFFFEBE54 , 32'h0001E5AE , 32'h000024F6 , 32'hFFF9B3FE , 32'h00021566 , 32'hFFFBDF5F , 32'hFFFDD9CE , 32'hFFFE1EB6 , 32'hFFFB0418 , 32'h000443A5 , 32'hFFFD4ED4 , 32'h0000D4A3 , 32'hFFFA6BBC , 32'h00019F1D , 32'hFFFBDA62 , 32'h000049A2 , 32'h0002F5AA , 32'hFFFAF0A3 , 32'h00010ACD , 32'h0003B112 , 32'hFFFE4E8D , 32'h00004843 , 32'h0002CCD7 , 32'hFFFCDF36 , 32'h000126D0 , 32'h00004681 , 32'hFFFE91A6 , 32'hFFFE6D42 , 32'h0006546F , 32'hFFFD37F9 , 32'hFFFAD38E , 32'hFFFDC286} , 
{32'h0002468C , 32'h0000CFCD , 32'h0002A978 , 32'hFFFF2D10 , 32'hFFFFCDEB , 32'hFFFF3B0B , 32'hFFFF9593 , 32'h000520F8 , 32'hFFFC7FFD , 32'hFFFE1E87 , 32'hFFFDF074 , 32'h00026DA5 , 32'h000217A1 , 32'hFFFEB258 , 32'hFFF99541 , 32'h000305ED , 32'h0000920A , 32'h00000344 , 32'hFFFE67B9 , 32'h0003BCAD , 32'h00013791 , 32'h00023B50 , 32'h00018A99 , 32'hFFFF6BA0 , 32'h0002E689 , 32'hFFFEF015 , 32'h000167D7 , 32'hFFFBD3CF , 32'h00028218 , 32'hFFFEB2C2 , 32'h0001EF57 , 32'hFFFFF15D , 32'hFFFD77C2 , 32'h000190F7 , 32'hFFFE33F5 , 32'hFFFEC551 , 32'hFFFF4BC9} , 
{32'hFFFF805C , 32'h00017906 , 32'hFFF80814 , 32'hFFFAB8C1 , 32'hFFFC9948 , 32'h000414BC , 32'hFFFBC686 , 32'h000311C5 , 32'hFFFF758B , 32'h0005F0ED , 32'hFFFBDE58 , 32'h00005A65 , 32'hFFFC586A , 32'h0002CCDD , 32'h00017466 , 32'hFFFFF048 , 32'h00066123 , 32'h0003CC00 , 32'h0001027A , 32'h0003369D , 32'hFFFE3358 , 32'h00027622 , 32'hFFFFEB68 , 32'h00050B32 , 32'h0000F8EE , 32'hFFFC9A69 , 32'h0003D876 , 32'hFFFB6F28 , 32'hFFFD0DB8 , 32'h00041CED , 32'h0005CBA0 , 32'h0005D547 , 32'h0006B9FF , 32'hFFFD0F08 , 32'h00002B9B , 32'h000100DA , 32'h00027120} , 
{32'hFE247FC0 , 32'hFA697280 , 32'hFCBD2C74 , 32'h05DBAAB8 , 32'hFEA7C95C , 32'hFF64AC49 , 32'hFE45C8B0 , 32'h0336EA04 , 32'h07189318 , 32'hFE5B7574 , 32'h00F13BA1 , 32'h05B067E8 , 32'hFE9ABA80 , 32'hFE39158C , 32'h013CAA44 , 32'hFA2D8578 , 32'h020F4A28 , 32'h014EC9B8 , 32'hFAE276F0 , 32'hF8FB7128 , 32'h05B89FD0 , 32'h006A9B38 , 32'hFEEDB354 , 32'h088AC240 , 32'hFFE0ADF3 , 32'h044F8BD8 , 32'h08563110 , 32'h022E6404 , 32'h01DBDA04 , 32'h00E51720 , 32'h00861F91 , 32'hFC953948 , 32'hFAC83D50 , 32'h0346B34C , 32'hFBC1A4F8 , 32'h02D77B3C , 32'hFD4B011C} , 
{32'h000106BF , 32'h00018AEC , 32'hFFFCFE15 , 32'h0001AA84 , 32'hFFFD3BC8 , 32'h000281BA , 32'hFFFFF568 , 32'hFFFDE01C , 32'h00039D15 , 32'hFFFF9B06 , 32'h000005C6 , 32'hFFFD9263 , 32'hFFFB107F , 32'h0003FFE4 , 32'h0001B971 , 32'hFFFE31BD , 32'h0000DB23 , 32'hFFFFE0D9 , 32'h000172DB , 32'h00008B08 , 32'h0001EAE1 , 32'h000112B0 , 32'hFFFEA91F , 32'hFFFDAA4C , 32'h00019F37 , 32'h00036E3E , 32'h0001E86C , 32'hFFFFC582 , 32'h0001481F , 32'hFFFECFD1 , 32'hFFFF14A4 , 32'h00014489 , 32'h0001D070 , 32'h0001CFE7 , 32'h00054658 , 32'hFFFF150A , 32'h00007CBB} , 
{32'hFDE3D4C4 , 32'hF9AB4250 , 32'hFC4F0E0C , 32'h06A4A1A0 , 32'hFE78DBD0 , 32'hFF50D926 , 32'hFE0F7A9C , 32'h039E26D0 , 32'h080C0BB0 , 32'hFE25A030 , 32'h01113E40 , 32'h066E6C58 , 32'hFE6EAE70 , 32'hFDFCA1E0 , 32'h016918F0 , 32'hF96527B8 , 32'h02593F84 , 32'h017C82EC , 32'hFA2DD8B8 , 32'hF80AEBF8 , 32'h06736558 , 32'h007B8040 , 32'hFEC824AC , 32'h09B208C0 , 32'hFFDBEFC6 , 32'h04E13838 , 32'h0976CCE0 , 32'h027D97CC , 32'h0219AC3C , 32'h0103E398 , 32'h009632A4 , 32'hFC21A53C , 32'hFA112E80 , 32'h03B9D8E8 , 32'hFB332DD0 , 32'h033C18CC , 32'hFCECC124} , 
{32'hF13A90C0 , 32'h0B17D060 , 32'h05B1D000 , 32'hFB37F2F0 , 32'h049728A8 , 32'hF1D7FAF0 , 32'h07026730 , 32'hFC65FCC0 , 32'h0F57B7A0 , 32'hFE40F220 , 32'hEFBDCA20 , 32'h04CC4690 , 32'h0ABA76D0 , 32'h03F3C898 , 32'h04847268 , 32'h0262BC6C , 32'h06C0BD80 , 32'h00DA4FC4 , 32'h009E04E6 , 32'hFD806F94 , 32'hFE0E18B8 , 32'hFE2D79C8 , 32'hFBB64FB0 , 32'hFFD90273 , 32'hFD0ECC48 , 32'hFC8644FC , 32'h0B6C2710 , 32'hF5B38F50 , 32'h006E6B80 , 32'h07160860 , 32'hF7A47A20 , 32'hFBC63B80 , 32'h06AB7528 , 32'hFC2A4608 , 32'h02402C54 , 32'h02A10760 , 32'hFEABE414} , 
{32'h079C9ED0 , 32'hF1D7BBD0 , 32'hFF128DB6 , 32'h02C2C928 , 32'hFC9E5D64 , 32'hFCBD3050 , 32'hFAEB6878 , 32'h08FBA260 , 32'h0FF77CE0 , 32'h00417313 , 32'hFF055B82 , 32'h0B25BB90 , 32'h000607DD , 32'h07E75B90 , 32'h043E4D68 , 32'hF2F60B00 , 32'h0475B360 , 32'hFE983610 , 32'hF180E790 , 32'hF4F112D0 , 32'h02201A7C , 32'h049FDE08 , 32'hFD23EFA4 , 32'h06D50410 , 32'h05CBA450 , 32'hFE2E61B4 , 32'h09040D90 , 32'hFCC10FDC , 32'h01DEA260 , 32'hFDAFE6B0 , 32'h01701A28 , 32'hF8A30EC0 , 32'hFEA83BE4 , 32'h0F613F40 , 32'hF991E988 , 32'h02CBF754 , 32'hFC7148B0} , 
{32'h16B7E4A0 , 32'hF545C6C0 , 32'hFAC6D438 , 32'h02C45D68 , 32'h00222629 , 32'hFF18F7E6 , 32'h0869B900 , 32'hFB0287E0 , 32'h056E4648 , 32'h05434F38 , 32'hFCCAA950 , 32'hFE4F9594 , 32'h02586848 , 32'h1B69F380 , 32'hFCE0F178 , 32'hFA0A83C8 , 32'h08716C40 , 32'h07CE0728 , 32'hF262E2A0 , 32'hFE69581C , 32'h0032F70C , 32'h067106F8 , 32'h0D459BA0 , 32'h03F1236C , 32'h05873730 , 32'hFC431A28 , 32'hFB4A23D8 , 32'hED07D380 , 32'h03DF3AF8 , 32'hFB234E68 , 32'hF04C9690 , 32'hFCEC65D0 , 32'h0C62EA80 , 32'h098797D0 , 32'hFB5EDA90 , 32'h01A057EC , 32'h0142A070} , 
{32'hFDB0A960 , 32'hF689C9F0 , 32'hFAB30140 , 32'h09EE08B0 , 32'hFDC175D8 , 32'hFCAF4518 , 32'hFB568910 , 32'h0B9991E0 , 32'h09D66E10 , 32'h0082B32C , 32'h018A0C2C , 32'h0A0C3870 , 32'hFD374F7C , 32'hFBBFFE50 , 32'h04D15E90 , 32'hF434CFB0 , 32'h06608BD8 , 32'h035C5B10 , 32'hF8527BC0 , 32'hF14D2300 , 32'h0805FCE0 , 32'h0437FEF8 , 32'hFF43BC10 , 32'h112D8F40 , 32'hFF8F9B49 , 32'h0614FD98 , 32'h142A1480 , 32'h033FCA6C , 32'h07C83EB0 , 32'h0554FCD8 , 32'h05F1BED0 , 32'hF9EEB6E8 , 32'hF3D54920 , 32'h07886BB8 , 32'hF73BAA10 , 32'h0400DD68 , 32'hFFAFD6C8} , 
{32'h05AA6470 , 32'hFADE9128 , 32'h008AE22B , 32'h004B501E , 32'hFC244A54 , 32'hFD899AE0 , 32'hFECA8D48 , 32'hFDF8A228 , 32'hE7332520 , 32'hFA91C1C0 , 32'h024A380C , 32'hF60CF300 , 32'hF00130E0 , 32'hFA549E50 , 32'hF7666700 , 32'hEC0BE500 , 32'h0CAA45B0 , 32'hFD496008 , 32'h0C1F6EA0 , 32'h06877190 , 32'h00916F22 , 32'h0AA31190 , 32'h0BD4E000 , 32'h06E82F88 , 32'h087EC3A0 , 32'hF6A2F0D0 , 32'hF8E9F168 , 32'h01466944 , 32'h03079E3C , 32'hFC1232A8 , 32'h0A2D9800 , 32'hFF93090C , 32'hF73D4390 , 32'h05613350 , 32'hF0B6BEA0 , 32'hFDBBB308 , 32'h01FB3B28} , 
{32'hFE306CF0 , 32'h00F1190B , 32'hFF48171E , 32'h0143732C , 32'hFED9C490 , 32'h003B1C4D , 32'hFF6C6058 , 32'h0059D4B6 , 32'hFF30F7B6 , 32'h02825944 , 32'hFE90478C , 32'hFF235019 , 32'hFE3D5098 , 32'hFFB7CD6B , 32'h00CFFC7D , 32'hFFD31D03 , 32'h009FCF7A , 32'hFE3E3F68 , 32'hFCB8079C , 32'hFFBB62C8 , 32'hFD5C7620 , 32'h0361B3B8 , 32'hFF5B928E , 32'hFEF72EF0 , 32'hFF13EA4C , 32'hFEE98BE8 , 32'hFECC4A0C , 32'hFF9D7EEB , 32'hFF4ACA37 , 32'hFF228F76 , 32'hFE7E207C , 32'hFDE6C80C , 32'h0064E02C , 32'hFFB0D417 , 32'h013A3CB0 , 32'h00D88309 , 32'h0036334D} , 
{32'hFF6691C3 , 32'h020A78E4 , 32'h058B4228 , 32'h00C92D8B , 32'hFEDC857C , 32'hE685DE40 , 32'h06296358 , 32'h0996C780 , 32'hE6AC7C60 , 32'hF9613510 , 32'hFD3366C4 , 32'hFBBD8948 , 32'hFF84143B , 32'hFFBDB402 , 32'h01980A34 , 32'hEF5ADA40 , 32'h0D055D90 , 32'h0458C848 , 32'h0B41D7B0 , 32'hFEA49698 , 32'hF8FFBE78 , 32'h14C60420 , 32'h03BA62E8 , 32'h07E81F68 , 32'h08392030 , 32'hFDC9E668 , 32'h01A968B0 , 32'h0BF85D30 , 32'hFEFA0BEC , 32'hFBCA2808 , 32'h02228114 , 32'h01AF1568 , 32'h02F1B980 , 32'h03D5CBB8 , 32'hF19592C0 , 32'hF80D9980 , 32'hFBA4F2D8} , 
{32'h0773D208 , 32'hFCB75D88 , 32'h07311AD0 , 32'hED1A4DC0 , 32'h033F826C , 32'hFD201604 , 32'hFC59B0D8 , 32'hEDBE76A0 , 32'h07369D00 , 32'h1C5615A0 , 32'h0A3D85F0 , 32'hFF863705 , 32'hF0FAB4A0 , 32'hF874B9F8 , 32'hF9AA7210 , 32'hF0879070 , 32'h08C28A00 , 32'h0561B4A8 , 32'hF5AD5E60 , 32'h063FF1A8 , 32'hFA68CD60 , 32'hFC82BBB4 , 32'hEA1BC540 , 32'h064FC0A8 , 32'hF7CB5080 , 32'hEF7D8640 , 32'h04DB4B58 , 32'h165C7F00 , 32'h0C788230 , 32'hFB4F5E40 , 32'h00DF0EE7 , 32'hFFF2864D , 32'hF9757CE8 , 32'hF4BE7D80 , 32'h0B252900 , 32'h06192D28 , 32'hFFE1C0AD} , 
{32'hF09D18C0 , 32'h077D5020 , 32'hF95FAC38 , 32'h0AB34B30 , 32'h00B6112C , 32'h0724AE90 , 32'hFEA59D0C , 32'h06FC2ED0 , 32'hF63673C0 , 32'hFB8C0108 , 32'h01169BB8 , 32'h01D97E64 , 32'hFF969884 , 32'hF2654A30 , 32'hF9B09A30 , 32'h03806F5C , 32'hFCDAE604 , 32'h01A01238 , 32'h023C1E08 , 32'hFFEE1BD2 , 32'h0410E868 , 32'hFB16E888 , 32'hF9E2FF28 , 32'hFF5837F7 , 32'hFD4E8264 , 32'h00B564C6 , 32'hFFF2BC14 , 32'h0CD9B7C0 , 32'hFE3DA400 , 32'h000A48C7 , 32'hFDF461C4 , 32'h031184CC , 32'hF8747430 , 32'hF4C05490 , 32'h07AAE440 , 32'hF97ABD08 , 32'hFC02CC30} , 
{32'hF9873C88 , 32'h0432E1A8 , 32'hFDB30820 , 32'h019DB7B0 , 32'h00162BF5 , 32'h03970DC0 , 32'hFFD46F8F , 32'hFF58AADA , 32'hFBA912C0 , 32'hFD483D68 , 32'h003490F1 , 32'hFF1706B7 , 32'hFE8B8BD4 , 32'hF883A440 , 32'hFD7EEAE0 , 32'h02561350 , 32'hFD9F49CC , 32'hFFCE74E6 , 32'h044A4EC0 , 32'hFF2347FE , 32'h02F8F07C , 32'hFBAAFE18 , 32'hFF0B7CE5 , 32'hFF60FD63 , 32'hFDF6FF68 , 32'h0187E5E8 , 32'h01687D28 , 32'h069A5ED8 , 32'hFF0449E4 , 32'h008D253B , 32'hFFCAA492 , 32'h00CECCE3 , 32'hFD4DC2C0 , 32'hFC50A2EC , 32'h017E2470 , 32'hFFDBDB07 , 32'hFF59A262} , 
{32'hF2DB1500 , 32'h0885D600 , 32'hFB4B1480 , 32'h0343120C , 32'h002DB94A , 32'h07461E18 , 32'hFFAA5E9E , 32'hFEA6A068 , 32'hF731D3F0 , 32'hFA831F30 , 32'h0067C7AC , 32'hFE1DA508 , 32'hFD107B0C , 32'hF0D1EA70 , 32'hFAF07A70 , 32'h04BC20E8 , 32'hFB2F6DF0 , 32'hFF9F09B5 , 32'h08B86030 , 32'hFE3CAFC4 , 32'h060513C8 , 32'hF7392B50 , 32'hFE120E40 , 32'hFEBC70B8 , 32'hFBDB0BC8 , 32'h0315EAA0 , 32'h02DAE610 , 32'h0D60AD80 , 32'hFE08FF08 , 32'h0121CA70 , 32'hFF92B05A , 32'h01A13D90 , 32'hFA899210 , 32'hF8816400 , 32'h03083198 , 32'hFFB319BE , 32'hFEAE2258} , 
{32'h000262D6 , 32'h0000116D , 32'h00012F47 , 32'h0001D5CF , 32'h0006DC7B , 32'h00016690 , 32'hFFFFB54E , 32'h0000E871 , 32'h0002A6A8 , 32'h0000C1A1 , 32'h0000CD3A , 32'h0000D804 , 32'hFFFE7EAB , 32'hFFFF5CBE , 32'hFFFDE6BA , 32'h0000B166 , 32'hFFFFF7F8 , 32'hFFFC9586 , 32'hFFFCE566 , 32'h00038F29 , 32'hFFFF97CE , 32'hFFFEF338 , 32'h000318F0 , 32'hFFFEB293 , 32'h0002CF18 , 32'hFFFFDBC2 , 32'h00008C39 , 32'hFFFFEEB2 , 32'hFFFF73E4 , 32'hFFFFA39C , 32'hFFFF4E54 , 32'hFFFD3992 , 32'h0000EBEF , 32'h00002DAD , 32'hFFFE828F , 32'hFFFFDFEA , 32'hFFFBB512} , 
{32'h00008C52 , 32'h0003E8E8 , 32'hFFFFE1C2 , 32'h00020F51 , 32'h00006E7F , 32'hFFFFEAF9 , 32'hFFFA93A3 , 32'h000578A1 , 32'h000269E5 , 32'hFFFEC601 , 32'hFFFC4DCA , 32'hFFFF4BEC , 32'h00076F6A , 32'h000404AE , 32'h00035043 , 32'hFFFE81F4 , 32'hFFFD2B90 , 32'hFFFEEF35 , 32'h0002886C , 32'hFFFC5E51 , 32'hFFFC0437 , 32'hFFFF46E0 , 32'h0003A025 , 32'h0000C382 , 32'h00000D3F , 32'hFFFCC0CA , 32'h0000A200 , 32'hFFFF561B , 32'hFFFF54D3 , 32'hFFFDAF6B , 32'hFFFBE702 , 32'hFFFFEC10 , 32'hFFFF315E , 32'hFFFC3EE4 , 32'hFFFE12F3 , 32'hFFFE0CA5 , 32'hFFFED788} , 
{32'h0000F678 , 32'hFFFD0220 , 32'h00011336 , 32'h00039FD9 , 32'h0002F026 , 32'hFFFBCA8D , 32'hFFFFDF43 , 32'h0003ACCC , 32'h00023697 , 32'hFFFE0D87 , 32'hFFFE0C4D , 32'h00029725 , 32'hFFFB5442 , 32'h0002E929 , 32'hFFFFBA7F , 32'h00030D0D , 32'hFFFF8182 , 32'h0001E87C , 32'hFFFFF72D , 32'hFFFE4B49 , 32'h00018722 , 32'h0003D818 , 32'h0003496C , 32'h0005566E , 32'h0000D05F , 32'hFFFD1545 , 32'h0003B24F , 32'h0002D12F , 32'h00024A0C , 32'hFFFE5590 , 32'h00030A73 , 32'h0001798F , 32'h000320F3 , 32'hFFFDD5EB , 32'h0002073C , 32'hFFFAF85C , 32'hFFFC7F21} , 
{32'hFFFEDFC3 , 32'hFFFE9185 , 32'h0001E202 , 32'h000383E0 , 32'hFFFEC41D , 32'h00008738 , 32'h000593F4 , 32'h00025A61 , 32'hFFFDBFDC , 32'hFFFF2C66 , 32'hFFFEB027 , 32'h0000BD97 , 32'hFFFB0B99 , 32'hFFF8F485 , 32'h0001F795 , 32'h0002786B , 32'h000311C2 , 32'hFFFB2A95 , 32'hFFFF3552 , 32'h00073530 , 32'h00023089 , 32'hFFFE0359 , 32'h0005FF4D , 32'hFFFCEBCC , 32'h0001ADD6 , 32'hFFFF7B4F , 32'h0000D66A , 32'h0002BCF5 , 32'h0001F1EB , 32'h00021BE3 , 32'hFFFF3054 , 32'h0001EBBE , 32'h00014F89 , 32'h000492CE , 32'h00024AFB , 32'h00004250 , 32'hFFFDEFB6} , 
{32'h00007DB5 , 32'hFFFD4F0A , 32'h00038E24 , 32'hFFFEDB0B , 32'hFFFF7644 , 32'h0002143A , 32'hFFFE3463 , 32'h0002B8ED , 32'h0004BBCE , 32'h0002ABAB , 32'h00019122 , 32'h00025FAD , 32'hFFFAF9DE , 32'h0000BD42 , 32'hFFFAB2BB , 32'h0000C572 , 32'hFFFAB04E , 32'hFFFFBE59 , 32'hFFFFA38C , 32'h0002548C , 32'h000194AE , 32'h00000495 , 32'h00003409 , 32'hFFFADE85 , 32'hFFFCD753 , 32'h00011646 , 32'hFFFE73A3 , 32'h00002FDA , 32'h00060737 , 32'hFFFA9E63 , 32'h00046553 , 32'hFFFEB2A1 , 32'hFFFEFBBA , 32'h00043E28 , 32'hFFFB4493 , 32'hFFFA2BC8 , 32'hFFFE1151} , 
{32'h0000B928 , 32'hFFFBE7CA , 32'h00029C87 , 32'h0004686C , 32'h0000B0DA , 32'hFFFD01A5 , 32'h00027245 , 32'hFFFDDF72 , 32'hFFFD1C16 , 32'h000365E2 , 32'h00057B9C , 32'h0000D8FA , 32'hFFFEA4D0 , 32'hFFFDB96E , 32'hFFFDA357 , 32'hFFFFD682 , 32'hFFFC21E2 , 32'h000219BD , 32'h00036F0F , 32'h000565A1 , 32'hFFF94A2A , 32'hFFFE1EDE , 32'h000567DB , 32'h0002DAF8 , 32'h00033AE2 , 32'h00025D23 , 32'h00020D79 , 32'h0003BB6E , 32'h0000E82A , 32'h0000D57D , 32'hFFFCB5C8 , 32'hFFFF529E , 32'h00034AA0 , 32'h00033C59 , 32'h0002A9AD , 32'h0003FAEC , 32'hFFFE9969} , 
{32'h0003751B , 32'hFFFF21C7 , 32'hFFFACABC , 32'hFFF98B7B , 32'hFFFC1188 , 32'h000223EE , 32'h0000326E , 32'h00065660 , 32'hFFFA7A50 , 32'hFFFE97E7 , 32'h0004639A , 32'hFFFC9957 , 32'hFFFFEC49 , 32'h00014F44 , 32'h00004942 , 32'hFFFEBD90 , 32'hFFFD8317 , 32'h00073197 , 32'h00076255 , 32'h0000AA93 , 32'h0000AADB , 32'hFFFD904F , 32'h0000DB55 , 32'h00006F0E , 32'hFFFFCCA3 , 32'hFFFB043E , 32'h000276D8 , 32'h0003BFA7 , 32'h0000E9CD , 32'h00054E15 , 32'h00044AE0 , 32'h00071F6B , 32'h0006268F , 32'hFFFD772F , 32'h0005C7FA , 32'h0002CBC4 , 32'hFFF96D6E} , 
{32'h00030CD4 , 32'h00004113 , 32'hFFFFFCBD , 32'h000030F8 , 32'hFFFF91FC , 32'h00009D14 , 32'h000358D8 , 32'hFFFAED6E , 32'hFFFF9899 , 32'hFFFD72A0 , 32'hFFFF82A8 , 32'h000215A5 , 32'hFFFEE465 , 32'h00025426 , 32'hFFFD8CA4 , 32'hFFFBE20F , 32'h0001D070 , 32'hFFFFDD79 , 32'h0003B4BC , 32'hFFFF2C08 , 32'h00032FBC , 32'hFFFE486D , 32'hFFFBD0C6 , 32'h0001E6BE , 32'hFFFDE688 , 32'hFFFF2BC8 , 32'h000088DA , 32'hFFF97B9F , 32'h00012449 , 32'h0009E7B0 , 32'h00004A50 , 32'h0000310C , 32'h0000CE9B , 32'h0003D11A , 32'h00027847 , 32'hFFFFCFCF , 32'h0001B4DB} , 
{32'hFFFFB079 , 32'h00025AF6 , 32'h000046DA , 32'hFFFEB843 , 32'hFFFD3932 , 32'hFFFFEB87 , 32'h00016ADD , 32'h00028C71 , 32'hFFF9F04B , 32'hFFFB8971 , 32'h00006C54 , 32'h00029DA8 , 32'hFFFDEF6D , 32'h000405A4 , 32'hFFFA6923 , 32'hFFFFC812 , 32'hFFFC3597 , 32'hFFFFFB6B , 32'h00054C26 , 32'h00074FA8 , 32'h00046B34 , 32'h00018827 , 32'h0004B663 , 32'hFFFF4D4F , 32'h00010255 , 32'h0005C322 , 32'hFFFF531B , 32'hFFFDD204 , 32'hFFFFD70D , 32'hFFFE912A , 32'h0000B262 , 32'hFFFD12AC , 32'hFFFC5336 , 32'hFFFE54EA , 32'hFFFF594E , 32'h000477F5 , 32'h00030773} , 
{32'hFFFD6F10 , 32'h0001AA4F , 32'hFFFF4B89 , 32'hFFFECD49 , 32'hFFFEC7E7 , 32'hFFF98D49 , 32'hFFFCBF33 , 32'h00010569 , 32'hFFFD1D9F , 32'h000257D7 , 32'h00013877 , 32'h000323CF , 32'h00062F3B , 32'h0001FD81 , 32'hFFF7EC94 , 32'hFFFE335D , 32'hFFFEED0A , 32'h00012C44 , 32'hFFFEEBDB , 32'hFFFD6DE4 , 32'h0000FE7C , 32'hFFFE72A9 , 32'hFFFBD644 , 32'hFFFF38A8 , 32'hFFFF36A2 , 32'h00008D07 , 32'h0001D2D8 , 32'hFFFEC4D0 , 32'hFFFF8CFF , 32'h00054624 , 32'h000271E4 , 32'hFFFE2E35 , 32'hFFFF79DA , 32'h0002E5F7 , 32'h00016DE0 , 32'h000216D6 , 32'h00009AA1} , 
{32'hFFFFA1EF , 32'hFFFF528A , 32'h000112EF , 32'hFFF66F52 , 32'hFFFE8922 , 32'h00012564 , 32'h0004841F , 32'hFFFD0F04 , 32'h00050770 , 32'hFFFE5C16 , 32'h0001E220 , 32'hFFFA80CE , 32'h00047F4D , 32'h00020CA4 , 32'h000092E3 , 32'hFFFD0EF5 , 32'hFFFD13EB , 32'h0006C8FE , 32'h00002972 , 32'hFFFBF220 , 32'h000026E7 , 32'hFFFD824D , 32'h00033DD8 , 32'hFFFD045E , 32'h00018630 , 32'h00011DF8 , 32'hFFFE7959 , 32'hFFFF3CBB , 32'hFFFC0ED4 , 32'h0000B635 , 32'h0004B01D , 32'h000365C1 , 32'h000239C0 , 32'h0002D6E2 , 32'hFFFF437A , 32'hFFFC475A , 32'h0002269D} , 
{32'hFFFE0007 , 32'hFFFED3BF , 32'h00036B6F , 32'h0003DA5E , 32'h00036286 , 32'h0001DF0F , 32'hFFFF52F2 , 32'hFFFE945F , 32'h0000741F , 32'h00044833 , 32'hFFFE016C , 32'h0000231F , 32'h00030DFC , 32'h00013B3B , 32'hFFFEBBE8 , 32'h0000465B , 32'hFFFF44DE , 32'h00004F50 , 32'h00005EC8 , 32'h00008DFE , 32'hFFFC0BF7 , 32'hFFFF4AA6 , 32'h00023580 , 32'hFFFA60BD , 32'h0002F410 , 32'h000083C3 , 32'h00043BCA , 32'h00017949 , 32'hFFFD97E2 , 32'hFFFC71AE , 32'h00025331 , 32'hFFFCF6B5 , 32'hFFFC6946 , 32'hFFFDB230 , 32'hFFFFE33C , 32'hFFFDC8BB , 32'hFFFFD08C} , 
{32'h0025FAA0 , 32'hFFF4A14A , 32'h0000ECD4 , 32'hFFF825D3 , 32'hFFEAD67A , 32'hFFFB445C , 32'h0002FE44 , 32'hFFE6F46B , 32'h000E1A61 , 32'h0008CB87 , 32'hFFE15B23 , 32'hFFF8DE89 , 32'hFFD1970C , 32'h0014812E , 32'hFFF921AF , 32'h0009CA75 , 32'h001BCE26 , 32'hFFFB92AE , 32'hFFE2802B , 32'h000E8904 , 32'hFFE6831F , 32'h0005EB26 , 32'h000F142D , 32'h00156915 , 32'h000757D2 , 32'h00086BEA , 32'hFFFFB556 , 32'hFFE4C89D , 32'h0007B345 , 32'h00021F66 , 32'hFFF4E921 , 32'hFFF63544 , 32'h000DFEA7 , 32'h0015C381 , 32'hFFE420DD , 32'h0004F220 , 32'hFFFA5F1B} , 
{32'hFA4028E0 , 32'h046ED590 , 32'h02E840F8 , 32'hFFDB47D0 , 32'h0367DCB0 , 32'hF8D27140 , 32'h04004B10 , 32'hFE5AE168 , 32'h087248C0 , 32'hFEFF74D0 , 32'hF982A810 , 32'h0190AD9C , 32'h055990D0 , 32'h0157D3AC , 32'h03D6D244 , 32'h05E4DB08 , 32'h023D777C , 32'h01241370 , 32'h004022BA , 32'hFA16B9A8 , 32'hFE8952AC , 32'hFEB21E24 , 32'hF9E96678 , 32'h00A068B9 , 32'h00631C36 , 32'h0009C81F , 32'h0720A520 , 32'hFF2B2BFC , 32'hFF4A9A14 , 32'h01637DD8 , 32'hFC050190 , 32'h01F0705C , 32'h08481090 , 32'hFDEC0D58 , 32'h041FDAE8 , 32'hFF81CABD , 32'hFE34687C} , 
{32'h01ED0EDC , 32'h057D1548 , 32'h03BE3A80 , 32'h05412448 , 32'h030AF544 , 32'h00FD3A5D , 32'hF8263290 , 32'h01761A24 , 32'h0193FF54 , 32'hFEB87E44 , 32'h0234CF74 , 32'h05237C90 , 32'hFD2E6F84 , 32'h0A02DCA0 , 32'hFC14B43C , 32'h0183098C , 32'h0709B3A0 , 32'hF5A7E280 , 32'h05BCB050 , 32'h04EA6968 , 32'hFBB0C970 , 32'hFBD621F0 , 32'h00DC5F03 , 32'h01A2C5E8 , 32'hFE2D4310 , 32'h0421CD90 , 32'h05E55FE8 , 32'h04BE3D78 , 32'h02E58C9C , 32'hF85222E0 , 32'hFE35E1C4 , 32'hFED5FA10 , 32'h03254354 , 32'h0029D425 , 32'hFDC18694 , 32'h0246DA88 , 32'hFF25324E} , 
{32'hFD0A0A48 , 32'hF7B1C970 , 32'hFB24D488 , 32'h07F4C738 , 32'hFD77C620 , 32'hFED4C53C , 32'hFE0FF6F4 , 32'h04CEE340 , 32'h0A5608E0 , 32'hFD677D50 , 32'h017CCF1C , 32'h08020AE0 , 32'hFE057FC0 , 32'hFDC58F5C , 32'h01C5044C , 32'hF79BC0A0 , 32'h02E62970 , 32'h020EC418 , 32'hF8DC3A40 , 32'hF5FB4A90 , 32'h08288360 , 32'h00FC2688 , 32'hFE995FC4 , 32'h0C38AF20 , 32'hFFB5B304 , 32'h060D53F8 , 32'h0C45DF30 , 32'h03BD60C0 , 32'h0192D044 , 32'h0162CFC4 , 32'h014FD454 , 32'hFAE29598 , 32'hF868BB00 , 32'h044C15F0 , 32'hF99B74F0 , 32'h0452A630 , 32'hFC57DA14} , 
{32'hEFA08FA0 , 32'h029F58B0 , 32'hF24D5E60 , 32'hFFCB0630 , 32'hFC56BF08 , 32'h3499DF40 , 32'h0986DC40 , 32'h00FB8218 , 32'h3D96D740 , 32'hC88D1C80 , 32'hE594EE20 , 32'h0EB78AD0 , 32'h0D264C80 , 32'h2372B640 , 32'hEC366C80 , 32'hE6A569A0 , 32'h040F9B98 , 32'h180B5260 , 32'hDF355800 , 32'h0C0A5000 , 32'h0A18B9D0 , 32'h00673944 , 32'h19045440 , 32'h1F3A39C0 , 32'hF91AF7D8 , 32'hF7207F80 , 32'hECA915C0 , 32'hFC5A0418 , 32'h024C9DF8 , 32'h138A92E0 , 32'hE2B88BC0 , 32'hF4030760 , 32'hFC44E6A0 , 32'h00EC7333 , 32'h15569E60 , 32'h126AB440 , 32'h0EFFA580} , 
{32'h00434DE1 , 32'hF93A76B8 , 32'h09BAE5A0 , 32'h06216C78 , 32'h00B9E54B , 32'hEDB497E0 , 32'h02B4F520 , 32'h094668E0 , 32'h082D4750 , 32'hF06A6CD0 , 32'hFAB841F8 , 32'h0A15D910 , 32'h064D39B8 , 32'h0A7CE3B0 , 32'h020E5480 , 32'hF6077000 , 32'h0E715340 , 32'hFFD737B6 , 32'hF09B9A40 , 32'hFCE7C808 , 32'hFDF90E00 , 32'hFA53AB28 , 32'h044F73D0 , 32'h070AE160 , 32'hFDAEF0E0 , 32'hF7B60F70 , 32'hF4CCA480 , 32'hF98E7E10 , 32'hFE9A4BD4 , 32'h08133710 , 32'hFBC355A0 , 32'hFF85125A , 32'h093D0A20 , 32'h021F0AFC , 32'h0A1D16B0 , 32'h058C4C98 , 32'h06C0BA80} , 
{32'h093DAA40 , 32'hF969ADA0 , 32'hFE715C2C , 32'hF79667E0 , 32'hF8851F90 , 32'hFDF6C05C , 32'h016CE14C , 32'hFFD74E18 , 32'h111200E0 , 32'h0E6114D0 , 32'hEE9C60C0 , 32'h09B16CC0 , 32'hF6D1E8F0 , 32'h2186C440 , 32'hF8EB2710 , 32'h02CC8884 , 32'h0CC63400 , 32'h1117B3E0 , 32'hE96C2180 , 32'h09A86060 , 32'hF64B9FD0 , 32'hF5401350 , 32'h1D80EF40 , 32'h0BC23F60 , 32'hFD8D1EA4 , 32'h05908E68 , 32'hF1F0FD90 , 32'hF047AB10 , 32'h00190FC3 , 32'hF8967198 , 32'hEFB3B980 , 32'hFF8B1F06 , 32'h076BD4E0 , 32'h0D0B97C0 , 32'hEB42DDC0 , 32'h052983A8 , 32'h02F81DB4} , 
{32'h0F1FBC60 , 32'h07BC6DA8 , 32'hF102C7A0 , 32'hF6BA7F60 , 32'h026FAFF0 , 32'hE5766120 , 32'h060563C0 , 32'h1280DFA0 , 32'hF61DCF00 , 32'h1BEC85A0 , 32'hFD9C8570 , 32'h072EE3D0 , 32'hEB3DB000 , 32'h16F11BA0 , 32'hF4B6C0C0 , 32'hFF022013 , 32'h178B5960 , 32'h061E04C8 , 32'hED89CB20 , 32'h10D96860 , 32'hF473D820 , 32'hE24C8920 , 32'h146E8D00 , 32'hFE1AD9F0 , 32'hFEF8FC08 , 32'h08B7FA40 , 32'h01DC6740 , 32'hF23A0210 , 32'hEB18B200 , 32'hF856DD90 , 32'hFDA11464 , 32'hF9D27840 , 32'h1628ADA0 , 32'h131EA340 , 32'hF8E934D0 , 32'h039EAABC , 32'h04369690} , 
{32'h041B0BC0 , 32'h0853A050 , 32'h02A84C34 , 32'h006D99C3 , 32'h08CE8050 , 32'hE602AA60 , 32'h11054200 , 32'hEE23C7E0 , 32'hF2423A70 , 32'h1C256680 , 32'h03B57BD4 , 32'hFF087B42 , 32'hEE6C2320 , 32'h00934950 , 32'hFA019480 , 32'hFC5DC0AC , 32'h03698BB8 , 32'h0259D55C , 32'hF3AE3FC0 , 32'hF38D20F0 , 32'hECBF1F80 , 32'h039C3DF0 , 32'h107EDF60 , 32'h05094528 , 32'h05E9A758 , 32'h09F4D9F0 , 32'h153A61E0 , 32'h019382DC , 32'hE4329DC0 , 32'h093B5A60 , 32'hF5385650 , 32'hF583E110 , 32'hED37D260 , 32'h069190D0 , 32'hF666BE20 , 32'hF38B1FF0 , 32'hFEE3F7EC} , 
{32'h010F7D44 , 32'h13FD3060 , 32'hEB7F9380 , 32'h0FABAD10 , 32'h04699318 , 32'hE5AF8100 , 32'h06CC0860 , 32'hEF5EE380 , 32'hF2480900 , 32'h0078D55D , 32'h02E99634 , 32'hDF900B00 , 32'hFDD9836C , 32'h049D8530 , 32'hFB45AB30 , 32'hEC770EE0 , 32'h049F01C0 , 32'h1659D780 , 32'h074A86D8 , 32'hFD7F3604 , 32'h03EA8608 , 32'h0CF3B580 , 32'h08115740 , 32'h1B1F3500 , 32'h12DF80A0 , 32'hE671B820 , 32'h03E6F54C , 32'h0E05FB80 , 32'hF376B110 , 32'h0331E30C , 32'hF4E700B0 , 32'hFF91577F , 32'h0C1FD080 , 32'h114D1460 , 32'hE62B9260 , 32'hFE3B5018 , 32'h006446BF} , 
{32'hF20ACFD0 , 32'h1DCDF8C0 , 32'h02654CB0 , 32'h0468C338 , 32'h117B8640 , 32'hF21C4E40 , 32'h146BF9E0 , 32'hF0645830 , 32'hED3FEC80 , 32'h0F959840 , 32'hF2866370 , 32'hF63C4DD0 , 32'hEBD2C880 , 32'h0C55AF20 , 32'hF4E85640 , 32'hE6BB3E80 , 32'hF9D84488 , 32'h07325970 , 32'h15600D60 , 32'hF378C8E0 , 32'h01850408 , 32'h11483C40 , 32'h02D06C7C , 32'h1B604140 , 32'h189B5080 , 32'hE7DFA820 , 32'h037B59D0 , 32'h074AA448 , 32'h0BC1A520 , 32'hFAA0FF98 , 32'hF5F2CA10 , 32'h004F97D3 , 32'h0623CA78 , 32'h07937708 , 32'hE2BB5E60 , 32'hFA0D08A0 , 32'hF985DE80} , 
{32'hEC5484A0 , 32'h174B0320 , 32'hEF7C7080 , 32'h05108D48 , 32'h024D2D28 , 32'h1DA09D80 , 32'h103CE7C0 , 32'hF82677A0 , 32'h0EE02020 , 32'hFD20011C , 32'hFB808440 , 32'hEF31ABA0 , 32'h0C09F680 , 32'h13E896E0 , 32'hF6D69BA0 , 32'hED35DD80 , 32'hE7CFF620 , 32'h13B39C20 , 32'hFD472340 , 32'h04B1B8E0 , 32'hFD0C8790 , 32'h1B7825A0 , 32'hF4E4F760 , 32'h1D3DFC20 , 32'hFB0384E0 , 32'hFC2297B0 , 32'hFD163858 , 32'h149B4720 , 32'h0CD98760 , 32'h04A40828 , 32'hFF9AF2D5 , 32'hFE988C38 , 32'h11CC1F80 , 32'h07EE8CC0 , 32'hFD3CF608 , 32'hEEBAFF00 , 32'hF314F860} , 
{32'hFAF9DC48 , 32'h02E89144 , 32'hFBE67438 , 32'hF6E6B430 , 32'h02610300 , 32'h16904A00 , 32'h05984310 , 32'hF17E4CD0 , 32'h164BD5C0 , 32'h050A4DD8 , 32'hF7DA25C0 , 32'hF0CD3CE0 , 32'hF9E6F4A0 , 32'h0199C800 , 32'h0119A280 , 32'hEFE033A0 , 32'h018E306C , 32'h0200F2F0 , 32'h0D318B10 , 32'h06E15C80 , 32'h05710A08 , 32'h0C0A57B0 , 32'hF5C80E70 , 32'h0FEC4760 , 32'h09BDD510 , 32'hFC3D2B4C , 32'hF8B931D0 , 32'h06B98F08 , 32'h04238DA0 , 32'h0B774640 , 32'hFF99E840 , 32'h023B51C4 , 32'h0ACB3FA0 , 32'hFF5C8789 , 32'h0463E8B8 , 32'hFE1F2228 , 32'hFD761B88} , 
{32'hF21F9150 , 32'hFF82D294 , 32'h01566444 , 32'hF7515FF0 , 32'h022B6CE0 , 32'h04D28668 , 32'hF89536A0 , 32'h03BCF004 , 32'h01E54A70 , 32'hFC85E01C , 32'hFEAED0A0 , 32'h041AD688 , 32'hFB5A07B8 , 32'hFA8CB2E0 , 32'hFBF067B8 , 32'h025C638C , 32'hFD699208 , 32'h05C65E70 , 32'h01517154 , 32'hFB8D1C48 , 32'hFCFA427C , 32'hFDE3BB10 , 32'h08093F20 , 32'h0632D418 , 32'h001ACDD2 , 32'hFFC53E40 , 32'hFACD2258 , 32'h04F04618 , 32'hFCFB3CB0 , 32'hF8AF13D8 , 32'hFCE8215C , 32'h06CE1B40 , 32'hF9FACD30 , 32'hFED8B274 , 32'hFDDF7490 , 32'h00F7BA53 , 32'h01DB8C88} , 
{32'hFF1CCC69 , 32'hFFF0C068 , 32'hFEB5ED10 , 32'hFFCCD297 , 32'h0013FB7A , 32'hFEEFE538 , 32'hFF6C47D3 , 32'h020C3ACC , 32'h0046216E , 32'h00D6AC61 , 32'h02051B9C , 32'h0059A8B2 , 32'hFE7093E8 , 32'h008C8F55 , 32'hFF3F93CB , 32'h0065A5F1 , 32'hFFE7EF5D , 32'hFE618B6C , 32'h00797C30 , 32'hFF8ADDB1 , 32'h016AEAE4 , 32'hFFE3F87D , 32'hFF5C8A67 , 32'hFE6FFFB8 , 32'h00A90A3D , 32'hFF7B7F6A , 32'h01FD7270 , 32'hFE4B477C , 32'hFFFBA65C , 32'hFF479F24 , 32'h019A82D0 , 32'h00103743 , 32'hFD7464C8 , 32'hFE565994 , 32'h01865FD8 , 32'hFF96DDAC , 32'hFE518B34} , 
{32'hF2F75CA0 , 32'h0B670A10 , 32'hF632B5E0 , 32'h03CF35D4 , 32'h01315D70 , 32'h1A51F620 , 32'hFDDC83C8 , 32'hF7D24B60 , 32'h0F9DCE50 , 32'h088C4BB0 , 32'h026B9868 , 32'h01BA8C98 , 32'h005821BF , 32'h01E1A9B4 , 32'hFDBAF2D0 , 32'h0BC6E130 , 32'hEF1444E0 , 32'hFFBA2F8D , 32'hF0669040 , 32'hFD0FFF08 , 32'hFB6C61F0 , 32'hF28307D0 , 32'hFC9A1FAC , 32'hFB722660 , 32'hF3D53610 , 32'hFE815818 , 32'hFF0AD270 , 32'hF7CEDF60 , 32'h06C5CCF8 , 32'h02CABDF4 , 32'hFD1BE5B4 , 32'hFD24A7C8 , 32'hFD9CB074 , 32'h02698ABC , 32'h0BDA83C0 , 32'h0307D8AC , 32'hFD9A02C4} , 
{32'h03355CC8 , 32'h07FD15A0 , 32'h065A0238 , 32'h029DF5BC , 32'hF58FEDC0 , 32'hFEC97DE0 , 32'hFBE23780 , 32'hFF54C12A , 32'h009B3474 , 32'hFE1D399C , 32'hFEDCCD9C , 32'hFBA24700 , 32'h02D5C2CC , 32'hFD458790 , 32'hFE183AF4 , 32'hFD7AFB38 , 32'hFFE517B8 , 32'h04662F30 , 32'h00081D67 , 32'hFCD40CFC , 32'hFFC35592 , 32'hFFE35788 , 32'h002B70E0 , 32'hFF11AF8A , 32'hFFFD2D8F , 32'h01BDF088 , 32'hFF85A335 , 32'hFE3A0438 , 32'h03D09384 , 32'hFA2FD8D0 , 32'h00A8B6E6 , 32'h00B1A0B0 , 32'hFF7858DE , 32'h004B0917 , 32'h03AAE488 , 32'h04C891E0 , 32'h00CE691E} , 
{32'h00072812 , 32'hFFFA0B41 , 32'h000283FB , 32'hFFF4076B , 32'hFFF21539 , 32'hFFFC6D50 , 32'h0011CA58 , 32'hFFFD1523 , 32'h0004C6E6 , 32'h0000E7FC , 32'hFFF7517B , 32'hFFFDC9BD , 32'hFFF8BF80 , 32'hFFFCF5C5 , 32'h00000C6E , 32'h0000A73D , 32'h00029D92 , 32'h00051E83 , 32'hFFECB486 , 32'hFFFFC116 , 32'h00019310 , 32'h0007E24E , 32'h00012073 , 32'hFFFFD695 , 32'h0009FBC4 , 32'hFFFBB88A , 32'hFFFA9E93 , 32'hFFF37B2B , 32'h00014401 , 32'h0001CD4D , 32'hFFFFD7D7 , 32'hFFFFE904 , 32'hFFFD18BD , 32'h000245D6 , 32'hFFFD984F , 32'hFFFC434E , 32'h00006410} , 
{32'h0012757D , 32'h000E2BC7 , 32'h0038E2A1 , 32'h00200768 , 32'h0022B8C9 , 32'h001C8D1A , 32'hFFEC80FE , 32'h0007CD51 , 32'h001A308A , 32'hFFED9F4A , 32'h00027E2B , 32'h0012802B , 32'hFFF48ACA , 32'h00422FC4 , 32'hFFF31CCC , 32'hFFD93831 , 32'h002761E6 , 32'hFFBF0095 , 32'h002E7D55 , 32'h001F7599 , 32'hFFE67F0A , 32'hFFC97679 , 32'h00153A83 , 32'h000D84A9 , 32'hFFF402CB , 32'h000295F6 , 32'h001973BD , 32'hFFE9189F , 32'h000E9EF3 , 32'hFFDC2818 , 32'h000F24D5 , 32'h000ABBB8 , 32'h001ED919 , 32'h0027F98B , 32'hFFF08E26 , 32'h00080B81 , 32'hFFDD30C9} , 
{32'h0001CBF8 , 32'h0004FD48 , 32'hFFFA0A99 , 32'h0003D6CD , 32'h0002E377 , 32'hFFFF4194 , 32'hFFFFA89E , 32'hFFFE4BA7 , 32'hFFFA94B1 , 32'h0004A526 , 32'hFFFCC16D , 32'h00039150 , 32'hFFFEDB30 , 32'h0000692A , 32'h0000C920 , 32'hFFFFB444 , 32'h00000925 , 32'hFFFF22B0 , 32'hFFFE8B17 , 32'hFFFBB1CB , 32'hFFFD6816 , 32'hFFFFB934 , 32'h000168A1 , 32'hFFFEEDEA , 32'h0001881C , 32'hFFFC16C0 , 32'hFFFC4033 , 32'hFFFDBD22 , 32'h0001D137 , 32'hFFFFA035 , 32'h00032859 , 32'h0001B2D8 , 32'h0002F9BA , 32'h0005104A , 32'h0001D9F4 , 32'hFFFB551E , 32'hFFFDE8A3} , 
{32'h0000BBE7 , 32'hFFFC0BCA , 32'h00035C95 , 32'hFFFA6292 , 32'h0001DE2F , 32'h00023F52 , 32'hFFFC002F , 32'hFFFF1D84 , 32'hFFFD3163 , 32'hFFFC763C , 32'hFFFC6539 , 32'h0001EACF , 32'h0000A080 , 32'hFFF8F39E , 32'h0004519A , 32'hFFFC47B4 , 32'hFFFD2C6D , 32'hFFFD0049 , 32'h0003C00D , 32'hFFF8633C , 32'hFFFDD49F , 32'hFFFC73AE , 32'h00018B4E , 32'h0002A099 , 32'h0003CC90 , 32'hFFFD267A , 32'h0003C3D0 , 32'hFFFEF879 , 32'hFFFE13AC , 32'h00010890 , 32'h0004D93A , 32'h000564F6 , 32'hFFFF838B , 32'hFFFF7495 , 32'hFFFFCF29 , 32'hFFFCC442 , 32'hFFFF41DC} , 
{32'h0003DEDB , 32'hFFFE30A7 , 32'hFFFF631B , 32'h0000C02F , 32'h000121EA , 32'h00009B16 , 32'hFFFBF2A3 , 32'h00033D91 , 32'h0000EE7A , 32'h0006633C , 32'h00032557 , 32'hFFFD1564 , 32'hFFFD825C , 32'hFFFFA3F8 , 32'hFFFA9801 , 32'h00095597 , 32'h00055E31 , 32'h000361C7 , 32'hFFFF2C2C , 32'h00038467 , 32'hFFFDAC9B , 32'hFFFDF6D4 , 32'hFFFF64BA , 32'hFFF82D48 , 32'h0001C69A , 32'hFFFFA34C , 32'h000096F0 , 32'h00000165 , 32'h0001F5D9 , 32'h000246C6 , 32'h00013BF5 , 32'hFFFCE606 , 32'h00013B62 , 32'hFFFD331A , 32'h0002884D , 32'hFFFAE172 , 32'hFFFD24AF} , 
{32'h000796C8 , 32'h00055B9E , 32'hFFFE76A0 , 32'hFFFB5420 , 32'h00006A0F , 32'h000202DD , 32'hFFFD670D , 32'h000187A1 , 32'hFFF9E3B4 , 32'h00017CBA , 32'hFFFA2A52 , 32'h0003057C , 32'hFFFF740E , 32'h0003EEB4 , 32'hFFFDA9F3 , 32'hFFFA69D9 , 32'h00095E0D , 32'h0006E486 , 32'h00016981 , 32'h0000FFC7 , 32'hFFFFE309 , 32'h00038A04 , 32'hFFFF6B0B , 32'h00004D6E , 32'hFFFF3ABA , 32'h0000018C , 32'h00012433 , 32'hFFFEFA5F , 32'hFFFE502C , 32'h0000C79E , 32'hFFFC7208 , 32'hFFFEA006 , 32'hFFFA7B54 , 32'h0001A3DB , 32'h00003558 , 32'hFFFC190A , 32'hFFFB13D9} , 
{32'hFFFC370E , 32'h00069228 , 32'h000334A0 , 32'h0000C4A4 , 32'hFFFF43F1 , 32'hFFFD2EF2 , 32'h00025E3E , 32'h000313AB , 32'hFFFF4970 , 32'h000043A7 , 32'h00006D81 , 32'hFFFFF84E , 32'h00057346 , 32'h00020511 , 32'hFFFF1F95 , 32'hFFFF4AF5 , 32'hFFFE9222 , 32'h00009DF8 , 32'h00013FE1 , 32'hFFFF3E9A , 32'h00086A75 , 32'hFFFD1D38 , 32'h0000579A , 32'h0003F8A2 , 32'hFFFF8EF6 , 32'h0001815D , 32'h0001E870 , 32'hFFFA3C29 , 32'hFFFF82DF , 32'h0001F92E , 32'hFFF9D59D , 32'hFFFD8D3A , 32'h0002B43E , 32'hFFFD8DF1 , 32'h00048EEC , 32'hFFFDD0F2 , 32'h0000681E} , 
{32'h0005289F , 32'hFFFFD4C6 , 32'hFFFC30D7 , 32'hFFFE0967 , 32'hFFFE65DA , 32'hFFFDBDD9 , 32'hFFFFCB2B , 32'h0004F2D3 , 32'hFFF87364 , 32'hFFFDAFD7 , 32'hFFFCEDAD , 32'h000004A7 , 32'hFFFE0A5F , 32'hFFFE71CB , 32'hFFFF2A01 , 32'hFFFF53F8 , 32'h00019727 , 32'h0003DA66 , 32'hFFFC5A78 , 32'hFFF94019 , 32'h0005C6EA , 32'h0005A2A8 , 32'h0005D224 , 32'h0000E6AD , 32'h0004FDF9 , 32'hFFFF0917 , 32'hFFFE5C87 , 32'hFFFEF2B5 , 32'h000316F3 , 32'h000011F8 , 32'h00007928 , 32'h00006E50 , 32'h000357CB , 32'h0002E81B , 32'h00036FC0 , 32'h0004E0C2 , 32'h00018455} , 
{32'h00058BA6 , 32'h00008E03 , 32'h00009525 , 32'h00032C32 , 32'h0001149A , 32'h0005846B , 32'h0001E06F , 32'hFFF8C5DF , 32'h00026A99 , 32'hFFFDA162 , 32'h00070A1F , 32'hFFFD1F4A , 32'hFFFF3E5F , 32'hFFFEDFE2 , 32'h00030653 , 32'hFFF8A910 , 32'h000348A4 , 32'hFFFEE64D , 32'hFFFF2AB0 , 32'hFFF88647 , 32'h00027AFC , 32'hFFFE358D , 32'hFFFE9E15 , 32'h00020732 , 32'hFFFDF033 , 32'h0000EF41 , 32'hFFFAF498 , 32'h0000F8CD , 32'h00037852 , 32'h00028F17 , 32'h0002A49D , 32'h00051B1E , 32'hFFFDB2CE , 32'h00002182 , 32'h000039A8 , 32'h000142EB , 32'h00032BF6} , 
{32'hFFB21713 , 32'h004131F7 , 32'hFFCC1276 , 32'h002A663D , 32'h00057DC9 , 32'h0028081B , 32'hFFFC4F35 , 32'h00012852 , 32'h0000F202 , 32'h001E0AA6 , 32'hFFE19E62 , 32'hFFE553C2 , 32'hFFF8F58A , 32'hFFE78BAE , 32'hFFEB920C , 32'hFFFD315B , 32'hFFE39EA0 , 32'hFFF9422A , 32'hFFE4C6A9 , 32'hFFFEFEA1 , 32'hFFDD1E6D , 32'h00127A60 , 32'hFFF373BF , 32'h00001030 , 32'hFFFC06CC , 32'hFFE24A17 , 32'hFFF69B1C , 32'hFFF756C6 , 32'h002CCF9A , 32'hFFF13E4D , 32'hFFF955E2 , 32'hFFEC9EB3 , 32'h000BCCC7 , 32'h001D607F , 32'h0000E784 , 32'h00169251 , 32'hFFF00CEF} , 
{32'hF6C4B5A0 , 32'h07348E80 , 32'h02B6F55C , 32'h013742D0 , 32'h04F7CF40 , 32'hF589B550 , 32'h069B3560 , 32'hFE6F9E70 , 32'h0D53B790 , 32'hFE2DF510 , 32'hF5989B50 , 32'h01B4F648 , 32'h06B2C6F8 , 32'h02469754 , 32'h06EE6E70 , 32'h09366000 , 32'h0098B79C , 32'h03B14034 , 32'h00D51774 , 32'hF5AD1910 , 32'hFC7B9344 , 32'hFC3D1F7C , 32'hF702D7B0 , 32'h00A8126E , 32'hFE72D5F8 , 32'hFF36C274 , 32'h0992C6C0 , 32'hFE7B12F0 , 32'hFF2AD304 , 32'h037CCC94 , 32'hFA6A72C0 , 32'h0405CD88 , 32'h0C91A800 , 32'hFD438B6C , 32'h05AEA3B8 , 32'hFD67F5CC , 32'hFE2D78EC} , 
{32'hFFC0FB1D , 32'h009D0584 , 32'hFE8E6E4C , 32'h0162A8C0 , 32'hFFCDBA05 , 32'h0000015E , 32'h00C7BFDA , 32'h00987A12 , 32'h00FCF0EC , 32'hFFA39520 , 32'hFEB8BD98 , 32'hFF064160 , 32'hFE4494D0 , 32'h007DF77A , 32'h012B83AC , 32'h00922D46 , 32'hFE0F4E78 , 32'h0186E628 , 32'h0078FC38 , 32'hFEAE6B5C , 32'hFE6619B4 , 32'hFEA62AF4 , 32'h0037286D , 32'h0025BD96 , 32'hFE4BE200 , 32'hFF3929F8 , 32'hFF1627AA , 32'hFF3E2BEC , 32'h002CC2E8 , 32'h014311C4 , 32'hFFF2E4FA , 32'h01106CF4 , 32'h0096CCC8 , 32'h0090184C , 32'hFF38E371 , 32'hFEADAE18 , 32'h00B487B4} , 
{32'hF575B990 , 32'h05A877A0 , 32'h02FCA900 , 32'h0ACA3BD0 , 32'h004BB8D5 , 32'hF3E0DAA0 , 32'h0ACBC090 , 32'h013AE1D0 , 32'h0277EDE0 , 32'hEE3CCC40 , 32'hEE804E40 , 32'h09597A90 , 32'h116F9EA0 , 32'h06103278 , 32'h0B171AC0 , 32'h0D6828B0 , 32'hFFED8BB0 , 32'h02AC7B50 , 32'hF9FF8738 , 32'hF72161E0 , 32'hF96BDD90 , 32'hFBD51600 , 32'h0108DD5C , 32'h086031D0 , 32'h005C8C8E , 32'h08E6EA00 , 32'h0C1A1400 , 32'hFB73D510 , 32'hFABB2D00 , 32'hFAFE7EA8 , 32'hFE2393BC , 32'h08EDFB20 , 32'h08396C40 , 32'hF51A58B0 , 32'h019ADCA0 , 32'hFCBCDC0C , 32'hF94F5370} , 
{32'hF0DBAB80 , 32'h0AB7B2A0 , 32'h03491BA4 , 32'hFA5874E0 , 32'h00A2B307 , 32'hF29F6C20 , 32'h05B3E390 , 32'h00C8005F , 32'h0F66F8D0 , 32'h002C588F , 32'hE889BA20 , 32'h036823EC , 32'h068CCBE0 , 32'h02E4C4B8 , 32'hFEF10E68 , 32'hF91DD630 , 32'h07EF8810 , 32'hFF21A7E1 , 32'h02105700 , 32'h09422200 , 32'hFD73253C , 32'hFE7AD558 , 32'h03CB91CC , 32'hFF787938 , 32'hF98EE098 , 32'hF912C6A8 , 32'h07641C68 , 32'hED714C00 , 32'h037F9B88 , 32'h0A34DED0 , 32'hF8BD77C0 , 32'hF42843E0 , 32'hFC014DD0 , 32'hFBE62DF8 , 32'hFCEFD7E0 , 32'h0688C0B8 , 32'h020EBEA8} , 
{32'h01E01500 , 32'hFF687E25 , 32'hFCC7AA58 , 32'hFCDDD4F8 , 32'hFF00E231 , 32'h10F04A80 , 32'hFF9FFDEE , 32'hFC83061C , 32'h118C0900 , 32'hFC84E6B8 , 32'h0032B2E9 , 32'h023AB510 , 32'h03B9A110 , 32'h04D640B8 , 32'hFC8AF974 , 32'h04E8F630 , 32'hF88A3E58 , 32'hFD18BF90 , 32'hF7FDAC60 , 32'h069448E8 , 32'h01BD8BB8 , 32'hFBC206F0 , 32'hFF28E0F0 , 32'hFA5A8340 , 32'hFAC3B980 , 32'hFB373E00 , 32'h0119C3D4 , 32'hFCC653F4 , 32'hFDEE0810 , 32'h04D86180 , 32'hF9325588 , 32'hFA05FE00 , 32'hFE1F6F84 , 32'h02C8525C , 32'h0D906BE0 , 32'h06627678 , 32'hFFEA854A} , 
{32'hF6CB4880 , 32'h070DD2C0 , 32'hF8784540 , 32'h014A7490 , 32'hFEA4F0C4 , 32'h14790440 , 32'hFA64F370 , 32'h00AA06D1 , 32'h0A192F70 , 32'h0391B440 , 32'hFE8718D0 , 32'h04F51C40 , 32'hFF7FD219 , 32'h001194A0 , 32'hFD590E40 , 32'h02EF0D00 , 32'hF3337BA0 , 32'hFB56CF88 , 32'hF2678EB0 , 32'hF808D1A8 , 32'hFC178578 , 32'hF5800910 , 32'hF95F0C18 , 32'hF7BD35F0 , 32'hFC281950 , 32'hF7BA7F60 , 32'h00DA4582 , 32'hFF9D0EF6 , 32'h031A5F24 , 32'hFE1AE7DC , 32'hFEF19114 , 32'hFAFBC560 , 32'h007A3778 , 32'h0AFE1A10 , 32'h07D129E8 , 32'h009A6027 , 32'hFC3BAFA4} , 
{32'hF0A348E0 , 32'h14BCEC80 , 32'hF97FA330 , 32'hF457EFD0 , 32'h04280178 , 32'hF3702310 , 32'hFA50D010 , 32'h0AD22160 , 32'h11CF5540 , 32'hF88DE680 , 32'hEE912560 , 32'hFB1395B8 , 32'h07A0EC00 , 32'h056601A8 , 32'h132E9BC0 , 32'h079E7580 , 32'h09A17110 , 32'h01B8EE78 , 32'hFCA7ED1C , 32'hFB063C80 , 32'hFD4C2160 , 32'h019A16F8 , 32'h1412B0C0 , 32'hFDBF8400 , 32'hF937DB70 , 32'h0261C34C , 32'hF3530770 , 32'hF610DAD0 , 32'hF4851660 , 32'h06BAD8E0 , 32'hF65BA9C0 , 32'hFC6B59A0 , 32'h0044D2A1 , 32'h00F6D7FD , 32'hF03CBF00 , 32'h0E29F980 , 32'hFF611E18} , 
{32'hF86C6308 , 32'h0B307DC0 , 32'h0301FBE4 , 32'hF815B8B0 , 32'hFAAB2628 , 32'hDF94DF80 , 32'h0FFBCE90 , 32'h07754390 , 32'h13D65B60 , 32'h1B858B40 , 32'hEDFECB20 , 32'h0C1C75C0 , 32'h16DCDC60 , 32'h221B8080 , 32'h0B0A8000 , 32'h0C577970 , 32'h1E7000A0 , 32'h09CD5630 , 32'hFBC1EEB0 , 32'hFA1A4CC8 , 32'hFCEE891C , 32'h0494F638 , 32'h11C32740 , 32'hDC0B5880 , 32'h07468890 , 32'hE10F9EA0 , 32'h16B27560 , 32'hDB042240 , 32'h091106C0 , 32'hF9BF2C48 , 32'h0DAD93F0 , 32'hFAF122B0 , 32'hEEE38A60 , 32'h04D740D8 , 32'hFB49AFE8 , 32'h0D9C2450 , 32'h036FD1E4} , 
{32'hF60A4850 , 32'h159CB940 , 32'h14E247A0 , 32'h09D512A0 , 32'hFF94B31E , 32'hDD532000 , 32'h1AB9FFE0 , 32'h08BD35D0 , 32'h0573BD70 , 32'h095FA380 , 32'hE9AA0320 , 32'hFF48B3EB , 32'h170A4B00 , 32'h22498AC0 , 32'h03544680 , 32'h00E50F39 , 32'h0B74B4F0 , 32'h0E0864B0 , 32'hFC08B060 , 32'hE4D00800 , 32'hEF8976C0 , 32'h080B2710 , 32'h0AA99950 , 32'hF57AB8C0 , 32'h17345EA0 , 32'hE865CBA0 , 32'h18C20920 , 32'h0F405F90 , 32'hFC9CC2A8 , 32'h10E03C60 , 32'h1DCACB00 , 32'hFC66AD08 , 32'hF0AC6FB0 , 32'hFEDD5BB0 , 32'hE3B318E0 , 32'hF4BFEE70 , 32'h06DC7D40} , 
{32'hECD84C20 , 32'h0905CD40 , 32'h03E8F93C , 32'h01BAA0C0 , 32'h016EB488 , 32'hED6B9DE0 , 32'h0AB1A180 , 32'hFCC1540C , 32'hEF044700 , 32'hFFC9E6D6 , 32'hFF6878D9 , 32'h0067211C , 32'hFF93172E , 32'h12800880 , 32'h06F93B78 , 32'hEF4D9520 , 32'h09DF58B0 , 32'h082C5250 , 32'hFC329378 , 32'hF4659FA0 , 32'hF9FC64E8 , 32'h00541894 , 32'h0D86AA70 , 32'hEC1769E0 , 32'h22A4A200 , 32'hF6252920 , 32'h04213D78 , 32'h140D2180 , 32'hF9AC1E98 , 32'hFE20D138 , 32'h0AA43490 , 32'hEDF75D40 , 32'h0518F288 , 32'h0256E3C8 , 32'hE3F3D4E0 , 32'h05A049D8 , 32'hFCB15C60} , 
{32'hF3466210 , 32'h00A9F5B8 , 32'h05969118 , 32'h0D031660 , 32'hFAD16DC0 , 32'hD942AC80 , 32'h0CDE05C0 , 32'h10025720 , 32'hEB9687C0 , 32'hF017F710 , 32'hF62AF220 , 32'h04140E88 , 32'hF6EE7A60 , 32'h1D4D9700 , 32'hFECDFDA8 , 32'hF221BBB0 , 32'h0D64C670 , 32'h0D404EF0 , 32'h072C3370 , 32'hEA8C5820 , 32'hFD1D93E8 , 32'h01994A78 , 32'h0C6E57E0 , 32'hF722A660 , 32'h22849300 , 32'hEFB67CE0 , 32'hF5BB4B20 , 32'h22828400 , 32'hFDCF328C , 32'h042F20E0 , 32'h16130820 , 32'hEFDFD340 , 32'h05126500 , 32'hFA367218 , 32'hEB549020 , 32'h0E172C60 , 32'h0308BC4C} , 
{32'hDAE49BC0 , 32'h13C90520 , 32'hF5C8B280 , 32'hF65D83D0 , 32'hF700EC90 , 32'hF75C6C50 , 32'h065705A0 , 32'h0D2EB0F0 , 32'h0485DBC0 , 32'h165E8800 , 32'hFD7E01C4 , 32'hFC21BB20 , 32'hEFF76000 , 32'h28082C80 , 32'hFDECD320 , 32'hFE316058 , 32'hEDC4D8E0 , 32'h0DAE5430 , 32'hF9309DE0 , 32'hEDCE60A0 , 32'hF8FE9E60 , 32'h069EDD60 , 32'h02879D04 , 32'hFDE481E8 , 32'h11CA6680 , 32'hF4CADCF0 , 32'hE7388780 , 32'h0E242320 , 32'hFD791B80 , 32'hE95FC700 , 32'h05504738 , 32'hFD1DD81C , 32'h01771EA4 , 32'hFB010A70 , 32'hFA0BFE78 , 32'h190A5500 , 32'h09BE7800} , 
{32'hD855B640 , 32'h1AFAA200 , 32'hEEB9AB60 , 32'h01B3A9B4 , 32'h0093B32B , 32'h0F1FCB70 , 32'h19F00A80 , 32'hF7F98160 , 32'h248DACC0 , 32'h009B63AC , 32'hEB051AE0 , 32'hF5BB1850 , 32'h151C92E0 , 32'h1C4E9FE0 , 32'hFCB00128 , 32'hF0EFDE60 , 32'hF00A4090 , 32'h140E62A0 , 32'hF799DC10 , 32'hFB169F10 , 32'h065808F0 , 32'h17427020 , 32'hF7231C60 , 32'hFAD185F0 , 32'h12591E40 , 32'hFCD91D00 , 32'hFBD6FCD0 , 32'h0A433800 , 32'h10839B80 , 32'h08A0D040 , 32'h1DEE15C0 , 32'h0D2912E0 , 32'h09E8E6E0 , 32'hF17B7F60 , 32'h09F86750 , 32'hF65D0940 , 32'h01961508} , 
{32'hEF3E4C20 , 32'h0C6C91F0 , 32'hE4FB3A20 , 32'hF06A8380 , 32'hF750C100 , 32'h157B7BC0 , 32'hFBAB0018 , 32'hF222D0E0 , 32'h0F35DAD0 , 32'h2AB58600 , 32'hED7A7860 , 32'hDA106480 , 32'hEDAA92C0 , 32'h0CEADD10 , 32'hF5303BA0 , 32'h0F15FE30 , 32'hE612CD20 , 32'h0CFEB970 , 32'h27FF2980 , 32'hFE7281A0 , 32'hFC2B7264 , 32'h31E41C80 , 32'hE6349D80 , 32'h0E5C6750 , 32'h0D4F9130 , 32'h1DAA0EA0 , 32'h12D86740 , 32'h0DEE7230 , 32'h12290AC0 , 32'hE9A13900 , 32'h035481F0 , 32'h058D1760 , 32'hF0CBDCC0 , 32'hFF615295 , 32'hF96BF538 , 32'hFB289FD8 , 32'h0E462910} , 
{32'hE139DEC0 , 32'hFD6C3EEC , 32'hD9AA65C0 , 32'hFA231EE0 , 32'hE9766980 , 32'hF64D5500 , 32'h0B70D5C0 , 32'h0153EB1C , 32'h0035B1A7 , 32'h0A938960 , 32'h09F38C70 , 32'h065D8C70 , 32'h0247C118 , 32'h0F35F460 , 32'h02C12D04 , 32'hF5A6D410 , 32'h0C8BC8B0 , 32'hF3733FB0 , 32'h0FA6F5C0 , 32'h0983A410 , 32'h02F651E8 , 32'h0CA9F670 , 32'hFCA99E0C , 32'hFDB3F818 , 32'h02703694 , 32'h06EFD538 , 32'hFDEAA664 , 32'hEF035060 , 32'h121DE0A0 , 32'hF2ABB5C0 , 32'h104FF100 , 32'h1FD0CF40 , 32'hE9905F20 , 32'h074DC0C8 , 32'h0066BD19 , 32'hFF34C670 , 32'hFAF026A0} , 
{32'hF83BA4B0 , 32'h04722828 , 32'h03C10DCC , 32'hFAD2E1A0 , 32'h0F7C6BF0 , 32'hFDC679BC , 32'hF4D26A90 , 32'h020C56C8 , 32'h0509D330 , 32'h1B4D98E0 , 32'h06D716B0 , 32'hF6951D40 , 32'hF8AAA2B0 , 32'hFE8ECBE4 , 32'hF95BAE68 , 32'hFAD3FDD8 , 32'h06194C00 , 32'h05426DF0 , 32'h0627D520 , 32'hFDAC8798 , 32'hF90CC818 , 32'h04D80080 , 32'hE33D4520 , 32'h021308B8 , 32'hFDC1C58C , 32'h08C25BF0 , 32'hF8482DA8 , 32'hF99FDB78 , 32'hF8C09E40 , 32'h0FDD16D0 , 32'h0987A630 , 32'h0719B0E0 , 32'hF465C380 , 32'h021188F4 , 32'h00259DC3 , 32'h05A95E08 , 32'h096F6F90} , 
{32'hF823BA60 , 32'h07532BB8 , 32'hFBB87780 , 32'hF49B4F60 , 32'h003206ED , 32'hFD8390A8 , 32'hFBEE5BF8 , 32'h0452B788 , 32'h03DEB0C0 , 32'h13668C40 , 32'h0A7901C0 , 32'hF85C1630 , 32'hE80E71C0 , 32'hFE92F3CC , 32'h012AF660 , 32'h02A2A894 , 32'hF4AE5AE0 , 32'h015B3550 , 32'h11C01B60 , 32'hF637D370 , 32'h0DE03B20 , 32'hFCF6F45C , 32'hF0157360 , 32'hFD362000 , 32'h0086A6F9 , 32'hFCFBB978 , 32'hFC669030 , 32'h06D6BB58 , 32'hFCBA6C94 , 32'h0014B8FD , 32'hFAF15110 , 32'hFA96AF68 , 32'hF6D81F60 , 32'hFE026EA0 , 32'h08A528B0 , 32'h0F77CE20 , 32'hFE7E2BC8} , 
{32'h000856B2 , 32'h00515A15 , 32'hFFEBFF95 , 32'h0011A5AC , 32'h001AD2D8 , 32'h000A4AFF , 32'hFFCDD2D4 , 32'h000A2FC3 , 32'h0010002D , 32'hFFFC699E , 32'h00020C3B , 32'h005D6345 , 32'hFF8FA585 , 32'h0070E526 , 32'hFFD650DB , 32'h0003667B , 32'h009C3518 , 32'hFF692B18 , 32'h002ADD42 , 32'h0064FD04 , 32'hFFE00F8A , 32'hFFFB8D21 , 32'h001AE29D , 32'h0031F4EB , 32'h0044F428 , 32'h0076E17B , 32'h00351C24 , 32'hFFB280C5 , 32'h00301DED , 32'hFF98E8FA , 32'h002B8263 , 32'h003FAB1D , 32'h0030C38A , 32'h000A3F4A , 32'hFFE1221E , 32'h00465220 , 32'hFFAC0380} , 
{32'hF4ADF9B0 , 32'h09F4CCA0 , 32'hFDB39A90 , 32'h051444D0 , 32'hFDE48D84 , 32'h0495DA20 , 32'hFCB59784 , 32'hFD0A4174 , 32'hFBB667D0 , 32'hFA3C7B38 , 32'h05167F38 , 32'hFD2F9870 , 32'hFB8FC290 , 32'hF3E35460 , 32'hFA3804E8 , 32'h0362B5EC , 32'hFBCDE640 , 32'h00831D15 , 32'h06D2D228 , 32'hFE801178 , 32'h05047640 , 32'hF8700560 , 32'hFEFE3884 , 32'hFEA0EC58 , 32'h0061215D , 32'h03F0C9C4 , 32'h003EC3A2 , 32'h09B02240 , 32'hFB4095C8 , 32'h026D98DC , 32'h010C1888 , 32'h05700528 , 32'hFC5C0230 , 32'hFB4D8DA8 , 32'h011CCAE4 , 32'h028DCC50 , 32'hFD0BA438} , 
{32'h001DD8CB , 32'hFFEA8982 , 32'h0041E4FB , 32'h004D2CDB , 32'h0029565C , 32'h0029EDD2 , 32'hFFE17326 , 32'hFFF3DC35 , 32'h00070ACC , 32'hFFF80ECA , 32'h00115964 , 32'hFFC45F32 , 32'hFFFE9A70 , 32'h005EB48E , 32'hFFE8DE30 , 32'h00048C36 , 32'h0073F844 , 32'h0006AF5C , 32'h00081B86 , 32'h004244BD , 32'hFF9EAE4F , 32'hFFBB2FA6 , 32'hFF9510E5 , 32'h001931C1 , 32'h000B59E2 , 32'h00117B20 , 32'hFFD922D6 , 32'hFFB9838D , 32'h0003F045 , 32'hFF88F872 , 32'hFFDEB299 , 32'hFFD77053 , 32'hFFF42EEC , 32'h0015EDE2 , 32'hFFC5F6D5 , 32'h003B7D90 , 32'h00293AB2} , 
{32'h000B8F3E , 32'hFFFBF5EC , 32'h0003B328 , 32'hFFFE47AA , 32'h0003BF4E , 32'h0007C9E5 , 32'h00077FBA , 32'hFFE9808F , 32'h00096B99 , 32'hFFFF826A , 32'hFFF1DD7C , 32'hFFF08A5C , 32'hFFEEDF89 , 32'h0001E6FF , 32'hFFF096AB , 32'hFFFE74D7 , 32'h000D9C71 , 32'h0000028F , 32'h0001C6A3 , 32'hFFFEA2C5 , 32'hFFFB24B7 , 32'h00048586 , 32'h00098BCB , 32'h0006F12D , 32'h0000EA14 , 32'hFFF41633 , 32'h000416A9 , 32'hFFF13CC4 , 32'h0002771D , 32'h00002561 , 32'hFFF9485E , 32'hFFFC4699 , 32'h0003844D , 32'h0008FF44 , 32'hFFFDD5BA , 32'hFFFBE7B2 , 32'h0003375E} , 
{32'hFFFF26C9 , 32'hFFFAE0DF , 32'hFFFF0FCE , 32'hFFFF6FD2 , 32'h0005D137 , 32'hFFFF1494 , 32'h00004AD2 , 32'hFFFE3D73 , 32'h0000C2AD , 32'hFFFC1CF4 , 32'hFFFB892D , 32'hFFFE8B2D , 32'hFFFD98F7 , 32'hFFFCB7F8 , 32'h00015C6B , 32'h0003DB58 , 32'hFFFF06AA , 32'hFFFC9F52 , 32'h0005B421 , 32'hFFFE6BAC , 32'h0002C750 , 32'h00062210 , 32'h0004E285 , 32'hFFFA43C4 , 32'h00020F07 , 32'hFFFFBB48 , 32'h0008B159 , 32'hFFFD6E5D , 32'hFFFF0BF3 , 32'hFFFC2B63 , 32'hFFFA024A , 32'h0001E29E , 32'h00019E02 , 32'hFFFF022C , 32'h0001C847 , 32'hFFFD568B , 32'h0002E89F} , 
{32'hFFFCEAF3 , 32'hFFFDEA4A , 32'hFFFFF4BE , 32'h00001C39 , 32'hFFFC2F83 , 32'h000301EA , 32'h0003623A , 32'hFFFE0A42 , 32'hFFFA227E , 32'hFFFCF79A , 32'h0000281F , 32'h00019805 , 32'hFFFD5452 , 32'h00025534 , 32'h0002780E , 32'hFFFD5F28 , 32'hFFFAD98D , 32'hFFFEA8C3 , 32'hFFFB3F8C , 32'hFFFF8F41 , 32'h000276AA , 32'hFFF9C8F7 , 32'h00039FE9 , 32'hFFFCA1F9 , 32'h00074A47 , 32'hFFFF20BA , 32'hFFFC0222 , 32'hFFFFCBB5 , 32'hFFFC7FA4 , 32'hFFFDAFCB , 32'h00013507 , 32'h0000B51D , 32'hFFFE5DA8 , 32'hFFF9B7F9 , 32'hFFFA193E , 32'h00033F50 , 32'hFFFC4580} , 
{32'h00026F8D , 32'h0002C41F , 32'h0002A7BB , 32'hFFFF7907 , 32'hFFFB704F , 32'hFFFD9459 , 32'hFFFD65DB , 32'hFFFE2A46 , 32'hFFFCD9CA , 32'h0000B8F8 , 32'hFFFEAC6D , 32'hFFFFA98B , 32'h00054047 , 32'hFFFE8614 , 32'h0006FD95 , 32'hFFFFD56D , 32'h00004897 , 32'h0007A5FE , 32'h00048F42 , 32'hFFFCE7DE , 32'hFFFA2C1F , 32'hFFFDB596 , 32'hFFFFE5A0 , 32'h00010D7A , 32'hFFFFB17C , 32'h000188FF , 32'h0000AB5D , 32'h0002D8F1 , 32'hFFFE01F2 , 32'hFFFEBA84 , 32'hFFFEC422 , 32'hFFFD1A77 , 32'hFFFE0BFB , 32'h0003378F , 32'hFFFEC8B6 , 32'h0004D292 , 32'h00001525} , 
{32'hFFFFA548 , 32'hFFF89DE9 , 32'hFFFBC167 , 32'h0002FFAF , 32'h00008975 , 32'hFFFE4481 , 32'hFFF8CCA5 , 32'hFFFE3582 , 32'h0004062D , 32'h000037BD , 32'h0002D71E , 32'h0003DEEE , 32'hFFFDFC17 , 32'h0004A067 , 32'hFFFB9E9A , 32'hFFFEF6E6 , 32'h0001DABF , 32'h00037FDB , 32'h0002B361 , 32'hFFFB73B1 , 32'h00042D51 , 32'hFFFD837F , 32'h0002F417 , 32'h0000FA24 , 32'h00012DF5 , 32'hFFFD0695 , 32'h0002DF8D , 32'hFFFF546B , 32'hFFFB2615 , 32'h000A02AE , 32'h00000573 , 32'h000169FC , 32'hFFFCCA0C , 32'hFFFDCCEF , 32'hFFFF6568 , 32'hFFFD69EA , 32'h0003A7FF} , 
{32'hFFFE27E3 , 32'h0000664F , 32'hFFFD22D0 , 32'hFFFFAC56 , 32'hFFFB0AF4 , 32'hFFFC7F90 , 32'hFFFC852D , 32'hFFFEB01B , 32'hFFFFD451 , 32'hFFFC277E , 32'hFFFABD76 , 32'h0000D5EF , 32'h0004118C , 32'hFFF9F96E , 32'hFFFDD6AC , 32'hFFFDE07D , 32'hFFFF14DC , 32'hFFFC6B5E , 32'h0001D933 , 32'h0000CC8B , 32'hFFFFF2FC , 32'h0002C0E2 , 32'h000312BA , 32'hFFF660F4 , 32'h0002CA5D , 32'h0000B5A1 , 32'hFFFCA238 , 32'hFFFF2AA5 , 32'h00009288 , 32'h00009634 , 32'h00017D67 , 32'h000071EE , 32'hFFF96650 , 32'hFFFE6D32 , 32'hFFFFD561 , 32'hFFF9C4A3 , 32'h000142D9} , 
{32'h00033238 , 32'hFFFC6D1B , 32'hFFFAA85B , 32'h0000B730 , 32'hFFFB3F19 , 32'h0002282F , 32'hFFFC55CC , 32'h0000B03E , 32'h0001C4EF , 32'hFFFDC173 , 32'h0005632D , 32'hFFFD031F , 32'hFFFD2380 , 32'hFFFE856A , 32'hFFFBB69E , 32'hFFFBFC6A , 32'h00025A84 , 32'h0001FD3C , 32'hFFFF752F , 32'hFFFE20C7 , 32'h00020C18 , 32'h00000B0C , 32'hFFFFD051 , 32'hFFFEFC6D , 32'hFFFBD05F , 32'hFFFB78A9 , 32'hFFFC9C80 , 32'hFFFECAED , 32'h0001D326 , 32'hFFFAEFBF , 32'hFFFEF02C , 32'hFFFE26A0 , 32'hFFFEC64A , 32'h00016DDD , 32'h00002915 , 32'h00052EDF , 32'h000593E9} , 
{32'hFFFA17AF , 32'h0012A1E6 , 32'h00038F7C , 32'h0004EC05 , 32'h0000C857 , 32'h000D979F , 32'hFFFBEBDB , 32'h00003C3A , 32'hFFFE04C2 , 32'h00000E60 , 32'h0006C493 , 32'h0007DD0A , 32'hFFFDA78B , 32'hFFFD9F01 , 32'hFFFAF7C6 , 32'h0002D3B8 , 32'h0002CEF8 , 32'hFFFFADF6 , 32'hFFF5C21F , 32'hFFFAD2F8 , 32'h0000C711 , 32'h0005759D , 32'hFFFEDE31 , 32'hFFFC07D0 , 32'hFFF87908 , 32'hFFFE3C26 , 32'hFFFD2AC1 , 32'h0001A9F8 , 32'h0001F6E2 , 32'hFFF9A622 , 32'hFFFBAF2D , 32'h00011C9A , 32'h00045AB5 , 32'h000781E3 , 32'hFFFC36CB , 32'hFFF60E04 , 32'hFFF9AED5} , 
{32'hF7305210 , 32'h06BE9D90 , 32'h02F84F70 , 32'h00F49016 , 32'h04C74330 , 32'hF5C70AF0 , 32'h06478228 , 32'hFEAC2DAC , 32'h0CA321A0 , 32'hFE5C7D74 , 32'hF5FD2180 , 32'h01C9EA18 , 32'h069176E8 , 32'h022265F4 , 32'h06933868 , 32'h088BA300 , 32'h0133F86C , 32'h032D35EC , 32'h00C7E0D4 , 32'hF66AEAA0 , 32'hFD007EB8 , 32'hFCBF81E8 , 32'hF70C49C0 , 32'h009FC43E , 32'hFEDDC1F8 , 32'hFF2727FF , 32'h0951C4D0 , 32'hFEB02340 , 32'hFF31BDE7 , 32'h03068790 , 32'hFA912C58 , 32'h03CD43A4 , 32'h0C1C26A0 , 32'hFD1D6328 , 32'h05B006D8 , 32'hFDAFA96C , 32'hFDEE3494} , 
{32'hF5DE2190 , 32'h047B0790 , 32'h04FA0828 , 32'h01965AF4 , 32'h06CD4A00 , 32'hFB0A3758 , 32'h0216C8E4 , 32'hFFEC8E97 , 32'h0B65BB50 , 32'hFFD0E141 , 32'hF398FDF0 , 32'hFB455C08 , 32'h04970070 , 32'h02D75BDC , 32'h081F3520 , 32'h08ECE660 , 32'h052A0948 , 32'hFF981AD4 , 32'h01D5C448 , 32'hF6472600 , 32'h06B3B190 , 32'hFD59BA10 , 32'hFAA534A8 , 32'h01CC9468 , 32'h02269E8C , 32'hFE790030 , 32'h01E10494 , 32'h00024DE8 , 32'hFDC750B0 , 32'hFF58BA7D , 32'hFE8284EC , 32'h06C35E20 , 32'h0A709800 , 32'h05B54B98 , 32'h05E3A028 , 32'hFE1525E8 , 32'h042C9A10} , 
{32'hF371DD80 , 32'h030C7F50 , 32'hF7680A50 , 32'hFF2B6EF7 , 32'h0C5C7230 , 32'h193BA480 , 32'h0B61B570 , 32'hF40B5760 , 32'h30DD2C80 , 32'hFCA032EC , 32'hF3C12FA0 , 32'h04009330 , 32'h0C52D270 , 32'h11F82620 , 32'h024FE418 , 32'h13904BA0 , 32'hEF728CE0 , 32'h05F84FB8 , 32'hF5A0C820 , 32'hF7BFF930 , 32'h0151D11C , 32'hF59A2630 , 32'hF16998E0 , 32'hFE9B7374 , 32'hFE8ADC5C , 32'h074F0978 , 32'h07720D98 , 32'h03C916AC , 32'hFF501D18 , 32'h0D9581D0 , 32'h00B6B6BC , 32'h00A1193C , 32'h0CD055B0 , 32'hF841D778 , 32'h0B8547C0 , 32'hFBE8E4F0 , 32'hF8DB8590} , 
{32'hFF5FDCFA , 32'h083F7D40 , 32'hF57D9D90 , 32'hFA192E58 , 32'hFD764E78 , 32'h30A3E500 , 32'h09D05CD0 , 32'hEBF40140 , 32'h2A8CBFC0 , 32'hF0B0F730 , 32'hF538A3B0 , 32'h00238FC9 , 32'h02A304C8 , 32'h07517F60 , 32'hFF88FCF3 , 32'hFD7828F8 , 32'hEB9BC9E0 , 32'hFE9EA284 , 32'hFC3BD56C , 32'h076AF340 , 32'h076896C0 , 32'hF8744A60 , 32'hF9309C78 , 32'h032E4C00 , 32'hFB4FE260 , 32'h104C5680 , 32'hFD76F2C4 , 32'h032D316C , 32'h02F2D378 , 32'h0A8FB3A0 , 32'h054709F0 , 32'h00438562 , 32'h03255C10 , 32'h06A03798 , 32'h0AA19CE0 , 32'h08140DC0 , 32'h08251E70} , 
{32'hFF0C1D13 , 32'h15C0F280 , 32'hF8BB0940 , 32'hF8D4C988 , 32'hF2249C30 , 32'h2925D040 , 32'h18A88360 , 32'hFB620D80 , 32'h3F175F80 , 32'hE6B884C0 , 32'h01CEEA08 , 32'h09D25300 , 32'h0E076860 , 32'h0A4C81D0 , 32'h0D777D00 , 32'h194661E0 , 32'h015638C4 , 32'h0E91C370 , 32'hFE4A3444 , 32'h17A64F80 , 32'h0294B258 , 32'h10F6C9C0 , 32'hF42A1EF0 , 32'h0E6CC5E0 , 32'hF450B9A0 , 32'h019000A0 , 32'h079E5BC8 , 32'h00D916E0 , 32'h0228E938 , 32'hFE52B5AC , 32'h0ACB5870 , 32'hEE4FA240 , 32'h142381E0 , 32'hF9E6F8F0 , 32'h0D50C630 , 32'h02E30F34 , 32'hF827A5C8} , 
{32'hE3DC9E40 , 32'h2A800240 , 32'hFE53E954 , 32'hE112D2C0 , 32'hF2743AE0 , 32'h027E7120 , 32'h0736E7E8 , 32'h03172BD0 , 32'hFBF87140 , 32'h0E780DA0 , 32'hE5896800 , 32'h03CE5E20 , 32'h1DA67F60 , 32'h0BFB9FB0 , 32'h03341724 , 32'h103A4E80 , 32'h02860B98 , 32'hED46F060 , 32'hF06C3440 , 32'h0F2B4310 , 32'h05898908 , 32'hF6B87890 , 32'hF1061540 , 32'h0A02FFD0 , 32'h0BD12930 , 32'hDCA28C80 , 32'h0F7FD430 , 32'hDF37CFC0 , 32'h07E60298 , 32'h1F9250A0 , 32'hFF6BD0D4 , 32'hEDE171E0 , 32'hE7CAD640 , 32'hF33B6970 , 32'hE14596E0 , 32'h0F6FDF00 , 32'h0B13D430} , 
{32'hFF6D336B , 32'h12895B20 , 32'h05D381C0 , 32'hEF5CC900 , 32'hFC4E6690 , 32'hFC9C58A8 , 32'h00628F79 , 32'h0748F1D0 , 32'h06500588 , 32'hFCFBD5FC , 32'hE69C2F80 , 32'h01B38804 , 32'h09F40450 , 32'h095B0AA0 , 32'h0C316360 , 32'h155B9FE0 , 32'h002D6439 , 32'hE8883A40 , 32'hF0E7EB30 , 32'h0EAFBA90 , 32'hFD3FBB38 , 32'hF0FA4C20 , 32'hF1FC0B10 , 32'h03D6D050 , 32'hFA5E35A8 , 32'hFFD012CB , 32'h0C7A7660 , 32'hF0567ED0 , 32'hFBD823B0 , 32'h13CCF4A0 , 32'hFEF24410 , 32'hF0E71C00 , 32'hE9DCDF60 , 32'hF2B89170 , 32'hE67165A0 , 32'h104DC120 , 32'h0BB768F0} , 
{32'hF2EAE0A0 , 32'h2055F9C0 , 32'h064D68D8 , 32'hEA6F71C0 , 32'h08717B00 , 32'hE5D92BA0 , 32'hFF188B4B , 32'h0A541DB0 , 32'hF1A9AEF0 , 32'h0840A390 , 32'hEF611520 , 32'h102EA580 , 32'h05327638 , 32'hF8CBDF58 , 32'hF87B2EB0 , 32'hEBCF0880 , 32'h0115DA78 , 32'hF60AAFA0 , 32'h0673F2F8 , 32'h0C54C9D0 , 32'h039983E4 , 32'h020F2F94 , 32'h095D10C0 , 32'hF24BA640 , 32'hF227D930 , 32'hF74CDA80 , 32'h1B3A46C0 , 32'hED4170C0 , 32'hFECBC190 , 32'h073509D8 , 32'hE27458E0 , 32'hEE0F8BC0 , 32'hE86FE120 , 32'hFBBF73D8 , 32'hFBAFCCF8 , 32'h06378CF0 , 32'h05BFA328} , 
{32'hF33FD900 , 32'h190634A0 , 32'h11CAFFE0 , 32'hFA4AC628 , 32'hF42706E0 , 32'hDB6C99C0 , 32'hFFE13C4D , 32'h0F784650 , 32'hF22F79F0 , 32'hFA5A9D68 , 32'hEFDB3380 , 32'hFD503EBC , 32'h0818A550 , 32'hF86B2DE8 , 32'hFA2378B8 , 32'hE8FE2E20 , 32'h10EE1CA0 , 32'h061EB9A0 , 32'h0ED858B0 , 32'h060F2338 , 32'hF9F2D858 , 32'h0A23F7A0 , 32'h015ABB04 , 32'hF8BAB268 , 32'h00D7F143 , 32'hFCBFD9A8 , 32'h06C7C518 , 32'hFEF1D620 , 32'h0B4F7E00 , 32'h006BE417 , 32'h05A03DC0 , 32'hEF383EC0 , 32'hF37733F0 , 32'h09DF5B50 , 32'hEE296900 , 32'h00A6F510 , 32'h09C37420} , 
{32'hE95D0E80 , 32'h1EBE7180 , 32'hFA3FF5C0 , 32'hF4E57840 , 32'hF52C6550 , 32'hD8EE0640 , 32'h0B3E3950 , 32'h1AFF9720 , 32'hD92D4400 , 32'h02A12CA0 , 32'hED3FC640 , 32'h03C23E30 , 32'h03368528 , 32'h06A83938 , 32'hF6CF7EE0 , 32'hDF1A6080 , 32'h0D432B10 , 32'hFCA0CD44 , 32'h0F04EA30 , 32'h128C9BA0 , 32'h05EFE160 , 32'h214D4180 , 32'h1185A860 , 32'h0B689870 , 32'hFAF09130 , 32'h05E173F8 , 32'h09C4BA90 , 32'hFC7A6554 , 32'hF581A480 , 32'h0458EC60 , 32'h0A8D3A80 , 32'hFA016C50 , 32'h042B4050 , 32'h0BB53610 , 32'hF465E4B0 , 32'h00206335 , 32'hFA6A9BC0} , 
{32'hD4D40D80 , 32'h285A5AC0 , 32'hF92704C0 , 32'hF9B3A3F0 , 32'hFCB9FCF4 , 32'hE71F6520 , 32'h0C4CBDD0 , 32'hFCB0DA38 , 32'hD529F400 , 32'h0AFB4380 , 32'hE503DFC0 , 32'hF1A02390 , 32'h13E56A80 , 32'h17F45E40 , 32'hF4DD8F30 , 32'hECC16D40 , 32'h12FE1E40 , 32'h0835B840 , 32'h13434020 , 32'h1E37C140 , 32'hF61FD2C0 , 32'h1F24D1C0 , 32'h22492A80 , 32'h0368831C , 32'hE7F25540 , 32'h031272E4 , 32'hFD0015EC , 32'hE217FFE0 , 32'h0D973C00 , 32'h0796A458 , 32'h01950068 , 32'hFCC3579C , 32'hF5788790 , 32'hF2CD3E60 , 32'hFC115B4C , 32'hF3B51850 , 32'h1452E040} , 
{32'hE5FA2BE0 , 32'h0B374310 , 32'h02C8E944 , 32'hFC4777EC , 32'h0358723C , 32'h0E740CA0 , 32'h0FF709C0 , 32'hE9989C20 , 32'h1377B080 , 32'hF24EEB30 , 32'hE3B663C0 , 32'hF23E81D0 , 32'h0EADA6C0 , 32'h12D4C340 , 32'hF27998D0 , 32'hE466AC00 , 32'h0BEDAF80 , 32'h08C163F0 , 32'h0D3CDB50 , 32'h25B5A040 , 32'h0A4C3AD0 , 32'h12D22240 , 32'h051679E0 , 32'h046B8D00 , 32'h056351A0 , 32'h09E762A0 , 32'hF9466960 , 32'hFDC0D6E4 , 32'h09DF3D50 , 32'h0E179E70 , 32'h0E190DC0 , 32'hFA7F6B68 , 32'hF3511AE0 , 32'hEFBFE420 , 32'hF23B6320 , 32'h088D57C0 , 32'h0268D29C} , 
{32'hEC484700 , 32'h1856FA40 , 32'h0390E298 , 32'hF49B34A0 , 32'hF9368770 , 32'h10D78CE0 , 32'h04D0D4D8 , 32'hF6F4D900 , 32'hFE30C028 , 32'h00180119 , 32'hF5ED4510 , 32'hF2FFE200 , 32'h12A0F000 , 32'h09348AC0 , 32'hF7EFD8A0 , 32'hF264C4E0 , 32'hFB874C18 , 32'h12845340 , 32'h0DBFFF00 , 32'h22ECEDC0 , 32'h01391808 , 32'h0B903670 , 32'hFED1289C , 32'h0A5224E0 , 32'hFB340CF0 , 32'h08949600 , 32'hF2671BA0 , 32'h0DD383A0 , 32'hF95C4F48 , 32'hF992D870 , 32'hFC9341A8 , 32'h0BDFDCC0 , 32'h0A01F990 , 32'hFE564F08 , 32'hFA6052E0 , 32'h0720F638 , 32'hFF3E64CC} , 
{32'hD2D55A00 , 32'h334F2040 , 32'hEEE5E8E0 , 32'hF88E3ED0 , 32'h0377B628 , 32'h1B762740 , 32'h09BE2710 , 32'hEE102640 , 32'hE5B80220 , 32'h15B19520 , 32'hF6DF2EA0 , 32'hEDF9E000 , 32'hF470D060 , 32'hF62E3AC0 , 32'hE3159AC0 , 32'hFFFD03F0 , 32'hEC61CD40 , 32'h05789688 , 32'h116AE440 , 32'h12416900 , 32'hF92FCB10 , 32'hF1EDF600 , 32'h014D8340 , 32'hFE636418 , 32'hEAB2E5C0 , 32'hF0BB3F50 , 32'h05B02FA0 , 32'h0CA28DA0 , 32'hF775FF40 , 32'hFE545828 , 32'hF0143F60 , 32'h02E73B68 , 32'h12FE13E0 , 32'h0AC06E60 , 32'h126C23E0 , 32'hFD6F0274 , 32'hFBA9AB48} , 
{32'hF9124B60 , 32'h1617B760 , 32'hFC279B04 , 32'hEAEC7D20 , 32'h0623FF98 , 32'h0C089620 , 32'h01C56654 , 32'hF6FE1DC0 , 32'hFB45B470 , 32'h212ABF00 , 32'h08928BC0 , 32'hE7555460 , 32'hFE7D9EC8 , 32'hFDECB358 , 32'hFC4F5A68 , 32'h088A0680 , 32'hEE5550C0 , 32'h01A61A60 , 32'h1F504F80 , 32'h0DB0FCA0 , 32'hF2FFFB20 , 32'h18EC7D20 , 32'hFB8BFC78 , 32'hF4EB62C0 , 32'h064744B8 , 32'h03B885DC , 32'h0BB5D750 , 32'h068C5380 , 32'hFE8AC6D8 , 32'hF309E410 , 32'h060CD0D0 , 32'h16B904A0 , 32'hF8985B58 , 32'h005CD0C7 , 32'h04C5F110 , 32'hFE747D78 , 32'hF406C2F0} , 
{32'hEED618E0 , 32'h190927C0 , 32'hF3E730D0 , 32'hE8C2A260 , 32'h072416A0 , 32'h1838C260 , 32'hFD1F9FF8 , 32'hF87347E0 , 32'h0C622720 , 32'h2CDC2D80 , 32'h1034D100 , 32'hEE8BD720 , 32'hF2960220 , 32'hE6E03720 , 32'hFE6AE378 , 32'h0DA57040 , 32'hED067440 , 32'h07B53AA0 , 32'h1F9F83C0 , 32'h0A0C41E0 , 32'h0F4FE470 , 32'hFF1AC02F , 32'hF5200CD0 , 32'hF27EB460 , 32'hF0418050 , 32'h1A07F360 , 32'h0C9AAB70 , 32'h136010E0 , 32'hF10CA090 , 32'h08307140 , 32'hEFFFD5E0 , 32'hFA9E2790 , 32'hF4817B70 , 32'hF8DE2C68 , 32'h08E69470 , 32'h063672D8 , 32'hFA423B50} , 
{32'h063CFF50 , 32'h0A95F240 , 32'hFC22D4A0 , 32'hE71C2280 , 32'hFCB12EE8 , 32'hFD141520 , 32'h06BF7118 , 32'hFBF34A80 , 32'hFE410AF8 , 32'hFEEFCAC4 , 32'hFAE370E0 , 32'hFBEB8770 , 32'hFB0387E8 , 32'hFE83C860 , 32'h01297DAC , 32'hFF575922 , 32'hF7876D30 , 32'hF8802100 , 32'h0D566300 , 32'hFAE511D8 , 32'h007BDE96 , 32'hF871E918 , 32'h123DE1C0 , 32'hFF7C6AB0 , 32'hF8665CE0 , 32'h0CFD9FE0 , 32'h0BD60D80 , 32'h0119A9EC , 32'hF8D03230 , 32'h0329DECC , 32'h07B5F1A8 , 32'hF9DE72B8 , 32'h0FC71B30 , 32'h07943E98 , 32'hF57047D0 , 32'h119C1E80 , 32'h00FE28E5} , 
{32'h0381BCD4 , 32'h01F2BD58 , 32'h09349CB0 , 32'hF89C22E8 , 32'hFCEC9A88 , 32'hE55707A0 , 32'hFA2D4BF0 , 32'h0D54FCE0 , 32'hF3072C90 , 32'h11F75220 , 32'h130A3560 , 32'hFE8D9188 , 32'hF43997A0 , 32'h0EF6EC30 , 32'h0E2BF940 , 32'h0E19DAE0 , 32'hEB0CA160 , 32'hFC4BA508 , 32'h07282C48 , 32'hF2CCCF20 , 32'hFC0A0060 , 32'hF156FEE0 , 32'h05E9CD30 , 32'hF6533240 , 32'hF6E3E990 , 32'h0318A94C , 32'h0357DCA8 , 32'h02162720 , 32'hFAF1AE98 , 32'hF686E570 , 32'hFEE72B98 , 32'hF141EE50 , 32'hF991ADD8 , 32'h02450130 , 32'hF76797A0 , 32'h296817C0 , 32'h067AD688} , 
{32'h05CC89D8 , 32'hFE072868 , 32'hFD3CE350 , 32'hFE3435A4 , 32'hF9C48F48 , 32'hE2EBC360 , 32'h008414FA , 32'h13EA9880 , 32'hEE956480 , 32'h0E3D7430 , 32'h134DBD20 , 32'h11556780 , 32'hF99919C8 , 32'h0A363F40 , 32'h0AE573F0 , 32'h0E10EB80 , 32'hEAFAE0A0 , 32'h074C6510 , 32'hFCB10978 , 32'hF4661D60 , 32'hF16AA890 , 32'hF73E06F0 , 32'hFA770C08 , 32'hF402C000 , 32'hF9BFF698 , 32'h053ECC88 , 32'h00198995 , 32'hFFCF4041 , 32'hF7A6F6F0 , 32'hFB103EF8 , 32'hF5838F10 , 32'hF57427D0 , 32'hF8FD7708 , 32'hF6F2A3D0 , 32'hFCAF5E1C , 32'h15898820 , 32'hF8695850} , 
{32'h004B8B56 , 32'hFF93AA0D , 32'h006DB80F , 32'h0087A3DE , 32'hFFCF1FB9 , 32'hFFFCE706 , 32'hFFEB7294 , 32'h005C8AF4 , 32'h003AF75C , 32'h004A4B2D , 32'hFFF231EB , 32'hFFFA1B36 , 32'h00576093 , 32'h001D83A0 , 32'hFFEBE0A7 , 32'h008111A5 , 32'h000AF69F , 32'h005EFAFC , 32'hFFF17696 , 32'hFFDC212A , 32'h00019D53 , 32'h0040F1A3 , 32'hFF99B206 , 32'hFFB295BE , 32'hFFADB687 , 32'hFFF021B7 , 32'hFF4B15E1 , 32'h004BE8A8 , 32'h001ACB65 , 32'hFFB2A469 , 32'hFF6FB481 , 32'hFF16F2A6 , 32'hFFD9D4FC , 32'h001C28E1 , 32'hFFC0614F , 32'hFFB0E597 , 32'h00937CD7} , 
{32'h00479550 , 32'hFF8D4C27 , 32'h0097B05B , 32'h00A67F19 , 32'hFFB08741 , 32'hFFFE1335 , 32'hFFF11178 , 32'h00777FA5 , 32'h0044041B , 32'h006B39F5 , 32'hFFFB4A8A , 32'h00051AFF , 32'h007673CF , 32'h00225693 , 32'hFFF45F14 , 32'h00A4781F , 32'h0012D976 , 32'h00825011 , 32'hFFFCA2FC , 32'hFFBCA99C , 32'h0008044A , 32'h0050D538 , 32'hFFA1850D , 32'hFFB76C7B , 32'hFF744B71 , 32'hFFC7EE18 , 32'hFF39AEAB , 32'h009E2E56 , 32'h0015FAD8 , 32'hFFC522B0 , 32'hFF59E749 , 32'hFF0FCD1A , 32'hFFC44A5D , 32'h0027DA03 , 32'hFFC0398D , 32'hFF9C6063 , 32'h00ADA193} , 
{32'h0044F71B , 32'hFFC4690C , 32'h00552FAE , 32'h003F3011 , 32'hFFC3833F , 32'hFFF3F919 , 32'h000C9098 , 32'h004F9805 , 32'h0034FFC6 , 32'h0037960C , 32'hFFC5449D , 32'h0005C453 , 32'h0020AA17 , 32'hFFF6EB5E , 32'hFFF74747 , 32'h0041A6F1 , 32'hFFC5B3AD , 32'h00311457 , 32'h0012FE23 , 32'hFFAF79F1 , 32'h00243B63 , 32'h002F3451 , 32'h0005B5B1 , 32'hFFBEC99E , 32'hFFB4CEB9 , 32'hFFF1D130 , 32'hFFA10F49 , 32'h00451B6E , 32'h0019889A , 32'h00008547 , 32'hFF995FBE , 32'hFF5AF582 , 32'hFFFF6362 , 32'h00449E1A , 32'hFFE24357 , 32'hFF9BA02E , 32'h003AA6E3} , 
{32'h000397DF , 32'hFFFEDBCB , 32'h000072BF , 32'h0004E45B , 32'h00068943 , 32'hFFFFEADA , 32'hFFFE0F52 , 32'h00007B6C , 32'hFFFB0908 , 32'hFFFD0C53 , 32'hFFFEE07C , 32'hFFFE609E , 32'h00058104 , 32'h0004E539 , 32'hFFFF0FD3 , 32'h0000D91A , 32'hFFFB5BE4 , 32'h00066EFE , 32'h0000DCE5 , 32'hFFFC14C2 , 32'h0000AAC0 , 32'h00033062 , 32'h00030B17 , 32'h000138DB , 32'h00031579 , 32'hFFFE5044 , 32'h00017749 , 32'hFFFF77B8 , 32'hFFF8A827 , 32'h0000726B , 32'h00029A40 , 32'hFFFDEF8E , 32'hFFFE658C , 32'h0000C3B3 , 32'h0004D731 , 32'h0004A43C , 32'hFFFBF7C2} , 
{32'hFFFC20D1 , 32'h0000C406 , 32'h000759EA , 32'h000268FB , 32'hFFFE75F0 , 32'hFFFB9108 , 32'h00039B75 , 32'h0000265D , 32'h00008037 , 32'hFFFAEDEA , 32'hFFFBC763 , 32'hFFFCB5C6 , 32'h0000B335 , 32'hFFFF455B , 32'hFFFB8DA4 , 32'hFFFDAF04 , 32'hFFF89715 , 32'hFFFF47F6 , 32'hFFFDF23F , 32'hFFFA0ABF , 32'h00008B01 , 32'hFFFE1874 , 32'hFFFF46BC , 32'h00010A28 , 32'hFFFF62F0 , 32'hFFFDCB11 , 32'hFFFE0009 , 32'hFFFEE077 , 32'h0006C25A , 32'hFFFFD8C6 , 32'hFFFFB74B , 32'hFFFBBC39 , 32'hFFFC452C , 32'hFFFE6BCB , 32'h00031A74 , 32'hFFFE6C0A , 32'hFFFD000D} , 
{32'hFFFC461A , 32'hFFFD4AAC , 32'hFFFEECFC , 32'hFFFE565C , 32'hFFFE13BC , 32'hFFFCAE72 , 32'hFFFCA1BD , 32'h00053DA7 , 32'hFFFC55E8 , 32'h00006EF2 , 32'h00059BDF , 32'hFFFAAEBC , 32'h00009DFA , 32'hFFFF6FB3 , 32'h000300F0 , 32'h000065C0 , 32'h00069318 , 32'h0000D144 , 32'h0005A549 , 32'hFFF74496 , 32'h0005FA81 , 32'h0003B045 , 32'hFFFB9608 , 32'hFFFD48C7 , 32'h0000EB5C , 32'hFFF9BF51 , 32'hFFFD1097 , 32'h0007D228 , 32'h0003C217 , 32'h00016312 , 32'hFFFE292D , 32'h0001496E , 32'h0002F4C8 , 32'h00059AED , 32'h00031F91 , 32'hFFFB493A , 32'hFFFFF6A9} , 
{32'hFFFDD6E7 , 32'hFFFE20E4 , 32'hFFFC81BB , 32'hFFFC6344 , 32'h0004F4AC , 32'h000351F0 , 32'hFFFF8115 , 32'h00033EEA , 32'hFFFE1AB7 , 32'hFFFFC923 , 32'hFFFCFAAA , 32'h0007B785 , 32'hFFFE3BF1 , 32'hFFFDED05 , 32'hFFFA951D , 32'hFFFF0D37 , 32'hFFFFFD1D , 32'hFFFB26D0 , 32'h000250A9 , 32'hFFFE37C1 , 32'h0003F179 , 32'h000648B8 , 32'hFFFEAF04 , 32'hFFFF633C , 32'h00022762 , 32'h00018C8B , 32'hFFFF5828 , 32'hFFFD64EE , 32'hFFFEA147 , 32'hFFFC3DEB , 32'h0002AEE2 , 32'h0001EC61 , 32'hFFFF03BC , 32'hFFFE723A , 32'h0001237D , 32'h00013B78 , 32'h000146D9} , 
{32'h0000D612 , 32'h000056DF , 32'hFFFCE6C5 , 32'hFFFF8D0D , 32'hFFFD5013 , 32'h000454D9 , 32'hFFFEC259 , 32'hFFFE9A7E , 32'hFFFF38F9 , 32'h00001A63 , 32'hFFFF5491 , 32'h00024D94 , 32'h00016D7F , 32'hFFFDF82B , 32'hFFFCEB80 , 32'hFFFDC697 , 32'hFFFDADC7 , 32'h00044512 , 32'hFFFF7A49 , 32'hFFFF4373 , 32'h0001DD5E , 32'h0001300B , 32'hFFFF1925 , 32'h0001AB21 , 32'h0000F8A5 , 32'h0002FECA , 32'h0002CBE3 , 32'hFFFF9F13 , 32'h0003A6CB , 32'h000135BF , 32'hFFFE346F , 32'hFFFFBC59 , 32'hFFFD8FC5 , 32'hFFFCECE2 , 32'h0005D9BE , 32'h000439B1 , 32'hFFFC29CE} , 
{32'h0002A8D6 , 32'hFFFFC80D , 32'hFFFDAED7 , 32'hFFFBD3F0 , 32'h000256F7 , 32'h00051350 , 32'h00028D42 , 32'h00005054 , 32'hFFFF285A , 32'h00031BA5 , 32'hFFFE423A , 32'hFFFD5B9B , 32'h000613DF , 32'hFFF81FBC , 32'hFFFDBF27 , 32'hFFFE97C8 , 32'h00068E82 , 32'hFFFFECE5 , 32'hFFFDF1D6 , 32'h00066175 , 32'hFFFE6C61 , 32'h000511C0 , 32'h00039FE4 , 32'hFFFC88FF , 32'h000723FB , 32'h0003BB2B , 32'h00009E19 , 32'h0001F852 , 32'hFFFE8414 , 32'hFFFFD39D , 32'h000050CB , 32'h00078E8A , 32'h00021E4C , 32'h0000754B , 32'h00033B94 , 32'hFFFF3B09 , 32'h00026087} , 
{32'h028D6E58 , 32'h0211C030 , 32'hFC240D10 , 32'hFDA57C5C , 32'hFF5C4E72 , 32'h011B7874 , 32'hFDA146B4 , 32'h010CF3AC , 32'hFD6771B0 , 32'h0032FBBF , 32'hF7829690 , 32'h00FAD04E , 32'h04C841B8 , 32'h03B03B90 , 32'h037509E0 , 32'hFF255E98 , 32'h03C0475C , 32'h040508B0 , 32'h01B94D40 , 32'hFB262AD8 , 32'h02B52270 , 32'hFECBC0C4 , 32'hF9A7FD10 , 32'hFE895268 , 32'h0086713F , 32'h02ADB8AC , 32'h0B291DE0 , 32'h0333C044 , 32'h04551498 , 32'hFD9AF640 , 32'hFC4CEC90 , 32'h04DA0A50 , 32'h04555438 , 32'hFDD21EA8 , 32'h0265CCB8 , 32'h012DF15C , 32'h04A8C0A8} , 
{32'h00CDA3EF , 32'h0A846B40 , 32'h12E1A3E0 , 32'h051F2978 , 32'h11499640 , 32'h0138F0D8 , 32'hF927AAF8 , 32'h0FEDEE70 , 32'h0E15F9F0 , 32'h01364CB4 , 32'hF605F1F0 , 32'hFB895E90 , 32'h177C63E0 , 32'h081AA1F0 , 32'h02C6ABF4 , 32'h0C49EBB0 , 32'hFE19B04C , 32'h0064F817 , 32'h02744FA0 , 32'hF7777230 , 32'h026F5BBC , 32'hFAF6D9B8 , 32'h04BC9480 , 32'hFD3C3BE4 , 32'h069BF2D0 , 32'hF8018F30 , 32'h06A16318 , 32'h112441E0 , 32'h01E9ED44 , 32'hFF3F4F53 , 32'hFA4B1040 , 32'hFD094870 , 32'h138B3780 , 32'h0509ACB0 , 32'h03A4211C , 32'h03FD8068 , 32'h029E1354} , 
{32'h069CB020 , 32'hFDC9F55C , 32'h03A2B1E8 , 32'h028A0D80 , 32'h038B74FC , 32'h03FF2498 , 32'hFCD9605C , 32'hFF06D00C , 32'h08870450 , 32'h005D36DE , 32'h07397950 , 32'h10DE3100 , 32'h06373C40 , 32'hF9C9E090 , 32'hF3126990 , 32'hFE0A78C0 , 32'h14F37740 , 32'hF7F8BEB0 , 32'hF3CF91B0 , 32'h0A9D8BA0 , 32'h012A12E0 , 32'h0F5E7560 , 32'hFEA96BD0 , 32'h028D8478 , 32'hF7BCD470 , 32'hF688B9C0 , 32'hFF8E68C7 , 32'h045A9060 , 32'h0A11A120 , 32'h06604EF0 , 32'h06536528 , 32'h0C23CD90 , 32'h02DF05D0 , 32'hFDD952EC , 32'h098F6230 , 32'hF1497D90 , 32'hFA1ECD28} , 
{32'h0248B780 , 32'h0F1AEAD0 , 32'hFF9AEC19 , 32'hF7C64D90 , 32'hEE338B20 , 32'h24C68AC0 , 32'h145821A0 , 32'hFEC8A5A8 , 32'h1E0D12C0 , 32'hFC444A14 , 32'h0EC71090 , 32'hF8B51DF0 , 32'h02DD05BC , 32'hFE2EC95C , 32'h165D5060 , 32'h0C5453F0 , 32'hF9110BE8 , 32'h0D0CF9C0 , 32'h152A67A0 , 32'h139D4F80 , 32'h001D2788 , 32'h19E7BB80 , 32'hF860BC88 , 32'h041587E8 , 32'h0739B9C0 , 32'h069D8780 , 32'h0D54D930 , 32'hFC6784F4 , 32'h0D74CE00 , 32'hE8950B60 , 32'h1A113900 , 32'hF45A45D0 , 32'h005AF326 , 32'h0077CC8B , 32'hF1F23020 , 32'hE5D9B2E0 , 32'hF7C0D940} , 
{32'hF4734000 , 32'h0900F600 , 32'h069DCE28 , 32'hF56D6AB0 , 32'h05DA8290 , 32'h01FCC514 , 32'hF8F49878 , 32'hFAAB6E98 , 32'h189B4640 , 32'h01746694 , 32'hFE1E7240 , 32'hFAFFC668 , 32'h0EB02DB0 , 32'hEF8A51A0 , 32'h1566E480 , 32'h153A6040 , 32'hF2A235C0 , 32'hF4AA0930 , 32'h0C079510 , 32'hEF4E4C20 , 32'hFEB675F4 , 32'h161094C0 , 32'hE4B61C80 , 32'hED3CE8E0 , 32'h0222FCAC , 32'h08EAAD90 , 32'h16B089A0 , 32'hFB186B60 , 32'hFDB61FA4 , 32'h000EEF94 , 32'h0AB160F0 , 32'hFCE9A2AC , 32'hF7586050 , 32'hF7611FE0 , 32'hF462C840 , 32'hF50F7280 , 32'h057FEC18} , 
{32'hF3874690 , 32'h1BDEF160 , 32'h18ACDD80 , 32'hD61D8DC0 , 32'hF9F5A210 , 32'h0F2E3D60 , 32'hD36CD640 , 32'h335A3A00 , 32'hF84EFA98 , 32'h0096A878 , 32'hF87A90A8 , 32'h0E9CB3A0 , 32'h1C738D60 , 32'hF835EDD0 , 32'h1F3CD200 , 32'h12F562C0 , 32'hDA634140 , 32'hE573E8C0 , 32'hE244F0A0 , 32'hFF622A89 , 32'hFA8DBD10 , 32'h046B5198 , 32'hDDD27E00 , 32'hF575DA60 , 32'h18AC6840 , 32'hDB6FD2C0 , 32'h15630BE0 , 32'h083752E0 , 32'h04AE74A8 , 32'h2566CC80 , 32'h198ABEE0 , 32'hD7E79200 , 32'hEF6B0C20 , 32'hFF021AF3 , 32'hDDDA69C0 , 32'hF5980750 , 32'hFA72EAF0} , 
{32'hEBC6B2A0 , 32'h004F5CE4 , 32'h162E8A20 , 32'hEA137F20 , 32'hFABCC4D0 , 32'hE3E921A0 , 32'hF5495E90 , 32'h1D29EAA0 , 32'h117BE600 , 32'h08768040 , 32'hFB81ED10 , 32'h151CD660 , 32'h10EC35E0 , 32'hE94360E0 , 32'h2CF616C0 , 32'h11F92740 , 32'hFBBA77A8 , 32'hF72859B0 , 32'h021EC200 , 32'h02819440 , 32'hE9E21200 , 32'h07D59AD0 , 32'hD920BC40 , 32'hF26DC690 , 32'hFC9B8670 , 32'h02464AB0 , 32'h0D669660 , 32'h06F1F190 , 32'hF5336970 , 32'h0BDACEE0 , 32'h0C9C13B0 , 32'hFFD7C419 , 32'h0186EDAC , 32'hFB01B4C8 , 32'h031A1E80 , 32'h00C895B8 , 32'hF86F6E30} , 
{32'hF0D7AE20 , 32'h074DACF8 , 32'h13F23A20 , 32'hE8E03820 , 32'h06D8D9D8 , 32'hE8868500 , 32'hEBB20B80 , 32'h16E65B00 , 32'h05FB8D10 , 32'h153B90A0 , 32'h06925AE8 , 32'h0A4068D0 , 32'hF7764240 , 32'hDC33FAC0 , 32'h1AA4FC80 , 32'h0BB38B60 , 32'hFF6F00D9 , 32'hF71FD240 , 32'h0A76B720 , 32'hF3168A60 , 32'hF7E2E320 , 32'h04FBCDF0 , 32'hE9CECD20 , 32'hF9E5F3B8 , 32'hF8AC19D8 , 32'hF6B3E960 , 32'h0D5645E0 , 32'hFEF91B2C , 32'hFDCF5CC8 , 32'h121A4BA0 , 32'h1E19F640 , 32'h075F4A30 , 32'hF9785578 , 32'h039F5018 , 32'h14CBDBA0 , 32'hF3CA8480 , 32'h08267DA0} , 
{32'hF69F6C70 , 32'h0E634DC0 , 32'h14A82DA0 , 32'hD6BEC700 , 32'hF4376CE0 , 32'hC255C100 , 32'hF7B23C20 , 32'h1C08B300 , 32'hC15FADC0 , 32'hECD9C620 , 32'hF5620490 , 32'h07567BC0 , 32'hEF9A1920 , 32'hD686CF40 , 32'h27EB6940 , 32'hEFFFF080 , 32'h23A24EC0 , 32'hE7FC6060 , 32'h041D7F10 , 32'h0D6CB770 , 32'hF753CE10 , 32'h1656FBA0 , 32'hF3ECFC20 , 32'h0FEDF820 , 32'hF4E1EFF0 , 32'h001572A3 , 32'h130D02A0 , 32'hF0ADEB40 , 32'h11ADA0A0 , 32'hFD4C137C , 32'h0FA60B20 , 32'h01BD0604 , 32'h07B2C150 , 32'h1BAFACC0 , 32'hF7FCE4C0 , 32'h00B7901C , 32'h014CD63C} , 
{32'hDDE3F540 , 32'h19D1E140 , 32'h19C15900 , 32'hF307A030 , 32'h0227BB44 , 32'hD372CF00 , 32'h02E066C0 , 32'h0F705750 , 32'hDB684500 , 32'hDA962040 , 32'hF628C5D0 , 32'hFE2C4194 , 32'h022917AC , 32'hD8A5CA00 , 32'h0982CA00 , 32'hEC209E20 , 32'h116E7D20 , 32'hFB9DB600 , 32'h0F883AC0 , 32'h0BFBD6B0 , 32'h041F3AC0 , 32'h01028900 , 32'hF66A4E30 , 32'h08D08030 , 32'hF1AEEE10 , 32'hFDEACFF0 , 32'hE5B812A0 , 32'hFA10C000 , 32'h042F1800 , 32'h069DDAF8 , 32'h090FD380 , 32'hFD12F504 , 32'hFC425BA8 , 32'hF43B0560 , 32'h1097B320 , 32'hFBE0A948 , 32'h136E4A40} , 
{32'hDA8589C0 , 32'h1204EF80 , 32'h00F9E274 , 32'hEA76C780 , 32'hFA487E68 , 32'h04567608 , 32'h061EA5F0 , 32'hF8FCF680 , 32'hE42DC380 , 32'hE269C840 , 32'hF366EAA0 , 32'h03CAE184 , 32'h06D1E198 , 32'hE4E48460 , 32'hFC77C1BC , 32'hE6E601A0 , 32'h0752DCA0 , 32'h0092893D , 32'h15B9AF40 , 32'h3D42ECC0 , 32'h09A40FC0 , 32'hF81ABC80 , 32'hFAEF27A0 , 32'h0AD7E8F0 , 32'hD5A26380 , 32'h1BC6D880 , 32'hEC989D20 , 32'hF284DFB0 , 32'hFABA1C40 , 32'h0E5DEDF0 , 32'hFF33B592 , 32'hFC8A0544 , 32'hDCF00C40 , 32'hE913DC40 , 32'hF59FAD80 , 32'h06358F70 , 32'h11DC15C0} , 
{32'hE7B33120 , 32'h1DE92500 , 32'hFBFC7318 , 32'h06785588 , 32'hEECD4560 , 32'h0E4954F0 , 32'h0C093310 , 32'hF35CC520 , 32'hFC59CE60 , 32'hEC7C5820 , 32'hEC48A9E0 , 32'hF98B9CD0 , 32'h180F8A00 , 32'h07B47748 , 32'hF0C10870 , 32'hE9E711E0 , 32'hF12F0650 , 32'h09304A00 , 32'hFB726A10 , 32'h143C5EC0 , 32'hEF779E40 , 32'h11EB7C40 , 32'h00DC390B , 32'h1637BC60 , 32'hEEBECAE0 , 32'h16228A40 , 32'hEEAD5AC0 , 32'hFEBFD968 , 32'h09A19500 , 32'hF9E5EA80 , 32'hFAAFA958 , 32'hEE407A60 , 32'hFF2F49E5 , 32'hFDEE32E0 , 32'hFC57387C , 32'h02C13ABC , 32'h11D39B00} , 
{32'hEC0EDE00 , 32'h0BD0A0E0 , 32'hF62983B0 , 32'hF54728E0 , 32'h0540C2A0 , 32'h157B18C0 , 32'h02A59F90 , 32'hD9E2A3C0 , 32'h07D63D28 , 32'h0136C0C4 , 32'hF516C6F0 , 32'hF4CB9570 , 32'h0CE2DE00 , 32'hDC5AE840 , 32'hF80D9EA8 , 32'hFAF1FFC8 , 32'h067C0020 , 32'h0E0D5C50 , 32'h0146B3A8 , 32'h1407A780 , 32'hFE96E484 , 32'hEBCCD120 , 32'h11640D20 , 32'h16C027C0 , 32'h03BCF2C4 , 32'h0944E2D0 , 32'h06334AF8 , 32'h14E91D60 , 32'h091B0AF0 , 32'h08CB0860 , 32'h0502EF38 , 32'h0837D350 , 32'h04D6C780 , 32'h01D4C9AC , 32'hF84FBBA8 , 32'h1550B420 , 32'h00E4B873} , 
{32'hEA757680 , 32'h1FD1C8C0 , 32'h049AD0C0 , 32'hEA6C3520 , 32'h0822AE70 , 32'hFDA5891C , 32'h0B811370 , 32'hD8D65F80 , 32'hFCE75F68 , 32'h23BEF600 , 32'h066B6560 , 32'hF1A2A190 , 32'h0A72C900 , 32'h08DE6750 , 32'hF4174270 , 32'hEE62DA80 , 32'hFD97C128 , 32'hFB6D21A0 , 32'h12D44B20 , 32'h172802C0 , 32'h01091E14 , 32'h15734740 , 32'h0E8666B0 , 32'h158E8020 , 32'hF2928800 , 32'h0BAA1760 , 32'h10F27AA0 , 32'hF6CA3B00 , 32'hF05B6300 , 32'h00E46D6F , 32'hE999DC40 , 32'hF0387E10 , 32'hF4ACC7E0 , 32'h08D6CEA0 , 32'hF2921340 , 32'hF0100F50 , 32'h09D93580} , 
{32'h0765ACE8 , 32'h2605E680 , 32'hF7481B10 , 32'hC5493D40 , 32'hF65660F0 , 32'h06813660 , 32'h094D4C00 , 32'hC8D101C0 , 32'hFA6FE1A8 , 32'h2875D600 , 32'hEBBB5300 , 32'hE68819C0 , 32'hF86A6138 , 32'h0FC680E0 , 32'hFAF9BC48 , 32'h0ADD95A0 , 32'hEF2DC840 , 32'hFE1A7FCC , 32'h2D413180 , 32'h17D1DB60 , 32'hF919BBA8 , 32'hFDF99E10 , 32'h1DE2FC60 , 32'h05DD40B8 , 32'hF9943038 , 32'h15B02960 , 32'h265A4C00 , 32'hFBCCD7A0 , 32'hDD989440 , 32'hFE852718 , 32'h1D2E5860 , 32'h09D37A00 , 32'h2797A1C0 , 32'h03A13904 , 32'hDE12B3C0 , 32'h0C7CAFF0 , 32'h11AA8FA0} , 
{32'h06814B58 , 32'h17D643A0 , 32'h02EBC0B4 , 32'hD9EAEA40 , 32'h017558E8 , 32'h0EAAEFA0 , 32'hF98DC180 , 32'hD0469A80 , 32'h09050540 , 32'h19712B60 , 32'h1E1A8BA0 , 32'h0C720DC0 , 32'h0A880190 , 32'h01CB85D4 , 32'h0B4C2A60 , 32'h06B64CF8 , 32'h16F1F8E0 , 32'h0E4AFA80 , 32'h02849528 , 32'hFC881F74 , 32'h0B121100 , 32'hFCA49D1C , 32'hF636DF80 , 32'h0E64D4D0 , 32'hF1C0C6A0 , 32'hF25A6BA0 , 32'hF5AE99A0 , 32'h16249160 , 32'hF1123F40 , 32'h0DB45FF0 , 32'h1132AAC0 , 32'h160BC380 , 32'hF8D2A2C8 , 32'h0F8DF540 , 32'hF92ABE08 , 32'h335FE1C0 , 32'hE5676E20} , 
{32'h00731EBC , 32'h0ED21900 , 32'h0C03D7B0 , 32'hDFFDB2C0 , 32'h09F06E70 , 32'hFB2BB320 , 32'hFCE6EB90 , 32'hFDAD405C , 32'hF97E4578 , 32'h186E6DE0 , 32'h08D07150 , 32'hF04C3090 , 32'hFD681380 , 32'hFD8F0CEC , 32'hFE7B233C , 32'h08BB70C0 , 32'hF19A0980 , 32'hFD634FA4 , 32'h168C6E00 , 32'h1087A2C0 , 32'hE7B47900 , 32'h138ED780 , 32'hEA1FC060 , 32'hF47EF680 , 32'h0599E8F0 , 32'hF2E70A70 , 32'hF6BCF8F0 , 32'h094A1A30 , 32'hF48F4780 , 32'hFDE37F8C , 32'h0373F190 , 32'h116D01E0 , 32'h06C852B8 , 32'hFDED5020 , 32'h184DF1E0 , 32'h0590A048 , 32'hFE27DEC4} , 
{32'h0282C868 , 32'hFE51CD88 , 32'h06C46378 , 32'hF7AF9A10 , 32'h03AD87A0 , 32'hFEE66854 , 32'hF55407F0 , 32'h0A254630 , 32'hFAAEA310 , 32'h05F0E290 , 32'h190127E0 , 32'h12FF3A40 , 32'h2CCFAB80 , 32'h0961AF60 , 32'h08713260 , 32'h04A710B0 , 32'hF2F7EDA0 , 32'h06EFD160 , 32'hFF749529 , 32'hFF67CE2B , 32'h078568C8 , 32'hFBC1DA88 , 32'h055CC078 , 32'hF75E4190 , 32'hF5417060 , 32'h0C90F720 , 32'hF74BFE70 , 32'h0E615810 , 32'h04C36EB0 , 32'h01A30630 , 32'hF7041B10 , 32'hFD4BF6F0 , 32'h00B055AF , 32'h0ACAB710 , 32'hFFD2D97A , 32'hFBCBECB8 , 32'h06412AE8} , 
{32'h0515EB58 , 32'h0FBF14B0 , 32'h153B9880 , 32'hE260D1E0 , 32'h0B91D790 , 32'hF2A73280 , 32'hFE609B38 , 32'hE847FB00 , 32'hCE0EE740 , 32'h0BFE27E0 , 32'h21470FC0 , 32'h03DF10BC , 32'h08E23C40 , 32'h064746D8 , 32'h08F3EAC0 , 32'h1888B960 , 32'h03DE0D6C , 32'hF98060B8 , 32'h01B2DB00 , 32'h0083141C , 32'hF36DBBD0 , 32'hF7281820 , 32'h093B3C20 , 32'hD83E23C0 , 32'hFEBE3064 , 32'hEDD84B00 , 32'hF2EB9410 , 32'hF94A9A28 , 32'hEE385E40 , 32'hFA47A2C0 , 32'hF1899B30 , 32'h09492220 , 32'h0DD7FB70 , 32'hFDB46090 , 32'h034F30DC , 32'hFA0F0188 , 32'h0009D0D4} , 
{32'h036C6458 , 32'hFECF34D8 , 32'hFF5838F5 , 32'h0203A528 , 32'hFEBA1F24 , 32'hFBA5F470 , 32'hFC9F7DD4 , 32'h0D08D830 , 32'hFBBA30C8 , 32'h05BFC7C8 , 32'h07CA5D60 , 32'h09A48BD0 , 32'h0BD114B0 , 32'h034A8F14 , 32'h06E7E9B0 , 32'h05F99478 , 32'hF6C4C2E0 , 32'h02B7C320 , 32'hF6381240 , 32'h003856B6 , 32'hFF895DAB , 32'h01FCAE10 , 32'hFC53A48C , 32'hF89242C8 , 32'hFD2C1CD8 , 32'h0817D7E0 , 32'hFA8FE820 , 32'h062C6130 , 32'hFCDBB5F4 , 32'hFE5A5148 , 32'hF96D06F0 , 32'hFC9EBDAC , 32'h04726F88 , 32'hFEE6EE28 , 32'h00B01321 , 32'hFDCCA29C , 32'hFEA55420} , 
{32'h0047ED2A , 32'h002E3677 , 32'h006ABFF2 , 32'hFFA39C80 , 32'h00663F5C , 32'hFFE28520 , 32'h0003140D , 32'hFFBA1A78 , 32'hFF4D4618 , 32'h002EB65D , 32'h00D3D25A , 32'h00978FD0 , 32'h006EC446 , 32'hFFE1F6A6 , 32'h0013068E , 32'h005F360B , 32'hFFAFB5EC , 32'h004D8442 , 32'hFF91E0FB , 32'hFFD7D89E , 32'hFFD73C8C , 32'hFF8F60D8 , 32'hFFFAF261 , 32'hFF34792F , 32'hFFE4256F , 32'hFFE3A55B , 32'hFFA3B1BC , 32'h00654C11 , 32'hFFB24F03 , 32'hFFF36B3C , 32'hFF55F88E , 32'hFFDA624F , 32'h00D7A199 , 32'hFF9C18C8 , 32'hFFBBDF6F , 32'hFF793530 , 32'hFF861DDC} , 
{32'h0000E928 , 32'h00007D14 , 32'hFFF89905 , 32'h00010B72 , 32'h00033358 , 32'h0000E333 , 32'hFFFCD605 , 32'h0001CEAD , 32'hFFFE0CB0 , 32'hFFFC18E9 , 32'hFFFEBDB7 , 32'hFFFF494E , 32'hFFFB8B01 , 32'hFFFFF3A5 , 32'hFFFD2F16 , 32'h0001511F , 32'hFFFB13B4 , 32'hFFFF50C4 , 32'hFFFD90D0 , 32'hFFFCB7FE , 32'hFFFEC7EC , 32'hFFFFAB47 , 32'h000460C5 , 32'hFFFDB0C1 , 32'hFFFE0B6D , 32'h00032DD7 , 32'hFFFDB7BF , 32'hFFFA7288 , 32'h0000F583 , 32'h0008C7D2 , 32'h00003B59 , 32'hFFFE61E0 , 32'hFFFA8EA5 , 32'hFFFD73BC , 32'h0000BB74 , 32'h00013885 , 32'h00031F1E} , 
{32'hFFFCA19D , 32'h000062A0 , 32'h0000A5A8 , 32'h0000D76C , 32'hFFFE9A0D , 32'hFFFFCAE0 , 32'h000138F8 , 32'h0001449C , 32'h0000D54E , 32'hFFFCDFDC , 32'hFFFB58E4 , 32'h00004FFE , 32'hFFFFB9F1 , 32'hFFFF7369 , 32'h00010139 , 32'h0004026D , 32'h00004E9A , 32'hFFFFDBC1 , 32'hFFFCD37D , 32'hFFFFEFDD , 32'hFFFF57B4 , 32'hFFFB0509 , 32'h0003A295 , 32'hFFFEBBDB , 32'hFFFC7EC7 , 32'h00002C3A , 32'hFFF83A09 , 32'hFFF8A707 , 32'hFFFE6CF6 , 32'h00030B58 , 32'h0001E19B , 32'h00050C10 , 32'h00071BB4 , 32'h00011DBA , 32'h0005B5D1 , 32'h0000931D , 32'hFFFE8959} , 
{32'hFFFBD3BA , 32'h00014BA7 , 32'hFFF85F0E , 32'hFFFBEDA6 , 32'h00015916 , 32'h0000FE9C , 32'h0001464D , 32'hFFFB45F0 , 32'hFFFD5E9D , 32'h000051B7 , 32'h0000972C , 32'hFFFF41C3 , 32'hFFFE7184 , 32'h000140CD , 32'hFFFC05FB , 32'h000586E0 , 32'hFFFC6DC8 , 32'hFFFD1ED2 , 32'hFFFFC49E , 32'h00003D3D , 32'h0000209A , 32'h00005A59 , 32'hFFFCEFF1 , 32'h0000231E , 32'h000545DF , 32'h0004A4B8 , 32'h0006DC4C , 32'hFFFF8682 , 32'h0002CB8C , 32'h0002C81E , 32'hFFFF4FD8 , 32'hFFFD7309 , 32'hFFFE78C9 , 32'hFFFBAD81 , 32'h0000267D , 32'hFFFD894A , 32'hFFFE435E} , 
{32'hFFFBCEE9 , 32'h0007C796 , 32'h0001E259 , 32'hFFFF41CE , 32'hFFFEA519 , 32'h0004C89A , 32'hFFFFEB31 , 32'h00002EB5 , 32'h0000E1CA , 32'h0000C902 , 32'h000556AF , 32'h00028299 , 32'h00027FA3 , 32'h00008E6D , 32'h00046C81 , 32'hFFF82A5F , 32'hFFFFBAEA , 32'h0002AAAE , 32'h00023BD9 , 32'h0000C22D , 32'hFFFBE085 , 32'hFFFFDE78 , 32'hFFFB06DE , 32'hFFFF4487 , 32'hFFFECA5C , 32'h00036C72 , 32'hFFFDBDD7 , 32'h0000ED32 , 32'h0001038C , 32'hFFFD3349 , 32'hFFFBA9C4 , 32'h00028F9E , 32'h00033CA6 , 32'hFFFF767F , 32'hFFFD9FFD , 32'h0004445C , 32'hFFFC1C5D} , 
{32'h000140B7 , 32'hFFFDF79F , 32'hFFF9AA02 , 32'hFFFFA985 , 32'h0002A425 , 32'hFFFF76C2 , 32'h0003DDCA , 32'h00065EB3 , 32'hFFF89C19 , 32'h0004FD37 , 32'h0004A938 , 32'hFFFF698B , 32'hFFFF7613 , 32'hFFFCB7E0 , 32'hFFFF2616 , 32'h0004826B , 32'h000024C3 , 32'h00034ED9 , 32'h000041EB , 32'h0006B7EF , 32'hFFFD8585 , 32'hFFFE8E28 , 32'hFFFD4DB4 , 32'h0001BF05 , 32'h00016E47 , 32'h000401DC , 32'hFFF9E282 , 32'hFFFB353D , 32'hFFF83D00 , 32'hFFFB1EC0 , 32'hFFFF0796 , 32'h0001AF15 , 32'hFFFF79B7 , 32'h00077A82 , 32'h000426EC , 32'h00059828 , 32'hFFFD6D65} , 
{32'h000457DF , 32'hFFFFA0FC , 32'h0001B16F , 32'h0001C72D , 32'h000019BB , 32'h00006D57 , 32'h00036E14 , 32'h0001B6C6 , 32'hFFFE05BF , 32'h00001403 , 32'h0002D3DE , 32'h000029CD , 32'h00003DC8 , 32'hFFFE1657 , 32'h000073CB , 32'hFFFE5A6F , 32'h0002499D , 32'h0002A096 , 32'hFFFE3706 , 32'h000119B1 , 32'hFFFD6191 , 32'hFFFB9226 , 32'hFFFCE34B , 32'h0000E2CC , 32'h00002076 , 32'hFFFCB4DB , 32'hFFFDFCA0 , 32'hFFFF02A3 , 32'hFFFE80A5 , 32'hFFFD3E99 , 32'h000425CB , 32'hFFFCB1AA , 32'h0000B2DF , 32'h0001A2D8 , 32'h00041783 , 32'h00000788 , 32'hFFFCFB33} , 
{32'h00A7D599 , 32'h055CCF80 , 32'h0309B114 , 32'h04524300 , 32'h0341FCF0 , 32'h027E40D0 , 32'hF817F748 , 32'hFE8D3528 , 32'h039FE1A4 , 32'hFFB33A11 , 32'h00FC3022 , 32'h02A70EC0 , 32'hFD040A54 , 32'h0944B160 , 32'hFAADD460 , 32'h020204A0 , 32'h05FEC118 , 32'hF57D9F30 , 32'h062FD7A0 , 32'h03A21E0C , 32'hFAE52CA8 , 32'hFB12EC50 , 32'h002EE339 , 32'h0030E1FA , 32'hFEF28F80 , 32'h038EB534 , 32'h0844B5F0 , 32'h039FCA98 , 32'h039DEBD0 , 32'hF5CFD590 , 32'hFB81E6E0 , 32'hFEC1C0F0 , 32'h019BA428 , 32'h02755F20 , 32'hFD707908 , 32'h008234E0 , 32'h00157B2E} , 
{32'h004C4279 , 32'hFF0C8DB5 , 32'hFD8E5A54 , 32'hFFB43B8B , 32'h0260CA00 , 32'h0E2D0A30 , 32'hFD755488 , 32'hFB658D50 , 32'h0DC3DC40 , 32'h03B7D198 , 32'h02C38B94 , 32'h019FF794 , 32'h015355BC , 32'h0128435C , 32'hFF649344 , 32'h08D31140 , 32'hF9D575B0 , 32'h007CA302 , 32'hFA4CBBF8 , 32'hFFAB56FE , 32'h0018613C , 32'hF75043B0 , 32'hFE6C9594 , 32'hFBF5E238 , 32'hF9307998 , 32'h0221415C , 32'hFF9E8BB0 , 32'hFC529390 , 32'h004F7507 , 32'h01D63070 , 32'hFDF97200 , 32'hFD3C2A64 , 32'hFD8233B4 , 32'hFB568F58 , 32'h0900F660 , 32'h02F908DC , 32'h018AB2AC} , 
{32'h0A247570 , 32'h01686D34 , 32'hFAFB2698 , 32'h00C3EA16 , 32'h00F91E9B , 32'h09871360 , 32'hF56772B0 , 32'h018752B4 , 32'hF964D1A0 , 32'hFFBA2775 , 32'hF7E68A70 , 32'h04E9A518 , 32'h091EA300 , 32'h004A87A0 , 32'hFDAD0EDC , 32'hFA18BD60 , 32'h0F12F150 , 32'hFEA53CC8 , 32'hFFB5293D , 32'h03C8A34C , 32'h022592AC , 32'h000F1179 , 32'hFD54CB84 , 32'hFAC25930 , 32'hFF0FAF55 , 32'h0459E960 , 32'h131C2900 , 32'h06185700 , 32'h093FA240 , 32'hFAF54CB8 , 32'hFC9E337C , 32'h0985FFF0 , 32'h06237E78 , 32'hFEE4D994 , 32'h0091600E , 32'hF97309A8 , 32'h045BBB58} , 
{32'h07726490 , 32'h0C2706A0 , 32'h0428DFB8 , 32'hEC09C7C0 , 32'h00133B62 , 32'h10749380 , 32'hFCBE19FC , 32'h0FCE1D40 , 32'h09B91990 , 32'hFC2958BC , 32'hFE218F1C , 32'hF5E1E930 , 32'h05D552B8 , 32'h0C639460 , 32'hF73D9BE0 , 32'h07243280 , 32'hF8AD7070 , 32'hF6E5A490 , 32'hF358EFE0 , 32'h00042CE5 , 32'h0F7CCB50 , 32'hEE7DD1C0 , 32'hF6875550 , 32'h0B20DC10 , 32'hFFD3577B , 32'hEE577180 , 32'h03A39F04 , 32'hFBA29710 , 32'hF0501B80 , 32'hF9A3CF78 , 32'hFC58205C , 32'hFE90D6D8 , 32'hFA7E7560 , 32'hF0061890 , 32'hFA505898 , 32'hF78B07A0 , 32'hFF88EAD0} , 
{32'h075F7598 , 32'h045CDDB8 , 32'hFBD495D8 , 32'hF4A0C500 , 32'hFCFAD9EC , 32'h2E4E4E40 , 32'h0BA14280 , 32'h0E052C00 , 32'h13230B40 , 32'hC96CCE00 , 32'hFDAA049C , 32'h068E2710 , 32'h2097BD40 , 32'hFC405648 , 32'hFC383950 , 32'hE703C580 , 32'h0874A7D0 , 32'hF873E740 , 32'hF520B1C0 , 32'h28D76640 , 32'h0366E1DC , 32'h2C3BD400 , 32'hEB605000 , 32'hE0537600 , 32'h04A061B0 , 32'hE88805A0 , 32'h0E17A460 , 32'h0F761D60 , 32'h0289344C , 32'h0608F480 , 32'hED8FF5A0 , 32'h0539F870 , 32'hFE4212DC , 32'h1049E140 , 32'h10C92F00 , 32'h1245A700 , 32'h0EADA740} , 
{32'h076CDE40 , 32'hFF96E6CE , 32'hFC71D1FC , 32'hED4B8D00 , 32'hF7675340 , 32'h1C951F80 , 32'hED174840 , 32'h0620EAC0 , 32'h155478C0 , 32'hFB82CAA8 , 32'hF75ACFE0 , 32'hFF1936E6 , 32'h02CF4844 , 32'hF43B4E20 , 32'h0FE049E0 , 32'h1C316080 , 32'hED7AF180 , 32'hFB33A8C8 , 32'hF7D71E30 , 32'h08FE3440 , 32'hF22F8D80 , 32'hF60EC390 , 32'hE4E49440 , 32'hFE2D0094 , 32'hE5EA9CC0 , 32'h088B6790 , 32'h07BEAFB0 , 32'hEE0B9680 , 32'hFC820E3C , 32'h162E29C0 , 32'hFB7AD5A8 , 32'hFD6D4E38 , 32'hFDC4D254 , 32'hFC7AE5F8 , 32'hFB3ED270 , 32'h139D72A0 , 32'hF971D300} , 
{32'h029B427C , 32'h11DECD00 , 32'h126C2480 , 32'hF3EC6450 , 32'h0525D088 , 32'h114714C0 , 32'hEBB02260 , 32'h0A8B7FC0 , 32'h1EF4ECA0 , 32'hFD6D6E20 , 32'hEE48C780 , 32'hFEF38E74 , 32'hFCB937BC , 32'hE25EBAC0 , 32'h1B3F2100 , 32'h2187B640 , 32'h01303FF8 , 32'h049F8A40 , 32'hDCD9E7C0 , 32'h0E89C700 , 32'hF7323D10 , 32'h08564F80 , 32'hE7BBF580 , 32'hE705AB00 , 32'hE49ED8E0 , 32'h0D856D50 , 32'h07FD4928 , 32'h05AFA640 , 32'hEC3D6E20 , 32'hFD4DFC18 , 32'h0640D3E0 , 32'h14041BC0 , 32'h07043338 , 32'hF96A5D88 , 32'hE056CB80 , 32'h0A3C1D10 , 32'h13864C60} , 
{32'h02BD2D20 , 32'hFD390144 , 32'hF7248AA0 , 32'hEBC15420 , 32'h04A6EAE0 , 32'h0349EDE0 , 32'hE023D4E0 , 32'h037687C0 , 32'hF1BF8770 , 32'hEEC24820 , 32'hFF5979C4 , 32'hFEC06F68 , 32'hF6064350 , 32'hF1983430 , 32'h0B33EC80 , 32'hFEF6D85C , 32'h020FF6D8 , 32'hFB712368 , 32'hF620EDB0 , 32'h0ADE7650 , 32'hFF0A2B98 , 32'h020B4B40 , 32'hF9A383C0 , 32'h0B17E730 , 32'hFE44F78C , 32'h07D6C7C8 , 32'h02AF36E4 , 32'hE5594700 , 32'h142685C0 , 32'hFFF2114B , 32'hFA08D780 , 32'hFAA27D70 , 32'h0C3CF670 , 32'h042040A0 , 32'h0DAF32D0 , 32'hFE0BC060 , 32'hFA2391C8} , 
{32'h0C492DC0 , 32'h0645ABE0 , 32'hFC6AFAB0 , 32'hEF1C67E0 , 32'hFD80B9D0 , 32'hFEA634C4 , 32'hEE4988E0 , 32'h0D361C40 , 32'hE88DFAC0 , 32'h0C7BB1E0 , 32'h07D78FB8 , 32'hFE96BB40 , 32'hF67940F0 , 32'hE6F3C0E0 , 32'h0D34EC00 , 32'h136D20A0 , 32'hFE858A28 , 32'hFE112BF0 , 32'hFDBD4490 , 32'hF7630B90 , 32'hEF6580A0 , 32'h025D1BD4 , 32'hFAF71798 , 32'h064B4060 , 32'hED04D900 , 32'hED9815E0 , 32'hFA0037B0 , 32'hDD80EE40 , 32'h013C19D4 , 32'h0FDBEB40 , 32'hFA8BC548 , 32'h06C33428 , 32'h08EEB650 , 32'h0E1E49B0 , 32'h1801D060 , 32'hF3A5FD10 , 32'h06E85BC8} , 
{32'h19F2C400 , 32'hF23A4370 , 32'h01E0B334 , 32'hE6C43920 , 32'hF1C25350 , 32'hDB3F72C0 , 32'hFE8308D4 , 32'h10AAD2A0 , 32'hD5FFFC40 , 32'hECAEA6C0 , 32'hFDD6E7C4 , 32'h06218618 , 32'hF3272860 , 32'hF1006340 , 32'hFD5A2FF4 , 32'h086DB990 , 32'h0D1DD1F0 , 32'h02F80224 , 32'h17C06E60 , 32'h0D3C5CB0 , 32'hEF9F6AA0 , 32'h0C065710 , 32'hF734C7D0 , 32'h0B4D8420 , 32'hF72039A0 , 32'h06DF3EB8 , 32'h007F468A , 32'hFA11FF30 , 32'hF349A500 , 32'h00CD5505 , 32'hE2CF1400 , 32'h00004C45 , 32'h0B590FD0 , 32'hEF5CD460 , 32'hF8DC15E0 , 32'h0E2E5160 , 32'hFE59A958} , 
{32'h03418268 , 32'hF49F6620 , 32'h145E8920 , 32'hFB8DCC78 , 32'hFD18628C , 32'hE1768BC0 , 32'hFFC49F17 , 32'h2190FA80 , 32'hD1EBCC40 , 32'hC741A5C0 , 32'hF50B7FA0 , 32'h01775A8C , 32'h0D380090 , 32'hF98A9690 , 32'h0134E758 , 32'hECB9CEC0 , 32'h1911B3E0 , 32'h0AEAB150 , 32'h0098E458 , 32'h192D08E0 , 32'h09CDCA80 , 32'h04C9CC50 , 32'hF4FAD970 , 32'h0207A4C0 , 32'hF8B19E88 , 32'hF2BEB010 , 32'hDA043600 , 32'h05857C80 , 32'h0652A798 , 32'h15B97880 , 32'h16CA7B60 , 32'h0810C1B0 , 32'h14D08FC0 , 32'hE8F8B0A0 , 32'h0E06C880 , 32'h06141C38 , 32'hFC982B04} , 
{32'hFFB2BD4B , 32'h01CDA670 , 32'h146E0000 , 32'hE518F440 , 32'hFEC3E968 , 32'h04E829F8 , 32'hFE895FBC , 32'hE2D253E0 , 32'hE6389BE0 , 32'hC4071080 , 32'hF1DDCB30 , 32'h13AEB2C0 , 32'h1A2C73E0 , 32'h106CD940 , 32'hF1D9EFF0 , 32'hFFAD02EA , 32'hEDD1C260 , 32'h13705F20 , 32'hFBBA27D8 , 32'h1E224D60 , 32'h0262481C , 32'hFB411358 , 32'hF3B3F990 , 32'hF1A996D0 , 32'h0EA82150 , 32'h09451290 , 32'hEC745080 , 32'hF3A3A300 , 32'h0334E2D0 , 32'hEDCB8A40 , 32'h0A043320 , 32'hF3CAD210 , 32'h09906C70 , 32'hF2251240 , 32'hDFD25440 , 32'h0283F4B8 , 32'h04BC93F8} , 
{32'h12097420 , 32'hF1573FA0 , 32'h10623180 , 32'hE12F0440 , 32'h020AE7D4 , 32'h19AFDF80 , 32'h1316D940 , 32'hCA06FAC0 , 32'h06C99968 , 32'hD0DF8CC0 , 32'hF57D25B0 , 32'h0802F750 , 32'h2086B6C0 , 32'h0771AA38 , 32'h035B9D40 , 32'hF3F51FC0 , 32'hDC9C2800 , 32'h19917FC0 , 32'h058764B0 , 32'h07C00F30 , 32'h0D336BA0 , 32'h034CF8F8 , 32'hEDAC2A00 , 32'h1778CF20 , 32'hFBBE6498 , 32'h1137FD40 , 32'hD583EB00 , 32'h115D9DE0 , 32'hEC4AFD60 , 32'h0F8090F0 , 32'hFB8B9058 , 32'hF13A46F0 , 32'h15D01D40 , 32'h06E81300 , 32'h0060FD43 , 32'hD79D9740 , 32'h19577A80} , 
{32'h08026A50 , 32'h0C963450 , 32'h0E9BC1F0 , 32'hCF56EAC0 , 32'h02BBF450 , 32'h15E50EC0 , 32'hFFDAF35C , 32'hC2C81F80 , 32'hF93E4310 , 32'hEB299F60 , 32'h08B798F0 , 32'hFA46FFB0 , 32'hFE9FDCA4 , 32'h06FBED68 , 32'hFE339C2C , 32'h037CBEB4 , 32'h001D80A2 , 32'hFB905E28 , 32'h14281440 , 32'hF890AA38 , 32'hF5692010 , 32'hF102D670 , 32'h08026B70 , 32'hF36218C0 , 32'h01D710B0 , 32'hF068DB20 , 32'hF52747A0 , 32'hF901DFF0 , 32'hF3FE3BD0 , 32'hFE21DCE0 , 32'hFD4218DC , 32'hF757B700 , 32'h145C0B40 , 32'h06A489F8 , 32'hF6F511A0 , 32'hF341ECF0 , 32'h099EBA10} , 
{32'h0D999330 , 32'h1607ABC0 , 32'h18DC83C0 , 32'hC1358D40 , 32'h16132760 , 32'h113CA640 , 32'hF7164320 , 32'hBDC55E00 , 32'hFD243724 , 32'h269D29C0 , 32'h1B6CFB00 , 32'hFA5A5730 , 32'hF464BC00 , 32'hF153D830 , 32'hFFE88785 , 32'hFF8B87A7 , 32'hFCF9C3B0 , 32'h00ECFFC4 , 32'h1100E5C0 , 32'h076FB450 , 32'h01E23938 , 32'h046B6DE0 , 32'hF6DD8100 , 32'hED32E480 , 32'h085A6850 , 32'h00C12598 , 32'hFE0CC9EC , 32'h037E0F84 , 32'h05060928 , 32'hFBDD9518 , 32'hEFC8F960 , 32'hF6856D40 , 32'h05B85230 , 32'h0E8ED3C0 , 32'hF94CB230 , 32'hF9493F58 , 32'h07B5F200} , 
{32'h07215528 , 32'h0B66C590 , 32'h02C754DC , 32'hD8CECB40 , 32'h052579A8 , 32'h0D792510 , 32'hF9F9FEC8 , 32'hE8DC8240 , 32'h0131B438 , 32'h2117D200 , 32'h20395740 , 32'hFCB9F3A0 , 32'hFCE3374C , 32'h0795DF20 , 32'h06041010 , 32'hF45ABE00 , 32'hF46E5400 , 32'h02936740 , 32'h0D39B390 , 32'hFF403D91 , 32'h0DC4D640 , 32'h208EB200 , 32'hE6308500 , 32'hFDE26960 , 32'h06BDAD38 , 32'h00AC766E , 32'hFFD68511 , 32'h0E1CE680 , 32'hF90CC0B8 , 32'hFEA212B8 , 32'hF84AE8F0 , 32'hFD8C644C , 32'h0B622D40 , 32'h1B77B6A0 , 32'hF8163558 , 32'hF554C670 , 32'hFDCFDD0C} , 
{32'h0DC16470 , 32'h129AA1E0 , 32'h14E5FBC0 , 32'hE3BF4A00 , 32'h158BC640 , 32'h096E8EF0 , 32'hFF94F2BE , 32'hE3424300 , 32'hF357ADC0 , 32'hF088E2E0 , 32'h0FE54CD0 , 32'h1C23FFC0 , 32'h06149280 , 32'h0725A330 , 32'h0B5FA420 , 32'h0121A984 , 32'hFC9BBCAC , 32'h0B0D1980 , 32'hFFE06C86 , 32'hF8F0B5D8 , 32'h0E65ECC0 , 32'hFE632890 , 32'hFAC6D388 , 32'h021F2B54 , 32'h147F3900 , 32'h089955F0 , 32'hF8CC77B0 , 32'hF64EA6A0 , 32'h0BD37900 , 32'h04ECC108 , 32'hF94DDB40 , 32'h03A9F390 , 32'hFE1DDEF0 , 32'h0A0E4C20 , 32'hE82F4800 , 32'hF5AC7630 , 32'hF9E74058} , 
{32'h0604C460 , 32'h02DA1D40 , 32'h05A1A1D0 , 32'hF9813778 , 32'h07BE17B8 , 32'hEEBBED20 , 32'h0E969030 , 32'hF3F0DA50 , 32'hF3CC5B60 , 32'h13F8DFE0 , 32'h154FA920 , 32'h0CF94DB0 , 32'h0B207AC0 , 32'h0F067180 , 32'h015B3D60 , 32'hFDF3843C , 32'hFA112E88 , 32'h03751CD4 , 32'hF758B770 , 32'hF632B8D0 , 32'hF924D4B0 , 32'hFCCD7BC0 , 32'h0EB0E970 , 32'hFFB94674 , 32'hFD169E34 , 32'h0B3FAB30 , 32'h09712D40 , 32'h0C9DEE50 , 32'hED0FB300 , 32'hFE16A22C , 32'hE9728CA0 , 32'hFCF8E904 , 32'hFC6E3D30 , 32'h04ADF308 , 32'hF725B460 , 32'hFFD18888 , 32'hFFF32A4D} , 
{32'h089F8FC0 , 32'h1071A200 , 32'h0693B280 , 32'hD8E331C0 , 32'h0270B858 , 32'hFFC09A3C , 32'hFC5E38F4 , 32'hFB974CB0 , 32'hE6F4E780 , 32'h0739C818 , 32'hFA5E2628 , 32'hF54BB670 , 32'h0C4594A0 , 32'h0E4B53B0 , 32'hFD7A82F4 , 32'h05E1A6E0 , 32'hE8516D00 , 32'hF774AC30 , 32'h09CAF880 , 32'h07F02E00 , 32'hF145A750 , 32'h05E2C9D8 , 32'h00DC5B24 , 32'hFEC40E3C , 32'hFFFD7840 , 32'hFA77B648 , 32'h02C82970 , 32'h01541A78 , 32'hF4B00690 , 32'h0D1977A0 , 32'h07580AF0 , 32'h067C1010 , 32'h22129A00 , 32'h04573EE0 , 32'h046142F0 , 32'h067746F8 , 32'hE2F85960} , 
{32'h0D0CB450 , 32'h02833784 , 32'h0D1EA280 , 32'hEE7DB360 , 32'h0BDF6750 , 32'h04F407A0 , 32'h01C7FBA0 , 32'hEDC9B520 , 32'hF1B86B40 , 32'hFDAEC130 , 32'h18312A40 , 32'h07312760 , 32'h0AAA9DB0 , 32'hF8DB6B50 , 32'h11A0BE80 , 32'h0C9D58D0 , 32'hF61C6940 , 32'h043D02C8 , 32'hFE3CFE6C , 32'hF79BA240 , 32'h096AC910 , 32'h01E6AF84 , 32'h01046970 , 32'hF5DB2EA0 , 32'h047F7438 , 32'h0556BE50 , 32'hFE4F8C50 , 32'h0AA75AD0 , 32'h0C4DF730 , 32'hFBCF6598 , 32'hFD24C588 , 32'h077C7E50 , 32'h01DDCDCC , 32'h00F01243 , 32'hF2F094E0 , 32'hF5395CE0 , 32'hE52B3FE0} , 
{32'h05BF3920 , 32'h01D27250 , 32'h0AF5E090 , 32'hF765C370 , 32'h08F9D0C0 , 32'hFCA75628 , 32'hFD967BA4 , 32'hF6E3C800 , 32'hF36954C0 , 32'h02BBB01C , 32'h22754B80 , 32'h137B0D40 , 32'h216AB080 , 32'h0942BAE0 , 32'h08EBF220 , 32'h02CD8C8C , 32'hF2B774E0 , 32'h04040288 , 32'hF206FA20 , 32'hF68DAA00 , 32'h0323BD4C , 32'hF292BD10 , 32'h02246ED4 , 32'hF8AF4E78 , 32'hF8EF9270 , 32'h0646A8C8 , 32'hF71D3590 , 32'h154DD680 , 32'hF25785E0 , 32'h03ED5B24 , 32'hE89EC260 , 32'hF312E180 , 32'h10DADA80 , 32'h04B6C948 , 32'hF5DE6C70 , 32'hF8A67110 , 32'h02CD926C} , 
{32'h015E54D8 , 32'h00545C80 , 32'hFE2F3430 , 32'hFE6495A8 , 32'hFF85E47E , 32'hFDBD89E4 , 32'h0427A7B8 , 32'hFDEFCBA8 , 32'hFF91A606 , 32'hFED5E3E8 , 32'h07271C18 , 32'h07457958 , 32'hFE9D5F28 , 32'h000B9052 , 32'hFB4B0160 , 32'hFFA36DB3 , 32'hFD5B42D0 , 32'h05B22A28 , 32'hFF0F90C9 , 32'hFFCF8C26 , 32'hF6AB5560 , 32'h00E913A1 , 32'hFEFE2C5C , 32'hFD877FA8 , 32'hFDE6EF58 , 32'h035F6D28 , 32'h0122E9D4 , 32'hFE13233C , 32'hFDE607BC , 32'h02B35CB8 , 32'h02F5CA8C , 32'hFDBA2FE4 , 32'hFEDB03E4 , 32'hF9437E38 , 32'hFE87F3FC , 32'h066FA680 , 32'hF430E650} , 
{32'h00026075 , 32'h00047CCB , 32'hFFFF7ADE , 32'hFFFFE517 , 32'hFFFD9B74 , 32'hFFFFF39D , 32'h000137B4 , 32'h00051451 , 32'h0003405F , 32'h0000FCC5 , 32'hFFFEFAFA , 32'h000169E0 , 32'hFFFDC68C , 32'h00011D98 , 32'hFFFDE0AD , 32'hFFFE3576 , 32'h000073C9 , 32'h00026BC7 , 32'h000294E5 , 32'hFFF88DC0 , 32'hFFFFF1A4 , 32'h0001DE4F , 32'hFFF72855 , 32'h000103D7 , 32'hFFFCFEC3 , 32'hFFFE9D20 , 32'h0003975C , 32'h00022C9C , 32'h0001C7B6 , 32'hFFFE45CB , 32'hFFFACE10 , 32'h0002FDF2 , 32'hFFFC740C , 32'hFFFCA5AE , 32'h0000AD86 , 32'h0002C021 , 32'h00024A4C} , 
{32'h0000A046 , 32'hFFFFCDF0 , 32'hFFFED0A6 , 32'hFFFFB6C6 , 32'hFFFE0F2C , 32'hFFF8B8C5 , 32'h0007CB3E , 32'hFFFE5D34 , 32'hFFFEA5F1 , 32'h0002CC4C , 32'h00001162 , 32'hFFFFFF67 , 32'hFFFBB4D7 , 32'h0001B075 , 32'h0004EE34 , 32'h000269E8 , 32'h0003A5D2 , 32'h0002C9A5 , 32'hFFFE506D , 32'h00036296 , 32'h0000E2E5 , 32'hFFFC71B2 , 32'hFFF855A1 , 32'h00015601 , 32'hFFFBCF5E , 32'hFFFF4D31 , 32'h00019212 , 32'hFFFE23D9 , 32'h0006CAED , 32'h0003A5CC , 32'hFFFD35E8 , 32'h0001A286 , 32'hFFFBDE97 , 32'hFFFF291A , 32'h00059641 , 32'h000417B5 , 32'hFFFDE0A9} , 
{32'hFFFAB749 , 32'h0000C0C5 , 32'h0003983B , 32'h00048227 , 32'h0001F713 , 32'hFFFE1734 , 32'hFFFF4082 , 32'h00025130 , 32'h000749FC , 32'h00010972 , 32'hFFFF4CD7 , 32'h0001C49B , 32'hFFFE5431 , 32'hFFFEED19 , 32'h000161A1 , 32'hFFFDBC37 , 32'h0001E3C7 , 32'h00021E12 , 32'h0007B3D2 , 32'hFFFE89AD , 32'hFFFF1C9E , 32'h0003FCE0 , 32'h0002FA31 , 32'hFFF95BFE , 32'hFFFFC625 , 32'hFFFDFEB6 , 32'hFFFBC283 , 32'hFFFF2C94 , 32'hFFFF2385 , 32'hFFF9D52B , 32'h00052951 , 32'hFFF8983A , 32'h00042D7E , 32'h0001D76B , 32'h00064E20 , 32'hFFFFAAE6 , 32'hFFFCE1E4} , 
{32'h0005348B , 32'hFFFE080E , 32'h00015372 , 32'h00012FFA , 32'hFFFE0E10 , 32'h00004DCA , 32'hFFFE07CC , 32'h00015BC1 , 32'hFFFE1C3F , 32'h0002F809 , 32'h000684DB , 32'h00025C4B , 32'h00024161 , 32'hFFFE810A , 32'h0000C72C , 32'hFFFDEA29 , 32'hFFFEE7C5 , 32'hFFFE3821 , 32'h000481DC , 32'h0008FA1A , 32'h0009099D , 32'hFFF92D8A , 32'h000373D3 , 32'hFFFEE79A , 32'h0003BA37 , 32'h0001F935 , 32'hFFFBCEF6 , 32'hFFFB4C4F , 32'h00066E91 , 32'h000077BF , 32'hFFFFAF30 , 32'hFFFDD8C7 , 32'h00004D1C , 32'h00036BA1 , 32'hFFFE489A , 32'h0000E23D , 32'h00030A74} , 
{32'hFFFBDEE4 , 32'hFFFC4A11 , 32'hFFFF61A3 , 32'h00004ECF , 32'hFFFB2E62 , 32'hFFFF5BFE , 32'hFFFA35BF , 32'h0000EB16 , 32'hFFFEEC4D , 32'hFFFC0E82 , 32'h0000F9A9 , 32'h000204CA , 32'hFFFF6319 , 32'hFFF90A03 , 32'h00034F3E , 32'h0000DA72 , 32'h00024A18 , 32'hFFFDCC17 , 32'hFFFE63CB , 32'hFFFD3D3D , 32'h0004263D , 32'h0002002B , 32'hFFFD3493 , 32'h00007D25 , 32'h00039453 , 32'h0003A729 , 32'hFFFD54A7 , 32'h0000C8D1 , 32'hFFFD9068 , 32'hFFFD8832 , 32'h00007DEF , 32'hFFFEDF4F , 32'h00009ADF , 32'h000475B8 , 32'hFFFE08EA , 32'hFFFCC5B4 , 32'hFFFEBEE4} , 
{32'h0000A51E , 32'hFFFD14DA , 32'h00007BB4 , 32'hFFFAAE9F , 32'h0006305E , 32'hFFF42BCB , 32'h0002CF84 , 32'hFFFCF053 , 32'h000190BB , 32'h0003B54F , 32'hFFFF58B3 , 32'hFFFB5DD0 , 32'hFFFE14F4 , 32'hFFF75D25 , 32'h0001D50A , 32'hFFF95665 , 32'hFFFBAD10 , 32'h0005DC51 , 32'hFFFF8133 , 32'h0002D874 , 32'h0001E457 , 32'h00025BA9 , 32'h0000B652 , 32'h0006A1BB , 32'hFFFFAD3D , 32'hFFFE05A8 , 32'hFFFCC23F , 32'h00085B57 , 32'h0002A342 , 32'hFFFAD19E , 32'h0008DE76 , 32'h00022944 , 32'h0002862C , 32'h000153FB , 32'h0005CB96 , 32'h000474D8 , 32'h00055E25} , 
{32'h002FE18E , 32'hFFA78F43 , 32'hFFFEA13C , 32'h0007A7B9 , 32'h003B24A9 , 32'hFFF5D81D , 32'hFFDF11B4 , 32'h00276B06 , 32'hFFCDB138 , 32'hFFA9E261 , 32'hFFF44D01 , 32'h003FC9E9 , 32'hFFFE1F2E , 32'hFFD8351D , 32'hFFF1337C , 32'hFFD859F8 , 32'h006D712A , 32'hFFD83788 , 32'hFFBB8D66 , 32'h0017EC80 , 32'hFFD56533 , 32'hFFF2CCF3 , 32'hFFF537F4 , 32'h00487546 , 32'hFFD76D24 , 32'hFFB65F60 , 32'h00040C51 , 32'hFFF61670 , 32'h001EC161 , 32'h004C3CDC , 32'hFFF528EC , 32'h001345AC , 32'h00405BD4 , 32'h000559B7 , 32'h002BCF7F , 32'hFFEFB0D1 , 32'hFFD3003C} , 
{32'h089E5CA0 , 32'h0B7FD090 , 32'h086321B0 , 32'h05AEF190 , 32'h0C11D9F0 , 32'hFF928125 , 32'hF61E0D60 , 32'h0329B830 , 32'hFEA1F024 , 32'hFB92A9A8 , 32'hFC821E14 , 32'h0504E7A0 , 32'hFA9DC508 , 32'h08B508B0 , 32'h0167C6B0 , 32'h03AA7654 , 32'h0480F028 , 32'hEDE9DF60 , 32'h00701EDD , 32'h0A4C2A50 , 32'hF85F3B98 , 32'hFA2D8A58 , 32'h029B5648 , 32'h05A5E918 , 32'h02AB0B08 , 32'h07E73E18 , 32'h06348D38 , 32'h0F72F240 , 32'h0C3B7CE0 , 32'hF2278A60 , 32'hFB7A90D8 , 32'hFDCBCDA0 , 32'h078A1CB0 , 32'h0401C8C0 , 32'h0283FF88 , 32'hFB04F790 , 32'hF88A6170} , 
{32'h0529A320 , 32'h042F5678 , 32'hFF85D841 , 32'hFA260858 , 32'h01078F7C , 32'hFC053B30 , 32'h005B3498 , 32'h06382810 , 32'h0036EC0F , 32'hFAC8D568 , 32'h0563C6E0 , 32'hFAFC15E0 , 32'h0421A820 , 32'hFF239DB8 , 32'hF9A4BF58 , 32'hFFA770EF , 32'hFBBE2B80 , 32'hF9B28308 , 32'hFBED76B8 , 32'hFCF00760 , 32'h008766D2 , 32'hFDE02A80 , 32'h01E7AB18 , 32'h00DE1021 , 32'hFCB6C000 , 32'h03251934 , 32'h02C67E30 , 32'h077C1B00 , 32'h0F7FC660 , 32'hF59898D0 , 32'h0661C688 , 32'hF8095EB0 , 32'h035E1DB8 , 32'h012B5B30 , 32'hFD2239F0 , 32'h012ACEC8 , 32'hFF333645} , 
{32'h0FC51270 , 32'h0D1DF980 , 32'h03901F64 , 32'hFCF147F8 , 32'hFC928CD8 , 32'h0BE28DA0 , 32'hFF073757 , 32'h056A01D8 , 32'h0BEE5F50 , 32'hEEEE2C20 , 32'h04511278 , 32'h0D28C400 , 32'hFB8E1B88 , 32'hFFE8334D , 32'hF194DFA0 , 32'h13447CA0 , 32'h0F2428F0 , 32'hF15FF980 , 32'hF8D2F8A8 , 32'h0ACC9EF0 , 32'hFDEE9C88 , 32'h24F93F80 , 32'h02080844 , 32'h03F27E14 , 32'hFFAC5186 , 32'hF69D0BF0 , 32'hFD6D2438 , 32'h0C1C2910 , 32'hFFB9E0F0 , 32'h033505EC , 32'h005E0EE6 , 32'hEF6028E0 , 32'h0C82BAA0 , 32'hFFE189FB , 32'h09BAFD50 , 32'h07D95810 , 32'h04D5FCA8} , 
{32'h02FC41A8 , 32'h05B172F0 , 32'hFA742F18 , 32'hF94DF8C0 , 32'hF854BCA0 , 32'h15323640 , 32'h0047781D , 32'h042C1248 , 32'h090865D0 , 32'hEFB36C20 , 32'hF4A5C310 , 32'hF9950300 , 32'h0B01FE00 , 32'h045E5A88 , 32'hFF7A4DA0 , 32'hF8BC9590 , 32'hFEB037D4 , 32'hFE059040 , 32'hFA98EEE0 , 32'h09C3AA70 , 32'h0C2805D0 , 32'hFF5DB969 , 32'hEC4D5FE0 , 32'h0B8A5420 , 32'h045EE198 , 32'h01A000C8 , 32'hF932F078 , 32'h052F4C80 , 32'h067D36A0 , 32'hFD72F894 , 32'h039D231C , 32'h010DCC80 , 32'h00E47158 , 32'hFDC117A0 , 32'h0458E1C8 , 32'hFCC95218 , 32'hFEB19ED0} , 
{32'h0C1D0500 , 32'hFB4A02E8 , 32'hF74965A0 , 32'hFC3F6AA8 , 32'hFB76E9A0 , 32'h1E244E00 , 32'hF386B440 , 32'h0200714C , 32'h078B1AC0 , 32'hFFB29CCC , 32'h074C8290 , 32'h03227AF0 , 32'hFF9AA76C , 32'h01960F3C , 32'hFB928B10 , 32'h05069948 , 32'hF699A930 , 32'hFC26F158 , 32'hF7EB53B0 , 32'h089DD320 , 32'h006B9337 , 32'hFBA19000 , 32'hFBB3E000 , 32'hF259FA30 , 32'hF409DF90 , 32'hFAC670A8 , 32'hF892F400 , 32'hFCA6F8CC , 32'h048BE388 , 32'h063C8B10 , 32'h0907DFE0 , 32'hFB0B58C8 , 32'hF45D2C50 , 32'h025FEA98 , 32'h06A30BC8 , 32'h05580380 , 32'h039401D4} , 
{32'h31ECC780 , 32'hED7B0EC0 , 32'hF2CBD270 , 32'hF19BA6F0 , 32'hE27A45A0 , 32'h31C23840 , 32'hF30AD0B0 , 32'h1F808B60 , 32'hFB896830 , 32'hFAF14068 , 32'h2028A1C0 , 32'h07D0BC38 , 32'hF45F6020 , 32'hF87C7738 , 32'h2308C080 , 32'h102C56C0 , 32'hE3B8F300 , 32'h0261BF2C , 32'hE7CDB320 , 32'h2027F980 , 32'h062FDCB8 , 32'h1C566660 , 32'hF3D4DF70 , 32'h0A85E0D0 , 32'h02D89D40 , 32'h03420C2C , 32'hE11EE0A0 , 32'hF7B3FDF0 , 32'h20850C40 , 32'hFF8A119D , 32'h1D779300 , 32'hE46CF440 , 32'h02997C68 , 32'h11F79640 , 32'hE4EBCA20 , 32'hF5DE3950 , 32'h098AD9E0} , 
{32'h1CDFB200 , 32'hFA32F278 , 32'hEA598460 , 32'hFB825FE8 , 32'hF56F15A0 , 32'h21D86800 , 32'hE6B87D00 , 32'h07985FD8 , 32'hEB0CB140 , 32'h2248DEC0 , 32'h094B7750 , 32'hFC5E9780 , 32'hFEFCE1EC , 32'hFE757F4C , 32'h15655300 , 32'h261D91C0 , 32'hE132E3E0 , 32'h0FA33B40 , 32'hF2478800 , 32'hFA93E3D0 , 32'h0098B67C , 32'h090EF560 , 32'hF011F5F0 , 32'hF6A42AD0 , 32'hF8E98F20 , 32'h2C0142C0 , 32'h0987ACF0 , 32'h0D0A92F0 , 32'h0CD334A0 , 32'hF8063378 , 32'h122413E0 , 32'h10459BC0 , 32'hFE1BCCD4 , 32'hF7441E20 , 32'hE8D24E80 , 32'hFED2BC68 , 32'h10590540} , 
{32'h393A00C0 , 32'hFFE2A1B3 , 32'hFC39C830 , 32'hFD7778A8 , 32'hFACFDCE8 , 32'h1DBE2DC0 , 32'hDACD2F00 , 32'h1C566D20 , 32'hD575EF00 , 32'h1FC91BC0 , 32'hF653DC90 , 32'hF65D5BE0 , 32'hF7D60A50 , 32'hFDD6CC58 , 32'h251E3A40 , 32'h05B84698 , 32'hFABCFE70 , 32'h0B30C990 , 32'hF6DBAE10 , 32'hE4874C20 , 32'hF2D41280 , 32'h15DEBBE0 , 32'h07AC0800 , 32'h2F835680 , 32'hF1B79CF0 , 32'hFD62F150 , 32'h27463C40 , 32'hF653BA10 , 32'h1F101620 , 32'h1DEA8560 , 32'h04F54F58 , 32'h0163D718 , 32'h03817B78 , 32'h03001060 , 32'hFB78A840 , 32'hE7BE3B60 , 32'h36550D40} , 
{32'h4F3FDC00 , 32'hD85B0640 , 32'h0E1BD340 , 32'hFE13E740 , 32'hFF3F846B , 32'hF7A038B0 , 32'hEC1A5B80 , 32'h21FBF380 , 32'hBC7B7380 , 32'hF7BFDBA0 , 32'h0E87E3B0 , 32'hF5E9AA70 , 32'hF0F5A1B0 , 32'hEE9DB100 , 32'h0FFDFB60 , 32'hFF49FF97 , 32'h11C04580 , 32'h12C182A0 , 32'h16A2FFC0 , 32'hEF55C9E0 , 32'h128A1100 , 32'h0F5CA240 , 32'h049F8E80 , 32'h14C068A0 , 32'h1251F3C0 , 32'h093F4230 , 32'h07E0F198 , 32'h13BD2F40 , 32'hFFE40232 , 32'hFF6D9577 , 32'h1422CFE0 , 32'h1CF27020 , 32'h036255F8 , 32'hF695E7D0 , 32'hFC45C24C , 32'h000A719E , 32'h07D2C380} , 
{32'h52E2DA00 , 32'hD68ACA00 , 32'h22573D40 , 32'hFF78C719 , 32'h07509598 , 32'hD79A2FC0 , 32'hF0C5F120 , 32'h180749A0 , 32'hD5A18A40 , 32'hD6833240 , 32'h0607A928 , 32'h03C18F1C , 32'h11E749E0 , 32'hF289C610 , 32'h13400440 , 32'h0FA862E0 , 32'h0E8ABFC0 , 32'h14189840 , 32'h03409BE8 , 32'h09494EB0 , 32'h18D25780 , 32'hE14A1660 , 32'hEE0C4F60 , 32'h0180E294 , 32'h09622E80 , 32'h16321320 , 32'hFBFDE070 , 32'h25C189C0 , 32'hF2BE3E10 , 32'h0E224710 , 32'hFC09DB08 , 32'hFD05F580 , 32'h15FD4480 , 32'hEE92AFC0 , 32'h0BF2CDB0 , 32'hF8764FF8 , 32'hFCE7ECA4} , 
{32'h2A841A80 , 32'hDD680740 , 32'h09B59470 , 32'hF4AC64C0 , 32'h08EA84C0 , 32'hF8461FB0 , 32'h1260BC40 , 32'hF8385760 , 32'h02A99A90 , 32'hBEAAB600 , 32'hF2644C60 , 32'h058D0C00 , 32'h02AE331C , 32'h00345E12 , 32'hFE86023C , 32'h0DCF0830 , 32'hFD8D28F0 , 32'h0ABDA990 , 32'h1656C380 , 32'h15940B20 , 32'h0726E4B0 , 32'hDFF1E680 , 32'hF29589C0 , 32'h0C6F4120 , 32'h11E09940 , 32'h0E6BDE30 , 32'hFDEECFDC , 32'h04F6F1C0 , 32'hEEDBB880 , 32'hFBA42B90 , 32'hF96FB4B8 , 32'h11684BC0 , 32'hFC95A7AC , 32'hEB03F7E0 , 32'hDEE0EF40 , 32'hFD55D084 , 32'hF451E490} , 
{32'h3B74FD00 , 32'hD0A44700 , 32'h214A0DC0 , 32'hCC977C00 , 32'h0ADBB840 , 32'h02E3D7A0 , 32'h14B330A0 , 32'hDA2DC180 , 32'h2BFDCF80 , 32'hCCBF5540 , 32'hEC472D40 , 32'hEF6CB480 , 32'h03A59568 , 32'hF33D65B0 , 32'hE9142760 , 32'h110E65E0 , 32'h0815E2F0 , 32'h083D3E80 , 32'h2E9FC480 , 32'h00273763 , 32'h23AEE500 , 32'hD3CD83C0 , 32'h0F6C8080 , 32'hFF72ACAF , 32'h06FFBB58 , 32'h21CB3000 , 32'h156F3F80 , 32'h06AF9698 , 32'h05F97C80 , 32'h0B1ACCA0 , 32'h1791A320 , 32'h0862D190 , 32'hF14FECC0 , 32'hFD8BD198 , 32'hFD760534 , 32'hFF517094 , 32'h06FADD50} , 
{32'h58B97F80 , 32'hB8D7C200 , 32'h334EC200 , 32'hD0701A80 , 32'h092B78B0 , 32'hE58AC800 , 32'h02DE171C , 32'hCE7FA540 , 32'h2F44AC80 , 32'hDEC6D840 , 32'hF1BD0370 , 32'hF42341F0 , 32'hF4F29240 , 32'hF16E8950 , 32'hFCEF29E0 , 32'h096297A0 , 32'h167DB2C0 , 32'hF53CED90 , 32'h12DD3820 , 32'hF1FEB030 , 32'hF85C5DF8 , 32'hD4C8EE80 , 32'h08758490 , 32'h080D4CC0 , 32'hF383F960 , 32'h07D5B4D0 , 32'h0BA0BD90 , 32'hDD2D59C0 , 32'h18B19DA0 , 32'h07A911A8 , 32'h0353909C , 32'hF598A9E0 , 32'hE86CC640 , 32'h00E60C95 , 32'hF032CAF0 , 32'h063CBA58 , 32'h09E8D230} , 
{32'h3E61E9C0 , 32'hD543A840 , 32'h22BD0B00 , 32'hD4187C80 , 32'h0902D920 , 32'hE33DC6A0 , 32'hFE402C14 , 32'hE8042C20 , 32'h25609D00 , 32'h0E5D4070 , 32'h05FAE6D0 , 32'hF9F57738 , 32'hEB980820 , 32'hFEE8AE70 , 32'hF7D17350 , 32'h00E87982 , 32'h1ECC5EA0 , 32'hFCFDCA50 , 32'h1C9FDA00 , 32'hF75DE2E0 , 32'h0B8F6D20 , 32'h0114A828 , 32'h08F78B70 , 32'hF2EEFE90 , 32'h04168020 , 32'h009C0482 , 32'hFE0DF650 , 32'hF310AE10 , 32'h05007C48 , 32'h135C72A0 , 32'hF900E6F0 , 32'hE71DF8E0 , 32'hFDA357F4 , 32'h17636020 , 32'hF9A8DDE8 , 32'hF29A8B50 , 32'h1CB5A6A0} , 
{32'h4126F000 , 32'hC7C2A440 , 32'h28A43780 , 32'hCC132C40 , 32'h0F8121B0 , 32'hE27F3180 , 32'hF7B9CAE0 , 32'hF648D440 , 32'h36B193C0 , 32'h27BA1A80 , 32'h0C370AA0 , 32'hF51C14B0 , 32'hF81D8C60 , 32'h1BB60A80 , 32'h03D1F270 , 32'hD2EA8B80 , 32'h1204D3C0 , 32'h0E0087F0 , 32'hF8D78D60 , 32'h1C6B4100 , 32'h1902F740 , 32'h1D7BD040 , 32'hE4756420 , 32'hFD6A32C4 , 32'hEDFAD440 , 32'hFAFB1890 , 32'hFC8065CC , 32'h09D0C170 , 32'hF56E5E60 , 32'hF6767770 , 32'hEE2DB320 , 32'h00DFD2DB , 32'hF44F8C20 , 32'hF432B390 , 32'h11E907E0 , 32'hFE8F63DC , 32'hFC532CE4} , 
{32'h45799E80 , 32'hDB3B0600 , 32'h177D6FC0 , 32'hE0C41460 , 32'h056D74D8 , 32'hE42086E0 , 32'h05542598 , 32'hEB99E4E0 , 32'h1C155000 , 32'h3067E200 , 32'h161D0760 , 32'hF4837E10 , 32'h08E45650 , 32'h2E231FC0 , 32'h0327B3D4 , 32'hD5DB9E40 , 32'h0BFF9F90 , 32'hFC52336C , 32'hEBFE8FC0 , 32'h19066F20 , 32'hFF22E066 , 32'h23CD3800 , 32'hEE1CAF20 , 32'h09EB44A0 , 32'hFCFAA758 , 32'hEFF67340 , 32'h00908E30 , 32'hF4B31820 , 32'h0BD572B0 , 32'hFD486DDC , 32'h10ED41E0 , 32'h08457870 , 32'h01FC1D94 , 32'h08C27510 , 32'h11C9CC40 , 32'hFC875A78 , 32'hF6D19550} , 
{32'h45072B80 , 32'hD98028C0 , 32'h18C1F4C0 , 32'hE8A44B80 , 32'hFF462414 , 32'hE3266C80 , 32'h0ADA9570 , 32'hF9334DE8 , 32'h1ADA9580 , 32'hFB46E4B0 , 32'h0205756C , 32'h0115F100 , 32'h0A99F770 , 32'h24915600 , 32'h0D5038E0 , 32'hF5D37940 , 32'h132512C0 , 32'hFBB1CCB8 , 32'hFFAFFF98 , 32'h1002AAA0 , 32'h0122D6E8 , 32'h10D03640 , 32'hFF2110F6 , 32'hF95139D8 , 32'h10BCE3C0 , 32'h07F63140 , 32'h04AB2618 , 32'hEB414CC0 , 32'hF8ACC978 , 32'h0A3F6850 , 32'h07E1F808 , 32'hFAAFDD08 , 32'h038ED9B4 , 32'h06E5D038 , 32'h024244EC , 32'hFD618F74 , 32'h0B04F460} , 
{32'h2D880100 , 32'hDEE3DE40 , 32'h123DC2C0 , 32'hEB7711E0 , 32'hFB18D148 , 32'hF0F02D70 , 32'hF9A2E810 , 32'h03577F3C , 32'h18EB0B20 , 32'h00223820 , 32'hF69068B0 , 32'h035639E0 , 32'h067B0270 , 32'h1545CDA0 , 32'h0D2EFB50 , 32'h0D216CC0 , 32'h0D45B190 , 32'h064C5248 , 32'h0194BBEC , 32'h03582514 , 32'h00324F71 , 32'h0642FF60 , 32'h001423D1 , 32'hF77C1FB0 , 32'h0C6B5D90 , 32'h12A6D880 , 32'h0E087770 , 32'hFB3DF560 , 32'hEB5200C0 , 32'h069326D8 , 32'h01B53AD8 , 32'h056C2E58 , 32'hFEABC3B4 , 32'hF76EB890 , 32'hEF8E43E0 , 32'h0EF5A4C0 , 32'hF739AA20} , 
{32'h19DAFA20 , 32'hF44EB9C0 , 32'hFE02BFD4 , 32'hFE824CBC , 32'hF95C6630 , 32'hEA504440 , 32'h063EF980 , 32'h108D17A0 , 32'h098FCAE0 , 32'h0BE2C4A0 , 32'h120AEA80 , 32'h17CC3780 , 32'h11D9D2C0 , 32'h1AF16B00 , 32'h0624D1B0 , 32'hF47A1A20 , 32'hF1D28C00 , 32'h15E90200 , 32'hDD4318C0 , 32'h01B8536C , 32'hE004D7A0 , 32'h0E87FD70 , 32'hF7FC7940 , 32'hF57BFF40 , 32'h00D8722D , 32'h00D46890 , 32'h08C26650 , 32'hF791DA30 , 32'h0BEA32B0 , 32'h03308394 , 32'hFE96F9C8 , 32'hF994BBA0 , 32'h036BA9D8 , 32'hF6AFA9F0 , 32'hF4351B00 , 32'hFE59D2F0 , 32'hED8C8320} , 
{32'h13C6C5C0 , 32'hFB38AA10 , 32'h05B47098 , 32'hF6E86E00 , 32'hFEC44140 , 32'hF3CECFF0 , 32'h05EBD8F0 , 32'hF1A86600 , 32'hF5406DA0 , 32'hFFC86765 , 32'h12611120 , 32'h144776E0 , 32'hFE5E257C , 32'hF594F4A0 , 32'hF9EAE678 , 32'hF5F7C740 , 32'hF844A6B8 , 32'h0D9CE5F0 , 32'hE92A1FE0 , 32'h069143A0 , 32'hE888ED20 , 32'hED5363E0 , 32'hF1780210 , 32'h04372C90 , 32'hEE5B3F00 , 32'hF6B3E1C0 , 32'h03242788 , 32'h14B662C0 , 32'h060F4188 , 32'h094ACBA0 , 32'hF7359C00 , 32'hF247BBD0 , 32'h08FE18D0 , 32'hE20857E0 , 32'h01025784 , 32'hFF6C6A97 , 32'hF61A01E0} , 
{32'h00014627 , 32'h000251A9 , 32'hFFFD35CD , 32'h00006290 , 32'hFFFFA2AC , 32'hFFFF0555 , 32'h00013574 , 32'hFFFD129B , 32'h0000AAC8 , 32'hFFFC350F , 32'hFFFEAFD9 , 32'hFFFEF5BC , 32'hFFFDDC9C , 32'h00001A56 , 32'hFFFFDCA6 , 32'hFFF9EC0C , 32'h000294E8 , 32'hFFFFAD12 , 32'h0004E785 , 32'h0000DEDE , 32'hFFFFAD7B , 32'hFFFFEE57 , 32'h00038DF5 , 32'h0002E78A , 32'h0001C867 , 32'hFFFD13B4 , 32'hFFFB45B5 , 32'hFFFF327B , 32'hFFFCA3D6 , 32'h0003D8A7 , 32'h000210FA , 32'h00001124 , 32'hFFFE2F95 , 32'hFFFF7E85 , 32'h000174BE , 32'h0001F093 , 32'h000006C8} , 
{32'h00008038 , 32'hFFFBB357 , 32'h00022CFD , 32'h00015CD6 , 32'hFFFF1A3A , 32'hFFFE658F , 32'hFFF4BB2A , 32'h000090FE , 32'h00062C4F , 32'hFFFE725E , 32'h0001849B , 32'hFFFD1E6A , 32'hFFFFA5B1 , 32'h000311D4 , 32'h0000D7AE , 32'hFFFD329E , 32'hFFFB1643 , 32'h000186B9 , 32'hFFFDB283 , 32'hFFFBB75D , 32'hFFFE48CF , 32'hFFFF4524 , 32'hFFFED7C5 , 32'h0003BFFC , 32'h000264A4 , 32'hFFFE7D61 , 32'hFFFCD69A , 32'h000199AF , 32'h00002F9C , 32'hFFF9B3A9 , 32'h0001D6C4 , 32'hFFFF1714 , 32'h00030400 , 32'hFFF569E4 , 32'h000122EB , 32'hFFFD445E , 32'hFFFE7FA5} , 
{32'hFFFD1BD5 , 32'h0002C32D , 32'hFFFE1D71 , 32'h00013FF9 , 32'h0001A0AD , 32'h00002185 , 32'h0000ECA2 , 32'hFFFF3BDE , 32'h0002252D , 32'hFFFF491F , 32'hFFFF5400 , 32'h00014964 , 32'h0000BA4A , 32'hFFFEF00C , 32'h000146F1 , 32'h00047B5D , 32'h0003E0BF , 32'hFFFE1704 , 32'hFFFED5C4 , 32'h0000D827 , 32'h0005812A , 32'hFFFFCB58 , 32'h00005C19 , 32'hFFFE40FA , 32'h00055A19 , 32'hFFFFED9F , 32'h0000EC59 , 32'h00003C86 , 32'hFFFD5326 , 32'h00017F72 , 32'h0000086F , 32'h000295AE , 32'h00031D74 , 32'h0001032D , 32'h0001919C , 32'h00027F68 , 32'hFFFC1D23} , 
{32'hFFFF2860 , 32'hFFFF82CA , 32'hFFFD6D5E , 32'hFFFD55D5 , 32'h0005DE6B , 32'hFFF95734 , 32'hFFFCB686 , 32'h0003B221 , 32'hFFFA6495 , 32'hFFFE978E , 32'h0001889B , 32'h000093C5 , 32'h0001CA22 , 32'h0003D66E , 32'h00008FF9 , 32'h0003AC5B , 32'hFFFC5B19 , 32'h0000C80E , 32'h00004FF0 , 32'h0000580A , 32'h0000008C , 32'h0000902B , 32'hFFFE37C8 , 32'h0000DB60 , 32'h000167B1 , 32'h00027594 , 32'hFFFD3EDE , 32'h0003619F , 32'h000007B3 , 32'hFFFF434C , 32'hFFFEB7A4 , 32'hFFFC4247 , 32'h000458F2 , 32'h0002BE61 , 32'hFFFFA8D0 , 32'hFFFAFCCA , 32'hFFFD9847} , 
{32'h0002B11C , 32'hFFFB4573 , 32'h00046399 , 32'h0004829E , 32'hFFFEC439 , 32'hFFFE529B , 32'h00009D89 , 32'h00054F4B , 32'hFFFFB569 , 32'hFFFC5A39 , 32'h000276E8 , 32'h00029A0C , 32'hFFFD57C1 , 32'hFFFD3646 , 32'hFFFF96D1 , 32'hFFFC059B , 32'h000145B0 , 32'hFFFED091 , 32'h0000C552 , 32'hFFFE840A , 32'h0004C226 , 32'h00031DD6 , 32'h000067B8 , 32'hFFFE2D65 , 32'h00063B99 , 32'h000055AF , 32'h000402E7 , 32'h00004BCB , 32'h000554E2 , 32'hFFFE5EA2 , 32'h0004EE8F , 32'hFFFD93EB , 32'h0004C0C0 , 32'h0002B8EE , 32'h0000EF5F , 32'h00039E85 , 32'hFFFCFC11} , 
{32'h0001084F , 32'hFFFFE504 , 32'hFFFBC19D , 32'hFFFC8C66 , 32'h0001CCE1 , 32'h0003E4A7 , 32'h00019134 , 32'h00019A4A , 32'hFFFE5351 , 32'hFFFB0163 , 32'h00082F61 , 32'h00002C0E , 32'h00006870 , 32'h000210ED , 32'hFFF86DF0 , 32'hFFFABB96 , 32'hFFFAD875 , 32'h000113A8 , 32'hFFFBAB83 , 32'h00040CAE , 32'hFFFAEF74 , 32'h000794CD , 32'h0000E2EA , 32'h00056D4A , 32'hFFFEFC01 , 32'h0001973F , 32'hFFFF445C , 32'h0001ACE5 , 32'h0001453D , 32'hFFFEB3D6 , 32'h000216FF , 32'h00015140 , 32'hFFFD9DF3 , 32'h0003EC8C , 32'hFFFDEDE2 , 32'h0003992C , 32'h00052F13} , 
{32'h00009800 , 32'h000185BD , 32'hFFFD8043 , 32'h000858B5 , 32'h0001606F , 32'hFFF9D608 , 32'h0002087C , 32'h0005BA9F , 32'hFFFD5A2F , 32'hFFFA8F89 , 32'hFFFBDA0E , 32'hFFFE5276 , 32'h0004117E , 32'hFFFE4F68 , 32'hFFFF4B40 , 32'h0002B0C2 , 32'hFFF8E0C3 , 32'h00027077 , 32'h0005C856 , 32'hFFF8F0DD , 32'hFFFDFABC , 32'h000331C8 , 32'hFFFF5707 , 32'hFFF9C761 , 32'hFFFDE8AA , 32'h0005E367 , 32'hFFFFC8E6 , 32'hFFF948D3 , 32'hFFFC412C , 32'h00063462 , 32'h0003E22B , 32'hFFFBB1AF , 32'hFFFC086F , 32'h0003AEDB , 32'hFFFDD989 , 32'h0005459F , 32'hFFFB4439} , 
{32'h012C0848 , 32'hFF574C95 , 32'hFFC8694B , 32'hFF9E468B , 32'h004CE794 , 32'hFFAE2AC7 , 32'hFFA40900 , 32'h007AD680 , 32'hFEDAAB70 , 32'hFFDE5768 , 32'hFFB0B866 , 32'h00027E88 , 32'h001CBE78 , 32'hFF65A688 , 32'h007D5D76 , 32'hFF30641E , 32'h007DF107 , 32'hFFD6A994 , 32'hFFA4C0C5 , 32'h00848F5A , 32'hFF577E02 , 32'h00F1E7E5 , 32'hFF2144B2 , 32'h01DB6484 , 32'h00028D9B , 32'hFE71C43C , 32'h00DB4707 , 32'h00625319 , 32'h016127C4 , 32'h00B7CF66 , 32'hFFAE03E6 , 32'h00358930 , 32'h00B5D95E , 32'hFFCA4F51 , 32'hFF08D599 , 32'hFF12AF5D , 32'h0084A748} , 
{32'h086D5920 , 32'hFF5158D7 , 32'hF8E28CC8 , 32'hFF69FDE0 , 32'hFDD46EB4 , 32'h05657AA0 , 32'hFDA20940 , 32'h002A902D , 32'hF896BB60 , 32'h00D02CEF , 32'hF8E07438 , 32'hFF4D47EA , 32'h02A6C7B4 , 32'h06148560 , 32'hFF99A858 , 32'hFCCA82A8 , 32'h04400FB8 , 32'h04E00778 , 32'hFFDF2D06 , 32'hFC72F054 , 32'h0474BBC8 , 32'hFF94B7F7 , 32'hFE909644 , 32'hFFC1E8BA , 32'h01ACE6A0 , 32'h01C68740 , 32'h09D49E10 , 32'h027E0E94 , 32'h065876E8 , 32'hFBCAE9C0 , 32'hF992DF58 , 32'h036B6F1C , 32'h03460FD8 , 32'hFEFC25DC , 32'hFFC878EF , 32'h0249494C , 32'h054C5920} , 
{32'h44BA5E00 , 32'hF7D9D260 , 32'hE6AC74C0 , 32'h08306030 , 32'hF2D746B0 , 32'h18599FC0 , 32'hF11D0F30 , 32'hFF57DC4A , 32'hE92D6680 , 32'h03A4E2EC , 32'h040D4CC8 , 32'h07890BF0 , 32'hF577F290 , 32'h19E376E0 , 32'hF7DA6D60 , 32'hE2A48760 , 32'h0E703750 , 32'hFA1B9050 , 32'h07616B18 , 32'h0706F758 , 32'hEEEE0AA0 , 32'h0E31E670 , 32'h19ED94E0 , 32'h115EF8C0 , 32'h032E96EC , 32'hF0271F50 , 32'hECDF9F40 , 32'hE29BBD60 , 32'hF9A7C808 , 32'hF4752FD0 , 32'hF0A3F360 , 32'hEEF16E60 , 32'hFD745ADC , 32'h0F207330 , 32'hEED8C6C0 , 32'h08567370 , 32'hF0ECF500} , 
{32'h17992880 , 32'hF207E670 , 32'hF31F2D80 , 32'hFFCE9C78 , 32'hF4D27910 , 32'h1E1FBBA0 , 32'hEF7EFCA0 , 32'h06C5E8F8 , 32'hE591B960 , 32'hFF0222E1 , 32'h0E27CA80 , 32'hFC944114 , 32'hEFFBF4A0 , 32'h012D7578 , 32'hF6D50050 , 32'hF3EAACE0 , 32'hFA655870 , 32'h00930B36 , 32'hFE5CD8A4 , 32'h0F00B460 , 32'h053791D0 , 32'h031B7470 , 32'h0EAD19A0 , 32'hF97037E8 , 32'hFD6A5A60 , 32'hF9B7B6F0 , 32'hEE89A380 , 32'hFD3E2318 , 32'h034297F4 , 32'h029ACF5C , 32'h0DFC6A20 , 32'hFCFDF15C , 32'hEB580D80 , 32'h00100D8F , 32'hFA807358 , 32'h05B9E138 , 32'hFC3DAB30} , 
{32'h1C8DE780 , 32'hF8DA2850 , 32'hF1224E20 , 32'hFCA1FAEC , 32'hF608B2A0 , 32'h28E66B80 , 32'hFB8A9EA8 , 32'h058E0370 , 32'hEBF00020 , 32'h0776EE20 , 32'h18803340 , 32'hF9A64F88 , 32'hEBC2F600 , 32'hFDD7E144 , 32'hF7420920 , 32'hF168CE80 , 32'hF176A7F0 , 32'hFB0100F0 , 32'h022993F4 , 32'h198CE560 , 32'hFE9B44D4 , 32'h04E4BAB8 , 32'h104E0340 , 32'hF02AF100 , 32'h08D1A630 , 32'hF504E0D0 , 32'hF5E46780 , 32'h028A7DD4 , 32'hF8F51630 , 32'hFE506F4C , 32'h0B250410 , 32'hF8A06070 , 32'hDD979240 , 32'h09662F60 , 32'hEE9B6D80 , 32'h04303858 , 32'hFF10171D} , 
{32'h3F634C40 , 32'hEA464640 , 32'hE79E8100 , 32'h046F1190 , 32'hF23416B0 , 32'h4E3CA980 , 32'h0442FA80 , 32'h0CC061B0 , 32'hF691AA80 , 32'hEBEDCA20 , 32'h2BC5A540 , 32'hFAD0A288 , 32'hDCC18840 , 32'hF59BFEC0 , 32'h05180310 , 32'h05C13378 , 32'hEFFBA4E0 , 32'h0229D634 , 32'hF813ACE8 , 32'h17566640 , 32'h00430955 , 32'hF13FF3B0 , 32'h144FB5A0 , 32'h01907FEC , 32'h02045AB8 , 32'hEE1F2A40 , 32'hF3F54DD0 , 32'hFB08F598 , 32'hFE0CA454 , 32'hF37CEC60 , 32'hFF8E394B , 32'h0283DE1C , 32'hF04C7C10 , 32'h13A88FA0 , 32'h042A29F8 , 32'h0E8FD480 , 32'hF30A1080} , 
{32'h43C85E00 , 32'hF6E28460 , 32'hE3123060 , 32'hF800D158 , 32'hF098AF50 , 32'h4690B300 , 32'hECF08520 , 32'hFB30A800 , 32'hEC486E80 , 32'h1077A260 , 32'h08CF9830 , 32'hFEB2AEC8 , 32'hF70DB600 , 32'h149E18C0 , 32'hFB671338 , 32'h1781F220 , 32'hDCF38400 , 32'hFD740EFC , 32'hF1A0FED0 , 32'h102AE320 , 32'hFB6FB1E8 , 32'hF9FA5B10 , 32'h104CF680 , 32'hE9DE67C0 , 32'h015110F4 , 32'hF6FD3450 , 32'hEF32FDA0 , 32'hFCE19520 , 32'hFBA53CE8 , 32'h18E0E280 , 32'h0D25B570 , 32'hFBD635A8 , 32'hE9B9E9E0 , 32'hEFA3D320 , 32'hF39F1E00 , 32'h13133A20 , 32'h036A8918} , 
{32'h42DF8700 , 32'h0B1D8010 , 32'hDDE1EEC0 , 32'h1F2B00C0 , 32'h07A5FC88 , 32'h44999300 , 32'hF21C4CA0 , 32'hED3941C0 , 32'hF4B22AA0 , 32'h19EF9000 , 32'hFA5336A0 , 32'hF6802D90 , 32'hF71A40C0 , 32'h1EFB6C00 , 32'h0198316C , 32'h1921CF00 , 32'hF5FD96A0 , 32'h171F4880 , 32'hED1912C0 , 32'hD7A4D580 , 32'h0A15BD10 , 32'hF7C63580 , 32'h2B078540 , 32'h02D8367C , 32'hEFE2F720 , 32'hFA4D5100 , 32'h12453000 , 32'hE89704C0 , 32'hFEC02F4C , 32'h148DFE80 , 32'h006A1D10 , 32'hFAD9F798 , 32'h13FE7CC0 , 32'hE1518360 , 32'h1AA3D540 , 32'hFFDC19FA , 32'hFB41FEA0} , 
{32'h254CA900 , 32'hEFE972E0 , 32'hE3D904E0 , 32'h08B9DD10 , 32'hF69390B0 , 32'h1C338CE0 , 32'hEE79BE00 , 32'h017BC8DC , 32'hDBE130C0 , 32'h0F2DD9D0 , 32'h061EB338 , 32'hEF1D06A0 , 32'hF9E26A40 , 32'h10411640 , 32'hF7C8FD70 , 32'h0BBDBA70 , 32'hFF2C4E8E , 32'h12F1A440 , 32'h025D7884 , 32'hE851FFA0 , 32'h060089B8 , 32'h06BBB160 , 32'h1F7F1D00 , 32'h0590F360 , 32'hE98660C0 , 32'hFFA03740 , 32'h0D825970 , 32'hFE1B7D90 , 32'h085CF340 , 32'h0B0A0270 , 32'h12C41180 , 32'h07A4B808 , 32'hF6A7DD10 , 32'h033E3244 , 32'h0C616450 , 32'hF2BBA930 , 32'h0D306590} , 
{32'h38173300 , 32'hFB828888 , 32'hFFA01E59 , 32'h3E7E3300 , 32'h22A34140 , 32'hED9ADB80 , 32'h07F90D68 , 32'hFAAB3D50 , 32'hC365A6C0 , 32'h058B7040 , 32'hE8A1F120 , 32'hEF0F41A0 , 32'hF4F54640 , 32'hFD61C474 , 32'hECE61460 , 32'h13CF8760 , 32'hFCB2FBBC , 32'h0FFC50B0 , 32'hFE3618F0 , 32'hF3DF7200 , 32'h0F2A4180 , 32'h1349B8E0 , 32'hE69C50E0 , 32'hE5E5A060 , 32'h0FB2CC50 , 32'hF1F0D560 , 32'hF967FEF0 , 32'hFD65A7D8 , 32'hEDDD09A0 , 32'h0DACE8A0 , 32'hE8A99280 , 32'h174B0320 , 32'hF2987B10 , 32'hFC013E18 , 32'h137804C0 , 32'h0A0FF3E0 , 32'h09AB5BA0} , 
{32'h1BEFD260 , 32'hD9AA0500 , 32'hECE5F560 , 32'h46230A80 , 32'hF6DB08C0 , 32'hDD78C600 , 32'h387C4A00 , 32'hFB2AF1E0 , 32'hDEAD7300 , 32'hD7979800 , 32'hFD94E2AC , 32'hCD267C40 , 32'hF193FA60 , 32'h0EB1FF20 , 32'hF4387150 , 32'h0D972C70 , 32'h0639B1F8 , 32'h058E4728 , 32'h09509E20 , 32'h10073500 , 32'h0C6CB930 , 32'h188FABE0 , 32'hD2C59600 , 32'hF9000FF8 , 32'h0727C380 , 32'hEBCF0840 , 32'h1389A020 , 32'h2525E380 , 32'hE9A92D40 , 32'hF15DC550 , 32'h1502F4A0 , 32'h02A4AFC8 , 32'h10254C60 , 32'hEC56E700 , 32'hE941AE20 , 32'h06810940 , 32'hEA88B3A0} , 
{32'h1EBA08E0 , 32'hD6074280 , 32'hF0453B90 , 32'h199381A0 , 32'hF6DDEA40 , 32'hFF172DAA , 32'h0D4BFBE0 , 32'h10A92F60 , 32'hFB0BD390 , 32'hD3B7AE40 , 32'hF0A28280 , 32'hE758EE00 , 32'h0421FEC8 , 32'hF1C9C340 , 32'hDC59E500 , 32'h35B672C0 , 32'hE84B2B20 , 32'hF56B28C0 , 32'h14057C80 , 32'hF97EB7D0 , 32'hCB845C00 , 32'h03011FA8 , 32'hFCD0117C , 32'h1D0AE4C0 , 32'h0F97E260 , 32'h0B7C6090 , 32'h056E6C60 , 32'h14089220 , 32'h01966E7C , 32'hECDF5740 , 32'h040085C0 , 32'h0692BF80 , 32'h07DB9F00 , 32'h0DE4E7F0 , 32'h021F5E30 , 32'hF24E8D70 , 32'h0335E8C0} , 
{32'h241DAC40 , 32'hE4463A40 , 32'h01577A88 , 32'hFD22F4F4 , 32'h02F5B184 , 32'h13B8B9A0 , 32'h074725C8 , 32'hE28A6BA0 , 32'h20755640 , 32'hE2CE3160 , 32'hDC2C93C0 , 32'hD8F47900 , 32'hD9C48AC0 , 32'hE7C3A380 , 32'hEDBBEF00 , 32'h0F59EA00 , 32'hFA0914E8 , 32'hF0E72540 , 32'h1304CDE0 , 32'hF6245020 , 32'hEA10CA80 , 32'hFC6D26D0 , 32'hEA7C0A40 , 32'h1315EE60 , 32'h17813A40 , 32'hE93B1AA0 , 32'h06BDB9A0 , 32'hEBDB7E80 , 32'h18D25AC0 , 32'hF9A7C148 , 32'h01B390BC , 32'h026E9188 , 32'h098E4A70 , 32'h155489C0 , 32'hEC730FC0 , 32'hEF82DFA0 , 32'hFBC40BA0} , 
{32'h06CF0A40 , 32'hFD486510 , 32'hFA20F3F0 , 32'hFD73F49C , 32'h01AF7E48 , 32'h0D262050 , 32'h05638428 , 32'hF450AF90 , 32'h28883500 , 32'h0110CD20 , 32'hDB0DBA40 , 32'hEB9C1F80 , 32'hEDB373C0 , 32'hEB798860 , 32'hEF55D3A0 , 32'hFF8F2D79 , 32'h0A2421E0 , 32'hF90FCEA0 , 32'h1BEA46C0 , 32'h04CA5270 , 32'hEFCA3560 , 32'hDF6986C0 , 32'h04180B08 , 32'h03F5BF10 , 32'h04D3AE88 , 32'hE88F3260 , 32'h0F705EB0 , 32'hEE5564E0 , 32'h0E6A6320 , 32'h0D9177E0 , 32'h052D3F78 , 32'hFB8CEBC8 , 32'hF991AF40 , 32'hFBAB3878 , 32'hFA202BD0 , 32'h036BB668 , 32'h092D1270} , 
{32'h2B889B40 , 32'hD9ED8CC0 , 32'h0AB586B0 , 32'hEBAE1160 , 32'hFF5A0091 , 32'hE1A07A80 , 32'hFD0F17A8 , 32'h17825A40 , 32'h308118C0 , 32'h0C6314B0 , 32'hE86ACB60 , 32'hED851E80 , 32'hE535DC40 , 32'hF1024EB0 , 32'hF1653A50 , 32'hF9828548 , 32'hFF6337EA , 32'h001E2272 , 32'h1B6E1900 , 32'h05899360 , 32'h0FC77F30 , 32'h066050E0 , 32'hF89B2560 , 32'hE01A3940 , 32'hFA64FA00 , 32'hF8810F88 , 32'hFEAF5CFC , 32'h09735E00 , 32'hFFA36FDE , 32'hFBF91EF0 , 32'hE3F29BC0 , 32'hF2831EF0 , 32'hF703CC00 , 32'hE964B620 , 32'h04355580 , 32'hFCCB2978 , 32'h038E2144} , 
{32'h36AEA4C0 , 32'hCF165C80 , 32'h143C0FE0 , 32'hF2FB4CF0 , 32'h0B34AB20 , 32'hD5C80600 , 32'hF7B42DF0 , 32'h1AF8D5C0 , 32'h299D7DC0 , 32'h214DB180 , 32'hF7E5E3D0 , 32'hF3FC3BA0 , 32'hFB6F05C8 , 32'h04FF0BF8 , 32'hF44D7EB0 , 32'h0156D1EC , 32'h0415A6F0 , 32'hFDC82E5C , 32'h17594D80 , 32'h08546D70 , 32'hF9F8E118 , 32'h04ACBDC0 , 32'h07805BD0 , 32'hF326E6F0 , 32'h015CE464 , 32'hF6A75750 , 32'h068C63C0 , 32'hEF6030C0 , 32'hF8D9C828 , 32'hFDC08A94 , 32'hF9B389B0 , 32'hFA4B5AE8 , 32'hEFCC0E60 , 32'hF5354E10 , 32'hFE8739EC , 32'h06A2DFD8 , 32'hFEDF87E8} , 
{32'h2ECD3780 , 32'hDB788780 , 32'h134147C0 , 32'hFBEA1680 , 32'h02CEA6BC , 32'hDECE4200 , 32'hF9802888 , 32'h1EBFD180 , 32'h1A719AA0 , 32'h1D13A420 , 32'h0AC52A00 , 32'h148D1AC0 , 32'h38D43040 , 32'h20C7A5C0 , 32'h07A06700 , 32'hF9724A10 , 32'hE4296A40 , 32'hFC09AA78 , 32'hFEA04B20 , 32'h0CE20370 , 32'h02F23D50 , 32'h12A04FC0 , 32'h0C83B480 , 32'h082B7D20 , 32'hF60E21A0 , 32'h093BBD60 , 32'hEED361C0 , 32'hF4A3F190 , 32'hF09C6220 , 32'hEF18DDE0 , 32'hF52EB8A0 , 32'hFAEC1220 , 32'h157D6FA0 , 32'h078AE678 , 32'hFBF4FDE0 , 32'h048A8B20 , 32'h1B906380} , 
{32'h2BD31880 , 32'hEDC9B320 , 32'h0EB903D0 , 32'hF839EEE8 , 32'h020E2434 , 32'hE44198C0 , 32'hFC419448 , 32'h213D7E80 , 32'h0ACC2E00 , 32'h08356CD0 , 32'h09F95CC0 , 32'h15898D40 , 32'h15E1B5E0 , 32'h1A145AC0 , 32'h1C2B28A0 , 32'hFEB44A1C , 32'hFA7D85A0 , 32'h08CDFA30 , 32'hEA56E000 , 32'h0FAF4440 , 32'hFF63FEF8 , 32'h162FBE60 , 32'h09575FD0 , 32'hFF4832E8 , 32'h03EC7BC0 , 32'h24843B40 , 32'hFB2E6CD8 , 32'h06DFF9F8 , 32'hEDB9F280 , 32'hF4F3C050 , 32'hF8D1A488 , 32'h02CD720C , 32'h02B98340 , 32'hFE4B5AFC , 32'h04BE8008 , 32'hFAF4AC08 , 32'hF6AB4ED0} , 
{32'h1B71B6A0 , 32'hEE5231C0 , 32'h0345166C , 32'h0F1E5300 , 32'h0189C93C , 32'hE1BD91E0 , 32'h007E0F91 , 32'h0FA098B0 , 32'hFFC09F04 , 32'h06A7C1B0 , 32'hE16877E0 , 32'hF3D68360 , 32'h0094DBC6 , 32'h0F1DF960 , 32'hF5FE26B0 , 32'hE991EC20 , 32'h0539ACE0 , 32'hF2D03640 , 32'hFE66FE9C , 32'h028B0174 , 32'hF5808570 , 32'h1491D2E0 , 32'hF8F96020 , 32'hFE7398B8 , 32'h0943BBA0 , 32'hF83259F0 , 32'hF96C4328 , 32'hF66E9AE0 , 32'h08109D80 , 32'h0A581A50 , 32'hFE668494 , 32'hFCB9F670 , 32'h08E132F0 , 32'h09258730 , 32'hFC273E98 , 32'hFF38225B , 32'h082161B0} , 
{32'h1F88B740 , 32'hFEEEEE64 , 32'h095D1A10 , 32'hF2BFD380 , 32'h0B9BBBC0 , 32'hF28BDBC0 , 32'h078F34F0 , 32'h06ACDB08 , 32'hFDAD299C , 32'hFCCF44BC , 32'hFDF3BCAC , 32'h0222E358 , 32'h16DB3BE0 , 32'h1E88AE00 , 32'h0294AC70 , 32'h051B5800 , 32'hF9706248 , 32'hF9BA8018 , 32'hEF6B13A0 , 32'h0B6B69B0 , 32'hD7A49740 , 32'h11B1CBA0 , 32'h026333B0 , 32'h0E716A30 , 32'h13040240 , 32'hF5BD9E50 , 32'hFEF878BC , 32'hF5EDA340 , 32'h09AF7670 , 32'h0766A0F0 , 32'h16A16900 , 32'h1864EB20 , 32'h068EEDC0 , 32'h12516A40 , 32'h10D91260 , 32'h0D7BBB10 , 32'hF4C2FE30} , 
{32'h0925FF90 , 32'hF9E56D88 , 32'h00C4D852 , 32'hFEC52400 , 32'h04628960 , 32'hF97AAC20 , 32'hF8234F40 , 32'hF4DD7060 , 32'hF8FC7550 , 32'hFF251355 , 32'hF87F9DE8 , 32'h0527E0B8 , 32'h02515434 , 32'hFED5EF20 , 32'hF5C77660 , 32'hFCE14228 , 32'hF38489B0 , 32'hFA9834B8 , 32'hF4D2A140 , 32'hF7AB2BF0 , 32'hF6612250 , 32'hF3D2E030 , 32'hF49839D0 , 32'hFACE0D20 , 32'hF70B20B0 , 32'h06E96648 , 32'hFBDD3118 , 32'h0B38F630 , 32'hFA8B6568 , 32'h10CAE1A0 , 32'hF070D0E0 , 32'hFF3B04D3 , 32'h047826D0 , 32'hF8F6C640 , 32'hF74F4420 , 32'h048223D8 , 32'h0375DBEC} , 
{32'h046E3018 , 32'hFD19E140 , 32'h02B984C4 , 32'hFEBB15E0 , 32'h013282A8 , 32'hFEE541B8 , 32'hFFCD51D7 , 32'hFCBA3220 , 32'hFF70ED0C , 32'hFC6E8B50 , 32'h01E3C3EC , 32'h011E13B8 , 32'hFF7AB41B , 32'hFC904DC0 , 32'hFFE68703 , 32'h00652F0C , 32'hFD934A18 , 32'h01E692DC , 32'hFB2CB180 , 32'hFF0CCB11 , 32'h0021415B , 32'hF73BA980 , 32'hFD4D9EC0 , 32'h00E07EC1 , 32'hFC9C7E14 , 32'hFEB83E38 , 32'hFDA104C4 , 32'h061097C0 , 32'hFC81A4D4 , 32'h0284CE60 , 32'hF9AE50F8 , 32'hF9F37800 , 32'h0663E228 , 32'hFF787088 , 32'hFFB2218A , 32'hFE621F1C , 32'h01F56FD0} , 
{32'h000560EA , 32'h00020B70 , 32'h0001C463 , 32'hFFFE0792 , 32'h0000706E , 32'h0001E263 , 32'h00002EE8 , 32'hFFFF6675 , 32'h0001ADB6 , 32'hFFFB3348 , 32'h0000F0A4 , 32'hFFFB5F31 , 32'h00008CA4 , 32'h0001E482 , 32'hFFFFECBF , 32'h0000DC35 , 32'h00050E48 , 32'h000444FB , 32'hFFFEE0EE , 32'hFFFDD5FD , 32'hFFFF6C4F , 32'h00005537 , 32'h00035BD6 , 32'hFFFFC014 , 32'hFFFD2DF1 , 32'hFFFC91A0 , 32'h00005CCF , 32'h0000B80A , 32'h00013795 , 32'h00011FE6 , 32'h00002C67 , 32'hFFFD0239 , 32'hFFFF0368 , 32'hFFFE7BEE , 32'h00003373 , 32'h0004D7F3 , 32'h0001FF97} , 
{32'hFFF98935 , 32'h000074B0 , 32'h00010D9A , 32'hFFFBE906 , 32'h0003F87F , 32'hFFFF073C , 32'h0004DFD1 , 32'hFFFDFC1C , 32'h00010F3B , 32'h0002C19A , 32'hFFFE3CF1 , 32'h00008EFD , 32'hFFFF6475 , 32'h00046A54 , 32'hFFFEB41C , 32'hFFFE4B88 , 32'hFFFF3C91 , 32'hFFF9DE6D , 32'h00004326 , 32'hFFFEF38B , 32'h000116FE , 32'h0003ADD2 , 32'hFFFC9D9D , 32'hFFFF4C8B , 32'hFFFDA94E , 32'hFFFEBB9C , 32'h00002A35 , 32'h000100E9 , 32'hFFFF0268 , 32'hFFFE8B46 , 32'hFFFCF70F , 32'hFFFC43F3 , 32'h00038B41 , 32'hFFFE3FF9 , 32'hFFF9FE5E , 32'hFFFA00F3 , 32'h0002B348} , 
{32'h00044410 , 32'h00022011 , 32'h000388FE , 32'h0007F475 , 32'h00045E36 , 32'h00028229 , 32'h000698CA , 32'hFFF77ED3 , 32'h00028BF9 , 32'h0005B2C5 , 32'h0000C940 , 32'hFFFF3430 , 32'h0004FF49 , 32'hFFFCE78D , 32'hFFFAA3E9 , 32'h0000A0CE , 32'h00069D87 , 32'h0006AE36 , 32'h0005B8FD , 32'h0004EB3F , 32'h0002B319 , 32'hFFFADC8B , 32'h0000F61A , 32'h0002CCAF , 32'hFFFE07AE , 32'hFFFC5818 , 32'hFFFC5583 , 32'hFFF98B5F , 32'h00016AE0 , 32'hFFFD4881 , 32'hFFFCA56B , 32'h00029C8B , 32'hFFFE6841 , 32'hFFFD5F5A , 32'h000702CD , 32'hFFFB6A0D , 32'hFFF9E38C} , 
{32'hFFF98D39 , 32'h000238CA , 32'hFFF9F06F , 32'h000077D9 , 32'h000288E8 , 32'h000054CC , 32'h00015E04 , 32'hFFFCE3B9 , 32'hFFFDFA26 , 32'hFFFEBCC8 , 32'hFFFBC81C , 32'hFFFCFED6 , 32'h00006A43 , 32'h0003231F , 32'hFFFFC3C9 , 32'hFFFCAD67 , 32'hFFFEDDD0 , 32'hFFFC04E1 , 32'h0006EE72 , 32'h00029B01 , 32'hFFFD0932 , 32'h000458CB , 32'h00015939 , 32'hFFFFDB3E , 32'hFFFE31B7 , 32'h00008A2D , 32'h0000F05A , 32'h0001AB48 , 32'h0000EC4C , 32'hFFFA7D3D , 32'h000240D5 , 32'hFFFEED88 , 32'hFFFC665D , 32'h0003DF27 , 32'hFFFD7198 , 32'h0001E018 , 32'hFFFCCA24} , 
{32'h0005BC99 , 32'h00040998 , 32'hFFFDB9E3 , 32'hFFFFA405 , 32'h0000B5A4 , 32'hFFFCCDBF , 32'hFFFE0D96 , 32'hFFFF29AE , 32'hFFFF2F24 , 32'h0004CB2A , 32'h00006830 , 32'hFFFE15BE , 32'h000183F7 , 32'hFFFEDB86 , 32'h00027FFF , 32'hFFFA2B55 , 32'hFFFD377A , 32'hFFFAD42F , 32'hFFFA54F9 , 32'h0002146C , 32'hFFF7FF52 , 32'hFFFFA1FF , 32'hFFFEA6D5 , 32'h000057AA , 32'hFFFFFDD0 , 32'h0000D705 , 32'h00013BC9 , 32'h0001EB69 , 32'h0002D8A6 , 32'hFFFDF979 , 32'hFFFEA022 , 32'h000343DE , 32'h00015CB6 , 32'h00004A09 , 32'h00000EB4 , 32'hFFFC3570 , 32'hFFFD849E} , 
{32'h045A8188 , 32'hFD2A38E4 , 32'h0263776C , 32'h00B7276B , 32'h023DF2F4 , 32'hFD86764C , 32'h00CB6716 , 32'h02056FA0 , 32'h038B7BC0 , 32'hFFAC26C4 , 32'hFDF26F08 , 32'hFCF0B604 , 32'hFE7D8274 , 32'hFEB58FD4 , 32'hFCB6C264 , 32'h003A2130 , 32'hFC3AABD8 , 32'h0012643B , 32'hFFFD4553 , 32'hFBBE4FA0 , 32'hFD6BA91C , 32'h020968A8 , 32'h00510DB7 , 32'hFDCC5EAC , 32'hFF211851 , 32'hFF2BEFB9 , 32'hFDB83610 , 32'hFFB49802 , 32'h01BB0720 , 32'hFF3DC928 , 32'hFC9C4BE8 , 32'hFAA45120 , 32'h00A2655E , 32'h00F7940C , 32'h0311C77C , 32'hFD373618 , 32'h01BA16C8} , 
{32'h0C9BFC90 , 32'h06E171C8 , 32'hFE8AF350 , 32'h0EF51560 , 32'h051DD918 , 32'h072A2F70 , 32'hF8C92570 , 32'hFCAB26DC , 32'hFDE6A6E8 , 32'hFEBAB554 , 32'h011CABD0 , 32'h036D7414 , 32'hFAB8DC40 , 32'h1826E820 , 32'hF3344C50 , 32'h010B0A34 , 32'h0DC7F600 , 32'hF5AAF320 , 32'h030ABE10 , 32'h0511BA90 , 32'hFE531608 , 32'hF8276C38 , 32'h0B0F8C30 , 32'h064FFEE0 , 32'hFED01680 , 32'h04685130 , 32'h08516EA0 , 32'h0232E948 , 32'h08F33DE0 , 32'hF236B390 , 32'hEFF56160 , 32'hFD499178 , 32'h0A291570 , 32'h01B3ECF0 , 32'hFB2EC520 , 32'h05F750D0 , 32'hFE34A81C} , 
{32'h24EF1180 , 32'hF7827D30 , 32'hEF119B20 , 32'h13407280 , 32'hF2C13170 , 32'h141C6FA0 , 32'h060748F0 , 32'hFA4BB568 , 32'hE5205520 , 32'h000BE3E2 , 32'h0E993160 , 32'hF2B252F0 , 32'hF9389150 , 32'h09AC6EB0 , 32'hF3C38490 , 32'hEF49C960 , 32'h004BC881 , 32'hF6BC5440 , 32'hFC6972AC , 32'h1609BB80 , 32'h0E698040 , 32'h05096F30 , 32'h08F59C30 , 32'hF667D240 , 32'hFFFA2918 , 32'hFC331CFC , 32'hF9231108 , 32'hFD188248 , 32'h06C4BBD0 , 32'h06121128 , 32'h0060772C , 32'hEDAFB540 , 32'hF8100958 , 32'h0719C9F0 , 32'hFBE26948 , 32'h055D8FD0 , 32'hFF44B4E8} , 
{32'h1DEE0B80 , 32'hF385A1B0 , 32'hF2A12420 , 32'h033E62D4 , 32'hFA0087D8 , 32'h1F5CE720 , 32'hF47F9650 , 32'h06F61CA8 , 32'hE493D000 , 32'h01D6E7CC , 32'h0DB566A0 , 32'h03E77CF4 , 32'hF2A9E720 , 32'h0296FFC8 , 32'hFB5044D8 , 32'hF46A5150 , 32'hF539BB50 , 32'hFB2B5180 , 32'h04F6E840 , 32'h09CD3B60 , 32'hFF3A9184 , 32'h02D93194 , 32'h1026A560 , 32'h042435F0 , 32'hFC787B88 , 32'hF3551420 , 32'hF5CC1E70 , 32'hF4DD49F0 , 32'hFB8A4C60 , 32'h0A639330 , 32'h03F0DFC0 , 32'hFDC9ADC8 , 32'hF1C3FE30 , 32'h044492A8 , 32'hFA4C6E30 , 32'h06DAD2B0 , 32'hF0CC8110} , 
{32'h30CA2980 , 32'hFA682910 , 32'hE8149600 , 32'h13DB1700 , 32'hF3459A70 , 32'h1D2DBF00 , 32'h0196F9A8 , 32'hF807BAF8 , 32'hE03741C0 , 32'h04C06F88 , 32'h138F3A40 , 32'h02475C78 , 32'h033D1E14 , 32'h00FD4691 , 32'hEEF5C980 , 32'hECAE3120 , 32'hFE0D8F10 , 32'hF9BE1F10 , 32'hFB6FF6D8 , 32'h195250E0 , 32'hFD34A724 , 32'h051B2330 , 32'h06ECB5E8 , 32'hE80AC5A0 , 32'hF9726860 , 32'hF9FC8840 , 32'h0E8FE700 , 32'hF94BC340 , 32'h036A2464 , 32'h1C4E11C0 , 32'h0DC195E0 , 32'hF1A2C270 , 32'hF5946070 , 32'hED01ECC0 , 32'hFFBD15DA , 32'hF8022F18 , 32'hE7C13DE0} , 
{32'h154C1EC0 , 32'h07CB70F8 , 32'hEA13A8A0 , 32'h0FA7D8B0 , 32'hF1539CB0 , 32'h1B3141C0 , 32'h062A29B0 , 32'hF2173310 , 32'h07CC93B8 , 32'hFC9BBEF8 , 32'hFFB90298 , 32'hFF20E9C0 , 32'h0A76ECF0 , 32'h0B905B50 , 32'h00F29C02 , 32'hEE4225A0 , 32'hFCD0BFB8 , 32'hF2193AD0 , 32'h0839C7E0 , 32'h0AD60E80 , 32'hFB6DEE20 , 32'h0059B8B0 , 32'hF98440F0 , 32'hFD622DC0 , 32'h01B3DEA8 , 32'hFCC52AD4 , 32'hF7251A00 , 32'h025C3858 , 32'hFE452C40 , 32'h0A919730 , 32'h0CA1C880 , 32'hF37F8460 , 32'hFBB8D030 , 32'hF5186450 , 32'h02AD4E88 , 32'hFFA556F3 , 32'hEC5392A0} , 
{32'h19A524E0 , 32'h0E25BEE0 , 32'hF2EB6850 , 32'h19D914E0 , 32'h0650DF98 , 32'h19E0F480 , 32'h14CC2F40 , 32'hFF43F600 , 32'hFEA7C968 , 32'hFD180F08 , 32'h077C0878 , 32'hFFA35CD1 , 32'hF6F576F0 , 32'h02A09370 , 32'h0408DD20 , 32'hE9838760 , 32'hF644FFC0 , 32'hE8E98E60 , 32'hF803FA28 , 32'h13A0A4C0 , 32'h06ABAB58 , 32'hFF57770B , 32'hF6608BE0 , 32'hEDF9D940 , 32'h0A37BAD0 , 32'hFAE1BBD0 , 32'hFC98CB98 , 32'h0762B4C8 , 32'hF54526A0 , 32'h0150690C , 32'h0BAFCC60 , 32'hF9618118 , 32'h130AC0E0 , 32'h02555460 , 32'h08CD1CE0 , 32'h094A0B50 , 32'hE83794E0} , 
{32'h1DB71D40 , 32'h0FF7B1D0 , 32'hF1272FE0 , 32'h1F4F9B40 , 32'hFE8CD6F0 , 32'hFE0B43B0 , 32'h26AA7DC0 , 32'hF1D8F9B0 , 32'hFE314EE8 , 32'h0A18DAD0 , 32'h085E6580 , 32'hF96D1C90 , 32'h063BEB20 , 32'h03177F48 , 32'h06407698 , 32'hFCE7F1E0 , 32'h04EEE0C8 , 32'hFB41CB70 , 32'h02C72B58 , 32'h032C2480 , 32'h06DAA8C0 , 32'hFE3DD054 , 32'h00B43544 , 32'hFB2F05B8 , 32'hFFD285B8 , 32'h038B7410 , 32'h064B7E00 , 32'hFB4B53C8 , 32'hFE820510 , 32'h027C459C , 32'hFBC3BBA0 , 32'hF0D29D00 , 32'h03819FC4 , 32'h00958821 , 32'h02E6847C , 32'h02AF3F84 , 32'hFDDC2E28} , 
{32'h32FF8880 , 32'h2694DD00 , 32'hFBF3EB88 , 32'h316D8D00 , 32'h19153C80 , 32'hF56B9290 , 32'h37A83CC0 , 32'hE33051C0 , 32'hED168780 , 32'h1049C2E0 , 32'hFC96ADF4 , 32'hFD340A2C , 32'hEB563220 , 32'hFD5AB8E4 , 32'h0D4C1CF0 , 32'h01138450 , 32'h0133E554 , 32'h02BF4B48 , 32'hF3C02580 , 32'hFF752E85 , 32'h0E35D000 , 32'h0CE3B510 , 32'h03B4E360 , 32'h08E093B0 , 32'h06580708 , 32'h158F20C0 , 32'hF8E83288 , 32'hEC1B7340 , 32'h03FD1A50 , 32'h167FABA0 , 32'hFD7EB5B0 , 32'hFB29E658 , 32'hFDB05F7C , 32'hE6914060 , 32'h02AF4F88 , 32'h067F4FF8 , 32'hF6D0F270} , 
{32'h11FA38E0 , 32'h24F27580 , 32'hEE82FE20 , 32'h45050300 , 32'h160E6A60 , 32'hE90327A0 , 32'h44419C00 , 32'hE27DB700 , 32'hF270E8B0 , 32'h11598EA0 , 32'hFD2D5478 , 32'hE4FFE5E0 , 32'h155B7580 , 32'hFE137C2C , 32'h13EC4280 , 32'h191B5560 , 32'h01639CEC , 32'hF904AED8 , 32'hFF44BBA4 , 32'hFE76D67C , 32'h055DBAF8 , 32'h057193F0 , 32'hEFCD6980 , 32'hFFB5AC0F , 32'hEC556860 , 32'h1A898680 , 32'h0E8BBA90 , 32'hEBA88A00 , 32'h1712B8E0 , 32'h1A171420 , 32'h041ABAB8 , 32'h01218CE0 , 32'h0FDAFD90 , 32'hED1EA920 , 32'h08287C30 , 32'h0874BCB0 , 32'h045AFC78} , 
{32'h14919300 , 32'hEDCA3440 , 32'hEF5DD400 , 32'h3C9A1080 , 32'h083108C0 , 32'hF7A528F0 , 32'h250B4940 , 32'hEA209820 , 32'hEC00DE00 , 32'hF42689F0 , 32'hFE8A7B24 , 32'hDD180340 , 32'h0C95FD70 , 32'h0C8DAF80 , 32'hF5A1B1B0 , 32'h1CC05AE0 , 32'h07C08D18 , 32'h08103890 , 32'hDD5A2E00 , 32'h0B040A20 , 32'h19ECA4C0 , 32'hF43CBC10 , 32'hF6CBA860 , 32'hF314E730 , 32'hDC5F3FC0 , 32'hE895E0A0 , 32'h19B6A360 , 32'h04039FE0 , 32'h08905150 , 32'hFA5538A0 , 32'hEA2ABE80 , 32'h0E95E6A0 , 32'h0C21F540 , 32'h1673D6C0 , 32'hF07C3B20 , 32'hF4B95210 , 32'h0965D730} , 
{32'hFD792DF4 , 32'hDB80A440 , 32'hE7795D60 , 32'h222C7CC0 , 32'hE60197E0 , 32'hF0CB0990 , 32'h1613F5C0 , 32'hEA146300 , 32'hF95D77F8 , 32'hE06A55C0 , 32'hF57DCB90 , 32'hD543A7C0 , 32'h19ABA940 , 32'h0AC36840 , 32'h0DF28A50 , 32'h02E7C6E4 , 32'hF368F0C0 , 32'hEFBE9B40 , 32'h0322F200 , 32'h1FB6A020 , 32'hF759B820 , 32'hF3B3F7F0 , 32'hEE427000 , 32'hEBEFEF60 , 32'hF7505990 , 32'hE2887420 , 32'h1EE27960 , 32'h0BD37DB0 , 32'h0D684740 , 32'hFB65D308 , 32'hFD63C990 , 32'hEB7897A0 , 32'hF9D2B158 , 32'h1CBB1540 , 32'h02C5F508 , 32'hF37AB3E0 , 32'h053826C0} , 
{32'h028D779C , 32'hE930F960 , 32'hDD00CB40 , 32'h0ECCBB10 , 32'hF19DCD60 , 32'h038F698C , 32'h02BA0938 , 32'hE01F4300 , 32'h0FA88F80 , 32'hD9692680 , 32'hE3260FE0 , 32'hDD1AF900 , 32'hF3612050 , 32'h09665FC0 , 32'hE3AB3920 , 32'h0EB4ED40 , 32'hFE244B48 , 32'hE4C6F7E0 , 32'hE2675940 , 32'hFB8A53E8 , 32'hF7ABEAA0 , 32'h0DF8C380 , 32'h0959C520 , 32'hFCC4E92C , 32'h08E6D860 , 32'h0B27AA10 , 32'hF7D27910 , 32'hFFF6EA03 , 32'hF24EA1A0 , 32'hE91AD6E0 , 32'hF4A86100 , 32'hFF7EC10D , 32'h0E6D02B0 , 32'hFFD375C3 , 32'hFD188580 , 32'hF7207970 , 32'hF47A8EC0} , 
{32'hEE635D40 , 32'h0284DF58 , 32'hEFF166C0 , 32'h0B88BFB0 , 32'hF9E5D7D0 , 32'h045D2B58 , 32'h0D4017F0 , 32'hF23126F0 , 32'h0864F800 , 32'hECC58DE0 , 32'hE7A68D80 , 32'hEBAA87A0 , 32'hD1ABB5C0 , 32'hF3A01C30 , 32'hFAE9CAD8 , 32'h073F9858 , 32'h0DBDC640 , 32'hEEA48FE0 , 32'hF08B5300 , 32'hFFD54829 , 32'hF21C5DA0 , 32'h0357B808 , 32'hFF0533BB , 32'h0215E58C , 32'h06D59730 , 32'hF04232A0 , 32'h0303FE54 , 32'hE8185E00 , 32'h07E160B8 , 32'hFC24ED08 , 32'h02ADCA40 , 32'h019171E4 , 32'hFC11C288 , 32'hEC55CDA0 , 32'h00459059 , 32'h0EB0A620 , 32'hF01E9610} , 
{32'hF76E8860 , 32'hFF5D5C10 , 32'hF47F4A50 , 32'h12625DC0 , 32'hF3BA4870 , 32'h044A16F8 , 32'hF1181750 , 32'h19623780 , 32'h1CC0AD60 , 32'h1E1ABA00 , 32'hE9B95E40 , 32'hE105B620 , 32'hDDFB1F80 , 32'hEB933E20 , 32'h08D179A0 , 32'hFA02FD68 , 32'h15E761C0 , 32'hEEAE08E0 , 32'h01C33CEC , 32'h02506338 , 32'h1E5FC860 , 32'h06FEA468 , 32'hF5666A30 , 32'hE84DA300 , 32'h03065874 , 32'hF7C87810 , 32'hF22C0440 , 32'hFF610936 , 32'hF66F23A0 , 32'hF9F9C2D8 , 32'hF2F9E690 , 32'hFE02B25C , 32'h13000900 , 32'hF2324F20 , 32'hFB544F78 , 32'h0D463800 , 32'h0A48FE50} , 
{32'h059F1B00 , 32'hF169D710 , 32'hF5D548B0 , 32'h12B902E0 , 32'hE56A7A40 , 32'hEC27C860 , 32'hF1873B00 , 32'h1E27A4E0 , 32'h2C847800 , 32'h3A9A2540 , 32'hD0E7E280 , 32'hEAB46020 , 32'hCF8097C0 , 32'hE1084AA0 , 32'hF9B1DA88 , 32'hF801A1E8 , 32'h035DF8E4 , 32'hF5D97D70 , 32'h039D7C74 , 32'h128A9560 , 32'h2C15FDC0 , 32'hF363D760 , 32'h09223810 , 32'hEAFCFF00 , 32'hE2EF7A20 , 32'hF72E4470 , 32'hEBE78620 , 32'h08ABB0B0 , 32'h0F9A1820 , 32'h05B4D3B8 , 32'h0247F424 , 32'hF92A8F28 , 32'h11D083C0 , 32'hEF0096C0 , 32'hFB5AA388 , 32'hF2DCD3A0 , 32'hF318D230} , 
{32'h156E8FC0 , 32'hEBF8C460 , 32'hEB68B3A0 , 32'h18999360 , 32'hF91D8548 , 32'hEA883F40 , 32'h0184ED18 , 32'h3FB77D80 , 32'h1FAC69A0 , 32'h20CFDFC0 , 32'hD50B5C00 , 32'hF3CDB210 , 32'hFD03C578 , 32'hF1360C80 , 32'hEC606F20 , 32'h073E9450 , 32'hEA8C19E0 , 32'h14767460 , 32'h132ADDC0 , 32'h19640CA0 , 32'hE7E072C0 , 32'hFEF7EE80 , 32'h03B5C1D4 , 32'h07D30850 , 32'hF68E3E90 , 32'hF8EF2B38 , 32'hEC6C7FC0 , 32'h06D2E4F8 , 32'h025600E0 , 32'h01A8B48C , 32'h0CA25960 , 32'hFE516A0C , 32'hF8DFE600 , 32'hF332A940 , 32'h02117F30 , 32'hF76D3230 , 32'h00269A59} , 
{32'h151AC620 , 32'hED318D20 , 32'hF2A70800 , 32'h1C17DE20 , 32'hF8BE45B8 , 32'hF80A07B8 , 32'hF22CF900 , 32'h40DDC280 , 32'h19B05DE0 , 32'h23E78280 , 32'hEAFC8820 , 32'hFF42352E , 32'h13D02260 , 32'hFBF4AE68 , 32'hE96EA560 , 32'h04297E38 , 32'hE22F4DC0 , 32'h09B33500 , 32'h19D62660 , 32'h2190BBC0 , 32'hF4682250 , 32'hFB513238 , 32'h0B7DF620 , 32'h06B94E98 , 32'hFEE84118 , 32'h06DD2698 , 32'hED9705A0 , 32'h17AF31C0 , 32'h04449068 , 32'hF9FF7438 , 32'hF408DE90 , 32'hFCB0AE2C , 32'h01FAEE64 , 32'h0018EA79 , 32'hFF7CC206 , 32'hF2FB3F40 , 32'h07D3E960} , 
{32'h05EEC8C0 , 32'h04FAA588 , 32'hF8694898 , 32'h09974BA0 , 32'hFE61E09C , 32'hFF03B71B , 32'h09010E70 , 32'h0ECD88B0 , 32'h09F43590 , 32'h1D09EB00 , 32'hEE902540 , 32'hF4E720D0 , 32'hFCAC61F4 , 32'h051D96D0 , 32'hF9EF8A58 , 32'hFAA03590 , 32'hE8D24480 , 32'hFF37324C , 32'h04EA0570 , 32'h0AC08FE0 , 32'hF9697490 , 32'h082C5B00 , 32'h02BD7FB4 , 32'h11449440 , 32'h0BA76070 , 32'hF8267308 , 32'h0C9143A0 , 32'h0B13A060 , 32'h0003AF86 , 32'h09DACD40 , 32'h00D8BE5E , 32'hF78DB040 , 32'h01176514 , 32'h0000982C , 32'hF22ED3C0 , 32'hFA9C6940 , 32'h0A350C10} , 
{32'h0B4C34C0 , 32'hFAFD5750 , 32'hFEEE2808 , 32'h06A41C80 , 32'hF8AAB6B8 , 32'hF580FA90 , 32'hFCA6FA40 , 32'h181CF060 , 32'hFBEEB5D8 , 32'h063E0DB8 , 32'hFD4DCF3C , 32'h0129E208 , 32'h1285ECE0 , 32'h01471370 , 32'h0DA446F0 , 32'hFB2EC8D8 , 32'hE3FF0820 , 32'h0377BDBC , 32'hF1BBB810 , 32'h04E5CE20 , 32'hF83EAF38 , 32'hFDBC8038 , 32'hFA2A8D20 , 32'hF5911140 , 32'hFE59EEF0 , 32'h08D13D60 , 32'h040DB0B8 , 32'h053D6F98 , 32'h0302C460 , 32'hFA455860 , 32'hE9A3A600 , 32'hF22482A0 , 32'h0079021F , 32'hFEB6DCB0 , 32'h01B72904 , 32'hED2D99E0 , 32'h09A69750} , 
{32'h2BCE5000 , 32'hF1A92B20 , 32'h0F61D6C0 , 32'hF28CEEF0 , 32'h0A935E90 , 32'hE5D24880 , 32'h130C5840 , 32'h032D3E7C , 32'h116B04E0 , 32'h00650054 , 32'h0001476D , 32'hF6425D90 , 32'h0891CE00 , 32'h15D25920 , 32'h010603A4 , 32'hF7127C50 , 32'hF58813E0 , 32'h02C685C0 , 32'hF3EE9EF0 , 32'hFF864CAD , 32'hE2395B00 , 32'h14453C20 , 32'h06E8B7E8 , 32'h01440D88 , 32'h05524308 , 32'h059E6230 , 32'h01CCE518 , 32'hFD615DD0 , 32'hFA37E010 , 32'h01E41C78 , 32'h0401E640 , 32'h0D3EE9A0 , 32'hFD3F59D4 , 32'h01B4C120 , 32'h108FA7A0 , 32'h04DA9B58 , 32'h013DBADC} , 
{32'h0CD7A730 , 32'hF59E2140 , 32'h04BC31E8 , 32'hFC9EB4C8 , 32'h0BAC1930 , 32'hF0DD2AA0 , 32'hF7DB1DB0 , 32'hFB365758 , 32'hFF80BCA5 , 32'h06B4B9C8 , 32'hEAE4DF20 , 32'hF91FD120 , 32'h00AACFF9 , 32'h11063000 , 32'hF07823F0 , 32'hF489C7F0 , 32'hF428A1F0 , 32'hF2EB0310 , 32'hF4CB6350 , 32'hF0367B50 , 32'hF4B38F60 , 32'h07EECDB0 , 32'hFB745770 , 32'hF92A8E50 , 32'h03A700B0 , 32'h03068B74 , 32'hF36523A0 , 32'h00BB5390 , 32'h041191D8 , 32'h1022C140 , 32'hFDABFF48 , 32'h0B0C1720 , 32'h004EF0F0 , 32'h06A251D0 , 32'h069300A8 , 32'hFE01C974 , 32'h0A71CAC0} , 
{32'hFFFF9A22 , 32'hFFFF7BA4 , 32'h000319BE , 32'h00000D81 , 32'hFFFC5019 , 32'h00008477 , 32'hFFFF246F , 32'hFFFD6770 , 32'h0000F1B8 , 32'h000240B1 , 32'hFFFDC79B , 32'hFFFD36A7 , 32'hFFFCF703 , 32'hFFFED7B7 , 32'hFFFCE053 , 32'h00001D35 , 32'hFFFF1A65 , 32'hFFFE2FE8 , 32'h0002C92B , 32'h0000EDDC , 32'h00019633 , 32'hFFFE7708 , 32'hFFFF543B , 32'h00016B6E , 32'h000448CB , 32'h0001E351 , 32'h00013CAC , 32'hFFFE1B6D , 32'hFFFD4632 , 32'hFFFDA70A , 32'h000151A3 , 32'h0002E3F4 , 32'hFFFF3432 , 32'h00009C51 , 32'h0000B71A , 32'hFFFCED1E , 32'hFFFF17AB} , 
{32'h00017781 , 32'hFFFD5CB5 , 32'h00040185 , 32'h0000C6E7 , 32'h0004821F , 32'hFFFCAE3A , 32'h00010BF1 , 32'hFFFA5F09 , 32'hFFFFA1F1 , 32'h0000607A , 32'h0003DACE , 32'h0000E78E , 32'h00005646 , 32'h0001025F , 32'h0000E790 , 32'h000223C7 , 32'hFFFE026A , 32'hFFFD9999 , 32'hFFFEFDC7 , 32'hFFFD63AE , 32'h00058CFB , 32'h0000D1D9 , 32'h0000E6C5 , 32'h0006E7F3 , 32'hFFFF7E64 , 32'hFFFD0A25 , 32'h000056B3 , 32'hFFFE4B83 , 32'h0003D1AB , 32'h0004889B , 32'hFFFE6644 , 32'hFFFFA5B6 , 32'h00001CEB , 32'h000195B3 , 32'h00056764 , 32'h00007570 , 32'hFFFCF143} , 
{32'h0008B27C , 32'hFFFDCE1D , 32'h0004BDBB , 32'h0001CEA3 , 32'h000050DB , 32'hFFFB2941 , 32'h00007056 , 32'h0002717C , 32'hFFFBAEE1 , 32'h00063A1C , 32'h000323D7 , 32'hFFF67AF7 , 32'hFFFC8E1E , 32'h00014E78 , 32'hFFFCF871 , 32'hFFF96CD7 , 32'h0002B52E , 32'h000143D4 , 32'h000193C1 , 32'h0003E001 , 32'h00051AC3 , 32'hFFFB249B , 32'hFFF92BE3 , 32'hFFFB9D4B , 32'h00001C99 , 32'hFFF8A96A , 32'hFFFFC402 , 32'h0003F367 , 32'hFFFED355 , 32'hFFFB5C81 , 32'h000066BD , 32'hFFFC2076 , 32'hFFFADB4A , 32'hFFFCAFF3 , 32'h00014B9C , 32'h00003E5B , 32'hFFFE9703} , 
{32'hFFFFB3EF , 32'h0004475A , 32'h00032DBA , 32'h0000C25F , 32'hFFFC0584 , 32'hFFFEB92F , 32'h00015C55 , 32'hFFF81CD8 , 32'hFFFF0ABA , 32'hFFFE3889 , 32'hFFFDE2CF , 32'h000296BB , 32'h00057C49 , 32'h0000840A , 32'hFFFE70F5 , 32'h00002182 , 32'hFFFD6323 , 32'hFFFB8AD6 , 32'h0001025F , 32'hFFFF63B5 , 32'h0001C29A , 32'h000068C9 , 32'h00032DB8 , 32'hFFFEC2F1 , 32'h00000C49 , 32'hFFFEABA7 , 32'hFFFBEE2D , 32'h0006A48B , 32'hFFFCE0A3 , 32'h00013D69 , 32'hFFF33AFB , 32'h0003454A , 32'h0005DA2F , 32'hFFFB713A , 32'h000499C5 , 32'h0002A3BD , 32'hFFFE1A21} , 
{32'h00008F77 , 32'h000559D6 , 32'hFFFB820B , 32'h00016934 , 32'h000315AD , 32'hFFFDDDFF , 32'hFFFA7700 , 32'h00047C54 , 32'hFFFD50B5 , 32'hFFFB4B88 , 32'h0000D04D , 32'h000090B6 , 32'h0000BC8C , 32'hFFFE8431 , 32'hFFFBAB70 , 32'h00010281 , 32'h0004DA1A , 32'h0000AA5F , 32'hFFFFBF9C , 32'h000138D1 , 32'h000143AD , 32'h0002BB2B , 32'hFFFE77D1 , 32'hFFFE9699 , 32'hFFFFE985 , 32'hFFFD0C90 , 32'hFFFE96B1 , 32'h00001896 , 32'hFFFFB652 , 32'hFFF922E7 , 32'h00036DDA , 32'hFFF70217 , 32'hFFFF370A , 32'hFFFF82FB , 32'h00022769 , 32'h00007DEA , 32'hFFFCE3EA} , 
{32'hFFFD8164 , 32'hFFFF5521 , 32'hFFFBDBE4 , 32'hFFFFA679 , 32'h0001DA12 , 32'hFFFE6313 , 32'hFFFDC825 , 32'h0007241E , 32'hFFFADAE6 , 32'hFFFEA5A9 , 32'hFFFF49D5 , 32'hFFFB3540 , 32'h000197CA , 32'hFFFE6B3D , 32'h0005B22A , 32'hFFFB6E48 , 32'h0003E312 , 32'hFFFEFB73 , 32'h00002A17 , 32'hFFFF9E3D , 32'h00028B34 , 32'hFFFDA0F7 , 32'hFFFF4578 , 32'hFFFF9372 , 32'hFFFB85AB , 32'hFFFA4064 , 32'hFFF8DD7C , 32'hFFFF165F , 32'hFFFD28CB , 32'h0000D780 , 32'hFFFFB939 , 32'h00012B1B , 32'h000248E5 , 32'hFFF904CD , 32'hFFFEBCCF , 32'h00006E6F , 32'hFFF9022B} , 
{32'hFFFA56C9 , 32'hFFF9652C , 32'hFFFFF490 , 32'hFFFF1A9B , 32'hFFFA7DA7 , 32'hFFFE5E28 , 32'hFFFCE98D , 32'hFFFF3348 , 32'h000416CA , 32'hFFFC535F , 32'h00041BCD , 32'hFFF9D145 , 32'hFFFBCE71 , 32'h00045F89 , 32'hFFFE6CCB , 32'h00089E43 , 32'h0001968E , 32'h0004D728 , 32'hFFFF738C , 32'h0004D3DD , 32'h00031619 , 32'hFFFCDF2F , 32'hFFFE90F1 , 32'h0000D0B5 , 32'hFFFF9E05 , 32'hFFFD41FF , 32'h000237C2 , 32'h0002C895 , 32'hFFFE55F3 , 32'h0000A975 , 32'h00030779 , 32'hFFFD6C2D , 32'h00061B9A , 32'h00054DCC , 32'h0002C239 , 32'h000111CB , 32'h000017F5} , 
{32'h14DBD920 , 32'h0A036110 , 32'hFAD5CA08 , 32'h08B9A040 , 32'hF844C9B8 , 32'hFC514954 , 32'h0D5F9AB0 , 32'hFE394C20 , 32'hF4187C40 , 32'h04FA0488 , 32'h023A2AC4 , 32'hF1F4CC70 , 32'h0DC229C0 , 32'h0427F078 , 32'h02EBB330 , 32'h02B44DD4 , 32'h03FB8794 , 32'hEB3040E0 , 32'hFADB73D8 , 32'h0745A7B8 , 32'h104D1940 , 32'hFB3029F8 , 32'hE9BEBB80 , 32'h006CB3C2 , 32'h02D38C14 , 32'hFBE05C88 , 32'h0AF81F20 , 32'hFE219848 , 32'hFF45809F , 32'h09CC75B0 , 32'h0335850C , 32'hF3546430 , 32'hFF900445 , 32'hFA32AD48 , 32'h040B2258 , 32'hF7CC46F0 , 32'hFC1E4518} , 
{32'h19ABF880 , 32'h0E08A810 , 32'hFCF3DF74 , 32'h0B1C2CA0 , 32'h0BA772C0 , 32'h06B63DC0 , 32'h22D87780 , 32'h0226B8A4 , 32'h0407F9F8 , 32'h045DF5A8 , 32'h14D09E20 , 32'hF09B6E50 , 32'h0CBE9260 , 32'hF688FDE0 , 32'h09E352F0 , 32'hF52969C0 , 32'hF5A078F0 , 32'hE07CA6C0 , 32'h12CB8620 , 32'h04D33038 , 32'h0A5C80E0 , 32'h02199644 , 32'hF37EB370 , 32'hF244E570 , 32'hF8740948 , 32'hFEC8AA20 , 32'h0B9999B0 , 32'hFE20267C , 32'h0D9C0B60 , 32'h057652F0 , 32'h0E5BCEB0 , 32'hF6B782E0 , 32'h0A79BC30 , 32'h09C8FBA0 , 32'hF43D96B0 , 32'h03903780 , 32'hF7B2DC70} , 
{32'h19B31DA0 , 32'h019EAB40 , 32'hF58FB200 , 32'h0DC6B700 , 32'hFDFA39C8 , 32'h0D6D1A70 , 32'h111E9FA0 , 32'h0122583C , 32'hF2ECA690 , 32'h017D0F00 , 32'h11FF66A0 , 32'hF8E74670 , 32'hF966F550 , 32'hF9C86DF8 , 32'hFFD27B99 , 32'hE9CE38A0 , 32'hFCC7A7BC , 32'hE9A7CE00 , 32'h003D2350 , 32'h09F3D6D0 , 32'h07FF5C40 , 32'h00617416 , 32'h04D19430 , 32'hF6504610 , 32'hFD250494 , 32'h02F5BE68 , 32'hFDA53828 , 32'h067D5F30 , 32'h06E2A860 , 32'hFE04B3B0 , 32'h0FE4BCF0 , 32'hFA709318 , 32'hF54F88B0 , 32'h0921E400 , 32'hF831F0D0 , 32'h064AC6C0 , 32'h0F488870} , 
{32'h28584D40 , 32'h19DB7120 , 32'hEE4F2A20 , 32'h1EE8D780 , 32'hF8757DE8 , 32'hF88DD608 , 32'h1B0279C0 , 32'hF4E57750 , 32'hFE1AE468 , 32'h0AB12960 , 32'h0AF22270 , 32'h0B5978C0 , 32'h0FE9C190 , 32'hF582F5B0 , 32'h05290400 , 32'hED5181A0 , 32'h01802DC8 , 32'hF9447BF8 , 32'h0759A4F8 , 32'hFD55D578 , 32'hF13FC3E0 , 32'hF820D558 , 32'hE8BE5740 , 32'hF445D700 , 32'hF96B5418 , 32'hFB46C5B8 , 32'h085A3D60 , 32'hF4777630 , 32'hFB35DB38 , 32'h1488E9E0 , 32'h12C31980 , 32'hEF581420 , 32'hF9349C38 , 32'hF631AC50 , 32'hFEDA4E84 , 32'hF8BBC250 , 32'hF93AEA40} , 
{32'h31512280 , 32'h17C596A0 , 32'hEAAE4320 , 32'h2D15A080 , 32'h0AF831B0 , 32'hF3DB23F0 , 32'h3BF31440 , 32'hEDBD4A60 , 32'h00D0530E , 32'h0FC112D0 , 32'h0F7A3D80 , 32'hFB9BEF88 , 32'h13AE0600 , 32'hFA285280 , 32'hFA7188F0 , 32'hF1F4E000 , 32'hFA88D2E0 , 32'hED5D4F20 , 32'h065380F0 , 32'hF3C0BB00 , 32'hF6F912B0 , 32'hF97AEEC8 , 32'h03D13510 , 32'hFD967264 , 32'h0050FD17 , 32'h0BCE30B0 , 32'hFEDD404C , 32'hFFAD665B , 32'h05A4AAC8 , 32'h0496A198 , 32'hFC542FD0 , 32'hEDAAFD80 , 32'hF988E068 , 32'hFC2DA9EC , 32'hFD73BEB4 , 32'h02F26900 , 32'h06AD2AD0} , 
{32'h255A8800 , 32'h210098C0 , 32'hFE868368 , 32'h30A77DC0 , 32'h0FC8EEB0 , 32'hF9D09590 , 32'h512CDA80 , 32'hF19DC9D0 , 32'h0A363B50 , 32'h0AEBC610 , 32'h18382140 , 32'h0AD99160 , 32'h0595F280 , 32'hE67008E0 , 32'h16F11500 , 32'hEBF7E2A0 , 32'hF582B190 , 32'hE9988B20 , 32'h0A85C070 , 32'h077AF050 , 32'h05B47658 , 32'hFFE49BA1 , 32'hFA9C0828 , 32'hFD72C620 , 32'h0AA93F60 , 32'h06E925E0 , 32'hF917EBC0 , 32'h05C50FD0 , 32'hF76CD8B0 , 32'hF8C983B0 , 32'h03CA19E8 , 32'hF2B4E700 , 32'hE94090C0 , 32'h0B0F4840 , 32'h133262C0 , 32'h09FD4A40 , 32'h04221A18} , 
{32'h0599A588 , 32'h2560EA80 , 32'h0DE100B0 , 32'h21DC0600 , 32'h1E50F720 , 32'hE0C0B7C0 , 32'h392F25C0 , 32'hEC1F8560 , 32'h0E0E3A50 , 32'h1B09F8E0 , 32'h0B606750 , 32'hFC8787DC , 32'h065F5F48 , 32'hF04E0E60 , 32'h1F35F800 , 32'h01721720 , 32'hFE656B20 , 32'hEAB5D9A0 , 32'hF36FB590 , 32'hE78557E0 , 32'h05086450 , 32'hFC532640 , 32'h06EAD920 , 32'h0B9A1D20 , 32'hFACA7658 , 32'h1FBFB300 , 32'h08B19200 , 32'h005156F1 , 32'h074CF138 , 32'hFAA3B0E0 , 32'hFE19A150 , 32'hFBBD4BB0 , 32'h0341C4E4 , 32'h0DAFC960 , 32'h0B11A8C0 , 32'hF1B68F40 , 32'h17188B60} , 
{32'hF68049C0 , 32'h1C238480 , 32'h0214C724 , 32'h379B9840 , 32'h2A910900 , 32'hE2128120 , 32'h213CA4C0 , 32'hE5220520 , 32'h0CBEDD30 , 32'h14A60E20 , 32'h1E5A6260 , 32'hE6CEC440 , 32'h04D68B70 , 32'hF3A782C0 , 32'h1DC65300 , 32'h32557540 , 32'h06658588 , 32'h2135D880 , 32'hFE87C73C , 32'h06383E28 , 32'hF1182D70 , 32'hFBAD39D8 , 32'h0600A4D8 , 32'h2E185AC0 , 32'hFC7068D0 , 32'h03CFD158 , 32'hF20B39F0 , 32'hE5D45600 , 32'h055730C8 , 32'h0D9A8A20 , 32'h0B7C4560 , 32'h078FF360 , 32'hF00F2B70 , 32'hF1F86BA0 , 32'hF9ECC6C0 , 32'hF307A8C0 , 32'h102470C0} , 
{32'hC95C6300 , 32'hF6A887C0 , 32'h16E4C6E0 , 32'h144B38E0 , 32'h09128120 , 32'hC0C9BDC0 , 32'h0E800A50 , 32'hFA405700 , 32'h1782D800 , 32'hFC705F2C , 32'h33F4F800 , 32'hDD1A9080 , 32'hE8CE70A0 , 32'hFF2CB5DD , 32'h1BF0A9E0 , 32'h41BCE280 , 32'h03EC4CBC , 32'h23502180 , 32'hFDE13DEC , 32'h217658C0 , 32'h0F8BCFB0 , 32'hFEA772A4 , 32'h0F3847D0 , 32'h16BFA140 , 32'hF3A8AD20 , 32'hF99AC070 , 32'h04532188 , 32'hE7A8D240 , 32'h162D4AE0 , 32'hF3B0E810 , 32'hED78DEA0 , 32'hE77BDD20 , 32'h07C36220 , 32'hF2ED9C90 , 32'hF7164E40 , 32'h0D3707D0 , 32'hE32CA340} , 
{32'hBA521400 , 32'hA8163D00 , 32'h067DAA40 , 32'h0C98E070 , 32'hE27782E0 , 32'hD2B4C900 , 32'h0E483E10 , 32'hEDA92740 , 32'hFCA825B0 , 32'hFCC03DC4 , 32'h2C9E32C0 , 32'hBAA76080 , 32'h1260CD20 , 32'h0A0D3780 , 32'hEFF38440 , 32'h1623EE80 , 32'h01BCE670 , 32'hEEF78020 , 32'hF00C18E0 , 32'h12F210C0 , 32'hFD833794 , 32'hFEB7B9F0 , 32'hF3349D40 , 32'hEC80A520 , 32'hDD50C280 , 32'hF9263FE0 , 32'hFDF8FAF0 , 32'hF97FF610 , 32'h03F75F1C , 32'h0182BCC8 , 32'h0296C4D4 , 32'hFA3E3E40 , 32'hF9668E60 , 32'h21BEA840 , 32'h07F11B20 , 32'h1B1D29C0 , 32'hF7C2CF50} , 
{32'hEEAC7E20 , 32'hCB39B580 , 32'hD5844EC0 , 32'h0DDA1A80 , 32'hDC5B9E80 , 32'hE9133700 , 32'hF7D9C100 , 32'hE44603C0 , 32'h001C1927 , 32'hEFF9DBA0 , 32'hEF5F5FA0 , 32'hF1DB0E30 , 32'h08B3FA80 , 32'h094F4AB0 , 32'h0BC33960 , 32'h0CF5D130 , 32'hF8AEBA70 , 32'hED479500 , 32'hE82242C0 , 32'hE8DFBFE0 , 32'hF9306798 , 32'h0D4B5700 , 32'h00F8D89F , 32'h05BD4EF0 , 32'hED1B28A0 , 32'h010B464C , 32'h028F2618 , 32'h119EDC80 , 32'h07AEE698 , 32'h07AA55C8 , 32'h05C36648 , 32'h1AE1CEC0 , 32'hF7A780E0 , 32'h0E9449B0 , 32'hF77111A0 , 32'hF3F26DA0 , 32'h01A7CDF0} , 
{32'h034F653C , 32'hF59497B0 , 32'h05738ED0 , 32'h0F4F12B0 , 32'hF11A6080 , 32'hFB0388A8 , 32'hE15F5FA0 , 32'hD5C8D180 , 32'hF5C50ED0 , 32'hEDB34820 , 32'hBF009600 , 32'hFCF2AD98 , 32'hF3C39B40 , 32'hF0A94B10 , 32'hFAB94DC8 , 32'h28C591C0 , 32'h0DF1F9B0 , 32'hD2150980 , 32'hBFBDD480 , 32'hFAA92960 , 32'hD4968BC0 , 32'h140CA400 , 32'hFDE74E14 , 32'hDF259F80 , 32'hFBA1C560 , 32'h2261C600 , 32'hF32D5390 , 32'h01083148 , 32'hE995DFA0 , 32'h05D6B328 , 32'hF27EC500 , 32'h0947B740 , 32'hE5085280 , 32'h0C846C40 , 32'hEFCBA600 , 32'h0470B308 , 32'h07948F40} , 
{32'hF37CE3E0 , 32'h0199F70C , 32'hE27C0C60 , 32'h0B83D5B0 , 32'hDD37E7C0 , 32'hFF60FE4C , 32'hFABF0FF8 , 32'h00552564 , 32'hFA3B10D0 , 32'h114B6A00 , 32'hE1F79F80 , 32'hF7687920 , 32'hC1E57B40 , 32'hF82F7058 , 32'h0500A158 , 32'hEFB578E0 , 32'h14AD5160 , 32'hF6626C10 , 32'hE0076E00 , 32'h05A41EB0 , 32'h0B2210E0 , 32'h279EC240 , 32'hFA700E58 , 32'hF2F14780 , 32'h05224240 , 32'h13454B40 , 32'hEC388F40 , 32'h04D154C0 , 32'hEFDFDE20 , 32'hEBF71DC0 , 32'hF0EC37A0 , 32'hCE06F9C0 , 32'h0370C9FC , 32'hE1DEC560 , 32'h0083C6FD , 32'hF5C36BA0 , 32'h1883B5E0} , 
{32'hF820D590 , 32'h049A0F98 , 32'hF017F3E0 , 32'h0FE07A00 , 32'hEEAD7C40 , 32'h130DB0E0 , 32'hEC7183C0 , 32'h1943A280 , 32'h08368150 , 32'h16907B20 , 32'hECD82780 , 32'hF7FE7070 , 32'hDCF558C0 , 32'hEC500BC0 , 32'h0C1FF720 , 32'h0A90F1A0 , 32'h19A6CB40 , 32'hE1210AA0 , 32'h0D417AD0 , 32'h012DD300 , 32'h38DD9700 , 32'h00A5048B , 32'hE2956D80 , 32'hE3CA1340 , 32'h1DA68F60 , 32'hF23F3B70 , 32'hEF7A6260 , 32'hFA4F7C10 , 32'hF3346670 , 32'h038EA308 , 32'h019A0F34 , 32'hEEDE2260 , 32'h25522700 , 32'h213727C0 , 32'h02C95664 , 32'hFEB7FC0C , 32'h0E791580} , 
{32'hF1A18A80 , 32'h06B34DF0 , 32'hF5A24C30 , 32'h0DFB0280 , 32'hFB5677A8 , 32'h0C1FFCE0 , 32'hF7603280 , 32'h038C3210 , 32'hFEF73360 , 32'h05A4D140 , 32'hFE4B5F80 , 32'hFD014B94 , 32'hFB650E30 , 32'hF15AAFE0 , 32'h05CEE900 , 32'h06B0E040 , 32'h0B827940 , 32'hF6064C70 , 32'h0E0DE0F0 , 32'hFF992B4B , 32'h168020C0 , 32'hF29D45D0 , 32'h06F3B7F8 , 32'hF7A4C1B0 , 32'h061136A8 , 32'hFDA5F3C8 , 32'hFC558BDC , 32'hF1315FA0 , 32'hFC6FFB2C , 32'h0054C6E6 , 32'hFA921100 , 32'hEDDF38A0 , 32'h192EBD20 , 32'h02B750D8 , 32'hE2F01E00 , 32'h0BED6520 , 32'h07571A70} , 
{32'h14430420 , 32'h0248AB40 , 32'hEF9B25E0 , 32'h301B4440 , 32'hED9F1500 , 32'hF0B3A130 , 32'h10001540 , 32'h41884B00 , 32'h0ADB15F0 , 32'h23183AC0 , 32'hF0CB6620 , 32'h0D4FB970 , 32'h1BBD66A0 , 32'h03175480 , 32'h148FBA00 , 32'h15BA7620 , 32'hEE92B5A0 , 32'hFB8A35A0 , 32'h03F33208 , 32'h1E1B9700 , 32'h128EFFA0 , 32'hFE5768C0 , 32'h032C0980 , 32'hFA114E80 , 32'hF45B1F10 , 32'h39117900 , 32'hE7636200 , 32'h04F43CB0 , 32'hFB631CF8 , 32'h1E4A9900 , 32'hFD96D428 , 32'hF2E58690 , 32'h0FF11BE0 , 32'h13B79240 , 32'hFA85E828 , 32'h0D34FCA0 , 32'h0294E88C} , 
{32'h007EFB12 , 32'hECF37CE0 , 32'hEEBC33E0 , 32'h29DA6780 , 32'h0D6157B0 , 32'h005C5D72 , 32'hF945AE08 , 32'h413D2A00 , 32'h1A319AE0 , 32'h214FF640 , 32'hE92D9080 , 32'hF3D96AF0 , 32'h310E72C0 , 32'hDE4F1440 , 32'hD9943C40 , 32'h10679440 , 32'hF5DD1B90 , 32'h07B8E968 , 32'h161DAD60 , 32'h206CB1C0 , 32'hEC881220 , 32'hECF74D40 , 32'h1C5444E0 , 32'h0A624120 , 32'h0AF18780 , 32'hE7A131A0 , 32'hFE95B4F4 , 32'h08F51200 , 32'h0AB0B9F0 , 32'h007D999E , 32'hFB984688 , 32'h19CFB320 , 32'hFD4BD1A0 , 32'hEFF7A4E0 , 32'h0096210B , 32'h0D43F810 , 32'hF440AE80} , 
{32'h0B9D3F10 , 32'hFC514168 , 32'hF899E6C0 , 32'h0DABA220 , 32'hF66EF450 , 32'hFA669AD8 , 32'h041F07F8 , 32'h1E234780 , 32'h0D87E4C0 , 32'h0586C2E8 , 32'hE5CD7160 , 32'hF83B95F8 , 32'hF8BAA480 , 32'hF1DF13A0 , 32'hF755D130 , 32'hF9244250 , 32'hF269B6E0 , 32'hF732DB20 , 32'h05FB1AD0 , 32'h0BD29000 , 32'hF3968A00 , 32'hF9FB09F0 , 32'hFE432D40 , 32'h0878DCA0 , 32'hFA709A30 , 32'hF9EB2F78 , 32'h04FDB070 , 32'hFE1ECBA8 , 32'h0A53C620 , 32'h01706A0C , 32'hFBD9F488 , 32'h00F0192B , 32'h000CABA0 , 32'hF56CCD90 , 32'hFE596D28 , 32'hF606AAC0 , 32'h0E82E450} , 
{32'h18E9AA80 , 32'hF5D18A90 , 32'h0403E880 , 32'h04A7A520 , 32'hF3744EA0 , 32'hF6CD37E0 , 32'h00335D12 , 32'h17C62980 , 32'h0E134550 , 32'h00B35D71 , 32'hEF2AA5A0 , 32'hFCC4F398 , 32'hFF532399 , 32'hF86A5000 , 32'hFDBA2174 , 32'hFCFC2E58 , 32'hF2333FB0 , 32'hF4A1EF40 , 32'h095F0E20 , 32'h19976B80 , 32'hF399DD30 , 32'hF3E9A470 , 32'hFD3D2B70 , 32'h09E512F0 , 32'h0D486E10 , 32'hFD830EA4 , 32'h0E2C9720 , 32'h04B239A0 , 32'h02164108 , 32'h08613030 , 32'hFECB9074 , 32'h0ED6F4F0 , 32'hF7089ED0 , 32'hF1C1AF50 , 32'h03949834 , 32'h013B7E68 , 32'h0E286640} , 
{32'h062BE158 , 32'h0E018500 , 32'h0ADE3150 , 32'hECE3BF00 , 32'hEF9DB3E0 , 32'h04A69A48 , 32'h12061C40 , 32'h158EF7A0 , 32'hF5561C10 , 32'h08E2B460 , 32'h0375A67C , 32'hF30AA9F0 , 32'h0DAF45B0 , 32'h08856DD0 , 32'hE92F2C60 , 32'h015B6754 , 32'hF2D55D10 , 32'hDAED98C0 , 32'hE8189B20 , 32'hFB1DA030 , 32'hFDE37EE8 , 32'hF5BE57D0 , 32'hF4044620 , 32'h1A459980 , 32'h10C187C0 , 32'hF63F0A30 , 32'h08564510 , 32'hF69308F0 , 32'hEFAD6940 , 32'hF7F5AAB0 , 32'hFA670F70 , 32'h1703D0C0 , 32'hF8BB7F98 , 32'hF2DEFA70 , 32'hFD2BC9B8 , 32'hFEEA31A8 , 32'hFD46E40C} , 
{32'hF98C8210 , 32'hF5D04CC0 , 32'h045565E0 , 32'h02795520 , 32'h01395584 , 32'h017893A4 , 32'h01DAE3A4 , 32'h02FD9C8C , 32'hF5C9E7E0 , 32'h02C834AC , 32'hF1BDC7E0 , 32'hE940FAE0 , 32'h05047D78 , 32'hFB448F00 , 32'h136BC560 , 32'hE8599D60 , 32'hE8E52AA0 , 32'h10E92780 , 32'hF8447588 , 32'h03EE8DC4 , 32'hF9F1C688 , 32'hE76DB5E0 , 32'h019C517C , 32'hF0549630 , 32'h11DEEEA0 , 32'h062633B8 , 32'h0DCF7920 , 32'hF6756890 , 32'hFA3AFB98 , 32'hEF4052A0 , 32'hF5F29F00 , 32'hF9B1A0D0 , 32'hF5F3D8E0 , 32'h0C7E3530 , 32'hFEE9A014 , 32'hF2683CB0 , 32'hFB9A9CC8} , 
{32'h0000AC24 , 32'h00014649 , 32'h00018DA6 , 32'h000363C0 , 32'hFFFF7885 , 32'hFFFD9889 , 32'hFFFDCB3E , 32'h0000332E , 32'hFFFE3924 , 32'h00002AF2 , 32'h00019B00 , 32'hFFFFFB43 , 32'hFFFF13BE , 32'h0000BBB6 , 32'h00012E79 , 32'h00003D12 , 32'hFFFDB03D , 32'hFFFF5759 , 32'hFFFF5A53 , 32'hFFFDB786 , 32'hFFFDAA18 , 32'hFFFCA94B , 32'hFFFF6595 , 32'h00043B65 , 32'h000057A2 , 32'hFFFE0CB2 , 32'hFFFD6659 , 32'h00039155 , 32'hFFFE2CCB , 32'h0000C001 , 32'hFFFFBA0E , 32'h00012264 , 32'hFFFE8994 , 32'h0004B27C , 32'h00027228 , 32'hFFFC11A8 , 32'h0000DAA5} , 
{32'h000B3C53 , 32'h00044624 , 32'hFFF2B640 , 32'h000B12C2 , 32'hFFFBC0DC , 32'h00025BEE , 32'h0002B34C , 32'hFFF3CC10 , 32'hFFFC7661 , 32'hFFF9BFE5 , 32'hFFFEBE3D , 32'hFFF84293 , 32'hFFFDFCDC , 32'h0006BA8A , 32'hFFF33FEF , 32'hFFFBFCCD , 32'h0001D319 , 32'h0003DBF2 , 32'hFFF90169 , 32'hFFFFC12F , 32'h00020A93 , 32'hFFFCB042 , 32'h000E1F82 , 32'hFFFC2984 , 32'hFFFF2DCD , 32'h00010FDF , 32'hFFFEC9CA , 32'hFFF70DA9 , 32'hFFFB2A9C , 32'hFFFE10BB , 32'hFFF073EB , 32'h00009473 , 32'h00090B9F , 32'h00012CC6 , 32'hFFFBF3DD , 32'h00043949 , 32'hFFFB49BF} , 
{32'h000117BB , 32'h0000CD36 , 32'hFFFBE9E7 , 32'hFFFEB2CA , 32'h000020CB , 32'hFFFE502B , 32'hFFFBA30B , 32'hFFFDCEA0 , 32'h0000C21A , 32'h00043995 , 32'h00022E27 , 32'h00054DE5 , 32'h00043C94 , 32'hFFFE4B7B , 32'hFFFFFF72 , 32'hFFFE6937 , 32'h00028A8E , 32'h0003A3FF , 32'hFFFF2BD0 , 32'hFFFB7615 , 32'h00018440 , 32'hFFFF0B48 , 32'hFFFD40AB , 32'h0003FE25 , 32'h00053394 , 32'hFFFC945F , 32'h00034B7D , 32'h000086D4 , 32'hFFFC1E93 , 32'h00038D55 , 32'h00003D9A , 32'hFFFEFB16 , 32'hFFFF6DF1 , 32'hFFFFD634 , 32'hFFFBA08A , 32'hFFFD225C , 32'h00040F30} , 
{32'h0000E998 , 32'hFFFF8D74 , 32'h000196F6 , 32'h000524D8 , 32'hFFFEFBEE , 32'h00019EF4 , 32'hFFFF6554 , 32'h00009B11 , 32'hFFFDA4A5 , 32'hFFFD504D , 32'hFFFB1564 , 32'h0001F00A , 32'hFFFACC4D , 32'hFFFFFF4C , 32'h0002AEDA , 32'hFFFC6A13 , 32'hFFFE8DC5 , 32'hFFFCD17B , 32'hFFFAAC2D , 32'h000686A0 , 32'h000813DF , 32'hFFFE481E , 32'hFFFDB565 , 32'h00052BBF , 32'hFFFB9A44 , 32'h00053AA5 , 32'h00007271 , 32'hFFF6AB6E , 32'h00005F4A , 32'h0003C921 , 32'h00032EC2 , 32'hFFFE57D8 , 32'h000163BD , 32'hFFFEE9A9 , 32'hFFFF9EAB , 32'hFFF6121A , 32'hFFFCE2C2} , 
{32'hFFFF0C75 , 32'hFFFFA53B , 32'h0001D301 , 32'hFFFF2A4D , 32'h000367F8 , 32'hFFFB6ADA , 32'hFFFF377C , 32'hFFFF96F9 , 32'h00010DD9 , 32'h00070826 , 32'hFFFFF364 , 32'h00015475 , 32'hFFFBEBA7 , 32'hFFFE3E33 , 32'hFFFDFA38 , 32'hFFFFB464 , 32'hFFFEBBC2 , 32'h00009D3A , 32'hFFFD53EE , 32'hFFFC5D02 , 32'h0001F0FB , 32'hFFF6EEBC , 32'h0002CF9B , 32'h00036D9B , 32'h000415F9 , 32'h000604B5 , 32'hFFFE248B , 32'hFFFDD53C , 32'h0002653A , 32'hFFFF7AE2 , 32'h00015265 , 32'h0002CBEE , 32'h00094943 , 32'hFFFBDFE0 , 32'h00004CE7 , 32'h0001B29A , 32'hFFFFF216} , 
{32'h0005877D , 32'h0005FFA4 , 32'h00093E78 , 32'h000130A5 , 32'h000BE082 , 32'hFFFE0D5C , 32'hFFFBB912 , 32'hFFFF8D7C , 32'hFFFF09E0 , 32'hFFFED705 , 32'hFFFC2962 , 32'h0008348C , 32'h0001A1E9 , 32'hFFFF8906 , 32'h000055EA , 32'hFFFFC6DA , 32'h00018FC8 , 32'h00047658 , 32'hFFFDA362 , 32'h00034FB2 , 32'hFFFAD602 , 32'h000273B8 , 32'h00032F3D , 32'h00075DC8 , 32'h0004F72D , 32'hFFFBFFD0 , 32'h00037F5F , 32'hFFFCEE85 , 32'h00003D33 , 32'hFFFCE998 , 32'hFFFE0381 , 32'h000164F8 , 32'h00020E6B , 32'h0000A9C5 , 32'h0000CC62 , 32'h00029B2B , 32'hFFF940A8} , 
{32'hFFFA4E53 , 32'hFFF6B7D6 , 32'hFFF89111 , 32'hFFFEAA63 , 32'hFFF6F68D , 32'hFFFC7024 , 32'hFFF80C68 , 32'h0000538A , 32'hFFF8FEA2 , 32'hFFFBD1E7 , 32'hFFFE6F4E , 32'hFFFBC49A , 32'h0003460E , 32'h0000B87E , 32'hFFF8D078 , 32'hFFFD1BE7 , 32'h000290CF , 32'h0002C608 , 32'hFFFFEDC0 , 32'h00064E96 , 32'h0003915C , 32'hFFFEA16C , 32'h00037C67 , 32'h0000F737 , 32'hFFF94DE2 , 32'hFFFCB8A1 , 32'h0001AF98 , 32'h00055B8E , 32'hFFFFFE36 , 32'h00027B10 , 32'h00008E69 , 32'hFFFEC386 , 32'h0001249F , 32'h000302AD , 32'h00033376 , 32'hFFFA0B26 , 32'hFFF952C8} , 
{32'h02BE8E0C , 32'h0209FB8C , 32'hFFB698C3 , 32'hFDF8310C , 32'h0439F1C8 , 32'h00D59874 , 32'h053EC460 , 32'h04B78FA8 , 32'h02634914 , 32'hFEF72F24 , 32'h08CBFF00 , 32'hF6BBA880 , 32'h048975A8 , 32'hFC65C968 , 32'h03434CB8 , 32'hFB1889A0 , 32'h029ADC7C , 32'hF908BDB0 , 32'h030AF544 , 32'hF997F370 , 32'hFF08AFB3 , 32'hFE9A24E0 , 32'h036D3BA8 , 32'h04056F70 , 32'hFFD68BCB , 32'h01C0436C , 32'hFE0A29F0 , 32'h043B0F60 , 32'h0AC048C0 , 32'hFE74BC94 , 32'h0657E8B0 , 32'hF86AEAC8 , 32'h07279D78 , 32'hF9E12088 , 32'hFAA9C058 , 32'h01D5DC64 , 32'h00C1261F} , 
{32'h24BAAAC0 , 32'hFFDA12BD , 32'hF6C00A80 , 32'h1FB59300 , 32'h070B6D38 , 32'h0AD11BA0 , 32'h1DA19620 , 32'h01D27908 , 32'hF296BBA0 , 32'h0896C800 , 32'h2A138AC0 , 32'hF813D5D8 , 32'hF691C290 , 32'hEE023460 , 32'hFBDB5B98 , 32'hF41DF870 , 32'hF554A5B0 , 32'hEE1B8F20 , 32'hFB196C18 , 32'hF9A38660 , 32'h0B005FB0 , 32'h01DACD24 , 32'h0BE37EF0 , 32'h02785090 , 32'hFEBC5370 , 32'h1487B900 , 32'hE33E0360 , 32'h166FA100 , 32'h12657780 , 32'hE4D29860 , 32'h15E21260 , 32'h07CA7960 , 32'hE6019EE0 , 32'h0B5C4270 , 32'hF83F8C58 , 32'h02009A6C , 32'h19246E40} , 
{32'h1A4F2E40 , 32'h1D160A20 , 32'h0078257A , 32'h14C50960 , 32'h2170EB00 , 32'hFF499E57 , 32'h39025100 , 32'h048477C0 , 32'h0A54CE90 , 32'h028802D0 , 32'h0746AB28 , 32'h15B5A340 , 32'hF5402340 , 32'hEFB0A0C0 , 32'h093BBBE0 , 32'hED4158E0 , 32'hEB8DC6E0 , 32'hE9A9E9E0 , 32'hFD360310 , 32'hF922AF50 , 32'h09C52040 , 32'h0033F4D4 , 32'h01244B1C , 32'hFFF9BCC8 , 32'hFBB09E60 , 32'h06A400D8 , 32'hF023B1C0 , 32'h00C5F9F5 , 32'h09211A00 , 32'hF06490A0 , 32'hFDDD1860 , 32'h1DE09160 , 32'hE5A90E40 , 32'h056371B0 , 32'hEB8FB640 , 32'h0A110D50 , 32'h1D311D00} , 
{32'h03D5C130 , 32'h16D11F00 , 32'h0AF4F900 , 32'h1FEDFD60 , 32'h0DF6EED0 , 32'hE6BE4540 , 32'h34650CC0 , 32'hF66B7860 , 32'h1A86A4E0 , 32'h037EDEEC , 32'h13D32D80 , 32'h06DD9CB0 , 32'h01FD7020 , 32'hE89F6DA0 , 32'h02FCE3AC , 32'hEA443920 , 32'hF335D550 , 32'hE1F07200 , 32'hFAEAA448 , 32'h0181B000 , 32'hFE44CEFC , 32'hF6C42A90 , 32'hFFF9E91C , 32'h00D19703 , 32'h0895E650 , 32'h09E46C70 , 32'hF8B18298 , 32'h0A0C4660 , 32'hF56CB3E0 , 32'hF65282D0 , 32'hF6EC46A0 , 32'h11F08160 , 32'hF30E3230 , 32'h1BE8F240 , 32'hF5E836B0 , 32'h056709F8 , 32'h19A763A0} , 
{32'h07A860F0 , 32'h1D4EC9A0 , 32'h19190C80 , 32'h15C097E0 , 32'h1A113020 , 32'hFE26574C , 32'h2FDB9100 , 32'h06F90CB0 , 32'h12B3FEA0 , 32'hFF34FC73 , 32'hFB47F4A0 , 32'h1F20E040 , 32'hFCCA1D4C , 32'hEFFAF9C0 , 32'h056F7940 , 32'hF259B750 , 32'hF942B0E0 , 32'hEF5D87C0 , 32'hFB0BC148 , 32'h02E31574 , 32'h02770374 , 32'hF9E91C80 , 32'hF1FD6CB0 , 32'hF9AEADB0 , 32'h0316C678 , 32'hFB198320 , 32'hFC0707D0 , 32'hFD7E9844 , 32'hFE9D4C28 , 32'h0AA109F0 , 32'hF5D78570 , 32'h0EFC79F0 , 32'hFAF83F80 , 32'h0FAF1410 , 32'h045C5D98 , 32'h13062F60 , 32'h00C598E7} , 
{32'hF51AE0C0 , 32'h12475100 , 32'h15F540A0 , 32'h13F34AC0 , 32'h0007F034 , 32'hED7B96A0 , 32'h1CDCD780 , 32'hFD3E4F8C , 32'h1E8D17A0 , 32'hF838AAC0 , 32'h1E5FDE60 , 32'h08E49350 , 32'hF13050A0 , 32'hE98563A0 , 32'h0F0F5AC0 , 32'h063B4338 , 32'hFA7CC120 , 32'hF948EFD8 , 32'hFC0B5A74 , 32'h118F8AA0 , 32'hF2058C80 , 32'hF4666E30 , 32'h08AF5880 , 32'h041BAE40 , 32'h114FE480 , 32'hF562DF00 , 32'hF1D6CF50 , 32'h021130C0 , 32'hFCCD8784 , 32'hF8760E28 , 32'h078AA198 , 32'hEF734180 , 32'h0311F3B4 , 32'h0B493BA0 , 32'hFDCD3E6C , 32'hF2AA1240 , 32'hF9997588} , 
{32'hF0B43F70 , 32'h0706D4F8 , 32'h2F761AC0 , 32'h17158220 , 32'h11A61AA0 , 32'hE6E88200 , 32'h02CF73C0 , 32'hF81189F0 , 32'h127B77C0 , 32'h03D2B298 , 32'h028F5C78 , 32'hF6F227D0 , 32'hF9A217D8 , 32'hE61D06C0 , 32'hFED18194 , 32'h0E5A59B0 , 32'hF7E495B0 , 32'hEC3B19E0 , 32'hFBB06A90 , 32'h02F886F8 , 32'hF12053C0 , 32'h02525DF0 , 32'h048EA760 , 32'h0DD77950 , 32'h01332D58 , 32'h05EF6458 , 32'hEF20CCE0 , 32'hFCB35814 , 32'hF26141E0 , 32'hFF83B548 , 32'h0CFBAA00 , 32'hE4673940 , 32'hFD4F07A4 , 32'h0590F488 , 32'h032D5B18 , 32'hFFFC2143 , 32'hF0F2B620} , 
{32'hD3480B80 , 32'hF2424190 , 32'h2B847C80 , 32'h21DA6CC0 , 32'h04709818 , 32'hE1532300 , 32'hFF9E8ECB , 32'hEF7757A0 , 32'h03E9A104 , 32'h092AC690 , 32'h1B1CB100 , 32'hD4914B40 , 32'hFCD09284 , 32'h0CCA54B0 , 32'h049FE400 , 32'h1DABE5E0 , 32'hFAEDDC38 , 32'h10AB3280 , 32'hEFFED260 , 32'h1F92C1A0 , 32'h0BD5DD60 , 32'h0034E47A , 32'h06B70AB8 , 32'h07588CB0 , 32'h0EA9A4E0 , 32'h15CD9E60 , 32'h031ACBE8 , 32'hF95C7558 , 32'h19ED4AE0 , 32'h041AF790 , 32'hF098D9B0 , 32'h044925C0 , 32'hF78D8CE0 , 32'hE9BD5F40 , 32'hF78922B0 , 32'hFBD92AA0 , 32'h0E8E4DB0} , 
{32'hDB04FE00 , 32'hDBC9A7C0 , 32'h23CEDD00 , 32'h0C2F2580 , 32'hF8A06570 , 32'hE6990660 , 32'hE7705DC0 , 32'hF8A57B70 , 32'hF26CACC0 , 32'h079AF3B8 , 32'h10A70D20 , 32'hE090A9A0 , 32'hF28EB2B0 , 32'h0C198A90 , 32'h198AB300 , 32'h106BDA20 , 32'hE55B26E0 , 32'h1CC089E0 , 32'hFD612064 , 32'h0D010670 , 32'hF88C8B18 , 32'hFA0DBF70 , 32'hF6ACC6B0 , 32'hFBB40408 , 32'h0FDAD2D0 , 32'h126C4360 , 32'h00283C27 , 32'hFB197A40 , 32'h14BCA080 , 32'h0CA93660 , 32'hF9FC5118 , 32'hF15299E0 , 32'hF2588590 , 32'hF79D9460 , 32'h061C7EC8 , 32'hFE2953B8 , 32'h03ADD360} , 
{32'hE5048EE0 , 32'hD9D30E80 , 32'hCBB023C0 , 32'hF5CBF9F0 , 32'hC25D4580 , 32'hDB999980 , 32'hF90BA660 , 32'hFB9BEE48 , 32'h0E4DE7B0 , 32'hF32DE940 , 32'h0728F7C8 , 32'hE2C8A100 , 32'h08FC96A0 , 32'h1A520420 , 32'h15B47D60 , 32'h0652F998 , 32'hFAA48BA0 , 32'hF7B4BC10 , 32'h086997A0 , 32'hF0F73740 , 32'h02F39F78 , 32'hFBEAC908 , 32'h024C7918 , 32'h117D7D60 , 32'hE4CF8E60 , 32'hF584A900 , 32'hFF6349AC , 32'h1330F2A0 , 32'hFF69D022 , 32'h134D86E0 , 32'h020C60D8 , 32'hF9058468 , 32'hEBBF1DE0 , 32'h1D86E540 , 32'h00000B0B , 32'h29515E40 , 32'hF71A9030} , 
{32'hE5A5F600 , 32'hE0C3D000 , 32'hE32AB840 , 32'hFACE0558 , 32'hC2A65C00 , 32'hF0F68550 , 32'hFE48475C , 32'hD1B8FD40 , 32'hFDF997FC , 32'hFF05712B , 32'h00BADF2C , 32'hF8BBF950 , 32'h0ACB8680 , 32'h14A70F80 , 32'h2F4C2AC0 , 32'hEA0061E0 , 32'h052B2EF0 , 32'hD768EA40 , 32'hF855EFD8 , 32'h1128B860 , 32'hEEF123A0 , 32'h040C63F8 , 32'h048FA9D8 , 32'hF92171F0 , 32'hEA68E3E0 , 32'hFFA8AD2C , 32'hFFDE01EE , 32'h21189A40 , 32'h0D19B3C0 , 32'hF67F4500 , 32'hDFF14980 , 32'h01B45914 , 32'hF48C1D00 , 32'hE8C03B80 , 32'h0274554C , 32'hF5942F60 , 32'hFDCB52A8} , 
{32'hF44F9C10 , 32'hFDAE2058 , 32'hF09124D0 , 32'hFE9D1AD4 , 32'hE46BE480 , 32'h099EF780 , 32'hFE2A1874 , 32'hEF086CE0 , 32'hFA16E2E0 , 32'h0A3575C0 , 32'hF3DA97C0 , 32'h07D9B6D0 , 32'hF7EF2220 , 32'h00EF7F87 , 32'h2AA5DFC0 , 32'h0394CF44 , 32'h0CE77C90 , 32'hFE25F3D4 , 32'hF1F22D20 , 32'h06AEF030 , 32'h017C9D78 , 32'h0D74E300 , 32'hFCE53550 , 32'h0AAD9900 , 32'h025A37C4 , 32'h12A3FBA0 , 32'h05BD9B80 , 32'h09188490 , 32'hEC379D60 , 32'hFA312508 , 32'hF697CAA0 , 32'h0DBDCFC0 , 32'hF4CD8F60 , 32'hE4131CA0 , 32'hF430B5D0 , 32'h0449FD28 , 32'hF9A0DD88} , 
{32'h005DA546 , 32'hFF0F1C45 , 32'hF3E55CA0 , 32'h150C1DE0 , 32'hF864C0E8 , 32'hFFE010C7 , 32'hF1854FC0 , 32'hE02E7BC0 , 32'hFAC658C0 , 32'hF33298B0 , 32'hEFFF3320 , 32'h088A9DF0 , 32'hE6C74880 , 32'hFBE2AF70 , 32'h11E6C400 , 32'h08A12690 , 32'h16FF9EC0 , 32'h05A952B8 , 32'hFE59E6F0 , 32'h070E8360 , 32'h06B40038 , 32'h09290840 , 32'hEF8D4D00 , 32'h0D30E070 , 32'h1C591700 , 32'h0F3B5F20 , 32'h031B43D4 , 32'h024040BC , 32'hE6BDE3C0 , 32'h01FC7B98 , 32'hFCF71644 , 32'h00734CC4 , 32'hF2037580 , 32'h04741298 , 32'h0B047190 , 32'hF199D740 , 32'hF5FB0820} , 
{32'hF0793550 , 32'hFFD85370 , 32'hFC19D58C , 32'h093464C0 , 32'hF4350030 , 32'h0FE77680 , 32'hF8A3AB58 , 32'h03A7E638 , 32'hF95297F8 , 32'h0ED40200 , 32'hF6384E20 , 32'hFD33F2A4 , 32'h011010D0 , 32'h007420E6 , 32'h1C5F9100 , 32'h0F1BCCE0 , 32'h1BD334C0 , 32'hEC58F460 , 32'h06179408 , 32'h08859830 , 32'h270A8940 , 32'hFD478680 , 32'hF6705CC0 , 32'h0FFE0D50 , 32'h25A58640 , 32'h033D3598 , 32'hEC626F60 , 32'hFC0708BC , 32'hF6DCAFE0 , 32'hFD3F3190 , 32'h04E35F28 , 32'h11BF5B00 , 32'hFD932B88 , 32'hFCBA88B0 , 32'hFEBA2A5C , 32'h04B880D8 , 32'h0BBEE200} , 
{32'hFA876598 , 32'hFEB6ABFC , 32'hFFDA9893 , 32'h0FE48A90 , 32'hFEFC02DC , 32'h02DBA480 , 32'hF8D596B8 , 32'h05C66E48 , 32'hFDCD5F8C , 32'hFF7ECD4B , 32'hFDE7C4CC , 32'h01FEE2F8 , 32'h08EB51D0 , 32'h042E3C00 , 32'h0C553E30 , 32'h0E6D5CD0 , 32'h067BDE58 , 32'h0431F0F8 , 32'h0AA19B10 , 32'h0655B378 , 32'h0F33E7D0 , 32'h06BCC320 , 32'h03F720E0 , 32'hFC68D33C , 32'h0E195D40 , 32'h0C2B6E20 , 32'hF8F1ACC8 , 32'hF911CD40 , 32'hF5943BC0 , 32'hFF9159E0 , 32'hFAAC50D0 , 32'h01C40E6C , 32'hFB910DC0 , 32'h0214361C , 32'h052DFFF0 , 32'h02CC10B8 , 32'hF9A49FF0} , 
{32'hFDA73668 , 32'h05EFFE00 , 32'hF69F6360 , 32'h13E5F6E0 , 32'hF8477FD0 , 32'h07DE7D40 , 32'hEDD70060 , 32'h374E7680 , 32'hFCBFAB84 , 32'h02958724 , 32'h126282A0 , 32'h07EE3CF0 , 32'h45587A80 , 32'h19008420 , 32'hFDC5D758 , 32'h194F2B60 , 32'hF6788A00 , 32'hE27549E0 , 32'h2777B900 , 32'h0D020250 , 32'h0D57F480 , 32'hE9947E20 , 32'h0B331AB0 , 32'h1382AA60 , 32'h073FD5E8 , 32'h0B19B610 , 32'hFFE8C029 , 32'h030F1844 , 32'hF11621D0 , 32'hFE32BC98 , 32'hE7F1E4C0 , 32'hFA29AA68 , 32'h045F4B08 , 32'h11A834C0 , 32'hF8096898 , 32'hFB57CFE0 , 32'h09934640} , 
{32'hFE0D6750 , 32'hF7F3DC50 , 32'hFB33F840 , 32'h1BC3C280 , 32'hF612E380 , 32'hFCED31A4 , 32'h0CF66E60 , 32'h08A026F0 , 32'hEE4B88C0 , 32'hE33E7B20 , 32'hFC3F54B8 , 32'hF62B7E10 , 32'h12A085E0 , 32'h0A4EAF50 , 32'h02DD42A4 , 32'h0C35F4C0 , 32'hFFF68B1A , 32'hF5F4A290 , 32'hFE394D1C , 32'h011F13A8 , 32'h034D831C , 32'hF9D986D8 , 32'h0A33E750 , 32'hFBA2AD68 , 32'hFAD23F60 , 32'h097C2950 , 32'h09178180 , 32'hF6A50AC0 , 32'hF6B34D50 , 32'h0BB97DE0 , 32'h067B8388 , 32'hFAA8E188 , 32'h0D30E330 , 32'h006DDEBC , 32'hFF093CC4 , 32'hFE2922B8 , 32'h0646F228} , 
{32'h05209468 , 32'h0BB30080 , 32'h0886CF90 , 32'h03D510C4 , 32'h0157622C , 32'hFFF730B4 , 32'hFC7DE078 , 32'h0F55CD80 , 32'h0320125C , 32'h0A0D9680 , 32'h036A0C80 , 32'hF5489CB0 , 32'h12D58360 , 32'h0AA9F510 , 32'hFBE0DB08 , 32'hEDFA2A20 , 32'h0070757B , 32'hEF38C760 , 32'hF65D5FE0 , 32'h079349C8 , 32'h118DC600 , 32'hF2B4F750 , 32'h06B32FA8 , 32'h0FC46420 , 32'hFED68BF8 , 32'hE337AD20 , 32'h0548A290 , 32'h0388A9A4 , 32'hF71D90A0 , 32'h05344CF0 , 32'hFE7BE66C , 32'h027AD928 , 32'h02105358 , 32'hFD173AE4 , 32'h0269EEA0 , 32'hF83C8DC0 , 32'hF7A2EF20} , 
{32'h03F18700 , 32'hFD35FE44 , 32'hFD40D540 , 32'hFA55F2B8 , 32'hFE679618 , 32'h054D5008 , 32'hFDA0BA40 , 32'h0B5DE220 , 32'h04E88E20 , 32'hF9380D18 , 32'h04FE8888 , 32'hFDEC1EB8 , 32'h0208FAC0 , 32'hF4AF6D90 , 32'hF4F8BB60 , 32'hFA365070 , 32'hFB8E0AA0 , 32'hED8D64C0 , 32'hF48A3150 , 32'hF57B0C20 , 32'hF4B887C0 , 32'h09F6A6F0 , 32'h002D2061 , 32'hFF9FE119 , 32'h06813678 , 32'h061FAE90 , 32'hFF6DA86E , 32'h0A312B00 , 32'h0190A184 , 32'hFA142018 , 32'hFD8ACED8 , 32'hF0384E50 , 32'h067CDF98 , 32'h01B63FE0 , 32'hFA9D9E88 , 32'hFD6DC384 , 32'h0839F810} , 
{32'hFEB4BABC , 32'hE67D0C60 , 32'hFCEB69E0 , 32'h1067B380 , 32'hF883BD60 , 32'h0EAEED30 , 32'h0AECBFA0 , 32'h28C8F7C0 , 32'h1184ABA0 , 32'hFB962D18 , 32'hDA5BEF00 , 32'hF703DB40 , 32'hF099D970 , 32'hEAFC01A0 , 32'h00281F5D , 32'hD17B4E00 , 32'hE3A80DC0 , 32'hF9212088 , 32'hF314D860 , 32'hF40E7CC0 , 32'hF2633F30 , 32'hE417A7E0 , 32'hF80F9950 , 32'hF0172360 , 32'h100A1660 , 32'hFA3B9370 , 32'h292BD880 , 32'hFE3143C0 , 32'hFD02750C , 32'hE674E9E0 , 32'hFAECF3E8 , 32'hFD5122F8 , 32'hF0293510 , 32'h1A91A6A0 , 32'hFE7309E8 , 32'hFCBF57E0 , 32'h03BD2A50} , 
{32'hFDC37220 , 32'hF8FA9150 , 32'hFBAE59D0 , 32'h07BD9828 , 32'hFE5DEBF0 , 32'hFF7074CD , 32'hFDC30960 , 32'h0414EE88 , 32'h08ED5460 , 32'hFE152348 , 32'h0110B6F4 , 32'h0716CD58 , 32'hFE6D19D0 , 32'hFDD10658 , 32'h01776130 , 32'hF8BEC888 , 32'h02DBBDCC , 32'h0181AB60 , 32'hF96A4460 , 32'hF6E14240 , 32'h0767C738 , 32'h01006034 , 32'hFED72F8C , 32'h0AED9950 , 32'hFFD4EE89 , 32'h051FB138 , 32'h0AB43860 , 32'h02EA64C4 , 32'h026C0904 , 32'h00ED07CF , 32'h0088DD95 , 32'hFBC46910 , 32'hF98AFFF8 , 32'h041041B8 , 32'hFA4C1438 , 32'h03C39560 , 32'hFCA7F70C} , 
{32'h0016393A , 32'h0011EA01 , 32'hFFD476B5 , 32'h003F1641 , 32'h002C64C6 , 32'h00424C23 , 32'hFFE5372E , 32'h001AF9F6 , 32'hFFF350E7 , 32'h002DFC67 , 32'hFFDCB9C4 , 32'hFFD41F65 , 32'h00394E56 , 32'hFFEDA794 , 32'hFFDA6476 , 32'h001C84AB , 32'h00468D95 , 32'hFFC55B36 , 32'hFFE51F07 , 32'hFFE3A775 , 32'h002D7E3D , 32'h006E3E83 , 32'h0036EE73 , 32'hFFFE964E , 32'hFFE86B39 , 32'hFFB64C47 , 32'h002AA634 , 32'h0032B19E , 32'h001038CD , 32'hFFB5846C , 32'hFFFCBFD6 , 32'h003244A1 , 32'h002EAC52 , 32'hFFF6D3C4 , 32'hFFADC11B , 32'h0011E6BE , 32'h00165A53} , 
{32'h0022F935 , 32'hFFECFC9F , 32'hFFC55D09 , 32'h005EB16F , 32'h0020DAC0 , 32'h002102E8 , 32'hFFFA6A16 , 32'h0016F42A , 32'hFFD57D16 , 32'h000AEB1A , 32'hFFE22BD5 , 32'hFFDFB944 , 32'h002AE2F7 , 32'h00124FF1 , 32'hFFDFAE1D , 32'hFFF2C0F8 , 32'h0066BEA9 , 32'hFFCD4DEA , 32'hFFD1AD2D , 32'hFFCAB72E , 32'h00329049 , 32'h00915B7F , 32'h00408114 , 32'hFFFA9C18 , 32'h000548AB , 32'hFFAD7944 , 32'h001FAD52 , 32'h002B4077 , 32'h001DCE13 , 32'hFFA66997 , 32'hFFE48EFC , 32'h001C102A , 32'h0040DA60 , 32'h00033AF8 , 32'hFF9C6797 , 32'h000E0A25 , 32'h000221FB} , 
{32'hFFF9D6ED , 32'h00006C04 , 32'hFFF7BF6F , 32'h0001D455 , 32'h000313E7 , 32'h0003C3C0 , 32'hFFFA4D51 , 32'h000221C7 , 32'h0005ECF8 , 32'hFFFCBB06 , 32'h0000C88A , 32'h00012619 , 32'h000522BC , 32'hFFF9A99B , 32'h00031ABD , 32'h00011651 , 32'h0005DD1C , 32'h00033C3A , 32'h000217DE , 32'h0002892E , 32'hFFFE88D0 , 32'hFFF9239A , 32'h0002BBF5 , 32'h00003DFD , 32'hFFFED046 , 32'h00001C77 , 32'h00065CA6 , 32'h000109FB , 32'h0008986F , 32'hFFFB13D5 , 32'h0001D397 , 32'hFFFFC52F , 32'h00027D52 , 32'hFFF8B6C5 , 32'h0002B9B4 , 32'h000805DD , 32'h00058134} , 
{32'h0000DA99 , 32'h00096F89 , 32'hFFFDCF8B , 32'h00048C65 , 32'hFFFDC8E0 , 32'h00033771 , 32'h0003E025 , 32'h00001BBF , 32'hFFFF54C4 , 32'hFFF81857 , 32'hFFFAAD9D , 32'hFFFC2010 , 32'h0005500F , 32'h0003AAA1 , 32'h0005FC07 , 32'h0002F219 , 32'hFFFD0C86 , 32'hFFFFECAF , 32'h0002C58C , 32'h00015DD4 , 32'h0000714F , 32'h00059922 , 32'hFFFD5CD8 , 32'h00007496 , 32'h0002DB0E , 32'hFFFDC34A , 32'hFFFEB137 , 32'h0000A55D , 32'hFFFE5B41 , 32'h0000300A , 32'hFFFF1200 , 32'hFFF6A91A , 32'hFFFC13A0 , 32'hFFFC0855 , 32'h0000BE94 , 32'hFFFADDEA , 32'h0000AA83} , 
{32'hFFFAFBAA , 32'h00041EBD , 32'h0000EB9A , 32'hFFFB81BD , 32'hFFFC048D , 32'h00041F7B , 32'h00045DBD , 32'hFFFE1963 , 32'hFFF9F1CD , 32'h00002702 , 32'h0002F321 , 32'hFFFD328E , 32'h000443F7 , 32'hFFFFB559 , 32'h000010BC , 32'hFFFEAFF1 , 32'hFFFB4F47 , 32'h00022139 , 32'h0006323D , 32'hFFFB2093 , 32'hFFFBAD6F , 32'h00021BA2 , 32'hFFFDC4C7 , 32'h0005BA8F , 32'h000450C3 , 32'h000189A0 , 32'h0002CACF , 32'hFFFA24EE , 32'h0003D96F , 32'hFFFDE116 , 32'h00006CF8 , 32'h0006EA07 , 32'hFFFF8921 , 32'h0003FC6B , 32'h0001480B , 32'hFFFFB464 , 32'hFFFD890C} , 
{32'hFFFBE433 , 32'hFFF9ED35 , 32'hFFF43159 , 32'hFFF8DC3B , 32'hFFF540FD , 32'hFFFA84C1 , 32'h0001B4BC , 32'hFFFCC9FC , 32'hFFFF486A , 32'hFFFB7E33 , 32'h000342F1 , 32'hFFFA110E , 32'h000301FE , 32'hFFFC7D30 , 32'h0000651B , 32'hFFFA39C5 , 32'h000CCE3A , 32'h0001DB43 , 32'h0004483B , 32'hFFFB3CF3 , 32'hFFF727A1 , 32'h0000C4EE , 32'hFFFE7CB1 , 32'hFFFF1F3C , 32'hFFFC04A4 , 32'hFFF85E69 , 32'hFFFFB953 , 32'hFFFCFE96 , 32'hFFF2169B , 32'h0005D6EB , 32'h000B5280 , 32'hFFFBBEDB , 32'h0003F6E2 , 32'hFFFDD4D9 , 32'h00004F47 , 32'hFFF8EE02 , 32'h0000D636} , 
{32'hFFFD6639 , 32'h0005D173 , 32'h000214DC , 32'h0001F37B , 32'hFFFFA56B , 32'h000160E1 , 32'h00013AA2 , 32'hFFFEA941 , 32'h0004BB9A , 32'hFFFB21C1 , 32'hFFFBFC9B , 32'hFFFCC022 , 32'hFFFB4F37 , 32'h0001063B , 32'h000268B3 , 32'hFFFEA842 , 32'h000079C1 , 32'h000156C2 , 32'hFFFAC111 , 32'h0000B525 , 32'h00022FE3 , 32'h0000F8AC , 32'h0000E4DC , 32'hFFFFDC7A , 32'hFFFC2170 , 32'hFFFE37CC , 32'hFFFFDDC4 , 32'h0003D72B , 32'hFFFF4113 , 32'h0005258A , 32'hFFFD2267 , 32'hFFFD5ED4 , 32'h00008938 , 32'h0001CF7A , 32'h000212D5 , 32'hFFFFE0AD , 32'hFFFD9722} , 
{32'h00081034 , 32'h00108683 , 32'hFFFB11E3 , 32'h00247691 , 32'hFFC1340F , 32'hFFC67D02 , 32'hFFE62FEA , 32'hFFFD1C75 , 32'h00149682 , 32'hFFEB109F , 32'h00240938 , 32'hFFFCB9A0 , 32'hFFD37A2A , 32'h000852C4 , 32'h001E9EB1 , 32'hFFF76484 , 32'hFFD3A122 , 32'hFFEC9871 , 32'h0000A87E , 32'hFFE973FE , 32'hFFE8104A , 32'hFFE83923 , 32'hFFFCB501 , 32'h001EEE11 , 32'h004588E0 , 32'hFFE1C2FF , 32'h0015BBE6 , 32'h0009A776 , 32'h000B82D3 , 32'h0032B8B5 , 32'hFFE756B7 , 32'h001E1326 , 32'h0009A08C , 32'hFFFC2BAF , 32'hFFD8CBA6 , 32'hFFF328BC , 32'h002CB21A} , 
{32'hEF21BAC0 , 32'hEB92D5E0 , 32'h143CFBC0 , 32'h11ED02E0 , 32'h194EDAE0 , 32'h02F7755C , 32'h4873EF80 , 32'h0113B174 , 32'h0CCC2110 , 32'h1313F560 , 32'h1A535C80 , 32'h189BE220 , 32'hEEFBE9E0 , 32'hF8809DC0 , 32'hEE2B45E0 , 32'hFB055360 , 32'hEBCB83C0 , 32'hD1768AC0 , 32'hFBBD7890 , 32'h03054B6C , 32'hF14F5790 , 32'hFEF25158 , 32'h0B64D5F0 , 32'hFD15DDE8 , 32'h0AE62C40 , 32'h0064D734 , 32'hEFE60DA0 , 32'hF676BF50 , 32'hE1472820 , 32'h100E1A20 , 32'hF940F318 , 32'hF756F5A0 , 32'hFE8C6ECC , 32'hFF6B1072 , 32'hF10F7E90 , 32'hEDCC1CA0 , 32'hF6F89AF0} , 
{32'hE58F3C80 , 32'hF4AB3330 , 32'h1C55E8E0 , 32'h0E8CB310 , 32'h010E42FC , 32'hFA2E6A68 , 32'h1B8CB5C0 , 32'hFDEC87C0 , 32'h0DAFBED0 , 32'h0448BE38 , 32'h0A188230 , 32'h0F3B9EA0 , 32'hF8F44FB0 , 32'hFB23C080 , 32'hF3A8B330 , 32'hFF3096F4 , 32'hFA18CDA0 , 32'hFD539C6C , 32'h00AAE0B1 , 32'hFD1A8440 , 32'hF27BA260 , 32'h04EA3A90 , 32'h08ACC930 , 32'hEAF075A0 , 32'h05B806A8 , 32'h06FEF678 , 32'hF694BC30 , 32'hF9AB7D38 , 32'hFE587E20 , 32'h04F57D18 , 32'h0AFAF9A0 , 32'hFDE5F230 , 32'h0C139600 , 32'hF515B7F0 , 32'hFF6FA5EC , 32'hF734AFC0 , 32'h0176B9BC} , 
{32'hD6F1CB40 , 32'hF525ED00 , 32'h24CDEF80 , 32'hF431D880 , 32'h15770400 , 32'hFBB86328 , 32'hFE2055C4 , 32'h0D98E6C0 , 32'h20BA3D80 , 32'hF2BBCBD0 , 32'h183A1300 , 32'h0D939E60 , 32'hED4DE5C0 , 32'hE1FBDEC0 , 32'h01D85C94 , 32'hF9BB0220 , 32'hE855B220 , 32'hFDDEA094 , 32'h07950AA0 , 32'h00A89C52 , 32'hDD0AFD80 , 32'h0CB67E30 , 32'h11D3C140 , 32'h01397B0C , 32'hF8B7D988 , 32'hFC4A0B6C , 32'hDFD6AAC0 , 32'hFC09FEF0 , 32'hEC24CC80 , 32'h06B56220 , 32'h23687E00 , 32'h1113BB20 , 32'hF8C08E40 , 32'h0A8F1B40 , 32'hF746C620 , 32'h0C21B430 , 32'hF7DE1EE0} , 
{32'hEB0ED5A0 , 32'h07079598 , 32'h24EE3E40 , 32'h0B294660 , 32'hFA762C90 , 32'hF22AED20 , 32'hFE118168 , 32'hF9EC4ED8 , 32'h18475440 , 32'hEACB1380 , 32'h2069FE00 , 32'hF827E7B8 , 32'hEC589F20 , 32'hEE923B20 , 32'hF18088A0 , 32'hEBCAF4E0 , 32'hF1B19530 , 32'hE909E980 , 32'h0824E3A0 , 32'h094E0F90 , 32'hF583D270 , 32'hF99986D8 , 32'h0E092A20 , 32'h12BEBA40 , 32'h0B0750F0 , 32'hEB2E2E80 , 32'hEB82B020 , 32'hF5CE6DA0 , 32'hEAA395E0 , 32'h1D75E640 , 32'h113291A0 , 32'hFFFCEA77 , 32'h018CA688 , 32'hFC9450DC , 32'h04A67310 , 32'hF45C4C50 , 32'hF9083170} , 
{32'hD3561B40 , 32'hFB8E3B10 , 32'h31683740 , 32'hF63F81F0 , 32'h1B8D3DA0 , 32'hEE6C4BC0 , 32'hFA9317C0 , 32'h133FDFA0 , 32'h1BFCB3C0 , 32'hF583F600 , 32'h17A01B20 , 32'h0BDB9870 , 32'hED35A720 , 32'hE3FEF960 , 32'h10E49940 , 32'hF94C7CE8 , 32'hEC90A780 , 32'hEAD47980 , 32'hF8216CD8 , 32'h08561450 , 32'hEFF2B480 , 32'hFE3D0F30 , 32'h07172788 , 32'h0BE6E490 , 32'h04725020 , 32'hFB42D518 , 32'hE3594AC0 , 32'h03134FF4 , 32'hFBD01968 , 32'hF4C40620 , 32'h19DD7660 , 32'h085B9420 , 32'hF2302C20 , 32'h1379BCC0 , 32'h148BA760 , 32'hDE90F480 , 32'hEF4DBEE0} , 
{32'hD6795480 , 32'hE7AE8840 , 32'h323C74C0 , 32'h189AC460 , 32'h0A027890 , 32'h0243E4C4 , 32'hF78B7260 , 32'hFA36AF48 , 32'hFCC48FE8 , 32'hF7F3CB30 , 32'h30DB2E80 , 32'hE16EAAA0 , 32'hF46B3EC0 , 32'h0CF9C780 , 32'h089956B0 , 32'hFBC250C0 , 32'hE88EC980 , 32'h02FF11D0 , 32'hF4DCC540 , 32'h142D3320 , 32'h0A499F00 , 32'hF8ED8E98 , 32'hFF269EA6 , 32'h0C59C600 , 32'h2AA0B380 , 32'h097AD5F0 , 32'h01418870 , 32'hF9C02FE8 , 32'h0167A0B4 , 32'h0DAE6680 , 32'hED093960 , 32'hFFBDE03A , 32'hF3149A10 , 32'hF5F5A900 , 32'h02C4F424 , 32'h0A496A10 , 32'h076AAF60} , 
{32'hD41EE740 , 32'hE6A4D720 , 32'h332EBFC0 , 32'hF286A970 , 32'h06CD1D48 , 32'h0BEBFE90 , 32'hD4B837C0 , 32'h05FE8740 , 32'h053A5308 , 32'hF1413920 , 32'h235E29C0 , 32'hE81DE460 , 32'hE8FA12C0 , 32'h03D1F40C , 32'hF77990D0 , 32'hFD1A1DB4 , 32'hF2A7A810 , 32'h0995D6E0 , 32'hE8DA37C0 , 32'hFFD24C5C , 32'h0E750170 , 32'h166C6CC0 , 32'h13750900 , 32'h179DB4E0 , 32'h1DE02A20 , 32'hFE9096A8 , 32'h1421C600 , 32'h06C00FD0 , 32'hFEB08620 , 32'h030B3274 , 32'hE37F9DA0 , 32'hFED6BA48 , 32'h04669A58 , 32'hF075E1E0 , 32'hFC5779B0 , 32'h021F1DFC , 32'h108AFDA0} , 
{32'hE304C2E0 , 32'hD2DCD400 , 32'hFA0DCC90 , 32'h04A1EDB0 , 32'hC85113C0 , 32'hF89C4DA8 , 32'hF4C68630 , 32'hF5DFEDB0 , 32'h00F5B6E9 , 32'hFD1023A8 , 32'h1DA9C160 , 32'hC76DFA40 , 32'h10A5D780 , 32'h0471BDC0 , 32'h027D1CB4 , 32'hFF7DE097 , 32'hF670C9E0 , 32'h09CCEDC0 , 32'hFDAAB118 , 32'hF5FAC110 , 32'hED9AFEE0 , 32'hFC912150 , 32'h02A1E7F4 , 32'h0828C490 , 32'h02C3E53C , 32'hFB26DAF8 , 32'h05E26B90 , 32'hF40CECA0 , 32'hD3CF6F00 , 32'h1B120700 , 32'h1B3CD2A0 , 32'hF49AE520 , 32'h0867DE60 , 32'hF02F7DF0 , 32'h0469AAF8 , 32'hF4E9B530 , 32'h0D81E340} , 
{32'hD4F10900 , 32'hCF871C00 , 32'hE4BE0E00 , 32'hF8393B10 , 32'hB3399E00 , 32'hE3546660 , 32'hF37B71E0 , 32'hF4A75DE0 , 32'h15BBC140 , 32'h0999F630 , 32'h1CB63380 , 32'hF8AD8C68 , 32'h01372BF4 , 32'h10369E00 , 32'hFB9EED38 , 32'hEC5815E0 , 32'h02518A0C , 32'hEFAA1F40 , 32'hFE39639C , 32'h0124E42C , 32'hFDCB2574 , 32'h0825DCE0 , 32'h00FFEC9F , 32'h0380A960 , 32'hFA2A1B40 , 32'h07AB7D98 , 32'h069A69D8 , 32'h0E4D3B50 , 32'hE0B7C3C0 , 32'h08621350 , 32'h13D17380 , 32'hF4AED600 , 32'hFD345408 , 32'hEE000440 , 32'h07D0BA50 , 32'h07FC9C90 , 32'h25A45F00} , 
{32'hE9968300 , 32'hEFAC2000 , 32'hF17BDBF0 , 32'hF7D66930 , 32'hCD32F6C0 , 32'hF97306F0 , 32'hF908D728 , 32'hE74136A0 , 32'h05C2D378 , 32'h0958D180 , 32'hF3307DF0 , 32'h212720C0 , 32'hF8B62920 , 32'h1112A960 , 32'h13249800 , 32'h0A58F410 , 32'h0AC87F60 , 32'hFE66BD9C , 32'h09800AC0 , 32'h121C3440 , 32'h0DFB6600 , 32'hE80CD760 , 32'h10349260 , 32'hF5BEA190 , 32'hFEF39B30 , 32'h0C279C80 , 32'hF7563CE0 , 32'h13347060 , 32'h0C623EE0 , 32'h0EA68950 , 32'h0153B9C0 , 32'h0A2FA1F0 , 32'hEBF67900 , 32'h0718BA88 , 32'hFF05B5A1 , 32'hD690D680 , 32'hFE0BAC6C} , 
{32'hFDD0865C , 32'hFA359F40 , 32'h05D76030 , 32'h08AAA600 , 32'hF04DB170 , 32'h03BE2BAC , 32'hEFCEAA00 , 32'hECC9F7A0 , 32'h004858BB , 32'h0D5CE3A0 , 32'hEDE86360 , 32'h0F2D33F0 , 32'h02639154 , 32'h00AF7235 , 32'h0F647D50 , 32'h10296940 , 32'h048B0998 , 32'hF6A1B9A0 , 32'hF7450160 , 32'h0CE588D0 , 32'hEE82FF00 , 32'h04F72A18 , 32'hFFD688A5 , 32'hFC231794 , 32'h0013A8E9 , 32'h0C9E4DA0 , 32'h00214927 , 32'h0425F990 , 32'hF3099220 , 32'h01A5EE2C , 32'hFA0E4B60 , 32'hFE445914 , 32'hF5C7E2B0 , 32'h09831310 , 32'h0557BD10 , 32'h08421010 , 32'hFF627A5F} , 
{32'hFA1DDC70 , 32'hF4C41D20 , 32'h057A77F0 , 32'h05194188 , 32'hF0839F40 , 32'h03548964 , 32'hF62423D0 , 32'hFDE604D4 , 32'hFB454EE0 , 32'h045E4B20 , 32'hFA96B248 , 32'h19DD8400 , 32'hF8895150 , 32'h0999C4F0 , 32'h0FA25E50 , 32'hFFE9FBFD , 32'h0D923AF0 , 32'hFC74CFF0 , 32'h194E4520 , 32'h023E9FB4 , 32'h06315998 , 32'hF8B822F0 , 32'h034548FC , 32'h15D74C00 , 32'h1F0C9100 , 32'h13BFEDC0 , 32'h0BFC12C0 , 32'h03CD6FB4 , 32'hEF28E5A0 , 32'h09681F30 , 32'hF23DB3E0 , 32'hF0F13DB0 , 32'hEAC9C600 , 32'h061461A0 , 32'h1EBE05C0 , 32'h0904A6B0 , 32'hF948D510} , 
{32'hF6420020 , 32'h02352568 , 32'h0266B720 , 32'h0FBFAAD0 , 32'hFEFFD2C0 , 32'h09BFE140 , 32'hF1422F80 , 32'hFC052FB4 , 32'hFFCA31D8 , 32'h07E4A588 , 32'h02D4A5F0 , 32'hFE41C788 , 32'h00D46A7B , 32'h01CF63A0 , 32'h096634A0 , 32'h0553DBA8 , 32'h1AB3A460 , 32'hF8DD6310 , 32'h093570B0 , 32'h0E6752E0 , 32'h157D2960 , 32'hF1725250 , 32'hFFF8856C , 32'hF8E3E980 , 32'h0E9BB410 , 32'hFB675D70 , 32'hFF3D6753 , 32'hF9F09020 , 32'h0012DE2C , 32'h079A0C08 , 32'h0674DAF0 , 32'h04AA3B80 , 32'hFD443DA4 , 32'hFF718935 , 32'hFDBE2C74 , 32'h0B4DEF30 , 32'hFA9CF718} , 
{32'hFA3C1ED0 , 32'hF569BE20 , 32'h02A14C90 , 32'h1D3CF780 , 32'h0244E304 , 32'h16581260 , 32'hE8335DC0 , 32'hFB17E278 , 32'hF5DE2F40 , 32'h036D1320 , 32'h0F018EC0 , 32'hFE8B9218 , 32'h0C1CCBD0 , 32'hF05B0980 , 32'hF4060F30 , 32'h05416DC0 , 32'h162BD6C0 , 32'hF3E29450 , 32'hFCFC4B24 , 32'h137C8540 , 32'h08E70FD0 , 32'h065CB7C8 , 32'h096A9AF0 , 32'hFEE6EAA8 , 32'h0C225B50 , 32'hFAD66A10 , 32'hF556F730 , 32'hF7E56110 , 32'h0518E208 , 32'hF79E4FE0 , 32'hFE7194D0 , 32'hF7DD9E10 , 32'hEC8F7640 , 32'h05DEEE80 , 32'hF3E88520 , 32'hFF27B858 , 32'h0AFBDBB0} , 
{32'hF8ED4A10 , 32'h030DCC58 , 32'h02E1CE30 , 32'h0A1EB280 , 32'h137D7900 , 32'h185C37E0 , 32'hEDD84000 , 32'h14BD06C0 , 32'h02EF0DFC , 32'hF9DFC5C0 , 32'h1C274020 , 32'hFDB5499C , 32'h39B992C0 , 32'hE996E800 , 32'hF0601660 , 32'hFF3F43F8 , 32'h16F6D940 , 32'hE95D7560 , 32'h1DB1B960 , 32'h0853B540 , 32'hFE6AFED0 , 32'h041603E8 , 32'h0CF81C10 , 32'hF4EEBC60 , 32'h07D00C38 , 32'hFE08D3D0 , 32'h20410080 , 32'h083792C0 , 32'h00CECC7D , 32'h1A16D420 , 32'h0A27BBE0 , 32'h136CC980 , 32'hEA839660 , 32'h00CDF7D5 , 32'hF94CA820 , 32'h04E0C718 , 32'hF7C7EF40} , 
{32'hFA62FB98 , 32'h0C2D1E20 , 32'h0183588C , 32'hFE23D704 , 32'h08DF83D0 , 32'h0C097720 , 32'hF7AC8910 , 32'h198E0C00 , 32'h003B3F47 , 32'h02062120 , 32'h0DDCBF40 , 32'hF0A14FB0 , 32'h2DB396C0 , 32'hF8063FA8 , 32'hF980FDF8 , 32'h00C0D192 , 32'hFA361528 , 32'hECACE340 , 32'h102BB4A0 , 32'hFA293DF0 , 32'h1547DCE0 , 32'hEF543040 , 32'h09457010 , 32'h044A2320 , 32'hF9FD4AE0 , 32'hF5123E30 , 32'hFCE09A14 , 32'h08552500 , 32'hFF3E3AD1 , 32'hFD17ACD0 , 32'hF8C90690 , 32'hFDEEC72C , 32'hFB59C460 , 32'hF8D33430 , 32'hFC92AC74 , 32'hFDCC6438 , 32'h066394A8} , 
{32'hFCF28270 , 32'hFB10BF80 , 32'hFED69E54 , 32'h0D449040 , 32'hFDF8976C , 32'hFC0ECC3C , 32'hFE36A3A8 , 32'h12CBF920 , 32'h0064029E , 32'hDDDFDE00 , 32'h0EAA1320 , 32'hF3E76480 , 32'h1604AC60 , 32'h03307850 , 32'hF4B650C0 , 32'hF896D590 , 32'h00BA08EC , 32'hF5944F00 , 32'h01037480 , 32'hE8428F60 , 32'h08060970 , 32'h068D22F0 , 32'h0CFD3390 , 32'hF9DCEA18 , 32'hF0DE0970 , 32'hFD0F608C , 32'hFFAE627C , 32'hF927EFE0 , 32'hF4395DD0 , 32'h03969A3C , 32'h054A6F88 , 32'hF38905F0 , 32'h047DD428 , 32'h00350CCD , 32'h0B12BB30 , 32'h0DAE66A0 , 32'h0971F7C0} , 
{32'hFE44E044 , 32'hF8B03D28 , 32'hFC1F0D64 , 32'h0B34AEE0 , 32'hFFAF2512 , 32'hFECC1D10 , 32'h018F3B94 , 32'h0A5BDEA0 , 32'h0AB42E00 , 32'hF3A7CF60 , 32'hFE8B73DC , 32'h0DC83440 , 32'hFDA01098 , 32'hFF24A1F1 , 32'h00CB7219 , 32'hEFC96600 , 32'h05884378 , 32'hFE07BE68 , 32'hF3F3B4E0 , 32'hF4B531A0 , 32'h074B9608 , 32'hFBE67548 , 32'h02966DB4 , 32'h0ABF33F0 , 32'hFC4F77DC , 32'h00538156 , 32'h091AE070 , 32'h04A745B0 , 32'hFE7DCAA4 , 32'h06537E80 , 32'hFF51DB1A , 32'hFECAEC88 , 32'hF9D90900 , 32'h0648DED8 , 32'h00467B24 , 32'h0B51DBD0 , 32'h01327384} , 
{32'hFBC052C8 , 32'hF66233C0 , 32'hFFA042A7 , 32'h0BE2D630 , 32'h0F4051E0 , 32'h059C0598 , 32'hFF051D53 , 32'hF6D41620 , 32'h04B7DF78 , 32'hF0A7C1F0 , 32'h0400C560 , 32'h0B809260 , 32'hF7146B60 , 32'hF3B64AE0 , 32'h093214B0 , 32'hEDB309E0 , 32'hF70F3580 , 32'h0AA568B0 , 32'h11227E60 , 32'hF86423E8 , 32'hEED7A340 , 32'h18C3D440 , 32'h0775CB18 , 32'hE51A7FE0 , 32'hF7D25AA0 , 32'h04BCAF30 , 32'h0A41EB70 , 32'hFF978A0F , 32'h07E6F2E8 , 32'h04BC12B8 , 32'hFF2A7D61 , 32'h08D607C0 , 32'h0A225ED0 , 32'h090A0160 , 32'h026E5B4C , 32'h18880A80 , 32'h082B2F40} , 
{32'hFEC8CDEC , 32'hF9575668 , 32'h03EE5488 , 32'h0383A9CC , 32'h0431DEC0 , 32'h073A65D8 , 32'hFAA08A38 , 32'h003068C3 , 32'h04597F60 , 32'hFF7A12D5 , 32'hFAB05B28 , 32'hF6E28930 , 32'hFE2DA09C , 32'h00C8EED7 , 32'h08EFB630 , 32'h06EDC338 , 32'h05734FE8 , 32'hF924F338 , 32'hFE321C0C , 32'hF7E62F10 , 32'h0C1809F0 , 32'h008186C8 , 32'h008B42B8 , 32'h02852D64 , 32'h0AD75090 , 32'hFAB3E8E8 , 32'hF4B450C0 , 32'h024680D0 , 32'h02BE7508 , 32'hF9CC85B8 , 32'h06BAE410 , 32'h07DADAD0 , 32'h04368430 , 32'h0B66BBF0 , 32'h01B775E8 , 32'h0128641C , 32'h070BF5E8} , 
{32'hFFF61746 , 32'h000EBDA5 , 32'h000B54B8 , 32'hFFFA5111 , 32'hFFF8AA50 , 32'hFFFD667E , 32'h00042FD2 , 32'hFFF5B633 , 32'h00029F2C , 32'h000A4F09 , 32'hFFFFDD14 , 32'hFFF78A42 , 32'hFFFFF676 , 32'h0006130D , 32'h00051034 , 32'h00179F9C , 32'h0001C090 , 32'h00050CD2 , 32'h00089D33 , 32'hFFFF50E3 , 32'hFFF9CE0F , 32'h000FEBB5 , 32'hFFF7D33A , 32'h00088B2B , 32'hFFF57AB9 , 32'hFFFDD2F0 , 32'hFFF83B3C , 32'h000398BE , 32'h0013E4EE , 32'h0008CA3B , 32'hFFF611FD , 32'hFFF999EB , 32'hFFF87F58 , 32'hFFF67E97 , 32'hFFFFD268 , 32'h00061D4D , 32'h0003D157} , 
{32'hFFFB3EE1 , 32'hFFF7AB61 , 32'hFFFD70D0 , 32'h000069C5 , 32'h0005E06A , 32'h00018712 , 32'hFFFE3C0B , 32'hFFF64085 , 32'hFFF7FCCB , 32'h0001EC7D , 32'h000316ED , 32'hFFFD332B , 32'h000056E2 , 32'h0006FD1D , 32'h00058E5A , 32'h0000057F , 32'hFFFEA971 , 32'h00020965 , 32'h0001A272 , 32'hFFFF90B5 , 32'hFFFBE88C , 32'h000935FB , 32'h0000FBED , 32'h0006CF5F , 32'hFFFCAAEA , 32'hFFFB345D , 32'h00031A33 , 32'hFFF8E2EE , 32'hFFFDE8AE , 32'h000201C2 , 32'hFFF9E0D6 , 32'hFFFE7ADC , 32'hFFFED6D9 , 32'hFFF8D807 , 32'hFFFDD6E1 , 32'hFFFC279A , 32'h00017E42} , 
{32'h0001208A , 32'h0001D2CD , 32'hFFFEBD41 , 32'h0001DBC0 , 32'h00012D50 , 32'h000540E1 , 32'hFFFF48D8 , 32'h00007089 , 32'h00050D37 , 32'h000598D0 , 32'hFFFE5B72 , 32'h00005F44 , 32'hFFFAC6D0 , 32'h0004A5BB , 32'hFFFFAA5A , 32'h000571C2 , 32'hFFFD1CB0 , 32'h000321F0 , 32'hFFFC8538 , 32'hFFFE8ED0 , 32'hFFFADE74 , 32'hFFFF69C2 , 32'hFFFE1F0E , 32'h00025151 , 32'hFFFEB75D , 32'h0004380E , 32'h0005EC5A , 32'hFFFB4017 , 32'hFFFE85F8 , 32'hFFFF6B17 , 32'h00036DA8 , 32'h00017419 , 32'h0002F945 , 32'hFFFC2FAC , 32'hFFFF8252 , 32'h00003C89 , 32'h0000156E} , 
{32'h0000193A , 32'hFFF8B74B , 32'hFFF92762 , 32'h00020F50 , 32'h000137F9 , 32'h00042692 , 32'h00014EDD , 32'h00004EAD , 32'hFFFCC6FA , 32'h00033D1D , 32'hFFFE7ED5 , 32'hFFFD8F0A , 32'hFFFD63A7 , 32'hFFFC1D3D , 32'hFFFC396B , 32'h00043F75 , 32'h0004760B , 32'hFFF79401 , 32'h0006858E , 32'h000040E8 , 32'hFFFBE32B , 32'hFFFE6282 , 32'hFFFC08EB , 32'h00010096 , 32'hFFFD5727 , 32'hFFFC8DE1 , 32'hFFFFB882 , 32'h0001036B , 32'h000381C7 , 32'hFFFBE01E , 32'hFFFC7025 , 32'hFFFC4B77 , 32'hFFFF31DE , 32'h00010FFD , 32'hFFFEB8E0 , 32'h00014160 , 32'hFFFB5FE7} , 
{32'hFFFEA93A , 32'h000201AD , 32'hFFF95F49 , 32'hFFFFCAF1 , 32'h0000B47F , 32'h0004C51A , 32'h00030690 , 32'h0003BA38 , 32'h000CAA65 , 32'hFFFEBFA2 , 32'hFFFE87D4 , 32'h00012D69 , 32'h0005D21B , 32'h00011BCA , 32'h00047EF0 , 32'h0006694E , 32'hFFFB4DC7 , 32'h0000A603 , 32'hFFFFFFB8 , 32'h00004832 , 32'hFFFE8817 , 32'hFFFEB4E3 , 32'h0001F373 , 32'hFFFCDE40 , 32'h0000880A , 32'h0000B7FF , 32'hFFFE118B , 32'h000333B5 , 32'hFFFEED6E , 32'h0004CFBB , 32'h0002430D , 32'h0003D398 , 32'hFFFAED2E , 32'h000461B2 , 32'h0002C2F8 , 32'hFFFFED63 , 32'hFFFEF639} , 
{32'h0002C364 , 32'hFFFD8D4E , 32'hFFFE9663 , 32'h000929F9 , 32'h00071344 , 32'h0000A3C1 , 32'h000107D4 , 32'hFFFB1DFE , 32'h0000E223 , 32'hFFFF4705 , 32'h0007E752 , 32'hFFFFA933 , 32'hFFFE78D2 , 32'hFFFAEE39 , 32'h00038E23 , 32'hFFFFE007 , 32'hFFFB7E83 , 32'hFFFBF04A , 32'h00038511 , 32'h0001BB50 , 32'h00063F85 , 32'h00047BA3 , 32'h0003FE25 , 32'h00078953 , 32'hFFFF4660 , 32'h0000D497 , 32'hFFFC6A23 , 32'h00020123 , 32'h00040070 , 32'h0000B4F5 , 32'h0003AD91 , 32'hFFFA0A19 , 32'hFFFCBB8F , 32'hFFFB5BFF , 32'hFFFA4E29 , 32'h0005D3CA , 32'hFFFF90B4} , 
{32'h0000FB27 , 32'h00010509 , 32'h0001F90A , 32'h00036E94 , 32'h0000543E , 32'h0006165C , 32'h0002FE83 , 32'h00024424 , 32'hFFFA3B2F , 32'h000160B8 , 32'h0003BDF4 , 32'hFFFFA914 , 32'h0001EE86 , 32'hFFFCE6F6 , 32'hFFFFBCE3 , 32'hFFFF9CB6 , 32'hFFFC1F2A , 32'hFFFCF907 , 32'h000225AB , 32'h00039901 , 32'hFFFDCD19 , 32'hFFFD97F2 , 32'h00079511 , 32'hFFFDD58A , 32'h000229D2 , 32'hFFFD71BE , 32'hFFF7CDC6 , 32'h0003EABF , 32'hFFFFE632 , 32'hFFFB58C8 , 32'h0001F895 , 32'hFFFCD934 , 32'hFFF969D9 , 32'hFFFDCA1F , 32'hFFF89FC8 , 32'hFFFD38E7 , 32'hFFFE200B} , 
{32'h01D93AC4 , 32'h000FB087 , 32'h0441EB90 , 32'hFFC716CA , 32'h05D3E4C0 , 32'h0136D6AC , 32'h026FC870 , 32'h05FA0D40 , 32'h0389993C , 32'hFD66C4C4 , 32'h0502FD20 , 32'h01C130A8 , 32'h04B73E18 , 32'hFD8EACEC , 32'hFCCC51E8 , 32'hFA14A590 , 32'hFB9067B0 , 32'hFA35F020 , 32'h037CF0AC , 32'hFFE33C1C , 32'hFEE497AC , 32'hFC30E54C , 32'h03DBA1DC , 32'hFDDFEBA0 , 32'hFAC88788 , 32'hF8050F40 , 32'hFF98DCEF , 32'hFC7B7340 , 32'h001C2919 , 32'h02E8A7E8 , 32'h05FC2CE8 , 32'h0472E4B0 , 32'h00FE8D27 , 32'h081CE9B0 , 32'hFDF123E0 , 32'h018AECCC , 32'hF942F800} , 
{32'hEBDD04A0 , 32'hF293B900 , 32'h21340FC0 , 32'hFCBF0764 , 32'hF5B56880 , 32'h0310B9EC , 32'h10EBF8E0 , 32'h0A253CA0 , 32'h09B97E70 , 32'hFF2B182C , 32'h1C518500 , 32'hFF5C3B0D , 32'hF11B3B30 , 32'hF5880150 , 32'hF0281850 , 32'hF8BDF5F8 , 32'hE859DD60 , 32'hE826C420 , 32'hF97021D0 , 32'h020C5864 , 32'hEE791B80 , 32'h0A3C7200 , 32'h07B45BE0 , 32'h0BF64E40 , 32'h0B452790 , 32'h08DDD6E0 , 32'hEB4B1F80 , 32'hF4AB9F70 , 32'hEEBE1620 , 32'h10EE7180 , 32'h0493CA58 , 32'hF7FCC0F0 , 32'h0862D740 , 32'hE5F4FE60 , 32'hF621A650 , 32'hFBD466B8 , 32'h037CFFE0} , 
{32'hF0357AC0 , 32'hEC588540 , 32'h1C328980 , 32'hFC4C0728 , 32'hFDB90974 , 32'h10247B20 , 32'h0EF2A8A0 , 32'h0D7511C0 , 32'hF7930E90 , 32'hFCED2814 , 32'h0BD11600 , 32'h028B48C4 , 32'hFB348A70 , 32'h07937B10 , 32'hEDE6EAA0 , 32'h06A597A0 , 32'hF56A8BD0 , 32'hF1D508C0 , 32'hF86805F0 , 32'h06230BF0 , 32'h0109CB58 , 32'h092AB550 , 32'hFDE5D638 , 32'hFD0B68A4 , 32'h0762CC88 , 32'h09E0B250 , 32'h079C00C8 , 32'hFB31C800 , 32'h067174F0 , 32'h080D0720 , 32'h03BD985C , 32'h0A517250 , 32'h09CC0B40 , 32'hFE3B1FF0 , 32'hFE937D60 , 32'hFF851DF8 , 32'h04D621B8} , 
{32'hEFFC7D80 , 32'hF0D2BD10 , 32'h3755A500 , 32'hF85D1AE0 , 32'h00B3C474 , 32'h22709700 , 32'h1E9098E0 , 32'h13A855A0 , 32'hF4A44D00 , 32'hFCD43988 , 32'h14FFC940 , 32'h0B427480 , 32'hEEA4F680 , 32'h02C16004 , 32'hED6B0B20 , 32'hF1C068A0 , 32'hEDA9A5E0 , 32'hE6DE01A0 , 32'hF489B210 , 32'hF755E930 , 32'h01860FFC , 32'h09528B90 , 32'h034784C8 , 32'hFA19B8B0 , 32'h08961F70 , 32'h0DC38E50 , 32'h1325C5A0 , 32'hF67AE440 , 32'hF2B35700 , 32'h052DA648 , 32'hF977B030 , 32'h0AB95830 , 32'h145F1860 , 32'hE4DD8080 , 32'hF4DD4FC0 , 32'hFE8DFF44 , 32'h10BCDF80} , 
{32'hE1F624C0 , 32'hDA5D9380 , 32'h519DF200 , 32'h0BA231C0 , 32'hF5ED3090 , 32'h25AFC600 , 32'h2A7B4480 , 32'h1C4BDB00 , 32'hEE3EFFC0 , 32'h0A2039C0 , 32'h0CBEBED0 , 32'h04F51550 , 32'hF1935B00 , 32'h0A0F3050 , 32'hED3CF1E0 , 32'hE6AE67E0 , 32'hF2D502C0 , 32'hEAE2C200 , 32'hF4A1A680 , 32'h07188478 , 32'h0825B2C0 , 32'hFF3FEF03 , 32'hFBF62C10 , 32'hF8909438 , 32'hFDCCE260 , 32'h01824C88 , 32'h16DBFAC0 , 32'hEDB9EE40 , 32'h10383120 , 32'h06B52118 , 32'hFF86C390 , 32'h0DA27D30 , 32'h0FE266E0 , 32'hFA450A60 , 32'h0E0C2E80 , 32'hF1ED3920 , 32'hF7B386A0} , 
{32'hCE4EFD00 , 32'hD73C61C0 , 32'h5B3C1A80 , 32'hFCB22BF0 , 32'hEA78E520 , 32'h24F37CC0 , 32'h1B9E9740 , 32'h19939580 , 32'hF152BBD0 , 32'h0AABA330 , 32'h04CCFCB8 , 32'hF6764120 , 32'hED692B20 , 32'h119FF760 , 32'hECA8A300 , 32'hFFDF651D , 32'hF1288C30 , 32'h01DEC9A4 , 32'hEFCC4600 , 32'h0C723560 , 32'h0AAFEE00 , 32'h0966D730 , 32'h06027890 , 32'hFC7BFEA0 , 32'h069CA9E0 , 32'h0C725060 , 32'h1903E180 , 32'h04E4C410 , 32'h0AC177A0 , 32'h10343640 , 32'hF38F6D50 , 32'h0FFD1550 , 32'h0E8671A0 , 32'hF3327600 , 32'hF0C074A0 , 32'h005C413E , 32'h097A48D0} , 
{32'hE2429840 , 32'hE554DFE0 , 32'h3A885E80 , 32'hFCF5C850 , 32'hE03CE420 , 32'h2280DB00 , 32'hFB821180 , 32'h10DE59E0 , 32'hEB3C55C0 , 32'h03020134 , 32'h162C2E40 , 32'hEE8B98C0 , 32'hE5B61F20 , 32'h0C9CC190 , 32'hFD7E0C80 , 32'hEBBCAB60 , 32'hE89BDB00 , 32'hFE97AC98 , 32'hE9C7A080 , 32'h079E7700 , 32'hFFE8A3DA , 32'hEC857120 , 32'h0F97D750 , 32'hFB628190 , 32'h066A0648 , 32'h0BAF1540 , 32'h14BC1440 , 32'hE9C66D20 , 32'h09A8CE40 , 32'hFC8276AC , 32'hFD7A1CCC , 32'h1E4D8280 , 32'h02354554 , 32'hFDF64EA4 , 32'hFE03A610 , 32'hFC895808 , 32'h08E05230} , 
{32'hF8D54A80 , 32'hF94F20D0 , 32'h00103989 , 32'h0BAFC710 , 32'hDB451B80 , 32'h027CD5EC , 32'h0AF576A0 , 32'h04389718 , 32'h0970DAE0 , 32'hF5C181D0 , 32'h1CDD2340 , 32'hED12B5E0 , 32'hFF95D248 , 32'hF732ECF0 , 32'h0582A130 , 32'hF8172068 , 32'h0C2E21C0 , 32'h128BDBA0 , 32'h06800518 , 32'hFD0D9634 , 32'h026DF06C , 32'h01B843DC , 32'h0904C010 , 32'h083D5910 , 32'hF5E4A140 , 32'hF4230740 , 32'h0D43B7E0 , 32'hF774B440 , 32'hF4853D40 , 32'hEFF68180 , 32'h12B8B360 , 32'hF3DA8070 , 32'h0847E330 , 32'h03792ACC , 32'h120E4740 , 32'hFDB38194 , 32'hFD0EACF8} , 
{32'hF765CF50 , 32'hC7429640 , 32'hE3390680 , 32'h0B5DEEB0 , 32'hBC885680 , 32'hF23C6E40 , 32'h03E8B3F0 , 32'hF0A03EA0 , 32'hFE4AB3C8 , 32'hFBB66C30 , 32'h2CDE5F80 , 32'hDE4DA100 , 32'h08713E90 , 32'hF3CFBBD0 , 32'hF1CED2F0 , 32'hFB251AD8 , 32'hFF4F78BE , 32'h0A2BD300 , 32'h0C6EFBB0 , 32'hF55ECD40 , 32'hF272F920 , 32'hFDA78AB4 , 32'h05576740 , 32'hF575A360 , 32'hF96D5408 , 32'hF85329E0 , 32'hF9FBAEA8 , 32'h002009ED , 32'hE898C300 , 32'h0E503340 , 32'h0A945D90 , 32'h203A98C0 , 32'hFEAC6BEC , 32'h15276660 , 32'h0C229D60 , 32'h02B393FC , 32'h192C5200} , 
{32'hEB2DF400 , 32'hF24F84E0 , 32'hDE8D3B00 , 32'h0E45C950 , 32'h9F6E2200 , 32'hEF982620 , 32'hF769F6C0 , 32'hEADB5780 , 32'h08684520 , 32'h063450E0 , 32'h0C5B6B30 , 32'h1FE4F020 , 32'hEDD9EB40 , 32'h0561F8E8 , 32'h04B29550 , 32'hF845B378 , 32'h0579E9C8 , 32'hF4199330 , 32'h01D04080 , 32'h144A4400 , 32'h0E3F2E30 , 32'hCED16DC0 , 32'h011550EC , 32'h13BAEDA0 , 32'h0E830B30 , 32'h0B12B120 , 32'h082FC3F0 , 32'h04D83510 , 32'hF4EDFCD0 , 32'h0D665F20 , 32'h1591A740 , 32'h1E781D60 , 32'h1033C920 , 32'h216512C0 , 32'hF3991220 , 32'hE1FDC400 , 32'h175C4100} , 
{32'hF1F85350 , 32'h05A58E70 , 32'hFBECB6A0 , 32'h0E06F280 , 32'hE5106200 , 32'hFFB03E21 , 32'hF2F34700 , 32'h034D52C8 , 32'hFA216DE8 , 32'h1B88DB60 , 32'h03F3BB70 , 32'h16D6AEA0 , 32'hF2299D50 , 32'h17830940 , 32'h12AAFC60 , 32'h0BBDB590 , 32'h191365C0 , 32'hF46326B0 , 32'hFD5503DC , 32'h1CD3CD20 , 32'hED109CC0 , 32'hF0A4CD40 , 32'h0B6A3A70 , 32'h05807F88 , 32'hFB3F0DA8 , 32'h0314BC70 , 32'h023790F0 , 32'h0CDBA470 , 32'h05773BA8 , 32'hEF9B5120 , 32'hF9905380 , 32'h0E885E60 , 32'hF786D410 , 32'h00D731FC , 32'hFD144EF4 , 32'hF3753210 , 32'hEF956FA0} , 
{32'hF6F13340 , 32'hFD0AF328 , 32'h04F371F0 , 32'h0E571B40 , 32'hF960A660 , 32'h04FFD048 , 32'hF6BDA960 , 32'hEE96D940 , 32'hF86A6420 , 32'h03B03560 , 32'hED7E3160 , 32'h0B9488A0 , 32'hF66B1890 , 32'h0DEB3920 , 32'h051897B0 , 32'h06A72EA0 , 32'h03633814 , 32'hF78A9F60 , 32'hFB6EC288 , 32'h0DB7A9A0 , 32'hED251360 , 32'h04502E90 , 32'hFAC0BF70 , 32'hFE3638B8 , 32'hFFBB8FCE , 32'hFC0CFF30 , 32'h00DFAA4D , 32'hF722D570 , 32'hF1078D10 , 32'h00ABBAF9 , 32'hF9CA6DD8 , 32'h0D75ADD0 , 32'hF123C060 , 32'h0DAC54B0 , 32'h053F7530 , 32'hF74B6650 , 32'hFE1BB110} , 
{32'hF24528F0 , 32'hF8ED4060 , 32'h077A5D08 , 32'h10444E00 , 32'hFE090168 , 32'h01D8A87C , 32'hEEFDEC40 , 32'hF3BE4600 , 32'hFF303909 , 32'h0B8430F0 , 32'hEE4A0CA0 , 32'hFF87BEA8 , 32'hFECE8F38 , 32'h05B68A40 , 32'h016086F0 , 32'h18F395A0 , 32'h1A998AC0 , 32'h008F4165 , 32'h061D5D10 , 32'h078C28B0 , 32'h1BDE8E00 , 32'hFFDFC7B3 , 32'hFF677897 , 32'hFA58D0E0 , 32'h1B7B9040 , 32'h0135893C , 32'hEF7FA4A0 , 32'hFD6D9324 , 32'hF52D0890 , 32'h03AA6434 , 32'h0C9653E0 , 32'hFC793BC8 , 32'h0052A0BB , 32'h0F37F9A0 , 32'h17732120 , 32'hFF5EAF43 , 32'hFB3B2B40} , 
{32'hF9922C58 , 32'hED90CC40 , 32'h0581C408 , 32'h1BDD5CE0 , 32'h087377F0 , 32'h1DA9AE00 , 32'hE69621C0 , 32'hEEAFBA00 , 32'hFAE00308 , 32'h03D1B1A4 , 32'h0AA97040 , 32'hF6AB2F00 , 32'h09CFE5E0 , 32'hFAB71910 , 32'h1C1E6A00 , 32'hEA8BB9C0 , 32'h11557080 , 32'hEDC858A0 , 32'h0492BE98 , 32'h05AF6E10 , 32'h02E29E1C , 32'hFFFD29CD , 32'hFCD98854 , 32'hF30A7A50 , 32'h05828818 , 32'hE9EC7260 , 32'hEF89E420 , 32'hEEAD61A0 , 32'h0408CFF0 , 32'hF8E7B438 , 32'hF84224C8 , 32'h037D053C , 32'hEF55E120 , 32'hEDDA4680 , 32'hEEF2D860 , 32'h08DC3330 , 32'h0828C540} , 
{32'hF8D15FC8 , 32'hF5794AF0 , 32'h06D88DD8 , 32'h09980C80 , 32'h1388C000 , 32'h12630EA0 , 32'hE5ADB540 , 32'hF9CC44B0 , 32'h0282AF68 , 32'h00BE5E6A , 32'h1D46D1C0 , 32'h074EDA98 , 32'h24E0CC80 , 32'hF2DEFCD0 , 32'hFEE2388C , 32'hF9AB0B58 , 32'h05944488 , 32'hFEA368F8 , 32'h16D98BE0 , 32'hF8ED2178 , 32'h0EB6E060 , 32'h05DB7B28 , 32'hF6F16E20 , 32'hF61E7BE0 , 32'hFFC75153 , 32'hF3946C70 , 32'h09AC2C20 , 32'hFC1C7A94 , 32'hFB2AD390 , 32'h050E92E8 , 32'hEBB78CE0 , 32'hFADBAA88 , 32'h059815B0 , 32'h062AC4C0 , 32'hFD71AC7C , 32'h03A59B74 , 32'hFD6ADD0C} , 
{32'h02A6B4A0 , 32'hEF299FC0 , 32'hF9524C08 , 32'h0DC71830 , 32'h068525B0 , 32'h184F7E40 , 32'hE9E01BA0 , 32'h10EEEB60 , 32'hFCE84DA8 , 32'hFD370BB0 , 32'h2D438780 , 32'hE2A82620 , 32'h210C8B00 , 32'hFC511C28 , 32'h021A90D8 , 32'h00BFC21B , 32'h18FD8840 , 32'hE427FDC0 , 32'h18B7C240 , 32'hEA4427E0 , 32'hE5935D00 , 32'hF9425150 , 32'hF276A3D0 , 32'h0E806A80 , 32'hEC93C3E0 , 32'h0E7AD0A0 , 32'h0245C470 , 32'h0F39A9E0 , 32'hFD9C3724 , 32'hDE6DDAC0 , 32'hEFD9B720 , 32'hEF764DC0 , 32'h153A4100 , 32'hF9C63B90 , 32'hF3BE9EF0 , 32'h02FF6F60 , 32'h06A034A0} , 
{32'hFAFD5898 , 32'h019652E0 , 32'hFE01D87C , 32'h0FBB0F40 , 32'h0E6ACA00 , 32'h1D719960 , 32'hF8EC4688 , 32'h0FA50DE0 , 32'h0D4D0B50 , 32'hE3AF7580 , 32'hFAFDDD18 , 32'hDF68E700 , 32'h212B8A40 , 32'h05A8CE88 , 32'h0C4F1030 , 32'hF59BD870 , 32'hF123B4A0 , 32'hF087F0B0 , 32'h1C713A40 , 32'hF8BE5AD0 , 32'h0DE7FCC0 , 32'h33DE1F00 , 32'hFEFDBC84 , 32'h0AB4C2C0 , 32'hFBA2F8A0 , 32'h0F041F70 , 32'h02BC5538 , 32'hCC66D000 , 32'hF3C17890 , 32'hFC5D635C , 32'h03DA72B8 , 32'h15158560 , 32'hF229F640 , 32'h04B28A90 , 32'h03002734 , 32'hFD165820 , 32'hF07CAA00} , 
{32'h01693654 , 32'hFFFD334D , 32'h00FE75A3 , 32'h0616E820 , 32'h010665BC , 32'h06EB9CD0 , 32'hFCF3B884 , 32'h05819EC8 , 32'h06298E40 , 32'hF9A5C240 , 32'hFD807A34 , 32'hF43A4800 , 32'h0D05EC60 , 32'hFD8AF288 , 32'h02A1BAC0 , 32'hFE4336A8 , 32'hFEF1E560 , 32'hF8A84AA0 , 32'h00DA70AB , 32'hFE0FE4E4 , 32'h0E2526A0 , 32'h039D25E8 , 32'h04778170 , 32'hFF101530 , 32'hFBD5B800 , 32'h01A008F4 , 32'h02CA3790 , 32'hE4150C20 , 32'hF395F9B0 , 32'hFCCDDB34 , 32'hF78C1BA0 , 32'h10FC32C0 , 32'hFE69FA94 , 32'h046A2C38 , 32'h016CDA00 , 32'hF7A7BDD0 , 32'hF71EEF40} , 
{32'h03C9FBD4 , 32'hFC536468 , 32'hFD478E3C , 32'hFEC0D5FC , 32'h06C30B00 , 32'h0C0CFC30 , 32'h046D5D08 , 32'hFEC4604C , 32'h028F22D4 , 32'h03EE93D8 , 32'hFC6112E8 , 32'h04E9D120 , 32'h12CEF2A0 , 32'hE33EF720 , 32'hF69CC790 , 32'hF5BAF250 , 32'h0E7FC5E0 , 32'hFA279E08 , 32'hF0FE3F70 , 32'h0EA26380 , 32'hFB36B440 , 32'h04039CA8 , 32'h0EF30E70 , 32'hFB7B33C8 , 32'h07B686A8 , 32'h0034D4E2 , 32'h0B43BC80 , 32'h04A706A8 , 32'hFD743A64 , 32'h02AD277C , 32'h02243914 , 32'h0CB982A0 , 32'h0465B738 , 32'h05A7C200 , 32'h0107191C , 32'h0247A704 , 32'hFE279470} , 
{32'hF5F61460 , 32'h03B7AFE4 , 32'h030F0774 , 32'h0549E740 , 32'h0B9B98F0 , 32'hF8D45CC0 , 32'h0A771FC0 , 32'hFD34FC64 , 32'h114E6DA0 , 32'hF7E760B0 , 32'hF5A1D720 , 32'h0C848050 , 32'hFF28FBC4 , 32'hFCFBDD4C , 32'h0A917650 , 32'hFD0A20A8 , 32'hFF1C4288 , 32'h0518F560 , 32'h062F9E28 , 32'hF6736290 , 32'hF3D33D30 , 32'h03BA5184 , 32'hFC7C6F00 , 32'hF3401340 , 32'hF9C43030 , 32'h03695CD0 , 32'h0ED51630 , 32'h0292BDEC , 32'h0133934C , 32'h0496F020 , 32'hFB236278 , 32'h0A923920 , 32'h12D0AD20 , 32'h0762BA18 , 32'h06A1CEA8 , 32'h0C074F00 , 32'h03C9DAE8} , 
{32'hF99A1120 , 32'hF22B0E00 , 32'h002AD73F , 32'h0F52AE60 , 32'h07849FF8 , 32'hFE48153C , 32'hFB2C8940 , 32'hF4BEF1B0 , 32'h03E84BE4 , 32'hFA41B930 , 32'h01A48510 , 32'h0E7AA990 , 32'hF00E9440 , 32'hF94AFCF8 , 32'h08AEE2B0 , 32'hF6339740 , 32'hFB7DA2B0 , 32'h189DD2A0 , 32'h1072BB80 , 32'h00906978 , 32'hEB553360 , 32'h0E6DF0E0 , 32'h0B3373C0 , 32'hE8AEC440 , 32'hF5C50C70 , 32'h0C838480 , 32'hFFB0FB38 , 32'h00A97287 , 32'h0F490730 , 32'h08464EC0 , 32'h03509FE0 , 32'h04A6EFF8 , 32'h123F2160 , 32'h087C4430 , 32'hFFA43844 , 32'h0CA173B0 , 32'h00B95924} , 
{32'hFFEE7435 , 32'h000C23F0 , 32'h0002D29D , 32'h000326BC , 32'h0000CB8C , 32'hFFF54EA1 , 32'h000735BF , 32'hFFEFE113 , 32'h000CE6F4 , 32'h000376E9 , 32'hFFF86C83 , 32'hFFFC39FE , 32'h0002DF4A , 32'h0004213E , 32'h000353BD , 32'h0019622F , 32'h0008EA7C , 32'hFFFFBD0D , 32'h000B0736 , 32'hFFF74EFF , 32'hFFF8BC14 , 32'h001231C3 , 32'hFFEFE8E0 , 32'h000CCB0E , 32'hFFFBBDF0 , 32'h0004E1EB , 32'h0000E558 , 32'hFFFDCE0B , 32'h000BD144 , 32'h00056514 , 32'hFFF6761D , 32'hFFFFF389 , 32'h0003506E , 32'hFFF6A637 , 32'hFFF9C4AA , 32'h00084962 , 32'h0000CEC4} , 
{32'h00051478 , 32'h00021A84 , 32'hFFFEE5E5 , 32'h000242E5 , 32'h00044377 , 32'h00000638 , 32'hFFF79F7D , 32'hFFFECB91 , 32'h0005067F , 32'hFFFFFF00 , 32'h0000985D , 32'h0003DDF6 , 32'hFFFA86BA , 32'hFFFF72D1 , 32'hFFFEAB39 , 32'h000366E3 , 32'h0001C1B2 , 32'hFFFBBDBD , 32'hFFF75609 , 32'hFFFDB9EF , 32'h0002A712 , 32'hFFFDA682 , 32'h0000E4D9 , 32'hFFFC8547 , 32'h000021BE , 32'hFFFDB077 , 32'hFFFB7F8C , 32'hFFFC2BB1 , 32'hFFFD373E , 32'h000584AC , 32'hFFFE1E8A , 32'hFFFFF35D , 32'hFFFF9EBB , 32'hFFFC58B4 , 32'hFFFFD625 , 32'h00059C02 , 32'hFFFEE36A} , 
{32'h0005EE46 , 32'h00008024 , 32'h0004FB5B , 32'h0005C38B , 32'hFFFEDB5F , 32'hFFFD02F3 , 32'h0001D7B7 , 32'h0002C334 , 32'h0007DC80 , 32'h0001ADFD , 32'hFFFFDE63 , 32'h00055C6B , 32'hFFFFE7B9 , 32'hFFFA7594 , 32'hFFFF8721 , 32'h000636EF , 32'h0005753C , 32'h0000B6C3 , 32'hFFFB1FA9 , 32'h00014B78 , 32'hFFFFDC36 , 32'hFFFE43DC , 32'h0000A419 , 32'hFFFA5807 , 32'hFFFD36B4 , 32'h00018276 , 32'hFFFEC15C , 32'h00023B7B , 32'h0004BDA1 , 32'h000101B5 , 32'h0000E81C , 32'hFFFD8BF5 , 32'hFFFE834A , 32'h000196BE , 32'hFFFD14F3 , 32'hFFFD2854 , 32'hFFFDBFA7} , 
{32'hFFFF93C7 , 32'hFFFE3275 , 32'h000557C7 , 32'h0001DE7A , 32'h0000BF08 , 32'h00019DE8 , 32'h00017D16 , 32'hFFFCC086 , 32'hFFFD8976 , 32'h00072D29 , 32'hFFFA9661 , 32'h0004A5A2 , 32'h00037BE6 , 32'h000448BF , 32'hFFFEA562 , 32'hFFFF7303 , 32'hFFFB8F01 , 32'hFFFF2EEC , 32'h00013DA6 , 32'hFFFE18C1 , 32'hFFFA9D57 , 32'h0001A8E3 , 32'h00020A1C , 32'hFFFE8F17 , 32'h000134C4 , 32'h0001E731 , 32'hFFFB2333 , 32'h00031ED3 , 32'hFFF6FFAE , 32'hFFFF0314 , 32'hFFFD4B80 , 32'h00028EAB , 32'hFFFD99A0 , 32'hFFFF57A5 , 32'h000596D2 , 32'h0004CB94 , 32'hFFFF5C50} , 
{32'hFFFC8833 , 32'hFFFC2DAD , 32'h00044110 , 32'hFFF9293E , 32'hFFFD1CBD , 32'h0003F564 , 32'hFFF6F975 , 32'h00011962 , 32'h000115B2 , 32'hFFFE61A7 , 32'hFFFF6573 , 32'h00047FC2 , 32'hFFFB5592 , 32'hFFFF3A0E , 32'h0005535D , 32'hFFFDB313 , 32'h00007EE4 , 32'hFFFEF18A , 32'hFFFBCA4A , 32'hFFFD4E5C , 32'h00003FA0 , 32'hFFFCFBF2 , 32'hFFF69C13 , 32'h00013E39 , 32'hFFFBA670 , 32'hFFFE92B6 , 32'hFFFA6929 , 32'hFFFE45B1 , 32'hFFFDD73B , 32'h00031294 , 32'h00020F72 , 32'hFFFDD50E , 32'hFFFF3DC9 , 32'hFFFB0902 , 32'hFFFE3662 , 32'hFFFB88DB , 32'hFFFF16EF} , 
{32'h0009AA05 , 32'hFFFD40BE , 32'hFFFC3E5B , 32'h0008853E , 32'hFFFAF040 , 32'h000B6C76 , 32'h00020DA3 , 32'hFFF6FEEF , 32'hFFFAE5ED , 32'hFFFE57F0 , 32'h0004E3A8 , 32'hFFFD4999 , 32'hFFFAE294 , 32'h00024803 , 32'hFFF54BF3 , 32'h0000D2A8 , 32'hFFFEDB12 , 32'hFFFC77D8 , 32'hFFFBF9D2 , 32'h0003C4AE , 32'h00001B14 , 32'h000591BA , 32'h00018814 , 32'hFFFA3E9E , 32'hFFFBB064 , 32'h00023D5C , 32'hFFF51290 , 32'h00026254 , 32'hFFFE9179 , 32'h000036D4 , 32'h000212C2 , 32'h00038FD3 , 32'hFFF1DE29 , 32'h000374EF , 32'hFFFECC00 , 32'hFFFB7299 , 32'h0000ABCA} , 
{32'h00501A58 , 32'hFFCF7257 , 32'hFFD712AF , 32'hFFF1DDAB , 32'hFFCD94C2 , 32'h0060BC1C , 32'hFFD1A5A3 , 32'h001C5B40 , 32'hFF965A8D , 32'h000F768C , 32'h00641C84 , 32'hFFDE2534 , 32'hFFBF3493 , 32'hFFF27292 , 32'hFFCDBE38 , 32'hFFA751AB , 32'hFFEF6145 , 32'hFFDEA4F0 , 32'hFFFDD088 , 32'h0041682E , 32'h001A75EA , 32'h0001DEAC , 32'h005EC710 , 32'h0001BF81 , 32'h0001CE91 , 32'h000349DF , 32'hFF9E7563 , 32'h00053435 , 32'h001DB8D4 , 32'hFFE60B23 , 32'h0036ECC1 , 32'hFFEB609C , 32'hFFA1ABE2 , 32'h0013B0B5 , 32'hFFC6F3AE , 32'h00047D5E , 32'h001B0E27} , 
{32'hED210460 , 32'hEE98D0C0 , 32'h11CBCEE0 , 32'h010D9678 , 32'h0731F630 , 32'hFE658E14 , 32'h032C021C , 32'h05E5A6E8 , 32'hF95651D8 , 32'hFC5DEF44 , 32'h08BEE930 , 32'hF0E56870 , 32'hF64F6A20 , 32'h0A3FCCC0 , 32'hFBFEAC30 , 32'h0C7DBD00 , 32'hF9281CD0 , 32'hFD21E068 , 32'hF1674030 , 32'h101C78A0 , 32'h0ED7B830 , 32'h0447CD38 , 32'h017BB6F4 , 32'h00339359 , 32'hFE28585C , 32'h0658B4E0 , 32'h0D3DFFF0 , 32'h04905728 , 32'h112DDF00 , 32'h03AE3758 , 32'hF8877C38 , 32'h08693B80 , 32'h030D241C , 32'h0859B4A0 , 32'hFF15EA2E , 32'h03B61CFC , 32'h07333930} , 
{32'hE36D0080 , 32'hD8A40500 , 32'h11EEF920 , 32'hFB463508 , 32'h2B4D2CC0 , 32'h02E598D4 , 32'h00C4658E , 32'h0A206BE0 , 32'hF2DC3920 , 32'h06186940 , 32'hF552ABE0 , 32'hE79ECE80 , 32'hFCAB3AF4 , 32'h150B07C0 , 32'hF647C6C0 , 32'h0F1A1910 , 32'hFB28EE60 , 32'hECC65000 , 32'hF1B1BDF0 , 32'h066B41D0 , 32'h18DF4820 , 32'h08E18480 , 32'h0328D710 , 32'hFF95A5B4 , 32'hF41D4AD0 , 32'h02AFCA40 , 32'hFDBDA774 , 32'h0ABA7880 , 32'h0F2F7F80 , 32'h06226A78 , 32'hFD4FCA08 , 32'h1150C1E0 , 32'hFD7B3F04 , 32'h135E14A0 , 32'hFDEBF110 , 32'h04255318 , 32'h0E4197C0} , 
{32'hCDDFEF80 , 32'hC5E8A500 , 32'h0E774A20 , 32'hE12849A0 , 32'h4B1C5D80 , 32'h1AA3A420 , 32'h0EDB9FD0 , 32'h17FB8000 , 32'hF9A74C20 , 32'h084421B0 , 32'hEC4B3EA0 , 32'hF4EA4400 , 32'hF5F189E0 , 32'h16DE4F00 , 32'hFFF6EB3C , 32'h23277F40 , 32'h117459A0 , 32'hFA580EC0 , 32'hF57C2570 , 32'h013A2A9C , 32'h1FEBE260 , 32'h0CD9DDD0 , 32'h153EC0C0 , 32'h092DAB20 , 32'hEF09C6A0 , 32'hFF5E5A93 , 32'hEAB2E540 , 32'h0BBA3A50 , 32'h0102CF00 , 32'hE935F460 , 32'h13C386E0 , 32'h097E8A20 , 32'hF740FC00 , 32'h1DBD9BA0 , 32'hFF35AE19 , 32'h0B446DF0 , 32'h04DF3BC8} , 
{32'hDCFC44C0 , 32'hCCF72CC0 , 32'h1438D900 , 32'hF8337920 , 32'h43E7D700 , 32'h16323300 , 32'h250F14C0 , 32'h07766658 , 32'hE4633E60 , 32'hF7F2EC00 , 32'hF55F2C90 , 32'h05A7D5A0 , 32'hDF7C3580 , 32'h18169580 , 32'hFCC92788 , 32'hFA48FCA8 , 32'hFCB39B80 , 32'hF0F480E0 , 32'h0D7B56E0 , 32'h0FDCD460 , 32'h0E35F120 , 32'h006AEEF1 , 32'h08547840 , 32'h072DCD10 , 32'hF86D5240 , 32'h0586C110 , 32'h0E59DE80 , 32'h0E20B9B0 , 32'h193D43A0 , 32'h0C678CF0 , 32'hFEFD5AC4 , 32'h03B5BD40 , 32'h0120F224 , 32'h035D00BC , 32'h0ABDC820 , 32'hFD7086C4 , 32'h050DF2F8} , 
{32'hE2090DE0 , 32'hD1BC18C0 , 32'h17A62620 , 32'hF7F1F6A0 , 32'h2CEB9080 , 32'h1B5C5040 , 32'h1EF89E00 , 32'h15638720 , 32'hEA4BA4C0 , 32'h0394D82C , 32'hF65313F0 , 32'h035204C8 , 32'hF06BE9B0 , 32'h1FD07880 , 32'h033E18B0 , 32'h0CC8A310 , 32'hFFC32CDC , 32'hDFAC0A40 , 32'hF771A160 , 32'h16E43FE0 , 32'h06586688 , 32'hFB7790C8 , 32'hF9A3BFA0 , 32'hFA0685B0 , 32'hEDA901E0 , 32'h0BF834B0 , 32'h16EFB7C0 , 32'hFEE0F810 , 32'h0919ACC0 , 32'h02F6A9D4 , 32'h0D6DD9D0 , 32'h007A1A71 , 32'hFED5061C , 32'h0777C4D8 , 32'hFF7D543D , 32'hFA986158 , 32'hFA5134B0} , 
{32'hF5DD9DB0 , 32'hE5735360 , 32'h0DD83080 , 32'hF8439B40 , 32'h052B9000 , 32'h21A9FB40 , 32'h11602B80 , 32'h0F007320 , 32'hE3C659E0 , 32'h0C1CAEC0 , 32'hEBC23320 , 32'hF975BD08 , 32'h05A63AF0 , 32'h10149740 , 32'h15CF6D60 , 32'hE6F24620 , 32'h058F7AF0 , 32'hFF53651D , 32'h0459A3A8 , 32'hFA7246E8 , 32'hF7E4A600 , 32'hF00CCEE0 , 32'hF55749C0 , 32'hF8364FD8 , 32'h07FCDE90 , 32'h11BF5560 , 32'h15DAFEC0 , 32'hF836CDC0 , 32'h05BE19B8 , 32'hF67FB8F0 , 32'h00CE4AB3 , 32'hFD97ABE0 , 32'hF895A740 , 32'hF62A3510 , 32'h0F2A6920 , 32'hFB3CF498 , 32'hF74607C0} , 
{32'hEE4186E0 , 32'hD8A3C1C0 , 32'h25B90640 , 32'h03FA0240 , 32'hD5E954C0 , 32'h1D5750A0 , 32'h1618DA60 , 32'h07A8BF68 , 32'hEB42C800 , 32'h0B6A43A0 , 32'h025BE828 , 32'hF38CEFA0 , 32'h0668CC10 , 32'hFEA63308 , 32'hFC03022C , 32'hF7C57490 , 32'h01D35820 , 32'hFE44DFF0 , 32'hFE28250C , 32'hEEED4320 , 32'hF407E260 , 32'hF02440F0 , 32'hF411CD70 , 32'hFB8F3EB0 , 32'hE6DBFF00 , 32'h00C2C90E , 32'h108EE840 , 32'hFDF15670 , 32'hE743C820 , 32'h0B7F3CE0 , 32'hF0E1FFD0 , 32'hF1FD7D20 , 32'h1C24AAC0 , 32'h072FA478 , 32'h070FEB00 , 32'h070C6310 , 32'hF5406C50} , 
{32'hF81EA688 , 32'hC0CA6780 , 32'h15744940 , 32'hF88F64B8 , 32'hB4935D00 , 32'h21116940 , 32'h3E099780 , 32'h1474AFA0 , 32'hFC932858 , 32'h1EB1B260 , 32'h1D6007C0 , 32'h00729E5B , 32'h18D1DE00 , 32'hC0495AC0 , 32'hEE6B7F00 , 32'hF65C7F10 , 32'h0C25EF80 , 32'h2ADFD240 , 32'hF3EDD660 , 32'hED73E500 , 32'h10CC2160 , 32'h0D3AD100 , 32'h16795740 , 32'h03D056F0 , 32'h0A913660 , 32'hFA0DC680 , 32'h0F620430 , 32'hE675F3C0 , 32'hEF3A6000 , 32'h073540E0 , 32'h01D906CC , 32'hFC5A5EBC , 32'hFE79CB54 , 32'hF20C6460 , 32'hF3D2C570 , 32'h1A496480 , 32'h02274CF8} , 
{32'hEA2C4CC0 , 32'hEA00D800 , 32'h0B2B55B0 , 32'hF665BD90 , 32'hAE263680 , 32'h0ACDBBC0 , 32'h18C77B40 , 32'hF7354840 , 32'hF393B050 , 32'h14676820 , 32'h063A7008 , 32'h16DEFF60 , 32'h0B43B630 , 32'h0741E2C8 , 32'hED9A5F20 , 32'h07A30710 , 32'h015E18C8 , 32'h033BD8F0 , 32'h1DA9A400 , 32'hD726E300 , 32'hF3E86330 , 32'hF8B2E9B8 , 32'hEA57D8E0 , 32'h04655848 , 32'h128A53C0 , 32'h033FFB5C , 32'hF6941170 , 32'hE1A73920 , 32'h11C269A0 , 32'h06EAB608 , 32'hFA81E058 , 32'hF363B760 , 32'hFA45BB70 , 32'hFAE73968 , 32'h0A1B6780 , 32'hF7CCCE50 , 32'hF4F347C0} , 
{32'hFAE94260 , 32'h03E8D814 , 32'hE915A0A0 , 32'hF7395720 , 32'hB3912400 , 32'h13AC8400 , 32'h16168E40 , 32'hF6037F40 , 32'hFC3FC7A0 , 32'h0AAADA60 , 32'hFF83CF0E , 32'h35555000 , 32'h081A4BB0 , 32'h05D9BE58 , 32'h126C5FE0 , 32'h0028B77C , 32'h1B2E4F60 , 32'hEBB06660 , 32'h20E97B40 , 32'h02F7A70C , 32'hFDE55E34 , 32'h09EFF8A0 , 32'h0217D880 , 32'h02920848 , 32'h089E3ED0 , 32'h08ECBBD0 , 32'h0BD634E0 , 32'h05A5E6D0 , 32'h17E2AAC0 , 32'hFA5E6120 , 32'hFD853248 , 32'h214C0C00 , 32'hFED74134 , 32'hE8077A80 , 32'h01565F20 , 32'hFC7E9D40 , 32'hF42B3C80} , 
{32'hF6A03270 , 32'h0C3D7D60 , 32'h029DF5BC , 32'h0E1D7790 , 32'hF9E3DBE8 , 32'h01CAB59C , 32'hF6ABB890 , 32'h00DF637A , 32'hFE8917F0 , 32'h031571AC , 32'h019D8324 , 32'h0CA8E530 , 32'hF4CC7DD0 , 32'h1DDBB8E0 , 32'h010BC43C , 32'hFBC4FE68 , 32'h01D57404 , 32'hF71AF8E0 , 32'h101F66A0 , 32'h04D77590 , 32'h010EBFAC , 32'h0C2EEAF0 , 32'hF7709CB0 , 32'hFC7171F8 , 32'hF15984E0 , 32'h0209D4A8 , 32'h006977FB , 32'hF88402A8 , 32'h049FB148 , 32'hF3C80610 , 32'h004C7335 , 32'h0313E75C , 32'hF6887440 , 32'hFE8A9FE0 , 32'h03B35108 , 32'hFBD1C010 , 32'h02A0B2F4} , 
{32'hEDE59460 , 32'hF9AF7380 , 32'h03E40FA0 , 32'h1BAA2960 , 32'hFE65E43C , 32'h08AF4410 , 32'hF9C350B8 , 32'hEE4985E0 , 32'hFC058CD0 , 32'h01193DB0 , 32'hF9AD89F8 , 32'h18E48860 , 32'hF20E76A0 , 32'h09A43B00 , 32'h0D41DFC0 , 32'h02F85104 , 32'hF6E6B840 , 32'h08DC6970 , 32'h0F9E7AF0 , 32'hFE5888E4 , 32'hE3DCB340 , 32'h07588150 , 32'h06B6A178 , 32'hF29F48B0 , 32'h04433758 , 32'hF662DD70 , 32'hFDE9C1E8 , 32'hFA1AB050 , 32'h01384D60 , 32'hFCC779A0 , 32'hFA98AFA8 , 32'hFC96B2DC , 32'hF815C848 , 32'h0B887750 , 32'h0FC76660 , 32'h0BEBA120 , 32'hFBF3F230} , 
{32'hEEF8AA80 , 32'h041894B8 , 32'h0C4FC170 , 32'h1A433F40 , 32'h01D14368 , 32'hFF704B4C , 32'hE7637660 , 32'hED940F80 , 32'h05580FC8 , 32'h0AB84E30 , 32'hF920DD20 , 32'h04FBA240 , 32'h04667F00 , 32'h1D5FF2A0 , 32'hFAE26E38 , 32'h13354B60 , 32'h237D5B40 , 32'hFD9D6B78 , 32'h0D34ABA0 , 32'h041A8CC8 , 32'h144D9460 , 32'hF12019F0 , 32'h08897890 , 32'hF085B4E0 , 32'h177AA220 , 32'h01C4D3C0 , 32'h0126571C , 32'h0E1EF220 , 32'hFDF590B0 , 32'hF109FCC0 , 32'h11F0A720 , 32'hFA5AC768 , 32'h04E2ED50 , 32'hFAAB6A70 , 32'h0B0EEEA0 , 32'hFF5B9361 , 32'hF378A130} , 
{32'hFB2E2850 , 32'hF4B96B50 , 32'h0822E630 , 32'h1BD61620 , 32'h0DCADC50 , 32'h0BF6EE70 , 32'hEBC25C20 , 32'hF0F4FA20 , 32'h0CD775E0 , 32'h0609A5A8 , 32'h06286F00 , 32'h0CB52CA0 , 32'h0A743F60 , 32'hFA381ED0 , 32'h073E7450 , 32'hFDE383B4 , 32'h0DE6A060 , 32'h00105BE7 , 32'h17995F60 , 32'h0A890080 , 32'hE84A96C0 , 32'hFD7EA664 , 32'h10CF28C0 , 32'hEEAA0620 , 32'hF2143620 , 32'hFC964CD8 , 32'h095D4C80 , 32'h0689FEA8 , 32'h193B8280 , 32'hFB923C48 , 32'hFB780E98 , 32'h06F9AFB8 , 32'h0CFF7400 , 32'h000E4D1D , 32'hED3D0640 , 32'hFB378080 , 32'h0A210070} , 
{32'hF1BFEEB0 , 32'hEB953CA0 , 32'h07329BC8 , 32'h0CEFEF40 , 32'h113C0D40 , 32'h0423DD80 , 32'hDD450D40 , 32'h11CCDEE0 , 32'h00F0F082 , 32'h069369D0 , 32'h1256C4A0 , 32'hE940BB20 , 32'h317C55C0 , 32'h0C69F220 , 32'hF2E67830 , 32'hED2A54E0 , 32'h019A65B4 , 32'hF5395A20 , 32'h145E0960 , 32'hEB0F1100 , 32'hF3B83FE0 , 32'hFCE11814 , 32'hFDC1CF60 , 32'h0242B9A4 , 32'hF3E3C310 , 32'hE7A1DF40 , 32'hF0F5A820 , 32'h0B939CF0 , 32'h0FC4F300 , 32'h0C5519F0 , 32'h0030EAC0 , 32'h01866D58 , 32'hFE091284 , 32'hFA8C6FC8 , 32'hF5C81690 , 32'hF05D9570 , 32'h15503680} , 
{32'hF376F750 , 32'h038BD654 , 32'hFA3D2540 , 32'hE95655A0 , 32'h1345A780 , 32'h0E8C5AA0 , 32'hEBA719C0 , 32'h1248E560 , 32'h0E573B00 , 32'hED7937C0 , 32'h0B0B5C40 , 32'hD2087140 , 32'h08CE9D50 , 32'h05F3DCC8 , 32'h012263A0 , 32'hF88CBD18 , 32'h11FBDAE0 , 32'hF2D8D760 , 32'h083C9A90 , 32'hE3C00820 , 32'hF8B7CB00 , 32'h0AA04760 , 32'h0F1391F0 , 32'hF0CF4E30 , 32'h0695C790 , 32'h089E9C20 , 32'h0629D690 , 32'h05BDC5E0 , 32'h077001D8 , 32'hFCC47FEC , 32'hFC1E17C4 , 32'hFC29BE50 , 32'hF473F970 , 32'hF8BA3168 , 32'h00279A2F , 32'hED03E440 , 32'hFCFC2174} , 
{32'hF5D7A5A0 , 32'h1027DBA0 , 32'hEDF4ECE0 , 32'hFBFC7A78 , 32'h0CE26F50 , 32'h1B88CDE0 , 32'hEFD90900 , 32'h1CBABD60 , 32'h1124E7E0 , 32'hD248CA40 , 32'h03248448 , 32'hD2F29580 , 32'h16381AC0 , 32'h03BF338C , 32'h07600530 , 32'h05999758 , 32'h0A4F5750 , 32'hF69A6380 , 32'h1D440AA0 , 32'hE2FED7E0 , 32'hFDEF53B4 , 32'h1E3FBC20 , 32'h038C1F94 , 32'hEB3491A0 , 32'h1322FB20 , 32'h1F59ADA0 , 32'hFDDB30CC , 32'hF3399060 , 32'hFA001868 , 32'h26FABDC0 , 32'hF7FD2E30 , 32'hEF2ED8C0 , 32'hFAA9F488 , 32'hFC6F360C , 32'hF10DAD50 , 32'hF47D01B0 , 32'hE47B3180} , 
{32'hEDCA2920 , 32'h09E6B320 , 32'hF7CCB4D0 , 32'h0A03D910 , 32'h0932BCA0 , 32'h0FAA3720 , 32'hFC11FD24 , 32'h1BBBBC60 , 32'h070EE910 , 32'h0039E115 , 32'hFB53E120 , 32'hE8A452C0 , 32'hFF44A4CA , 32'h1D8D3C00 , 32'h0340FFE4 , 32'h14295840 , 32'h179F8940 , 32'h045C1038 , 32'h14BDB3E0 , 32'hE75012E0 , 32'h10097C20 , 32'h182922E0 , 32'h131AC420 , 32'hE99CA7A0 , 32'h168E0140 , 32'h18EDACA0 , 32'hF99364D8 , 32'hEDCD2BA0 , 32'hF7ABB7B0 , 32'h0C4E30C0 , 32'h156D5E60 , 32'h16735160 , 32'hF1480050 , 32'h148658C0 , 32'hF6A34200 , 32'h05C73D10 , 32'hEC09B160} , 
{32'h003147C2 , 32'h090A8F90 , 32'hFCEDC92C , 32'hFD265890 , 32'h0206CC08 , 32'h06DEB9D8 , 32'h08908E40 , 32'h169EDBE0 , 32'h056EE808 , 32'hF7C79900 , 32'h06792320 , 32'hF02CFA60 , 32'hFFC563E2 , 32'h08559B10 , 32'hFFDEB5BE , 32'h03B78120 , 32'h07689680 , 32'h055C4420 , 32'hFFB31742 , 32'hF22198D0 , 32'hF2197430 , 32'h06535F18 , 32'h08977F90 , 32'hF15C22B0 , 32'h053591B0 , 32'h0D26CD40 , 32'hFD9FB0A0 , 32'h08423F10 , 32'hFE1BBBBC , 32'h0DBB0AA0 , 32'hF409D290 , 32'h01FE4180 , 32'hF3B91E60 , 32'h055640C0 , 32'hFAB64058 , 32'hF87C69E8 , 32'hF78661C0} , 
{32'h0312C5EC , 32'hF8E2EC88 , 32'hF87096B0 , 32'h0AE9D450 , 32'hF87D0678 , 32'hFD442DB8 , 32'hFE58C500 , 32'h129590E0 , 32'h0C2D7630 , 32'h0463BC30 , 32'hEB087AE0 , 32'hFA34F228 , 32'hF5B13580 , 32'hF94A78F8 , 32'hF65B82B0 , 32'hFEDED498 , 32'hFDD45060 , 32'h007ABC35 , 32'h066E83B8 , 32'h06FAE8C0 , 32'hFA233B68 , 32'hFAFEDC80 , 32'hFF1458CA , 32'h02CA6184 , 32'h0156CAAC , 32'hFC0A103C , 32'h012946B8 , 32'hFFCC4683 , 32'h01A1C798 , 32'hFEDA07CC , 32'h04DAA278 , 32'h020194D8 , 32'hFE293290 , 32'hFAF340B8 , 32'h05A11188 , 32'hFFA47F3D , 32'h03D0CC2C} , 
{32'hFA5F5EC8 , 32'hF4207BB0 , 32'hFC5DB1E0 , 32'h0DCA9FF0 , 32'h0119F780 , 32'h00087D8C , 32'hFB11DEE8 , 32'hFFF625EF , 32'h08BF66A0 , 32'hFC330254 , 32'h02FB3648 , 32'h0C55B010 , 32'hF9D794C0 , 32'hF921D9C8 , 32'h04702180 , 32'hF6A4B010 , 32'h01B05D90 , 32'h09FDE310 , 32'h018DEB30 , 32'hF7B53FD0 , 32'h01342F20 , 32'h043AA868 , 32'h0226BD4C , 32'h01A5AD10 , 32'hFB039808 , 32'h0927B280 , 32'h08CA22C0 , 32'h019747F4 , 32'h06D1F598 , 32'h0261C980 , 32'hFE0EDB10 , 32'hFBB98158 , 32'h002FA40C , 32'h060771E0 , 32'hF81038D0 , 32'h085591F0 , 32'hFC8A0274} , 
{32'hFFC42D55 , 32'hFED66648 , 32'hFF2DBCD7 , 32'hFF450711 , 32'hFDBE2014 , 32'h00BBBBF4 , 32'hFE4F7420 , 32'hFFF724E4 , 32'h005CBAC3 , 32'hFF13627A , 32'hFF9EA311 , 32'h01D8047C , 32'hFF2A7F6F , 32'h00CEE888 , 32'hFE699360 , 32'hFF0562DB , 32'h00AD5906 , 32'h005AF3E3 , 32'hFFD400F8 , 32'hFF235CF6 , 32'hFF7B9771 , 32'hFEA5C188 , 32'h0024FFAC , 32'h0022F5AB , 32'h014EB1C0 , 32'hFE0119DC , 32'h008C0FFF , 32'h008A0A0F , 32'hFE088B34 , 32'h002DD52B , 32'h012A3790 , 32'h01523FE4 , 32'hFFE537E9 , 32'h0022E801 , 32'h007EB54F , 32'hFEE387A4 , 32'hFFC81F7C} , 
{32'hFFFFFC16 , 32'hFFFD292C , 32'hFFFE510A , 32'hFFFAC58B , 32'h000048E2 , 32'hFFFDCC1B , 32'h00027079 , 32'h00050575 , 32'h000066CB , 32'h00028891 , 32'h00038C19 , 32'hFFFE53EB , 32'hFFFE8D43 , 32'hFFF55314 , 32'hFFFFC9E3 , 32'hFFFD46A9 , 32'h00029A13 , 32'h0004DD52 , 32'h0001F7E5 , 32'hFFFA74A1 , 32'hFFFE52EF , 32'hFFFF2715 , 32'hFFFE197F , 32'h000454DC , 32'h000140F9 , 32'h0006237A , 32'hFFFDC09E , 32'hFFFF15B9 , 32'h0000D0C0 , 32'hFFFF0C32 , 32'hFFFFB67D , 32'hFFFF385C , 32'h0004207C , 32'h00039429 , 32'h0002A163 , 32'h0000ABCE , 32'h0000E2CE} , 
{32'h0005F456 , 32'h00057560 , 32'hFFFCFD32 , 32'hFFFFADC8 , 32'hFFFF1A1C , 32'h0000E4FC , 32'hFFFC513C , 32'hFFF9E2C6 , 32'hFFFDDC07 , 32'hFFFC975C , 32'hFFF9FF8D , 32'hFFFD4829 , 32'hFFFF2D3B , 32'h00035F24 , 32'hFFFC0D1C , 32'hFFFEB2A7 , 32'hFFFF005D , 32'h0004367A , 32'h00034C4C , 32'hFFFDDE41 , 32'h00027B6D , 32'hFFFFB31B , 32'hFFFA2A52 , 32'hFFFC6B69 , 32'h00072CCB , 32'h0001AE15 , 32'hFFFD352F , 32'hFFFF48A4 , 32'hFFF75A61 , 32'hFFFE866A , 32'h00065647 , 32'h00093B2D , 32'h00007106 , 32'h00000ECA , 32'h000004A3 , 32'hFFFE10FE , 32'h0000F2D0} , 
{32'h0003A3C0 , 32'hFFFF89BC , 32'hFFFE42A8 , 32'h00028748 , 32'hFFFE5D79 , 32'h0000ADA5 , 32'hFFFFB672 , 32'hFFFE5A7B , 32'hFFFEC796 , 32'h00016A06 , 32'h00010A5C , 32'h00012FAA , 32'h00024563 , 32'hFFFE4A58 , 32'hFFFAD128 , 32'h0001988B , 32'h00002A45 , 32'hFFF76E61 , 32'hFFF9EC2A , 32'hFFFDE313 , 32'h00017882 , 32'hFFFF2B4B , 32'h00020E2F , 32'hFFFFB8B5 , 32'h0006095C , 32'hFFFB7180 , 32'hFFFB62EB , 32'hFFFF42B2 , 32'h00047721 , 32'hFFFEB1B9 , 32'hFFFD1D50 , 32'hFFFD8B2E , 32'h00042BB6 , 32'hFFFECB1C , 32'hFFFE0941 , 32'h00027A0F , 32'hFFFEB160} , 
{32'hFFFE6FFE , 32'hFFFF88BA , 32'h000090AC , 32'h0002DE40 , 32'hFFFB0486 , 32'h0001A4F8 , 32'hFFFBB70B , 32'hFFFBD7DD , 32'hFFFC195B , 32'h0003E430 , 32'h0001FD00 , 32'h0005DC2C , 32'hFFFEEEAA , 32'hFFF7C9B7 , 32'h0001F73B , 32'hFFFFD262 , 32'hFFF964DF , 32'h00084D1C , 32'h00012D5F , 32'hFFFD3299 , 32'h00059C5C , 32'hFFFEBA0A , 32'hFFFDC593 , 32'h00025ACD , 32'h0001BFBA , 32'hFFFE7957 , 32'h00047411 , 32'h0004AF65 , 32'hFFFEB15D , 32'hFFFF58A8 , 32'hFFFFD452 , 32'hFFFCDB7F , 32'hFFF9537F , 32'hFFFC4EC2 , 32'hFFFBA527 , 32'hFFFC0644 , 32'h00014D0E} , 
{32'h0037174D , 32'hFFCF870A , 32'hFFEB333A , 32'hFFFD3600 , 32'hFFE1546E , 32'h00458478 , 32'hFFDE298F , 32'h000971DF , 32'hFFBCDFA1 , 32'h0010515A , 32'h003D0863 , 32'hFFEB97D0 , 32'hFFC58C3A , 32'hFFE9FDE0 , 32'hFFDD8C78 , 32'hFFBB3E06 , 32'hFFDF63D0 , 32'hFFFDA47E , 32'h000B21F4 , 32'h003A46C3 , 32'hFFFE4840 , 32'h0014D12D , 32'h003EA169 , 32'hFFF3AB11 , 32'hFFF26B70 , 32'h0003A6BD , 32'hFFA61B58 , 32'h000B7641 , 32'h0017CD07 , 32'hFFEE514F , 32'h0023CE47 , 32'hFFE6B21B , 32'hFFC29202 , 32'h00198D55 , 32'hFFD05BBF , 32'h000E5B5B , 32'h00133F2E} , 
{32'h0048977D , 32'hFFD441F4 , 32'hFFD844B2 , 32'hFFF22BB2 , 32'hFFCB6A9B , 32'h00623D13 , 32'hFFD47768 , 32'h001A1E41 , 32'hFF951255 , 32'h00121C06 , 32'h0066C7F3 , 32'hFFD4EB2E , 32'hFFBD28BF , 32'hFFEC86C1 , 32'hFFD37A12 , 32'hFFA7A813 , 32'hFFF36BB6 , 32'hFFE713F4 , 32'h00016916 , 32'h004B89AA , 32'h00169C03 , 32'h00061236 , 32'h0057147B , 32'h000665EE , 32'h0003D28B , 32'h0000EE50 , 32'hFF9C9520 , 32'h000B254D , 32'h00246507 , 32'hFFE22D9E , 32'h003A2A39 , 32'hFFE1739C , 32'hFFA6B3A0 , 32'h001352F6 , 32'hFFC5A1A8 , 32'h000D6C0F , 32'h0025F2FD} , 
{32'hFED45A38 , 32'hFABC4EE8 , 32'hFF620B4C , 32'h022008DC , 32'h08594900 , 32'hFAE01490 , 32'hF4522E90 , 32'hF9BBB0C0 , 32'hF7019500 , 32'h03EC073C , 32'hF216F9A0 , 32'hFE95B500 , 32'h02848740 , 32'h04BCCF50 , 32'hF2EA58E0 , 32'hF7CCD680 , 32'hF90A93E0 , 32'hF3D6E5E0 , 32'hFCB7E468 , 32'hF3907960 , 32'hFF764E24 , 32'hFED237E4 , 32'hF9C4D8E0 , 32'hFC2622D0 , 32'hFF923210 , 32'h055184A0 , 32'hF74A76E0 , 32'h04A7FCF8 , 32'h00270CD6 , 32'h0D15E1B0 , 32'hF99CB4A8 , 32'h0BD3D100 , 32'hFC236900 , 32'h00DB5474 , 32'hFD2D4138 , 32'h02FDFB00 , 32'h05B8FF90} , 
{32'hE11D7E80 , 32'hD1FE2C40 , 32'h081E2A20 , 32'hFB5D1668 , 32'h2BB16000 , 32'h049B47F0 , 32'h0A674470 , 32'h03F51160 , 32'hEBA98440 , 32'h03390A24 , 32'hF854C260 , 32'hFE01A20C , 32'hF349DBA0 , 32'h11A8DCC0 , 32'hFC266014 , 32'h0EBABFC0 , 32'hFC5F452C , 32'hF8D59FD8 , 32'hF6FC2F80 , 32'h0A712760 , 32'h0BCA8CB0 , 32'h09728230 , 32'h00E1C22E , 32'hF6C5F620 , 32'hEF897AC0 , 32'h0CDB7440 , 32'h07D0DE50 , 32'h0CBEB730 , 32'h16A08B00 , 32'h0D5DC9C0 , 32'hFD922D40 , 32'h0782F778 , 32'h036DD7EC , 32'h0BF00070 , 32'hFF253BDC , 32'h0828A710 , 32'h061B74C0} , 
{32'hED29EBC0 , 32'hE97937A0 , 32'hEB9838A0 , 32'hEC469600 , 32'h28A89A00 , 32'h0E7581E0 , 32'h0C2EDA40 , 32'h0878D200 , 32'hF2CAD880 , 32'h011B4754 , 32'hF1B40810 , 32'h0C226CA0 , 32'hFCEFD0B8 , 32'hFF245901 , 32'h01C452B8 , 32'h0C521A90 , 32'h06176BE0 , 32'hF9C56AE0 , 32'h0460CC08 , 32'hFEFA8D2C , 32'h02CBA584 , 32'hFD83C898 , 32'h060A0C10 , 32'h00A9CFBF , 32'hF3E8CE00 , 32'h03410670 , 32'hFE20D11C , 32'h06265990 , 32'h000D50AE , 32'hF3C21AA0 , 32'h0B2E6250 , 32'hF3D24B70 , 32'hF953A478 , 32'hF71EF760 , 32'h07838550 , 32'hFD3A8468 , 32'hFFD1E495} , 
{32'hED9DADC0 , 32'hDBCD9900 , 32'hF9789028 , 32'hFA7CC950 , 32'h28B27780 , 32'h24E021C0 , 32'h185800A0 , 32'h0B9E27A0 , 32'hEF4CD1E0 , 32'h08547710 , 32'hF6C07540 , 32'hEDC218C0 , 32'h1054B200 , 32'h117D3040 , 32'h09C46310 , 32'hF9E4C7F0 , 32'h20593200 , 32'hFA14F978 , 32'hFEB1A788 , 32'hF830D450 , 32'hDB79ED00 , 32'hF6930170 , 32'hE900A100 , 32'h01512490 , 32'hE205EC20 , 32'h0EE10B80 , 32'hFF4878FB , 32'hFF3C9089 , 32'hDD9D9700 , 32'hDB9F1D40 , 32'h24D5B740 , 32'hE516B2C0 , 32'hFB2ED788 , 32'h0C145AE0 , 32'h0D0E8350 , 32'h1C242520 , 32'hFD71EED8} , 
{32'hEEA2FCC0 , 32'hD34D7600 , 32'hFE55E72C , 32'hFAC53D28 , 32'h3DCAA000 , 32'h22679800 , 32'h14B63800 , 32'h09815890 , 32'hE6C9C160 , 32'h0BEAD5F0 , 32'hE43AB320 , 32'hFFF538B4 , 32'hFA4B9300 , 32'h23034300 , 32'h2488A440 , 32'hEF81C640 , 32'h05BA4CA0 , 32'hF8446E88 , 32'h0B86F230 , 32'h1857FA40 , 32'hFFDD38A4 , 32'hE8206600 , 32'hF9F69400 , 32'h016C936C , 32'hE0202E00 , 32'h0469BDB8 , 32'h095D3E90 , 32'h01030200 , 32'hEEB29320 , 32'h0B3B51F0 , 32'h21C1A1C0 , 32'hF4C448E0 , 32'hF0A646F0 , 32'hF9599EA0 , 32'hFED8A83C , 32'hF7349D10 , 32'hE9E7B2A0} , 
{32'hE507D000 , 32'hBDF87B00 , 32'hE4660E80 , 32'hEE2B9480 , 32'h30899E40 , 32'h16759EC0 , 32'h24A74580 , 32'h05F2BA88 , 32'hEC0CCEA0 , 32'h0E7A5300 , 32'hE8879CA0 , 32'hF0A088B0 , 32'h06134540 , 32'h01620DA4 , 32'h26F461C0 , 32'hF8845E18 , 32'hFE007EC8 , 32'hFDBF436C , 32'hFAFD42C8 , 32'h03C29ECC , 32'hF9F96E00 , 32'hF8E2DE18 , 32'hFC8DC7C8 , 32'hFD10AA3C , 32'hF75EC0E0 , 32'hFCC6C7B4 , 32'h040B74F0 , 32'hFF3FBE11 , 32'hE26C9420 , 32'h07AE4960 , 32'h0CAEFF70 , 32'hE3F6A0C0 , 32'hFCE2C5F0 , 32'hFF211195 , 32'h02618A84 , 32'hF0357D10 , 32'hF372F4A0} , 
{32'hE558D860 , 32'hCD26A600 , 32'hEF71FB00 , 32'hD1E55BC0 , 32'h1BFD8FA0 , 32'h18C0A780 , 32'h2B1660C0 , 32'h05555CA0 , 32'hE8E13AE0 , 32'h28228CC0 , 32'hD8950980 , 32'hF56C0BE0 , 32'h183BC040 , 32'hC6798380 , 32'h08B2F040 , 32'h013F15A8 , 32'hFE0A7F64 , 32'h2F55C6C0 , 32'hED142A60 , 32'hF784FBF0 , 32'h03960BCC , 32'hF86E1158 , 32'h191F5F60 , 32'h047176C0 , 32'h14D143A0 , 32'h01FD3510 , 32'hF5A4C5F0 , 32'hF9FBAB08 , 32'hFF534E7C , 32'hE1E31C60 , 32'h010202D8 , 32'hEFBAA5E0 , 32'hFCCCFB44 , 32'h00285C4E , 32'hFEDB447C , 32'h0CA8C0B0 , 32'hFC0375D8} , 
{32'hE308F6E0 , 32'hC05E9F80 , 32'hD8D83F80 , 32'hCC17FC00 , 32'hEEE1D240 , 32'h134800E0 , 32'h44751E80 , 32'h094823E0 , 32'hEC3521E0 , 32'h13C7D420 , 32'hEA7CB5C0 , 32'h1DF6C7C0 , 32'h1597B6A0 , 32'hDA850BC0 , 32'hEF0F3620 , 32'h0A428020 , 32'h06962D18 , 32'h24B4A900 , 32'hFE6F55D8 , 32'hD7D6DD40 , 32'h1436FBE0 , 32'h0DF958B0 , 32'hFBB430C0 , 32'hEE9EE660 , 32'h007D460C , 32'hF70E1040 , 32'hE0BBA960 , 32'hE68128E0 , 32'h0EAB8060 , 32'hFBB66400 , 32'hFC9C3F08 , 32'hFAFDD480 , 32'h035BC814 , 32'hFF71BF9D , 32'h02225620 , 32'hE592E3E0 , 32'h126876E0} , 
{32'hE8F4FFE0 , 32'hC5876140 , 32'hDDA4A680 , 32'hD9AD1CC0 , 32'hC3211B40 , 32'h091F3E10 , 32'h42F09280 , 32'h00F9C565 , 32'hF2DFD6A0 , 32'h012F7F9C , 32'h0860A040 , 32'h3303EE40 , 32'h0C0EA4F0 , 32'h0624D1F8 , 32'hCCF93680 , 32'h1B17FF60 , 32'h0F93BC00 , 32'hE25B2A00 , 32'h1CBDCA00 , 32'hEAE1F0A0 , 32'hE9F68720 , 32'h15DAC880 , 32'hDBC852C0 , 32'hED943880 , 32'h0E255B20 , 32'h115F9220 , 32'hF8905698 , 32'hF16FA830 , 32'h2984D500 , 32'hE88D4880 , 32'hF76AFD40 , 32'hF6FAA4C0 , 32'hFBC6FA80 , 32'hF18D2D10 , 32'h0DC48E60 , 32'h088E19E0 , 32'h076DC2F0} , 
{32'hF8E1ECE0 , 32'hF98BDB80 , 32'h118822A0 , 32'h0D626FC0 , 32'hF8624AA0 , 32'h161F6DE0 , 32'h179968E0 , 32'h14FA8B40 , 32'hEB7B35C0 , 32'hF93CF778 , 32'hEAA6E060 , 32'h21D67A80 , 32'h0B66FEB0 , 32'h177070A0 , 32'hF64105B0 , 32'h05FA3FB0 , 32'h14507100 , 32'hE642A360 , 32'h05734430 , 32'hFBBD0290 , 32'hF48DBE50 , 32'hF4AA0A90 , 32'h0A41F650 , 32'hFC14D9B4 , 32'h01FF9AB0 , 32'h04D9EE30 , 32'h0C056140 , 32'hEFAA26A0 , 32'h178F1FA0 , 32'hEECADEC0 , 32'h04927330 , 32'h0817D870 , 32'h06E7BCC0 , 32'hF9A15CA8 , 32'h02870524 , 32'hF4C5EF80 , 32'hFDEE55D0} , 
{32'hF7121A20 , 32'hFCE2CA1C , 32'h0AEE13C0 , 32'h04104E28 , 32'hF5A95AE0 , 32'h119E4500 , 32'h03464238 , 32'h112F1E00 , 32'h0120E0FC , 32'hF8465AC8 , 32'h073CC408 , 32'h0F306050 , 32'hF0F087C0 , 32'h1C4773C0 , 32'h0050DA8C , 32'h0896F880 , 32'h063E3200 , 32'h089A5410 , 32'h0B903700 , 32'hFF64DCD4 , 32'h0299EAB8 , 32'h0000AA30 , 32'hF6588470 , 32'hF3A9B980 , 32'h04860120 , 32'hF932EF08 , 32'h11E73340 , 32'hF4D4B980 , 32'hFD51F704 , 32'hEC6E1860 , 32'h0EAB8510 , 32'hFC23EF9C , 32'h08985DB0 , 32'hF215B320 , 32'h064F2B30 , 32'hE5CA98C0 , 32'hF3A03470} , 
{32'hFF2D5E89 , 32'hF6589B10 , 32'h1054C760 , 32'h2A380F80 , 32'h0B6A0140 , 32'h01213268 , 32'hE632A7E0 , 32'hF0007D10 , 32'hF77A5E60 , 32'h0E172990 , 32'hF503F9E0 , 32'h1D4472A0 , 32'h08BA16B0 , 32'h0FD927C0 , 32'hF6604B50 , 32'h2A7F1C80 , 32'hFD78D110 , 32'h0C5E9CE0 , 32'h149A2B60 , 32'h21597580 , 32'hF401D130 , 32'hFE22DE8C , 32'hEBF359A0 , 32'h13435C00 , 32'h16CB97E0 , 32'hE67A4FE0 , 32'h002AC74B , 32'hF1BBC8B0 , 32'hFFDFCFC2 , 32'hFD244ABC , 32'hFE3BF200 , 32'h025E413C , 32'hEB610DC0 , 32'h02346CBC , 32'hFB511DD0 , 32'hEE83E660 , 32'hFCFFD0D8} , 
{32'hEFEEC480 , 32'hF79109E0 , 32'h110CACE0 , 32'h1B44B880 , 32'h16D69800 , 32'h11529060 , 32'hE1E38C60 , 32'hD8FA08C0 , 32'h0EB1ABC0 , 32'h0D57A0D0 , 32'h159684A0 , 32'h0AF4A030 , 32'h254719C0 , 32'hFEFFC25C , 32'hF7D5E950 , 32'hF98B8450 , 32'h20D6BC80 , 32'h0B466210 , 32'h041FCCD0 , 32'h0B3DAAE0 , 32'h027BDCAC , 32'hF562C970 , 32'h10B98500 , 32'hD1563600 , 32'h10D0EDE0 , 32'hF0BBDF20 , 32'h09682410 , 32'h099965C0 , 32'h1D0DBB00 , 32'h0975C5C0 , 32'h02A7D368 , 32'hFAD043D8 , 32'h0BD78040 , 32'h09213730 , 32'h03FBAFB0 , 32'hF0B04350 , 32'h0BE61580} , 
{32'hF4026D10 , 32'hF7FBFD00 , 32'h07DA4D50 , 32'h15B11E40 , 32'h16561960 , 32'h0FC1F1D0 , 32'hF0814F80 , 32'h08AA5460 , 32'h08788C10 , 32'h0ADAF700 , 32'h128D82C0 , 32'hF68ECB80 , 32'h176CFC20 , 32'hFEDCE704 , 32'hFC6262BC , 32'h00487EDD , 32'h15B4C320 , 32'h0D394B20 , 32'h108C70C0 , 32'hF6DBF950 , 32'hFC74B1F0 , 32'hF3372430 , 32'hF717D7C0 , 32'hF7CB95F0 , 32'hFF0E31EF , 32'h063718C0 , 32'hED2CEB40 , 32'h011AC708 , 32'h06BED450 , 32'hF163D310 , 32'h03949494 , 32'hF30038E0 , 32'h057B4648 , 32'hFE9B45FC , 32'hF531F940 , 32'h070B9DF0 , 32'h1BE8CA20} , 
{32'h00798721 , 32'hEBDE3F80 , 32'h065FAA10 , 32'h1B494160 , 32'h1006A620 , 32'h06967910 , 32'hED5A4300 , 32'hF9D0EF00 , 32'h0E4E92D0 , 32'h058A89B8 , 32'h1CE494C0 , 32'hF4A0B7A0 , 32'h10306F60 , 32'hF99E24D0 , 32'h01B116B8 , 32'hFAA489B8 , 32'h17A82720 , 32'h04D31C48 , 32'h01A543A4 , 32'hEDA47C80 , 32'hF9731E10 , 32'h00F3BFE2 , 32'hFF659BD3 , 32'h079D4438 , 32'hF6399560 , 32'hFDE51054 , 32'hF93E1A30 , 32'h08A95390 , 32'h0E272570 , 32'hEEC5EF80 , 32'h025CDB0C , 32'h03BD70B0 , 32'hFC2FEEBC , 32'hE99E5CA0 , 32'h076A73D8 , 32'hEB7F0320 , 32'hFAFCF458} , 
{32'h1166F120 , 32'h16881A40 , 32'hE9382D20 , 32'hFC476E88 , 32'h0BFA7F50 , 32'hFE9A1A4C , 32'h023D895C , 32'h059601E8 , 32'h1654E7C0 , 32'hF6D49B20 , 32'h04158110 , 32'hF793AF60 , 32'h01CB36B0 , 32'hF78C23B0 , 32'h04DC7F50 , 32'hF05122C0 , 32'h05B6F460 , 32'hFAC3CFA0 , 32'h10232640 , 32'hD4ECAA40 , 32'hE5C29260 , 32'h00D1AA16 , 32'h190EB8A0 , 32'hF73EC0C0 , 32'hE044C300 , 32'hFD5016AC , 32'hFA7901F8 , 32'hF9D0F448 , 32'hDA919800 , 32'hEC8D1D40 , 32'h07B73890 , 32'h10A6B780 , 32'h00B1DAC1 , 32'hE3C9B360 , 32'hF55000E0 , 32'hD96C64C0 , 32'hFC9882E8} , 
{32'hF73A8140 , 32'h07D9DBE0 , 32'h06132038 , 32'hF9D577F0 , 32'h00755CC7 , 32'h07A4EF18 , 32'hFB37DCB0 , 32'hEF5E0580 , 32'hF5982EE0 , 32'hDF8B5180 , 32'h0F121550 , 32'h012E28CC , 32'h082B0A10 , 32'hF305BFC0 , 32'h00402E1E , 32'h0D9CAE80 , 32'h0203AD04 , 32'hF0F5A910 , 32'hF630E560 , 32'hEB9D0D80 , 32'hFDBB81F4 , 32'h0196F2A4 , 32'h01A60F5C , 32'hEF56CE40 , 32'h020CCD18 , 32'h07659B80 , 32'h04649588 , 32'hFE7ABA1C , 32'h00344BC2 , 32'hFE0F3EC4 , 32'h0638DAC0 , 32'hF70ABDB0 , 32'hE901DE20 , 32'hF5BEA1A0 , 32'hF55B1550 , 32'hF0C66BC0 , 32'h04E4DDD0} , 
{32'hFB32D7B8 , 32'h0332413C , 32'hF9FE1A40 , 32'h02DA07A4 , 32'hFEB73FBC , 32'h051D1618 , 32'h0615F5C0 , 32'h0CBE9570 , 32'h07268490 , 32'hF4336CE0 , 32'h0B11CC20 , 32'h078D7D28 , 32'hFC0DF374 , 32'h045CBE70 , 32'h008A1FDC , 32'hF5A97800 , 32'h0E770F90 , 32'h1063DEA0 , 32'hF9F54528 , 32'h0120FF64 , 32'h01F7DEF4 , 32'hFB0AC970 , 32'h01968030 , 32'hF9E0EAE0 , 32'h0146253C , 32'hFBA08728 , 32'hFF3BBF5B , 32'hF5D375F0 , 32'hF4340260 , 32'h0AE89500 , 32'hF700A290 , 32'h09E3CFE0 , 32'hFE48A16C , 32'hF9C5F3F0 , 32'h07A9BD80 , 32'h073C87C8 , 32'h10745E60} , 
{32'hFB9CE940 , 32'h0E17B260 , 32'hFFAFAEDA , 32'hFB3D5DF0 , 32'h11B49960 , 32'h0B161760 , 32'h0F6913D0 , 32'h05F8B500 , 32'h0D8F56E0 , 32'hE50332C0 , 32'h02A54CD0 , 32'h01A252C0 , 32'h0AB5E850 , 32'hF7FB9390 , 32'h0DEDEF50 , 32'hFAA8CF30 , 32'h01A5D8F8 , 32'hF984DB48 , 32'h03350CC8 , 32'hF3426A50 , 32'hFB5710F0 , 32'h16E0C780 , 32'hF86B6848 , 32'hF0C00B80 , 32'h0587B278 , 32'hF0717120 , 32'h1E770060 , 32'h027998E4 , 32'hF2738860 , 32'hFF14BA11 , 32'hEBE14F60 , 32'h0D4B58F0 , 32'hFACAA088 , 32'h012846F4 , 32'h0F931B10 , 32'h14BE2AC0 , 32'h1930C740} , 
{32'h001905EF , 32'hFF33530C , 32'hFE300538 , 32'hFDCE5A54 , 32'hFE983E44 , 32'hFEECF87C , 32'h025B6688 , 32'hFFF79982 , 32'hFF17C976 , 32'hFE4E5AEC , 32'hFF939113 , 32'h00C31482 , 32'hFDD736C4 , 32'h0147D71C , 32'hFD0C10A4 , 32'h0472DC98 , 32'hFE34D0BC , 32'h00A42B58 , 32'h01A3989C , 32'hFEA80F28 , 32'hFAF40C40 , 32'h045EB498 , 32'hFC6A7F04 , 32'h02F96F1C , 32'h009D846F , 32'h032CBDDC , 32'h00B8626E , 32'h02C4A908 , 32'h0090BE79 , 32'hFDF350E4 , 32'hFFCFC761 , 32'hFEC48218 , 32'hFE56DC7C , 32'h00AAB52A , 32'h019CD0D0 , 32'h00C36415 , 32'h0292BB04} , 
{32'hFFFB515C , 32'hFFFFC4B2 , 32'h00039281 , 32'h0004CFDF , 32'hFFFF7020 , 32'hFFFE03B7 , 32'hFFFF8B26 , 32'hFFFE38A8 , 32'h00012328 , 32'hFFFED40C , 32'hFFFC5408 , 32'h000049FD , 32'h00031F22 , 32'hFFFE259E , 32'h0003042B , 32'h00035F2A , 32'h00017F5F , 32'h0002F2E2 , 32'hFFFEF543 , 32'hFFFB29F7 , 32'h0001AC1A , 32'h00001605 , 32'hFFFB5F6D , 32'h0003E257 , 32'h0002BB1A , 32'hFFFD9BB7 , 32'hFFFE40C2 , 32'h00003BE3 , 32'h000546A8 , 32'hFFFE873A , 32'hFFFFFDBA , 32'h0002AE63 , 32'h00015E44 , 32'h00018AC7 , 32'hFFF9E34F , 32'h00017434 , 32'h0000D760} , 
{32'h0000353E , 32'h00018B57 , 32'h0003C746 , 32'hFFF91FD7 , 32'hFFFA778D , 32'h00049EBB , 32'hFFFD7317 , 32'h00017768 , 32'h0001CF54 , 32'h00008213 , 32'h000048A9 , 32'hFFFE8D11 , 32'h00009976 , 32'hFFFBBB42 , 32'h00028D18 , 32'hFFFFC762 , 32'hFFFFE362 , 32'h0000CBC9 , 32'hFFFCE422 , 32'h00005C1C , 32'h0000978C , 32'h00038638 , 32'hFFFB88D5 , 32'hFFFE4DAB , 32'hFFFF8A9D , 32'hFFFC0339 , 32'h0003FEE5 , 32'hFFFD5248 , 32'h0004504A , 32'h000656FF , 32'hFFFDB78C , 32'hFFFDFE3E , 32'h0002042D , 32'hFFFF4852 , 32'hFFFE4FE1 , 32'h0000E4A8 , 32'hFFFFCEED} , 
{32'hFFFA7C44 , 32'h00006A1F , 32'h0007942C , 32'hFFFEF33B , 32'hFFFF6072 , 32'h0003873F , 32'hFFFEF212 , 32'hFFFF1A88 , 32'h000397A3 , 32'h00060769 , 32'hFFFEE117 , 32'hFFFF5270 , 32'hFFFA93CE , 32'h0001FD9C , 32'h000116D1 , 32'hFFFDB21E , 32'h0001606C , 32'hFFFC1E7D , 32'h0001BD43 , 32'hFFFD19FF , 32'h00028F14 , 32'h0006173B , 32'hFFFDE029 , 32'hFFF64893 , 32'hFFFCE940 , 32'hFFFE477A , 32'h000110AC , 32'h00000101 , 32'hFFFCDCA2 , 32'hFFFDEABC , 32'h000093D7 , 32'hFFFC59C0 , 32'h0004A3BD , 32'hFFFDE31E , 32'hFFFF6C06 , 32'hFFFF0CAC , 32'hFFFB7C8F} , 
{32'hFFFE32E2 , 32'h0000F564 , 32'h0004FFE7 , 32'hFFF93E92 , 32'hFFFF2A35 , 32'hFFFE446E , 32'hFFFF733C , 32'h00045ABC , 32'h00016B0B , 32'h00074F79 , 32'hFFFEDD3D , 32'hFFFFC1EB , 32'hFFFDB12F , 32'hFFFA95F3 , 32'h00066B9F , 32'h00028988 , 32'hFFFF01EC , 32'hFFFDA1DB , 32'hFFFB0A51 , 32'h000238AF , 32'h0003D3CA , 32'hFFF9C713 , 32'hFFFEBB18 , 32'hFFFE1049 , 32'hFFFF12E2 , 32'h0000F03D , 32'h0000DE91 , 32'hFFFE9439 , 32'h0007C427 , 32'hFFFFCC0B , 32'hFFFECBC9 , 32'h000538CD , 32'h0002401C , 32'h000593D4 , 32'hFFFF4466 , 32'hFFFC0A2E , 32'hFFFCBDDD} , 
{32'h00020D15 , 32'h00008849 , 32'h00057332 , 32'h00079FFB , 32'hFFFACA47 , 32'hFFFD8F44 , 32'hFFFF18AC , 32'h00039AED , 32'hFFFB7186 , 32'hFFFBEB55 , 32'h0001F5A3 , 32'hFFFEADCE , 32'h000448CA , 32'hFFFD74B1 , 32'h0003EDCA , 32'h00009E28 , 32'h000187EC , 32'h00035AB5 , 32'hFFFD4238 , 32'h00004793 , 32'h000175BD , 32'h0001E002 , 32'hFFFDFBA7 , 32'hFFFF5876 , 32'hFFFCAFEA , 32'h0002DB9A , 32'hFFFF5956 , 32'hFFFD9503 , 32'hFFFEFE38 , 32'h0004123E , 32'h00001451 , 32'hFFFED6D8 , 32'h00014C10 , 32'hFFFEDD16 , 32'h0000439A , 32'h000B2C31 , 32'hFFFF5682} , 
{32'h00022F5D , 32'h00005A69 , 32'h0001C48B , 32'hFFFC55F6 , 32'hFFFE86A5 , 32'hFFFFC756 , 32'h0001A72D , 32'hFFFC9A71 , 32'h00022AEA , 32'h0002E155 , 32'h0003C033 , 32'h0000C620 , 32'hFFFF5896 , 32'hFFFE29EF , 32'hFFFF12C9 , 32'hFFFCFBDF , 32'hFFFA70A8 , 32'hFFFD2A4D , 32'hFFFCDC39 , 32'h000277E0 , 32'h00056D08 , 32'hFFFBC23A , 32'hFFFEDBE2 , 32'h0001F587 , 32'h00071ABB , 32'h00061F9E , 32'h00018AB0 , 32'hFFF9CAC4 , 32'h000314EB , 32'h0004BC32 , 32'h00009394 , 32'h0000AAF5 , 32'h00022D37 , 32'h0001F915 , 32'h00026C2E , 32'hFFFDF88A , 32'h00046423} , 
{32'h0003B6BF , 32'h0008A4FE , 32'hFFFC014B , 32'hFFFF2147 , 32'hFFF9C832 , 32'h00026B2C , 32'h000AFBC3 , 32'h000A274C , 32'h00035FDF , 32'h000723DD , 32'h00026911 , 32'hFFFF48A3 , 32'h000C907D , 32'h0000F5FD , 32'hFFF7EFE9 , 32'h0005BC22 , 32'h00010F8D , 32'hFFF7AB1E , 32'hFFFCFF34 , 32'hFFFDCE50 , 32'h00047929 , 32'hFFFFB0D7 , 32'hFFFE6D40 , 32'h00065153 , 32'h0004F153 , 32'h0000CBBE , 32'h0002D103 , 32'h0000D69C , 32'hFFFD10A5 , 32'hFFFF8E90 , 32'hFFFF376A , 32'hFFFD2601 , 32'h00042A1C , 32'h00025DD1 , 32'hFFFE94D0 , 32'hFFFDA81A , 32'hFFFE85EB} , 
{32'hFEE42BDC , 32'hFD807EBC , 32'hFE4012B4 , 32'hFE7E0FD4 , 32'h00A2C646 , 32'h0231FE48 , 32'h02031FB0 , 32'hFF472A26 , 32'h0043E1C4 , 32'h024D70AC , 32'hFDD73DE4 , 32'hFE4E7C2C , 32'hFF94C15D , 32'hFF372273 , 32'h070E0DD0 , 32'hFE92E2C0 , 32'h024EF758 , 32'hFD4D070C , 32'h0183A924 , 32'h00E97B7B , 32'hFDB057AC , 32'hFEDC9B7C , 32'h0031D2AE , 32'h02734794 , 32'h043FF6C8 , 32'hFE8FD18C , 32'hFE2EBABC , 32'h00CF334E , 32'hFF624800 , 32'h04336888 , 32'hFD045D50 , 32'h025CE494 , 32'h0340B458 , 32'hFCDF12C4 , 32'h000F230E , 32'h011F6278 , 32'hFFC6E249} , 
{32'hF8990C70 , 32'hF0735C50 , 32'hFDE112C8 , 32'h0C1E6760 , 32'h0746DDF8 , 32'h00EE62E2 , 32'hFE12AAD4 , 32'hF4FC1FC0 , 32'h03BF5DF8 , 32'hFD961E84 , 32'hFF055BCB , 32'h0AFC9A30 , 32'hF163C7D0 , 32'hF9230AE0 , 32'h1032CD00 , 32'hF58ECBA0 , 32'hFEDD9868 , 32'h12BF2860 , 32'h10762A60 , 32'h01B61D2C , 32'hEA9D4740 , 32'h0BAF8200 , 32'h0A3D6940 , 32'hEE1AB600 , 32'hFB6BC938 , 32'h097ED1F0 , 32'hFDC09868 , 32'h018318AC , 32'h0C97C9A0 , 32'h0C6C4090 , 32'hFF867EC5 , 32'h07085E98 , 32'h145FCE40 , 32'h03E144A4 , 32'h001CA916 , 32'h0CB85FA0 , 32'h00912D10} , 
{32'hEE25B1A0 , 32'hEF5A0EA0 , 32'hDFEE6840 , 32'hFE335A94 , 32'h14CA9F60 , 32'h0B041A90 , 32'hEAEFAAA0 , 32'h003C9871 , 32'hE9B39600 , 32'hF19BB7C0 , 32'h0E41F300 , 32'h07242AE0 , 32'hEA4817E0 , 32'hF48953C0 , 32'hFF5FAEF5 , 32'hF7D15C50 , 32'hEEEAE360 , 32'h00B75E11 , 32'h1871B140 , 32'h0EA6C870 , 32'hF8D5E768 , 32'hFBE52EB8 , 32'h0B8899E0 , 32'hF4F4E280 , 32'h03D9F86C , 32'h0B56FAE0 , 32'h05122388 , 32'h04C3F410 , 32'h0644D2C0 , 32'h106371A0 , 32'h0342D0C8 , 32'hF4F22EE0 , 32'h04278D90 , 32'hF2C8EBE0 , 32'h0F295030 , 32'h03A3C1A0 , 32'hFE73261C} , 
{32'hFA30B2D8 , 32'hFC4E9F0C , 32'hEBD2B320 , 32'h03ACC4B8 , 32'h1DFF2D00 , 32'hF43628A0 , 32'hE4AFDF20 , 32'hF77DDD90 , 32'hF7BC4770 , 32'hF8E4CDF0 , 32'hFF31518B , 32'hF5796730 , 32'h00E201CB , 32'h13380580 , 32'h12536220 , 32'hF05295C0 , 32'hF30C3340 , 32'hF5367740 , 32'h082B46B0 , 32'h08B3D2A0 , 32'hF9E2C3F8 , 32'hEF540620 , 32'hFFBE04C6 , 32'h072F4310 , 32'h09DBB600 , 32'h0B8FB3E0 , 32'h01F72B68 , 32'hFDD901B0 , 32'h046FC810 , 32'h07AA9458 , 32'h091D2440 , 32'hF9EB7BC8 , 32'hF2042EF0 , 32'hFE65DD5C , 32'h1A02E980 , 32'h08772F10 , 32'h04643E00} , 
{32'hF2508680 , 32'hEDEADB20 , 32'hE2ACF0E0 , 32'hE894F0C0 , 32'h2C485200 , 32'hF8293A28 , 32'hEA19DA80 , 32'hFFAFB642 , 32'hF21524D0 , 32'h03447C10 , 32'hEFFB40C0 , 32'hFA6D7290 , 32'h0E7390C0 , 32'hF9348E00 , 32'hEB488320 , 32'hFF420222 , 32'hF6872CA0 , 32'h02F6F88C , 32'hEF40FA60 , 32'hF6D79230 , 32'hF4AC6390 , 32'h03C494C4 , 32'h1514E5E0 , 32'h0E0EB2C0 , 32'h0BD6B8A0 , 32'h03F147B8 , 32'h04F2FFF8 , 32'h00B51298 , 32'hFE8C1FDC , 32'hFA1AE608 , 32'hFD4F2154 , 32'h1648B760 , 32'hFF91ED87 , 32'hEEF64180 , 32'h07AA9B60 , 32'h135575A0 , 32'h0B7CE230} , 
{32'hEDCCB040 , 32'hE33EB580 , 32'hE251AFE0 , 32'hEA0975C0 , 32'h3F2D8140 , 32'hFFBBFE7A , 32'hF42C7DD0 , 32'h0A6BFEA0 , 32'hFE16096C , 32'h05CF9A38 , 32'hFC89AF50 , 32'hF288D630 , 32'h0DFC38D0 , 32'hF3F9D160 , 32'hFF54CB95 , 32'hF5AB5440 , 32'hFB3CACD0 , 32'h0F18B250 , 32'hED8B0200 , 32'h0A772CF0 , 32'hE94589E0 , 32'hF04B6200 , 32'h0FEE5190 , 32'h08941810 , 32'h1045BB20 , 32'h04C57230 , 32'hFEEE3DAC , 32'hF9C0BE20 , 32'hE49C3DA0 , 32'hEAA827A0 , 32'h02F3ED34 , 32'hEED33AE0 , 32'hF9846940 , 32'hFD01C02C , 32'hF8646BD8 , 32'h05118E08 , 32'h042ABEE8} , 
{32'hE8A0ECC0 , 32'hD7B22BC0 , 32'hE6F51580 , 32'hDEFC34C0 , 32'h25BFA3C0 , 32'h069B4700 , 32'h27AF2500 , 32'h0B3079A0 , 32'hEDF20A80 , 32'h031A5FF4 , 32'hE7B5A140 , 32'hF7C4BD40 , 32'h008E51C2 , 32'hF6A91D40 , 32'h15947580 , 32'hED373140 , 32'hF17BDD90 , 32'h13E1BA20 , 32'hFB477970 , 32'hF7BBAD40 , 32'h08B3ED70 , 32'hFB096998 , 32'h06D892B0 , 32'h04D077C8 , 32'h08240560 , 32'hEF55FDA0 , 32'hFA82E0C0 , 32'hFDEFA774 , 32'hF1BC1BD0 , 32'hFF915273 , 32'hF969CF88 , 32'hF1C374D0 , 32'h03B57900 , 32'h071EE6B0 , 32'h02B8BB00 , 32'hE182E220 , 32'hF2014E20} , 
{32'hE5EF3680 , 32'hBC0EED80 , 32'hB5F09C00 , 32'hDBAE5600 , 32'h2714DE80 , 32'h020671CC , 32'h3A51F380 , 32'h06E26E38 , 32'hFB9F9658 , 32'h0E1B49C0 , 32'hF7A9C7A0 , 32'h13F28720 , 32'h059FD1F8 , 32'hF57C9BE0 , 32'h169B01C0 , 32'hF99DC0E8 , 32'h07334140 , 32'h0FCB6A50 , 32'hF8238B08 , 32'hF5729960 , 32'h16AC5560 , 32'hFFB9900E , 32'hF2A349F0 , 32'h105E1F80 , 32'hFD84BEF4 , 32'hEDA98D00 , 32'hF8258E38 , 32'h0498DFE8 , 32'h011056B0 , 32'h1346BBE0 , 32'hE9993D40 , 32'hFD551C14 , 32'h090E8D50 , 32'hFEC125C4 , 32'hEEF79E40 , 32'hF77CCA00 , 32'hFBF15F30} , 
{32'hE5B8F3E0 , 32'hBFCBB180 , 32'hB23A4C00 , 32'hDA89A840 , 32'h0118CAD4 , 32'hF02A2060 , 32'h2CD27800 , 32'hF61E3350 , 32'hFC732FF8 , 32'h1541F4C0 , 32'h12AD4B60 , 32'h12E6A580 , 32'h1603A500 , 32'hF0E9DDF0 , 32'hFE9563A4 , 32'h1CD1E320 , 32'h12DAFCE0 , 32'hF2E572C0 , 32'h0BC3DAB0 , 32'h02C62850 , 32'hF8F4BCD0 , 32'h00BC9F38 , 32'hFEA942FC , 32'h046AA6A8 , 32'h0A556290 , 32'hE9FE2560 , 32'hF2512F10 , 32'h011FD814 , 32'hFBD3B6D0 , 32'h232C5240 , 32'hF4959460 , 32'h15919320 , 32'h0065B08A , 32'h10CF1140 , 32'hFCB292CC , 32'hF2E0DAE0 , 32'h05F61E28} , 
{32'hFFCA1DA7 , 32'hD2C18C80 , 32'hE17EA5E0 , 32'hD4CFE900 , 32'h1EEA32A0 , 32'hFBF2A9F8 , 32'h201410C0 , 32'h0AFCA640 , 32'hFA9F9408 , 32'hFB9F4CD0 , 32'h027A7848 , 32'h29A79600 , 32'hFF5B8C0F , 32'h0B5EE960 , 32'hDE5C3F40 , 32'h379AE840 , 32'h14D30FC0 , 32'hFB74C300 , 32'h1863E2C0 , 32'h0055B7AF , 32'hF0F58C10 , 32'h1CA37260 , 32'hFA71F828 , 32'h150D8700 , 32'hF8507170 , 32'h00275B7A , 32'hFE07AD50 , 32'h1139E920 , 32'hF6E1A680 , 32'h077067C0 , 32'hFF871B52 , 32'hF4C419B0 , 32'hEF4B7C20 , 32'hF49162D0 , 32'hFACDC838 , 32'h0FE4A700 , 32'h06FFDE88} , 
{32'h0B09DAC0 , 32'hDA137080 , 32'h11046340 , 32'h0B2BC5E0 , 32'h130BB4C0 , 32'hFDAD06F8 , 32'h0390D3DC , 32'h0508BC58 , 32'hF93BF840 , 32'h0EAA3090 , 32'h06056548 , 32'h30499F00 , 32'hF1BD44E0 , 32'h16D909A0 , 32'hE9842460 , 32'h0E59C060 , 32'h06D01728 , 32'hE944D340 , 32'h28ECB940 , 32'h0D0A4C10 , 32'hFF795FF6 , 32'hF4AEDE20 , 32'h00A96FCC , 32'hFFB0911F , 32'h179EA780 , 32'h01DCBBE8 , 32'h140AF2E0 , 32'h02A6ABD8 , 32'hDD2AE380 , 32'hE7F55560 , 32'hF09219C0 , 32'h02D17044 , 32'h06B74B20 , 32'hEFB451C0 , 32'h0FA7A290 , 32'hF5898E20 , 32'h068E98D0} , 
{32'hF940F6B8 , 32'hDC609980 , 32'hF8D4E928 , 32'h29C91980 , 32'h17FE0460 , 32'h0C9755B0 , 32'hF302C670 , 32'hF92884B0 , 32'h0277DDB8 , 32'h07C3FB10 , 32'h05C5F000 , 32'h14220400 , 32'hF7529FC0 , 32'hFEB18350 , 32'h00B33993 , 32'h111877E0 , 32'hF8A71BC8 , 32'h0BF5C5F0 , 32'h179461E0 , 32'h0E8877B0 , 32'hF44E7CE0 , 32'h0B88DAE0 , 32'hF20E3460 , 32'h040F52A0 , 32'h017DC514 , 32'hE6ED6240 , 32'h046A5550 , 32'h036FDC14 , 32'hE5D78D00 , 32'h0ABF04C0 , 32'hE5B0D240 , 32'h04309C18 , 32'hEF296560 , 32'hFDEC28F0 , 32'hEA6FDD40 , 32'hEBB4BAC0 , 32'hFE977F00} , 
{32'hF24E6FD0 , 32'h004E26DF , 32'h0090E684 , 32'h27793EC0 , 32'h11075E00 , 32'h0D444C50 , 32'hE3869C60 , 32'hF51652B0 , 32'hF48A02B0 , 32'h0B6E96E0 , 32'h07F9D280 , 32'h06DC4B70 , 32'h11761AA0 , 32'h0308E100 , 32'hE6DA1E40 , 32'h04C82328 , 32'h0818F3D0 , 32'h036B0944 , 32'h02C3BE2C , 32'hF609A0D0 , 32'hF1595350 , 32'hF6F86620 , 32'hE06F18A0 , 32'h01C0FF9C , 32'h044109E8 , 32'hF6648160 , 32'hF2AB6F80 , 32'hEC9D7520 , 32'h0A83C780 , 32'hFC29BADC , 32'hF5C49420 , 32'hFC1B90F8 , 32'hEFC14A60 , 32'h08D2C1D0 , 32'hEE2F8AE0 , 32'h071D9950 , 32'h10E5FB20} , 
{32'hF116E450 , 32'hE45A9FC0 , 32'h0973CA60 , 32'h2B3F37C0 , 32'h099C4020 , 32'h04A2D3A8 , 32'hE5FEA5A0 , 32'hF076DFF0 , 32'h03590888 , 32'h09752590 , 32'h14BEDB20 , 32'h13F55340 , 32'h11A50D60 , 32'hF883FB58 , 32'h01C57A7C , 32'hFDFB8280 , 32'h0CB821E0 , 32'h1380F8A0 , 32'h15209080 , 32'h08CEFCD0 , 32'h0C4CFE70 , 32'hFEF3436C , 32'hEE171E80 , 32'hF6BB5640 , 32'hFA599A68 , 32'hF58ECD50 , 32'hF255B090 , 32'hF5661920 , 32'h114F6BE0 , 32'hFF9E24C8 , 32'hFA504830 , 32'hFDFB604C , 32'hFADE9DC8 , 32'hF7F64E80 , 32'hE92749E0 , 32'h17A237E0 , 32'h03A20EF4} , 
{32'h0ACF8E40 , 32'hF7478130 , 32'h0CFB7630 , 32'h0A0BE1A0 , 32'h163E0CE0 , 32'hFB81FDC8 , 32'hEBA42EE0 , 32'h05670F38 , 32'h11C208C0 , 32'h0E6A5B40 , 32'h0C76AF60 , 32'hFB6E2950 , 32'h1CCA82A0 , 32'h10E35900 , 32'hFC708BD8 , 32'hE57C35E0 , 32'h10EAB9C0 , 32'hE83DF220 , 32'h0A3CF980 , 32'hFFC4D9C2 , 32'hF7005CF0 , 32'hF5FA4C90 , 32'h0D389B70 , 32'h0059ACF6 , 32'hEA517DE0 , 32'hFED94F9C , 32'hF80D9488 , 32'hF4FB1C00 , 32'h14C81620 , 32'hEA6E6E40 , 32'h03E01314 , 32'h057C2908 , 32'h1808E880 , 32'hFD399654 , 32'hF05F5650 , 32'hFD936D8C , 32'hE95A98E0} , 
{32'h020694F8 , 32'h0EE966A0 , 32'h035ED960 , 32'hFE5CB514 , 32'h12E6F8A0 , 32'h0329427C , 32'hFCFD7218 , 32'h0AC8F590 , 32'h099F33A0 , 32'hF5F3E830 , 32'h050359E0 , 32'hF020CA00 , 32'hFFCA0288 , 32'hFBCEA610 , 32'hF7640B50 , 32'hFDD44308 , 32'h17685AE0 , 32'h07AF1860 , 32'hF4505040 , 32'hF54CAAF0 , 32'hF97870A8 , 32'h00F91580 , 32'hF5C86E70 , 32'hF00C0790 , 32'hFF80214E , 32'h0E2376C0 , 32'hF75DBF30 , 32'hFB48E408 , 32'h02FFBE8C , 32'hFF4C831B , 32'h05D27D58 , 32'h08265560 , 32'hF8CA9048 , 32'hFF1F441D , 32'hEE643A40 , 32'hEEA65340 , 32'hF8421CD0} , 
{32'hF5748CD0 , 32'h08EAA2B0 , 32'hF1778920 , 32'hE8502EC0 , 32'h06BFF540 , 32'h0C421ED0 , 32'h05D9B080 , 32'h20E69940 , 32'h118509E0 , 32'hF7B67C00 , 32'h118D6C80 , 32'hDE5B3AC0 , 32'hF5A320E0 , 32'h05A871E0 , 32'h089E9960 , 32'hF3FEDD90 , 32'h20826A00 , 32'hFC1CF840 , 32'hFA67B678 , 32'hE25E0360 , 32'hE45276E0 , 32'hFBF7DAB8 , 32'h0E6D6450 , 32'hF3273A80 , 32'hF776D260 , 32'h12259B00 , 32'hEF91E3C0 , 32'h11F06440 , 32'h09092400 , 32'h0A194F40 , 32'hDF73A680 , 32'h0F5E68A0 , 32'hF089E410 , 32'hEDF3E5A0 , 32'hE8746A80 , 32'hEC0CEC40 , 32'hE9F7CC80} , 
{32'hFEAB93CC , 32'h07B32D50 , 32'hF5847A30 , 32'hFC72C8EC , 32'h0550D7C0 , 32'h07C3DCC8 , 32'h0F3FF290 , 32'h0F217950 , 32'h0025311E , 32'hF69F3BD0 , 32'h0726E5F0 , 32'hF28541D0 , 32'hFADFB150 , 32'h03905248 , 32'h02CEFEBC , 32'h0233CCB4 , 32'h0F9C6A10 , 32'h0BD01B70 , 32'hFC219570 , 32'hFC7F1CEC , 32'hFC4C7034 , 32'h02F90A2C , 32'hFC9338EC , 32'hFB7DC3A0 , 32'h04F944B8 , 32'hF755A6F0 , 32'h0199F0F0 , 32'h08006A10 , 32'h018E5238 , 32'h0ADA48C0 , 32'hECCDC920 , 32'h057765E0 , 32'hFE0052D0 , 32'h015912AC , 32'hFC53D0A0 , 32'hF960C2B8 , 32'hFF6B099B} , 
{32'h03944CA8 , 32'h19CEDD20 , 32'hEF10EC80 , 32'hF8996AE0 , 32'hFB3E54F8 , 32'h1B9ED2C0 , 32'h145E37E0 , 32'h2C365580 , 32'h15736E80 , 32'hD6DBC980 , 32'h16AD7960 , 32'hF91AE258 , 32'hF4953560 , 32'hF7FA9730 , 32'h27905D00 , 32'h113157C0 , 32'h1A3E5920 , 32'h15684540 , 32'h077806C0 , 32'h16C67040 , 32'hFDFFAB28 , 32'h0B8710F0 , 32'h101C9FE0 , 32'hEC6DB880 , 32'h061C3450 , 32'hFA06A8C8 , 32'h0C636760 , 32'hFD74B4C8 , 32'hF67E4E60 , 32'hFE4F0CDC , 32'hF5756C10 , 32'h011D0314 , 32'hF69849B0 , 32'h1AF79F60 , 32'h0C888420 , 32'h071C2258 , 32'h0904E160} , 
{32'hF4ED99F0 , 32'h04B8A970 , 32'hFCB16AC0 , 32'hFF79DC30 , 32'h04F3A038 , 32'hF8ECE208 , 32'h0A6B6310 , 32'h0581CF10 , 32'h0A5FFE80 , 32'hF7F3C560 , 32'hF273C850 , 32'h028EB1CC , 32'h0C7C4330 , 32'h00FE5524 , 32'h0A504640 , 32'h0C42ABD0 , 32'hFE7216D4 , 32'h05112BB0 , 32'h08317C80 , 32'hF28A4C20 , 32'h0524BC58 , 32'h02604B94 , 32'hFA7F0938 , 32'hFC461620 , 32'h04D397C8 , 32'h04B51FB0 , 32'h02732AC0 , 32'hF422FB50 , 32'hF84C46C0 , 32'h06518A98 , 32'hF3872B30 , 32'h03824378 , 32'h10EC4780 , 32'h06062890 , 32'h03727B40 , 32'hF6B76DD0 , 32'hFE1644B4} , 
{32'hFDB97FB4 , 32'hF9F66838 , 32'hFC5AE864 , 32'h046E4B50 , 32'hFC26E998 , 32'hFE06D7BC , 32'h007EC3C9 , 32'h05E46BE8 , 32'h08071470 , 32'hFC77E578 , 32'h052C8B68 , 32'h0AB7CE80 , 32'hFBA888C0 , 32'h01A72758 , 32'hFF33C7F7 , 32'hF6BFA120 , 32'hFE2FAA18 , 32'h098B1F50 , 32'hF70728F0 , 32'hF4F3BF60 , 32'hFB00ADC0 , 32'h0056322E , 32'h036E40E0 , 32'h08D7EBE0 , 32'hFF2290BE , 32'h03523F10 , 32'h0DF152B0 , 32'h0DB85DC0 , 32'h0129B0E8 , 32'h060422C0 , 32'h033DE458 , 32'hFAF8FAE0 , 32'hF49343C0 , 32'h04067188 , 32'hFB3E6658 , 32'hFE1CC0B0 , 32'hFB926620} , 
{32'h0076AB73 , 32'hFF0230E2 , 32'hFF0F8FC7 , 32'hFF879E1D , 32'hFC6B621C , 32'h01E531A8 , 32'hFD57F170 , 32'h0082F823 , 32'h007682A1 , 32'hFF9F71FC , 32'h0144B594 , 32'h035B0C0C , 32'hFEF3ED54 , 32'h0194A534 , 32'hFDE6F1BC , 32'h00270395 , 32'hFFDDC03A , 32'h01AD9368 , 32'hFF968584 , 32'hFEE9B5E4 , 32'hFE88D4A4 , 32'hFD671890 , 32'h00E0D37A , 32'h004C3C5A , 32'h01256560 , 32'hFC7BD744 , 32'h0106C370 , 32'h00E48D4D , 32'hFE2FE9B4 , 32'h03399394 , 32'h0379EC14 , 32'h023CFA90 , 32'hFCF4075C , 32'hFEB6AE08 , 32'hFFC403CA , 32'h00B83555 , 32'h02199764} , 
{32'h000261EE , 32'h000262E4 , 32'hFFFC2E64 , 32'hFFFE0266 , 32'h00006F2F , 32'h0002A884 , 32'hFFFDD9EA , 32'h000129B1 , 32'hFFFF0C86 , 32'h00033EAC , 32'hFFFCFB64 , 32'hFFFDF9A6 , 32'hFFFBF78B , 32'hFFFE53E3 , 32'hFFFFA958 , 32'h0001C474 , 32'hFFFE13D0 , 32'hFFFBF36D , 32'hFFFDD3F1 , 32'h00036FFB , 32'h00029653 , 32'h00004A82 , 32'h00036F1B , 32'h0001DF13 , 32'hFFFD6E6C , 32'hFFFFEA6B , 32'h00044BCE , 32'h0002C5BD , 32'h00012F3B , 32'h00010D01 , 32'h0002FE0D , 32'h00023447 , 32'h00038EAC , 32'hFFFADE2F , 32'hFFFD1621 , 32'h00041C22 , 32'h0003F815} , 
{32'hFFFF4635 , 32'h0006C26C , 32'h00013E64 , 32'h000421EC , 32'hFFFC6F83 , 32'hFFFAFFA8 , 32'hFFFF7679 , 32'hFFFF6710 , 32'hFFFFDA9D , 32'hFFFF1E7A , 32'h000860B5 , 32'h000138E5 , 32'hFFFBA02C , 32'hFFFFC68C , 32'h0006DC30 , 32'h00001019 , 32'h0002E61F , 32'hFFFC52D7 , 32'h00064AE4 , 32'hFFFF0C14 , 32'h0002BC0D , 32'h00077D01 , 32'hFFFC6AEB , 32'h0006280A , 32'h00034CD0 , 32'h0008AFA1 , 32'hFFF86D36 , 32'hFFFA816F , 32'h0000385D , 32'h000078D9 , 32'h00031514 , 32'h00049DE7 , 32'h00040B29 , 32'h0003C5D5 , 32'h00053CAB , 32'hFFF8A9E8 , 32'h000023EF} , 
{32'h00023943 , 32'h0000A42F , 32'hFFFEC18D , 32'h0002191F , 32'h00013D8D , 32'hFFFCF6E8 , 32'h0003C974 , 32'hFFFBFE64 , 32'h0001FEB3 , 32'h00047141 , 32'hFFFB3305 , 32'hFFFC1AFC , 32'hFFFFAC00 , 32'hFFFDD185 , 32'h000479C6 , 32'h0005C295 , 32'h000380AE , 32'hFFF8F123 , 32'hFFF4A1E3 , 32'h00001A8F , 32'h000259B3 , 32'h00007E94 , 32'h0006511C , 32'h0008BD85 , 32'hFFFC9F95 , 32'h00051E7A , 32'h0000C616 , 32'hFFFEE4A1 , 32'h0000EF23 , 32'hFFFCBD85 , 32'h000453B9 , 32'h000418BB , 32'h0003C973 , 32'hFFFD7FE6 , 32'h0002847C , 32'hFFF7E9CD , 32'h0004B7E7} , 
{32'hFFFF1CD8 , 32'hFFFE407B , 32'hFFFB871F , 32'hFFFD782F , 32'h000116DE , 32'hFFFC482F , 32'h00084D4B , 32'h000786CB , 32'hFFFFCAD6 , 32'h0001BA8F , 32'h0004D2F2 , 32'h000A24D0 , 32'h0000FE3D , 32'hFFFEB72D , 32'h0002E43C , 32'hFFFF41DA , 32'hFFFE6BAC , 32'h0001F484 , 32'hFFFD95D6 , 32'h0000D502 , 32'hFFFFFB08 , 32'h0002FE68 , 32'h0005708E , 32'h00027E78 , 32'h00043BA1 , 32'hFFFFC550 , 32'h00009906 , 32'h000034A6 , 32'h0004B4BC , 32'h00046FF5 , 32'h00066DBD , 32'h000059F1 , 32'hFFFEF768 , 32'h00025673 , 32'hFFFC950D , 32'hFFFDB220 , 32'h0000CB6B} , 
{32'h00037FC6 , 32'h0001DB7F , 32'hFFFE3F9E , 32'h000339F7 , 32'h000566FB , 32'hFFFF64B6 , 32'h00011192 , 32'hFFFDF1B7 , 32'hFFFFE7D3 , 32'h0002E23A , 32'hFFFB2A8F , 32'h000702F8 , 32'hFFF99EAB , 32'hFFFF972F , 32'hFFFA5B88 , 32'hFFFC1689 , 32'h00038468 , 32'h00014A67 , 32'h00001E5B , 32'h0005BAF1 , 32'h0006D5FF , 32'hFFFF8CEE , 32'h0001D073 , 32'hFFFD3144 , 32'hFFFB109A , 32'h00018CA5 , 32'hFFFDA9BC , 32'hFFFB0130 , 32'h000090D9 , 32'hFFFEFC33 , 32'h0000AA0B , 32'h0001AE16 , 32'hFFFA984A , 32'hFFFF2D81 , 32'hFFFD2EA9 , 32'hFFFCFF62 , 32'hFFFFEBF5} , 
{32'h00016077 , 32'h000014DF , 32'h00000AFF , 32'hFFF93526 , 32'h0000137D , 32'hFFF94E93 , 32'hFFFB1CB2 , 32'h000053BF , 32'hFFFFB229 , 32'hFFFE6B3A , 32'h000023F0 , 32'hFFFBCB35 , 32'h000111E7 , 32'h00006DEC , 32'hFFFEFE74 , 32'h00081425 , 32'hFFFF04D3 , 32'h00059F74 , 32'h00042133 , 32'hFFFEC612 , 32'h0003EA22 , 32'hFFFE4122 , 32'h0004673F , 32'h00018EF9 , 32'hFFFD1AD5 , 32'h00012AC6 , 32'h0000F77E , 32'hFFFF8A7D , 32'h00018D02 , 32'hFFFC93F1 , 32'hFFFF7AA9 , 32'h0000FA72 , 32'hFFFC1C9D , 32'h0002C30F , 32'hFFFEAE18 , 32'h000260A9 , 32'hFFFB4259} , 
{32'h03DEACD8 , 32'h07D4A888 , 32'hF2ADC3A0 , 32'h00CA922B , 32'h07149FC8 , 32'hF58FC970 , 32'hF34EBAD0 , 32'hF9428A68 , 32'h050C91F8 , 32'hFB121EE0 , 32'hFF6DF265 , 32'hF7CCAA30 , 32'h0210E1EC , 32'h00272E53 , 32'h0A6878D0 , 32'h03510A5C , 32'h01A92C48 , 32'h07DA6260 , 32'hFFB9E44F , 32'h05A5C070 , 32'h01F71ADC , 32'hFF11DE8C , 32'h012161EC , 32'h054F1C68 , 32'hFD2FAE78 , 32'hFB2D3AB8 , 32'hFAE2C4A0 , 32'h08567F50 , 32'hFF7F13CC , 32'h00FA8535 , 32'h02A11F64 , 32'hFE6CBA38 , 32'hF9330168 , 32'h09735220 , 32'hFFEBF75F , 32'h06CB9920 , 32'hFF453DFF} , 
{32'hFFC1971F , 32'h00025525 , 32'hFF7857AE , 32'hFFE3B75D , 32'hFF6878B2 , 32'hFFDF15F4 , 32'h0013FA3F , 32'h0021CFC5 , 32'hFFC8C365 , 32'h0022AAD3 , 32'h00466822 , 32'hFFA16B35 , 32'h00537A5E , 32'h0000F35B , 32'hFFBEFA77 , 32'h000926AC , 32'h00351D65 , 32'hFF6848EA , 32'hFFB2EADE , 32'h0028A307 , 32'h001A5844 , 32'h002FB2B0 , 32'hFFEDC543 , 32'h0081CF13 , 32'hFF6BF56D , 32'hFFC8426E , 32'hFFD6443F , 32'h00016AAA , 32'hFF8D787B , 32'hFFDB49C6 , 32'hFFD0F186 , 32'hFFC2DF30 , 32'hFFE2F936 , 32'hFFE380C6 , 32'h005547ED , 32'hFFC572D1 , 32'h00A26302} , 
{32'h05A6AC28 , 32'h0291B678 , 32'hEC4A4200 , 32'h0C234300 , 32'h025658B8 , 32'hF2F2B620 , 32'hFA65F180 , 32'h0E4EF960 , 32'h0B2B8240 , 32'h000CA441 , 32'hEF2EFF20 , 32'hF2497610 , 32'hF6572E60 , 32'hFCAA177C , 32'hFAD8A558 , 32'h09EB77F0 , 32'hFE59B404 , 32'h0E410980 , 32'h05A837D0 , 32'h09E553C0 , 32'hF0A9B0F0 , 32'h04BBF7F8 , 32'hF0F293D0 , 32'h11BC6160 , 32'hFC0DDB04 , 32'hFCB09D04 , 32'hFCFCABEC , 32'h099636B0 , 32'h0333B2A0 , 32'h01E0C058 , 32'h0A8A28D0 , 32'hFC92B180 , 32'hF5D7DDB0 , 32'h063066C8 , 32'h040F0C00 , 32'h047F9B38 , 32'h0C4306D0} , 
{32'hFC06DEB0 , 32'hFAD21FA8 , 32'hF8E3FEC0 , 32'h0106B4E8 , 32'h0A04F7A0 , 32'hFFA3CC3F , 32'hF8F0E6A0 , 32'hFFD42187 , 32'hFDCDD398 , 32'hFD92AB50 , 32'h0156BCB0 , 32'hF9C2EFA8 , 32'hFE860FC4 , 32'h038EF87C , 32'h09FD5490 , 32'hF70D6220 , 32'hFAD6BE60 , 32'hF98AD9D8 , 32'hFE71DDF0 , 32'h05D3EB58 , 32'hFC3F95C0 , 32'hFA7E7CF0 , 32'h025128F4 , 32'hFE6872DC , 32'h02A18D30 , 32'h0648BB70 , 32'h04F98380 , 32'hF80C0C10 , 32'hFE7059B8 , 32'hFCA95EE8 , 32'h06F0C630 , 32'hFD01A5C8 , 32'h01147EB0 , 32'hF89A4300 , 32'h0936B6A0 , 32'hFD469E04 , 32'h03420D18} , 
{32'h035E5D80 , 32'h01714814 , 32'hD70A7FC0 , 32'hF8108228 , 32'h17F51280 , 32'hF387E150 , 32'hDC471740 , 32'hFF0F3F28 , 32'hFA172CB0 , 32'hF22C2600 , 32'hF75921D0 , 32'hEE48FAE0 , 32'h032ABE04 , 32'h057E59E0 , 32'h146BE0E0 , 32'hF27C0670 , 32'hFB4E6960 , 32'h0B532F80 , 32'hFEF6FEC8 , 32'h0AEC6EB0 , 32'hFEB5D224 , 32'hEEFD7220 , 32'hFF468FD1 , 32'hFCC7DC08 , 32'h0FC536E0 , 32'h08815110 , 32'h13466780 , 32'hFA7BCC18 , 32'hFEDC3E64 , 32'hF99648C8 , 32'h01DFCE98 , 32'hFC75C328 , 32'h04B10D08 , 32'hFFEE82CE , 32'h0DAF6BA0 , 32'hFFFAAD2D , 32'h0D66F5C0} , 
{32'h08A3E640 , 32'hFE98EFDC , 32'hC054B340 , 32'hE8093C20 , 32'h2C368680 , 32'hE142F860 , 32'hEAF39AE0 , 32'hFB699BD0 , 32'hF6F06DD0 , 32'hE79E3A40 , 32'h05BFE718 , 32'hE24EF280 , 32'h13A7E980 , 32'hEB9D79C0 , 32'h1E76DC80 , 32'hE4D75060 , 32'hE371B9A0 , 32'h14A86FC0 , 32'hF94F2410 , 32'hF67872F0 , 32'h0166BA20 , 32'hFC62F158 , 32'hFD9EFEF0 , 32'hEF28AF40 , 32'h16639220 , 32'hF070E070 , 32'h0DCBDFA0 , 32'hEC4DC260 , 32'hF09D4B70 , 32'hF0B38720 , 32'hFCA0AB88 , 32'h08758720 , 32'hF2C51070 , 32'hEF544160 , 32'h0F38BCC0 , 32'h03048F98 , 32'h0B332FE0} , 
{32'hF74F0F20 , 32'hF7748560 , 32'hB2249880 , 32'hEE3E0B60 , 32'h21F9A0C0 , 32'hD6677140 , 32'hE66A25E0 , 32'hF84B1EA0 , 32'h00D98A66 , 32'hED5F5200 , 32'h0F53C5F0 , 32'hEE750EA0 , 32'h02A62AD8 , 32'hFE551348 , 32'h0C6A2C80 , 32'hEEB9B6E0 , 32'hF563CEA0 , 32'h01D7256C , 32'hF61BA2C0 , 32'h135154A0 , 32'h03E0B630 , 32'hE71CADA0 , 32'h0813FC20 , 32'hF6D72850 , 32'h1CB11D80 , 32'h08E9C2A0 , 32'hFEAB87F0 , 32'hF0B2B540 , 32'h0EC325E0 , 32'hEF691820 , 32'h0613FD28 , 32'hFDBAFC18 , 32'hFB6A5570 , 32'h05E9A2D0 , 32'h136FB780 , 32'hF18F1560 , 32'h0B503B20} , 
{32'hE2AC9D60 , 32'hF01E9250 , 32'h80000800 , 32'hE310EFC0 , 32'h2CC2AEC0 , 32'hCF35B980 , 32'hF4BA56A0 , 32'h0415AB28 , 32'h0CE60BC0 , 32'hF59F6440 , 32'h30A23940 , 32'h0DCE0820 , 32'hF424BD90 , 32'h0ECD8C30 , 32'hF841FDF8 , 32'hF9625810 , 32'hEF0F9380 , 32'hE7D69F80 , 32'hF2AB37D0 , 32'h273CC940 , 32'h02D49408 , 32'hF39CB8C0 , 32'hFD9F1EE8 , 32'hEF5F2BA0 , 32'h14AF0BE0 , 32'h0969B5A0 , 32'h0EBE6D20 , 32'hD8F41100 , 32'h104BE660 , 32'hF6E159C0 , 32'h05842450 , 32'h0A55F010 , 32'h037B3300 , 32'hDCC9E900 , 32'hF94902A0 , 32'hF374B4B0 , 32'hF5C17700} , 
{32'hFBA7D2F0 , 32'hF21ED830 , 32'h9C108500 , 32'hE198AEC0 , 32'h18409440 , 32'hD40349C0 , 32'hF49E5EA0 , 32'h0C20ED60 , 32'h1F16AA80 , 32'hF9650830 , 32'h2792B700 , 32'h260F1040 , 32'hF8E307E0 , 32'h010270FC , 32'hF9632BF0 , 32'h07B75FA8 , 32'hFB3B9E40 , 32'hE46149A0 , 32'hF3F7D360 , 32'h09C0D7C0 , 32'h181B9FA0 , 32'h0A2CD5A0 , 32'hFFBAF345 , 32'h0598C5B8 , 32'h022A1998 , 32'h131D87E0 , 32'h068ACFA8 , 32'h06356EE0 , 32'h0DA36A40 , 32'h09237E50 , 32'h001A37D8 , 32'h060D1348 , 32'h0CAD2470 , 32'h0293AE04 , 32'hFF2B5106 , 32'h0215ED28 , 32'hF724FD10} , 
{32'hFFCD5067 , 32'h050F1EB8 , 32'hE6DEE400 , 32'hF1942AF0 , 32'h27928EC0 , 32'hF63C9030 , 32'h091793B0 , 32'hE3FAF480 , 32'hFDEA9A90 , 32'hF111A380 , 32'h2A94C880 , 32'h1A27E500 , 32'h0321AF18 , 32'h06867E58 , 32'hFDF7351C , 32'h160ABBA0 , 32'h05EB8998 , 32'hEEEA22A0 , 32'hF9A8E6C0 , 32'hF90AEEF8 , 32'h1E0CCA20 , 32'h24CEF600 , 32'h0426B6C8 , 32'h0E0D2B70 , 32'hF8C4DAD8 , 32'hE7358280 , 32'h020E6D68 , 32'h0F765D70 , 32'hFC012DEC , 32'h11EBCD20 , 32'hF99E3838 , 32'h0990C6A0 , 32'h01A15DDC , 32'hFCE5D780 , 32'hEDDA7620 , 32'h04E322C8 , 32'h04C67FB8} , 
{32'hF7FF6C80 , 32'hF4349A30 , 32'hF7DCC8C0 , 32'h02B9B51C , 32'h1DBA2BE0 , 32'h0227FFB0 , 32'hFB298F08 , 32'hFDA50534 , 32'h09F577F0 , 32'hFBC3FDC8 , 32'hF7756610 , 32'h1F6A0500 , 32'hEB4C0660 , 32'h162CE160 , 32'hEE091140 , 32'h18051AE0 , 32'hFAD5E2E8 , 32'hED2609E0 , 32'h133D5B40 , 32'h07C77260 , 32'hFBE28C90 , 32'h0943DF90 , 32'h053E6710 , 32'h0E9FF2F0 , 32'hEECA4560 , 32'hE8C28C40 , 32'hFBB55210 , 32'h0B963A80 , 32'hE8EDF540 , 32'h01468680 , 32'hF35F8E10 , 32'h112DBE20 , 32'hF8231878 , 32'hFB49C770 , 32'hEA3ED5E0 , 32'hF5722180 , 32'hFC68E744} , 
{32'hF0C44C70 , 32'hE6EF93A0 , 32'hF0FFF110 , 32'h2DB4F100 , 32'h2A7A0D00 , 32'h127652E0 , 32'hEF9CC840 , 32'hFD1BBAE0 , 32'hFD054484 , 32'h0A919060 , 32'h0DBA0750 , 32'h2EDBE8C0 , 32'h010275CC , 32'hFA1C1908 , 32'hE744F5A0 , 32'h0964B2F0 , 32'hFD153364 , 32'h203A2140 , 32'hF56289F0 , 32'h09E04A90 , 32'hFE4290A4 , 32'h02FDF6DC , 32'hD8518680 , 32'h030C6B20 , 32'hF90E16B8 , 32'hF565E3B0 , 32'h105630A0 , 32'hEA136320 , 32'hE5FB40C0 , 32'hF33F81A0 , 32'h0BAA9B90 , 32'hEAB9D520 , 32'hFED6DC90 , 32'h0D7D8FC0 , 32'hF5AD2CB0 , 32'hEA5B2FE0 , 32'h15CE31E0} , 
{32'hE9107860 , 32'hE9DA1E20 , 32'h020FDA70 , 32'h41161E80 , 32'h149103A0 , 32'h09165E10 , 32'hE1157F80 , 32'hEA3F2400 , 32'hFBEBE040 , 32'h01523B4C , 32'h140328E0 , 32'h12850EC0 , 32'h03CBCF2C , 32'hFB605AC8 , 32'hE0B1B3C0 , 32'h02620DAC , 32'h220C3900 , 32'h426B5600 , 32'hFE1F1F68 , 32'h0D2172E0 , 32'hEE0CC940 , 32'h12E82900 , 32'hD4EC6A80 , 32'hF2F08C10 , 32'hF4E4F290 , 32'h0ADBAAB0 , 32'hF843D788 , 32'hE67C2520 , 32'hF2D1AF50 , 32'hF85EA688 , 32'hFD718EE4 , 32'hFE360BEC , 32'hF752D950 , 32'hFEFAD2EC , 32'h0298CCBC , 32'hE8840520 , 32'hFDCC5C5C} , 
{32'hFC77DBA8 , 32'h08897FE0 , 32'h05E082E8 , 32'h0D577130 , 32'hFFE75CBF , 32'hFAB42DE0 , 32'hFD043BAC , 32'h014525F8 , 32'h061AA7E0 , 32'hFD6A8374 , 32'h0DFEC670 , 32'h0153F248 , 32'hF3DA2E70 , 32'h154DEF40 , 32'h0498E648 , 32'hED9C4D20 , 32'h03D1F5CC , 32'h12749740 , 32'h16AEB640 , 32'hF30BC2E0 , 32'h093C4380 , 32'hF250DFB0 , 32'hF02BD4A0 , 32'hFC7C1BDC , 32'hE312DA00 , 32'hF9DA6E70 , 32'hFBD01B08 , 32'hF1D94A90 , 32'hF701E3F0 , 32'hFC87D124 , 32'h048380A8 , 32'h0FEBD6A0 , 32'hFF6F4F7B , 32'h01CD6E64 , 32'h0542B8F8 , 32'hF63B02B0 , 32'hFC1602C0} , 
{32'hFF92BF89 , 32'hF9E25BF8 , 32'hF68EE600 , 32'hFCCBC4BC , 32'h0AA7C140 , 32'hF9989B20 , 32'h00D51CBC , 32'h085F2D60 , 32'h0E599C70 , 32'h09593A30 , 32'h144A2E40 , 32'h0244A57C , 32'hFB350178 , 32'h01515360 , 32'hFC5E182C , 32'hDEA82140 , 32'h0CDD6CC0 , 32'h0DE2D5E0 , 32'hED3E2B40 , 32'hEE65BE00 , 32'h043C9B08 , 32'hE1E26800 , 32'hE8055060 , 32'h18425BA0 , 32'hEF6DF2A0 , 32'hFDD625BC , 32'h09325F70 , 32'hFE736C84 , 32'h17E0A280 , 32'h08C18310 , 32'h0D3375D0 , 32'h0C42A9A0 , 32'hFFF90740 , 32'hF37B16A0 , 32'hF67C7D50 , 32'h052CD310 , 32'h03333370} , 
{32'hFFF29C15 , 32'h064A99A0 , 32'hF3424E60 , 32'hF653A940 , 32'h052F1378 , 32'h04D40078 , 32'h06D45598 , 32'h111BE160 , 32'h0B5F5DD0 , 32'hFBC3F228 , 32'h14466D60 , 32'hF5523440 , 32'hFD5CEC74 , 32'h03968884 , 32'hFC4A1D44 , 32'hF7109A90 , 32'h0F88DA10 , 32'h01988E40 , 32'h053A8B78 , 32'hF52D58D0 , 32'h033D3A68 , 32'hFF8E84D8 , 32'hFCFDDCDC , 32'hFE1D1908 , 32'hF8FBB288 , 32'h020A4FF4 , 32'hF9DF1890 , 32'h0162F188 , 32'h0DF175B0 , 32'h0B3084D0 , 32'hFCF93CF8 , 32'h081EA490 , 32'h02D80488 , 32'hF04E3E40 , 32'hF1C74760 , 32'h01CBA014 , 32'hFCE95A40} , 
{32'hFF0EA768 , 32'h07C74248 , 32'hFB8FD990 , 32'h01903758 , 32'hFD539BE4 , 32'h038E8314 , 32'h04B8BD48 , 32'h04E0CC60 , 32'h05840C30 , 32'h00223395 , 32'h089EB650 , 32'h05311F50 , 32'hF9E30060 , 32'hFFB6C341 , 32'h0032C9D7 , 32'h090D0970 , 32'h0B1B7680 , 32'hFCAF4980 , 32'hFFEB49BB , 32'h024CEA2C , 32'hFEF5F320 , 32'h070A6BF8 , 32'h01512318 , 32'h04A30950 , 32'hFF7A6B6F , 32'hF7674550 , 32'hFDAE0E40 , 32'hFF5E0040 , 32'hFE5CE124 , 32'hFD527618 , 32'h05039888 , 32'hFD38C200 , 32'h0B451DB0 , 32'hFA561C08 , 32'hFDE6C4E0 , 32'h08AB21B0 , 32'hFEFC7A74} , 
{32'h0968DAA0 , 32'h110869E0 , 32'hFD448FB0 , 32'h023DD880 , 32'h0AE412D0 , 32'h0A2CD5F0 , 32'h16707640 , 32'h099D7520 , 32'h0565C700 , 32'hF6A592C0 , 32'h02386AA4 , 32'h0ADAC0F0 , 32'hF7D302E0 , 32'hFA780CF0 , 32'h0B4F8700 , 32'hFCCAA740 , 32'h022753E8 , 32'h02CB5C78 , 32'hFA8CA628 , 32'h07AE71B0 , 32'hFD71E818 , 32'h04063010 , 32'h01FCA10C , 32'hF5E751E0 , 32'h0655ED18 , 32'hFD21E804 , 32'h03285114 , 32'h057C23D0 , 32'hFEF2C1E4 , 32'h00FDAF90 , 32'hF14AF020 , 32'h0C46F5D0 , 32'hF2604EF0 , 32'h08356DB0 , 32'h0450E120 , 32'h078630F0 , 32'h16466280} , 
{32'hF988A918 , 32'h11626640 , 32'hF54C7A90 , 32'hFA3715D8 , 32'hF6AA1070 , 32'h13A87F20 , 32'h11A05660 , 32'h0C750720 , 32'h0349A764 , 32'hF0D6C110 , 32'h142139C0 , 32'h0A330700 , 32'hF98F1098 , 32'h04A438A0 , 32'h1790C440 , 32'h05A24C38 , 32'h15F4B640 , 32'h12F6A7C0 , 32'h02506204 , 32'h19167BA0 , 32'h006A0B35 , 32'hFA013EB8 , 32'h03AB96AC , 32'h068A0508 , 32'h06AB59B8 , 32'hF71B52B0 , 32'h1327A600 , 32'hFD1CA914 , 32'hECB70B20 , 32'hF9BBC5B0 , 32'h047C4D98 , 32'h0D48B2F0 , 32'hFF1F7BBB , 32'hFE2F7524 , 32'hFCAE3CAC , 32'h03F4A24C , 32'h11D66A20} , 
{32'hFC44553C , 32'h11C0A000 , 32'h07145268 , 32'hFBF45A30 , 32'h05B3BC30 , 32'hFF34C499 , 32'hFE8DDD50 , 32'h0F19C590 , 32'h05DFE190 , 32'hF507BBE0 , 32'hEF157B40 , 32'h080ED3E0 , 32'h01B2B9F4 , 32'h0106FC58 , 32'h0DDDF680 , 32'h0E4F4D00 , 32'hFCB42140 , 32'h048223D8 , 32'h05FD0DE8 , 32'hFB35B160 , 32'h0DB12CE0 , 32'h03467718 , 32'hFEBB72FC , 32'hF5CEA4E0 , 32'h0ABE21A0 , 32'h02F42EF4 , 32'hF610CFA0 , 32'hECA37C60 , 32'h0BB38DB0 , 32'h01454B50 , 32'hF774D140 , 32'h0719E708 , 32'h06418340 , 32'h017EF618 , 32'hFF32FD3E , 32'h02A862A0 , 32'hF9ADD640} , 
{32'hFA9A7EE8 , 32'h05D882C8 , 32'h0033B364 , 32'hFF00D285 , 32'hF8DEC3A8 , 32'hF374C1D0 , 32'h05ACFB60 , 32'h058D6150 , 32'hFBFCB220 , 32'hF210F430 , 32'h064889E8 , 32'h0239F928 , 32'hD9F7F500 , 32'h32E8DCC0 , 32'h0BB544A0 , 32'h08BC8990 , 32'hDD817680 , 32'h01BD6AC4 , 32'h253E55C0 , 32'hE448F460 , 32'hFD0DFFE8 , 32'hFCC098DC , 32'hE1F273A0 , 32'h0C9F7ED0 , 32'hF8A512A8 , 32'h019D4678 , 32'hF2D98E30 , 32'h00386E61 , 32'h023988D4 , 32'hFDBE2998 , 32'hF65BABD0 , 32'hECE5D100 , 32'hF027CA70 , 32'h00F106BA , 32'h0863CE10 , 32'h085672E0 , 32'h0DF50AF0} , 
{32'hFFFF9355 , 32'hFFFFDE88 , 32'hFFFF54E9 , 32'hFFFDE5BE , 32'h00004445 , 32'h0004C81A , 32'h000214BE , 32'h0001ED1B , 32'h00031B7B , 32'h0002F953 , 32'h000056E5 , 32'h0003360B , 32'h00002B0A , 32'h0000163B , 32'hFFFF57E6 , 32'h0001395F , 32'hFFFB257B , 32'hFFFFD42C , 32'h00017F95 , 32'hFFFF3EA9 , 32'h00008443 , 32'h00031852 , 32'hFFFFF524 , 32'hFFFF7174 , 32'hFFFF468B , 32'hFFFDB088 , 32'h000413E8 , 32'hFFFB11E4 , 32'hFFFC7C68 , 32'hFFFC6175 , 32'h00006C77 , 32'hFFFE63A9 , 32'h00040F28 , 32'hFFFE076F , 32'h000116B0 , 32'hFFFFA614 , 32'h000239FD} , 
{32'hFFFF2EE9 , 32'h00008421 , 32'h00034EFC , 32'h0000AE60 , 32'hFFFE3652 , 32'hFFFB1891 , 32'hFFFFB48D , 32'hFFFF85E1 , 32'h00041AED , 32'hFFFCF8B6 , 32'h0002E69F , 32'h0003530E , 32'hFFFF17FC , 32'hFFFBFBCB , 32'h00028C72 , 32'h00009F97 , 32'hFFFE4C39 , 32'h000194C4 , 32'h0002DAB7 , 32'h0000689E , 32'hFFFF92DE , 32'hFFFB2F77 , 32'h0002E5EC , 32'h00033CE9 , 32'hFFFF6570 , 32'h0002EDAC , 32'h00015165 , 32'hFFFF15CC , 32'h0000AA8D , 32'h00011120 , 32'hFFFCB3AA , 32'h0001B858 , 32'h0000AC2D , 32'hFFFF3D14 , 32'hFFFFC743 , 32'hFFFF476C , 32'hFFFF5DB3} , 
{32'h0001C33A , 32'hFFFEBA13 , 32'hFFFFAB3B , 32'h00035BB3 , 32'h0002A14B , 32'hFFFEDDF8 , 32'hFFFA28B5 , 32'h00041908 , 32'hFFFC5570 , 32'h0002B34B , 32'hFFFAB5E9 , 32'h0000BD03 , 32'hFFFAE953 , 32'hFFFA248E , 32'h0003447E , 32'h00033C06 , 32'h00030333 , 32'hFFFECECB , 32'h0004F05C , 32'h000045A0 , 32'hFFFE0468 , 32'h0000C6A0 , 32'h000019B4 , 32'h00021208 , 32'h000146F7 , 32'h00029C0D , 32'hFFFF68A1 , 32'hFFFDEFF4 , 32'h00034079 , 32'h00029C51 , 32'hFFF978AC , 32'hFFFF2ECD , 32'h00004FF3 , 32'hFFFE01BB , 32'hFFFF6CC2 , 32'h0003BA7A , 32'hFFFF31BE} , 
{32'h00018D35 , 32'hFFFFDBF6 , 32'hFFFF8D1A , 32'h00071103 , 32'h00065B8A , 32'hFFFE93B9 , 32'hFFF8B946 , 32'hFFFEC9FD , 32'hFFFF4F4F , 32'hFFFF4110 , 32'h0001270B , 32'hFFFF0E11 , 32'hFFFC770C , 32'hFFFBC2E7 , 32'hFFFF0DB8 , 32'hFFFDD762 , 32'hFFFCDBA4 , 32'h00043393 , 32'h00006018 , 32'hFFFFE96B , 32'h0002AEF9 , 32'h0004E837 , 32'hFFFD6E25 , 32'hFFF8BE98 , 32'hFFFE69E7 , 32'hFFFE1E8D , 32'h00009BD1 , 32'hFFFF3477 , 32'hFFFD7476 , 32'hFFFBA24B , 32'hFFFCCF1E , 32'hFFFDAE9F , 32'h000024F5 , 32'hFFF9F209 , 32'hFFFBF1C8 , 32'hFFFF0E51 , 32'hFFF8C85D} , 
{32'hFFFF21F0 , 32'hFFFF5503 , 32'hFFFA57F6 , 32'h0000F06A , 32'h0001D683 , 32'h0002419A , 32'h0001B305 , 32'hFFF9A4CF , 32'h0004A9FA , 32'hFFFDD798 , 32'h00040AC9 , 32'hFFFD2D4C , 32'h00027012 , 32'h00082CAB , 32'h0000290F , 32'h00006D36 , 32'hFFF9AEA0 , 32'h00001A85 , 32'hFFFB9EF3 , 32'hFFFF2D31 , 32'hFFFDB164 , 32'hFFF97517 , 32'hFFF93DB0 , 32'hFFFE11F6 , 32'h0002872F , 32'hFFFEE11F , 32'hFFF8F549 , 32'h0001F1D8 , 32'h0004788E , 32'h00002DB8 , 32'hFFF6134D , 32'hFFFEFDD6 , 32'hFFFD0A69 , 32'hFFF9ACAD , 32'hFFFFFE37 , 32'h0004175B , 32'h0003DF1D} , 
{32'h0004C115 , 32'hFFFF8A2F , 32'hFFFEC603 , 32'h00022DC0 , 32'hFFFCAE35 , 32'h0003DBE5 , 32'h000335D6 , 32'hFFFFDF5E , 32'hFFFEF9BD , 32'hFFFBA879 , 32'h0006D885 , 32'hFFFD6757 , 32'h00009D08 , 32'hFFFD1A17 , 32'h0001FF4D , 32'h0002E989 , 32'hFFFF066A , 32'hFFFF51CC , 32'h000017B0 , 32'hFFFD66C2 , 32'hFFFC86FE , 32'hFFFE8298 , 32'hFFF93EAE , 32'hFFFE70B2 , 32'h000006DF , 32'h0004411F , 32'h0004369E , 32'hFFFCB97E , 32'hFFFE9D99 , 32'h00016F2A , 32'h00034704 , 32'h000027FB , 32'hFFFE4AF4 , 32'h000289DB , 32'hFFFD4EA1 , 32'hFFFA92E9 , 32'hFFFEC710} , 
{32'h00036780 , 32'hFFFA5641 , 32'hFFFC4C64 , 32'hFFFC8354 , 32'h00039E8E , 32'hFFFD4791 , 32'h000003FE , 32'hFFF99ECC , 32'h00025CBE , 32'h00010801 , 32'h00025579 , 32'h00035BF0 , 32'h00047598 , 32'hFFFDBD66 , 32'h00044F4C , 32'h00042158 , 32'hFFFEFA9F , 32'hFFFDE91A , 32'h000189FD , 32'h000519A7 , 32'h00056CE8 , 32'hFFFD4EF5 , 32'h0000E9B2 , 32'hFFFEF56F , 32'h00043163 , 32'h0002CE7F , 32'h0002811D , 32'h0001B5CD , 32'hFFFCB9D3 , 32'hFFFCBD78 , 32'h0000657D , 32'hFFF9FD33 , 32'h0000040A , 32'hFFFE9D70 , 32'hFFFED1A0 , 32'h0000B16E , 32'h0004D953} , 
{32'h0003DACE , 32'h00008AC6 , 32'h0004CA47 , 32'hFFFF6F33 , 32'h0000562C , 32'h0002FC21 , 32'hFFFCAFC5 , 32'h0000B520 , 32'h000245F4 , 32'hFFFE20DA , 32'h0005F3CA , 32'hFFFDEC5D , 32'hFFFFF141 , 32'hFFFDA407 , 32'h00025BAF , 32'h00031B43 , 32'h00032C35 , 32'hFFFEB1C2 , 32'hFFFF776C , 32'hFFFEC006 , 32'hFFFD7157 , 32'h0001C6CC , 32'hFFFE7608 , 32'hFFFDC271 , 32'hFFFF6C4D , 32'h00014BEA , 32'hFFFA1463 , 32'hFFFE65C0 , 32'h00028E8B , 32'hFFFF24AA , 32'h00004F0E , 32'h000547EA , 32'hFFFBA805 , 32'hFFFA6718 , 32'hFFFE81F1 , 32'h00003915 , 32'hFFFFE803} , 
{32'h0045D2F7 , 32'h00CEDE6F , 32'h0063B778 , 32'hFF326E4D , 32'h0236D9B4 , 32'hFF7E7BEB , 32'h000D5891 , 32'hFF6DE293 , 32'hFEA3B260 , 32'hFF52DBD8 , 32'h01152B8C , 32'hFE59EA08 , 32'h034C9210 , 32'h01963C68 , 32'hFF6D9B7B , 32'hFF25F785 , 32'hFDEAD18C , 32'hFFC9AB20 , 32'hFF1AB254 , 32'h007C6917 , 32'hFADAFC00 , 32'h0122BCAC , 32'hFF7F5FF2 , 32'h02250A88 , 32'h0078716A , 32'hFEF5ADC0 , 32'h025132BC , 32'h0002721F , 32'hFDFE90D4 , 32'hFEEFCA60 , 32'h00841CFE , 32'h04F66930 , 32'hFF073211 , 32'hFEC12D50 , 32'h0344B378 , 32'h05160BB0 , 32'hFCF1EF0C} , 
{32'hEF9C43A0 , 32'h0ADF3760 , 32'hFA1A4458 , 32'h04088F68 , 32'h01776D90 , 32'h089FD9D0 , 32'h00165F77 , 32'hFF4E3940 , 32'hF54C73D0 , 32'hFB5DD758 , 32'h01C968D8 , 32'hFE675B88 , 32'hFCDAD2AC , 32'hEFE961C0 , 32'hFCE98FAC , 32'h02593150 , 32'hF8F36680 , 32'h027A81A0 , 32'h0DEDA5A0 , 32'hFD97D500 , 32'h0A37D120 , 32'hEFCCDB00 , 32'hFC193FE4 , 32'hFF6E1A82 , 32'hF608EAF0 , 32'h0124D2EC , 32'h0368FBA8 , 32'h0F0EE860 , 32'hFD786F78 , 32'h0312F568 , 32'h0217AF34 , 32'h0640FF40 , 32'hF98BAFE0 , 32'hF6C578A0 , 32'h02C5AFB8 , 32'h006F2406 , 32'hFBAD6D70} , 
{32'h0AFC0B80 , 32'h1661E040 , 32'h019BD38C , 32'hE4944FC0 , 32'hFF8173FA , 32'hEF1E75A0 , 32'h0A6B7D60 , 32'hF7231A10 , 32'hF65E7190 , 32'h015C9434 , 32'hFB668678 , 32'hE36D1A40 , 32'hF2C7F0C0 , 32'h1F8673E0 , 32'hFF7141FA , 32'h0DFE3C30 , 32'hE75FF8A0 , 32'h04A7A5D8 , 32'h08BFB070 , 32'h09E40EF0 , 32'hE13C63E0 , 32'hFC58CF34 , 32'hFF4DC8D3 , 32'hF20D6200 , 32'h02D53C4C , 32'hF05A1080 , 32'hECBEE2A0 , 32'h093788C0 , 32'h046AFF10 , 32'h0A9F15E0 , 32'h10C37040 , 32'h12C81100 , 32'h08A473C0 , 32'h030E9808 , 32'h1879DE40 , 32'h00BD7302 , 32'h12A5F0C0} , 
{32'hFA968AC8 , 32'hF65AA3B0 , 32'hF19C37D0 , 32'hEFB10120 , 32'h025EBD44 , 32'h0362EF38 , 32'h05E5E630 , 32'h052D0B98 , 32'hF96DB6C0 , 32'hF1FE4A70 , 32'hFC8E7BEC , 32'hE8D7FAE0 , 32'h10FD6E80 , 32'h0C8BC6A0 , 32'hF3F60D80 , 32'hDCBFE200 , 32'h00778877 , 32'h1669C5A0 , 32'hFE8478B8 , 32'h159ED9E0 , 32'hFE1EC194 , 32'hE8C17F80 , 32'hD1392900 , 32'hE733D4E0 , 32'h168348C0 , 32'h15C767C0 , 32'h0CEBC1A0 , 32'hFDC4070C , 32'h029CF4B8 , 32'hDF65BAC0 , 32'hEF979CC0 , 32'h07D11AD0 , 32'h002C312B , 32'hFE297F54 , 32'hE633C660 , 32'h15B7CFC0 , 32'hFE609BAC} , 
{32'hFDA0FFDC , 32'hF5868040 , 32'hDE0FE200 , 32'hFA13E680 , 32'hF28E9F00 , 32'hF158E720 , 32'h09942830 , 32'h043A9310 , 32'hF981AAA0 , 32'h05412EA8 , 32'hFDA734F8 , 32'h0429FB10 , 32'h121D3B40 , 32'h02E0F844 , 32'h14C2A7C0 , 32'hFA007460 , 32'hF3031820 , 32'h1567C500 , 32'hFDAADEF4 , 32'hFA7BAAA0 , 32'h038B3584 , 32'hED22E060 , 32'hF43D3250 , 32'hEEE4C9E0 , 32'h01D14D94 , 32'hFEC3146C , 32'hFB363B28 , 32'hF5100500 , 32'h0E1687F0 , 32'hF7048FF0 , 32'hF04723D0 , 32'h0DF85D00 , 32'hFBD74038 , 32'h15D3E400 , 32'hFF3BE972 , 32'hF00A87B0 , 32'hFC20F5CC} , 
{32'hFF0573A8 , 32'h1428EF60 , 32'hDC3E9C00 , 32'hF59762C0 , 32'hFB12EAA0 , 32'hE94AA700 , 32'hF4FE4410 , 32'h1B0C1820 , 32'h061CCA80 , 32'hF66B1F50 , 32'h1E7D3D60 , 32'hFE225224 , 32'h0132FCF4 , 32'h00EF9762 , 32'hFD819A2C , 32'hECF98220 , 32'hE6B40A60 , 32'h00608DEC , 32'hF5109460 , 32'h070BB5B8 , 32'h08650B90 , 32'hF2B22C40 , 32'hFA08D420 , 32'hF2C77420 , 32'h17DF24E0 , 32'h16620B40 , 32'h00A8DAF1 , 32'hE711D420 , 32'h06C9D038 , 32'h07ADE2F0 , 32'hFC7414D4 , 32'h1737F8C0 , 32'h1FD15B40 , 32'hF996CE48 , 32'hF7701750 , 32'hFE96F2B4 , 32'h057EF168} , 
{32'hEF3FF6C0 , 32'h01785088 , 32'hF2B39EC0 , 32'hF202D880 , 32'h0475A2E8 , 32'hEDCBA540 , 32'hFBCE4250 , 32'h06C83C00 , 32'h01EBFE44 , 32'h02FC5814 , 32'h0723BEB8 , 32'h02656B08 , 32'h00C34538 , 32'hFE646E7C , 32'hF0A3E8B0 , 32'hF2594B80 , 32'hF9E67260 , 32'hF8BEFE58 , 32'hFAA43F20 , 32'hF487E270 , 32'h08798260 , 32'hFEB65A98 , 32'hF75E1CD0 , 32'hEF6EC7A0 , 32'h0DA29A70 , 32'h06EBF658 , 32'hF74584C0 , 32'hFDBC0250 , 32'h007E30DC , 32'hFE99420C , 32'h068E91C8 , 32'h04410620 , 32'hFEF9FE1C , 32'hF9264E68 , 32'h10F3A6C0 , 32'hFBBE8C90 , 32'h001CC471} , 
{32'h060EE358 , 32'h06A23460 , 32'hE5C1E6A0 , 32'h00273872 , 32'hF3615900 , 32'hDAEB0EC0 , 32'hF3DE6AB0 , 32'h02E5F090 , 32'h164BB6E0 , 32'hEF263340 , 32'h1C6AC640 , 32'h12409680 , 32'hF42C1580 , 32'hF2027520 , 32'hC4271480 , 32'h0C9D59D0 , 32'hDB2C7880 , 32'h05115D20 , 32'hF64B0DB0 , 32'hFC677C6C , 32'hF457DA80 , 32'h0E9B7DF0 , 32'h0075BFCE , 32'h06394870 , 32'h029B7A6C , 32'h029CAC04 , 32'h1B188E20 , 32'hF7BC8530 , 32'hFFE51DA3 , 32'hFBD58B40 , 32'hF49A1200 , 32'hFEA2E07C , 32'hFD3F4EA8 , 32'h09491310 , 32'hEAAA4BC0 , 32'h016F7E5C , 32'hE1594280} , 
{32'h02B303CC , 32'h09F15650 , 32'hEAA275A0 , 32'hEED1B500 , 32'h1219CF00 , 32'hC7755AC0 , 32'hF60E5960 , 32'h0A643910 , 32'hFD6269AC , 32'hEE4F6200 , 32'h201D9D80 , 32'h0EDDF570 , 32'hE0E90EC0 , 32'hF73D1FE0 , 32'hC2E9E500 , 32'h2A83CEC0 , 32'hEA047680 , 32'hFACC5068 , 32'hEB349C00 , 32'h05F3FD60 , 32'h30FED180 , 32'h13E32440 , 32'h1DDDFCE0 , 32'hF0BC27D0 , 32'hF2EBC350 , 32'hF4465410 , 32'h1F182700 , 32'hF9213590 , 32'h07CB9550 , 32'h06BF4A68 , 32'h02F5CB78 , 32'hFFF956AA , 32'h04648D98 , 32'h09134D30 , 32'h06363FB8 , 32'h09405BC0 , 32'hFAA9E8E8} , 
{32'h03D1A6A4 , 32'h03EF3E0C , 32'h08B26060 , 32'h09B10490 , 32'hFC75D72C , 32'hF9D592B0 , 32'hFA02F288 , 32'h09947C20 , 32'h000BEA2F , 32'hE93A2940 , 32'hFE1860E8 , 32'h0E1EFAE0 , 32'hF97602F8 , 32'h12809400 , 32'hF8A1DEC0 , 32'hFCB53558 , 32'hF9FF50B8 , 32'h00D393E9 , 32'hFD89D07C , 32'hF58CACB0 , 32'h034D0C9C , 32'h00DE312D , 32'hFE53084C , 32'hF83C2788 , 32'hEBC928C0 , 32'hF2124800 , 32'h00A99B89 , 32'h066D6BD0 , 32'hFA95F6D8 , 32'hFD357A30 , 32'hFFC636E0 , 32'hF73FF6D0 , 32'hF72E9E90 , 32'h0A3B9E80 , 32'h08E0B950 , 32'hF5FE8130 , 32'h00650AE4} , 
{32'hFB0B7720 , 32'h0061DB66 , 32'hFA0C2A08 , 32'h1B70F6E0 , 32'h0BC7DFE0 , 32'hF7674F20 , 32'hF3C67C70 , 32'h0D7BC930 , 32'h01509E38 , 32'hF7F477F0 , 32'hFE6EDDD4 , 32'h1E103D60 , 32'hF8BDF348 , 32'h0DB55040 , 32'hCF38CD80 , 32'hFCD09684 , 32'h1628D580 , 32'h194153E0 , 32'hED3B2620 , 32'hF601E900 , 32'h05E8BA98 , 32'hFFE13235 , 32'hE4FE5760 , 32'h0D3D1A70 , 32'h00FB81CE , 32'h01C9424C , 32'h03A8394C , 32'hFAE9B8C8 , 32'hDFE43900 , 32'h193CAFC0 , 32'h15D51F20 , 32'h07E53D00 , 32'hF9351ED8 , 32'h07FB04E8 , 32'h0C095D10 , 32'h01D066D0 , 32'h13C95940} , 
{32'hEDF52EC0 , 32'h0C324680 , 32'hF81AD990 , 32'h0B5D1FD0 , 32'h03A9975C , 32'h12E29880 , 32'hEB81E060 , 32'h0B6C1B90 , 32'hFF8EB387 , 32'h03ABFC50 , 32'h0AAD0A60 , 32'h0A8390A0 , 32'hFA4432F0 , 32'h1346FAE0 , 32'hF3D264C0 , 32'hFB7EA4A8 , 32'h186FE880 , 32'h09C3FE60 , 32'hF24367D0 , 32'hFFB63B21 , 32'hEC6C5DA0 , 32'hEB1F0280 , 32'hEC3E9200 , 32'h19E58B80 , 32'h01C48364 , 32'h04724188 , 32'h13118D80 , 32'hF6BF50C0 , 32'hF83152C0 , 32'hFBE07118 , 32'h1388BD00 , 32'hF966C010 , 32'h0B81FF30 , 32'h12F9CB20 , 32'hEF6C7860 , 32'h00DF6475 , 32'h09A6C070} , 
{32'hFDB3EDC4 , 32'h07012720 , 32'hFFCA349D , 32'h0515E138 , 32'h04C49048 , 32'h00E88D6C , 32'h0058B420 , 32'h09CEB7B0 , 32'hFB7F6528 , 32'h0537B3F8 , 32'hFBF43430 , 32'h04A48750 , 32'hF54F3F10 , 32'h1885C1A0 , 32'hFBC6CB28 , 32'h029CC824 , 32'h0E677240 , 32'h06B0CB08 , 32'hFD07CF94 , 32'h15B64160 , 32'hF0189200 , 32'hDD88D800 , 32'hEEC144C0 , 32'h06C35178 , 32'hFB548F00 , 32'h0F1C8C30 , 32'hF9EE9F38 , 32'hF841A5F8 , 32'hF6F631B0 , 32'h018C1D88 , 32'h1429DEC0 , 32'h03B4E514 , 32'h04D506F0 , 32'h0DC2E410 , 32'hF4DCC810 , 32'hF8C57C50 , 32'h0072DCF3} , 
{32'h01ACBF8C , 32'h09D03C70 , 32'hFA09F658 , 32'hFB6E9758 , 32'h0D1B8F50 , 32'hFC1DDA6C , 32'hFC067FD4 , 32'h0A57A3F0 , 32'h05472D48 , 32'h08065B20 , 32'h13E08F00 , 32'hFC07992C , 32'h04CF09D0 , 32'h01552B18 , 32'hDA568E80 , 32'hFC1592A4 , 32'h105CBB20 , 32'hF0DF3DC0 , 32'hFB6287F8 , 32'hF2A32B00 , 32'hF5FE8220 , 32'hF97702F0 , 32'hE26A8CE0 , 32'h0CC1DE70 , 32'hF77C94F0 , 32'h0D7CC1C0 , 32'hE36F1220 , 32'hF7414EC0 , 32'h12675FE0 , 32'h04C44F80 , 32'h1CE292A0 , 32'hF623A800 , 32'h1C3BB160 , 32'hF71482E0 , 32'hF1EB9D90 , 32'h0A16C080 , 32'h01BE2960} , 
{32'hFEBF0C00 , 32'h0F1F2A20 , 32'h09D39E40 , 32'hF8E99930 , 32'hE9A38D20 , 32'h02EECF58 , 32'h18A37CA0 , 32'h259A3E00 , 32'h05702D18 , 32'h00D9AB75 , 32'hFD5D5838 , 32'hE96ECA60 , 32'hEAF94080 , 32'h17B28660 , 32'hFE0EAE3C , 32'h09896F00 , 32'h2BAA5200 , 32'h16C5B4C0 , 32'hF2A19A10 , 32'hEFE68680 , 32'hEE1BB540 , 32'hE9888E20 , 32'h08C0EB10 , 32'hFAA93E00 , 32'hF621F8C0 , 32'h0CF22CD0 , 32'hDCF53F80 , 32'h1B69D740 , 32'h0BCC8AF0 , 32'h274C8C40 , 32'hECC91CA0 , 32'h05A4BFE8 , 32'hE450AAA0 , 32'h1093EA60 , 32'hF1B03610 , 32'hEF59A100 , 32'hDCA2F680} , 
{32'h0061A4A5 , 32'h11520080 , 32'hEF4708C0 , 32'hFEF2B358 , 32'hF5254990 , 32'h0AC4EAB0 , 32'h1A21ABC0 , 32'h21F3F480 , 32'h12357180 , 32'hFB97A908 , 32'h1E699640 , 32'h0FC65560 , 32'hE1B4B680 , 32'h0949ADA0 , 32'h15A379E0 , 32'h0CBFAE10 , 32'h18EE4420 , 32'h231651C0 , 32'hFB1B0220 , 32'h16D2B520 , 32'h04BC8860 , 32'hF02C86E0 , 32'hF960E1E8 , 32'h06169E08 , 32'hF8446008 , 32'hE6353F60 , 32'h03410B68 , 32'hFBC90700 , 32'hFFBD9BA4 , 32'hFEC79984 , 32'h06901298 , 32'h06782540 , 32'h0D94FB70 , 32'hFBFD3338 , 32'hEF9F2A60 , 32'hF2BE2050 , 32'h1584B5E0} , 
{32'h022B2198 , 32'h18092D20 , 32'h01865310 , 32'h00908061 , 32'hF1371800 , 32'h0D916CB0 , 32'h1C84D240 , 32'h2437F1C0 , 32'h0DC85CD0 , 32'hD8259E40 , 32'h1505F340 , 32'h010EA2AC , 32'hE88C9E60 , 32'h1B971400 , 32'h23E5A700 , 32'h13FB3D40 , 32'h02793388 , 32'h0F71A260 , 32'h14A9F900 , 32'h02B8CF68 , 32'h067515B0 , 32'hFEB0B6E8 , 32'h04621C68 , 32'hEC6598A0 , 32'hF5B666D0 , 32'hE6136EE0 , 32'h016CD958 , 32'hF0D4F240 , 32'hF4528820 , 32'hEE17DF00 , 32'hF9E742D0 , 32'h05C0D518 , 32'hFB72B2D8 , 32'h02BA50B8 , 32'hFEAFD594 , 32'hF230C510 , 32'h123C29A0} , 
{32'hEA0D4620 , 32'h1049C980 , 32'hF2EC8B60 , 32'h0A3180B0 , 32'hF9A80DB8 , 32'h084D1700 , 32'h080251A0 , 32'h0D0BAE20 , 32'h0257A844 , 32'hF402D6D0 , 32'hF7017690 , 32'hF42C35A0 , 32'hF94E95A0 , 32'h14DAF4A0 , 32'h09E072A0 , 32'h0CFE5540 , 32'hE0450FC0 , 32'h050E6310 , 32'h0F70A4F0 , 32'hEF1CF560 , 32'h070D42B0 , 32'h050CCE10 , 32'hFFA2EB85 , 32'h04F079B8 , 32'h063DBE78 , 32'h08CE3940 , 32'hECDA2FC0 , 32'hF043A260 , 32'hFD859138 , 32'h03833F5C , 32'hFC8566B0 , 32'hF444CA00 , 32'h03E51338 , 32'h0F560E10 , 32'hF9A26350 , 32'h0BEE4640 , 32'hFEDDFC98} , 
{32'h0135D6CC , 32'h08527CA0 , 32'h0277DE90 , 32'h07B881C0 , 32'hFF1808B9 , 32'hFACEB698 , 32'hFEB6A5DC , 32'h035D9F1C , 32'h010A7B1C , 32'hEE945D60 , 32'h06726758 , 32'hFE077BB0 , 32'hEA8053E0 , 32'h201E8C00 , 32'h071C5190 , 32'hFE2C6EF0 , 32'hF8960BA0 , 32'hFC6B2FE4 , 32'h0F351A90 , 32'hF5AA57B0 , 32'h0AC01530 , 32'h04747B50 , 32'hEA572940 , 32'hFB966040 , 32'hE94EAEE0 , 32'hF7C7C7E0 , 32'h00C518B9 , 32'hFDFF3D34 , 32'h015E984C , 32'hFF5D3411 , 32'hFAA1CC58 , 32'hFB262880 , 32'hFFC29CBC , 32'h009D88A4 , 32'hFBC855B0 , 32'hEBF37420 , 32'h05A7A678} , 
{32'hF32C51E0 , 32'h00D2A74D , 32'h089DD890 , 32'hF8DFDC90 , 32'h0205EF84 , 32'hFE9D93D4 , 32'hF3F61E10 , 32'h082B7950 , 32'h079064E8 , 32'hF27E2DF0 , 32'h034B0F00 , 32'h0D1A2E50 , 32'hE8496020 , 32'h1542A540 , 32'h01C2FB90 , 32'hFD8199D0 , 32'hF9CCF488 , 32'h04CD63E8 , 32'h05730E40 , 32'hF4AD44D0 , 32'hFA5A6A98 , 32'h0016F9FE , 32'hFECAD23C , 32'h00459266 , 32'hF67FAA10 , 32'hF893FE70 , 32'hF6265820 , 32'h04CE4D20 , 32'h031C715C , 32'hF6B158C0 , 32'hFCA9712C , 32'hFF5BDA0F , 32'hF783CA50 , 32'h04FA81F0 , 32'hFC6B75A8 , 32'hF24D96F0 , 32'h08701C70} , 
{32'hEFD364C0 , 32'hFB1C3E40 , 32'h049DCC08 , 32'hEFE125A0 , 32'h03CA27B4 , 32'h03E4AF7C , 32'hF4232350 , 32'h0691EC88 , 32'h0782AB90 , 32'hFCD74994 , 32'hFCFCE40C , 32'h07DF92D8 , 32'hF9E0E990 , 32'hFE80A3BC , 32'hFB6EE440 , 32'h01CD2070 , 32'hFE46DD24 , 32'h0A2C9710 , 32'hFD423550 , 32'hF909F590 , 32'hF8357750 , 32'h004ED67B , 32'h0E753C10 , 32'h0B1D0530 , 32'h01A72534 , 32'hFE100AB0 , 32'hF5B12E20 , 32'h01C95178 , 32'hFBE9EFF0 , 32'hF32574C0 , 32'hFA129C60 , 32'h0A64A770 , 32'hF98599A0 , 32'h01FC135C , 32'hFA917C68 , 32'h01D913C0 , 32'h0433E420} , 
{32'h00027C1B , 32'h0001B244 , 32'hFFFA3A76 , 32'h0002F1AD , 32'hFFFECE8C , 32'hFFFBF57B , 32'hFFFE3D5F , 32'h0002CB43 , 32'h000392B1 , 32'h00041DBA , 32'hFFFD9954 , 32'h0002E790 , 32'h0002F671 , 32'h0000092A , 32'hFFFA824B , 32'hFFFD90FD , 32'hFFFDD2A4 , 32'h0000F655 , 32'hFFFF5238 , 32'hFFFEFB78 , 32'h00017381 , 32'h00027474 , 32'h00066D1A , 32'hFFFCCCFB , 32'hFFFDDB56 , 32'hFFFF8D65 , 32'hFFFFF3BA , 32'hFFFC9B5A , 32'h00001A80 , 32'h0000D304 , 32'hFFFA6B0E , 32'h0002CCF7 , 32'hFFFFFDD6 , 32'h0001DFB1 , 32'h00033539 , 32'hFFFED71E , 32'hFFFAF4B2} , 
{32'h00022603 , 32'h00009C41 , 32'h0003C0F3 , 32'hFFFDE746 , 32'hFFFCC0E1 , 32'hFFFD5CCC , 32'hFFFD416E , 32'hFFFF1740 , 32'hFFFE59FE , 32'hFFFE810C , 32'h000045CE , 32'hFFFF4C59 , 32'h00037DA5 , 32'h00028E80 , 32'h0006506B , 32'hFFFC3D2A , 32'hFFFD5772 , 32'h0002C519 , 32'h0000298E , 32'h00015DF2 , 32'h0005736E , 32'h0002215A , 32'h0001D4A4 , 32'h0001BC34 , 32'hFFFC58B8 , 32'hFFFD40A2 , 32'hFFF9DBD4 , 32'h00074037 , 32'hFFFC055F , 32'hFFFEF61D , 32'h00026993 , 32'h0001A778 , 32'h00040DEC , 32'hFFFFB49F , 32'h0001434A , 32'hFFFEE1BF , 32'hFFFB14C4} , 
{32'hFFFFC9AA , 32'hFFFC1B89 , 32'h0005196C , 32'hFFFEA6A6 , 32'h0000A709 , 32'hFFFE3FF3 , 32'h0006AF1E , 32'hFFFF6B60 , 32'h000068B5 , 32'hFFFD7990 , 32'h00065101 , 32'hFFFB64B4 , 32'hFFFE1B73 , 32'h0002B218 , 32'h0003F7F4 , 32'hFFF90AC7 , 32'h0000F538 , 32'hFFFF3439 , 32'h0004A963 , 32'h0000AB9A , 32'h00006ACA , 32'hFFFFF28F , 32'hFFFB6624 , 32'hFFFC439D , 32'h0001D828 , 32'h0002EEDD , 32'h00024B8D , 32'h0000F13C , 32'hFFFA1494 , 32'hFFFD365A , 32'hFFFFDC77 , 32'h0002C156 , 32'hFFFEAC5F , 32'hFFFAC0B3 , 32'h00010D0A , 32'hFFFED5A4 , 32'h00016AF4} , 
{32'h00014F00 , 32'hFFF8FAE8 , 32'hFFF9A17C , 32'h00021908 , 32'h000036B9 , 32'hFFFDB7A2 , 32'h0002C822 , 32'hFFFFE69B , 32'h0002357E , 32'hFFFE59CA , 32'hFFFE65BD , 32'h00033735 , 32'hFFFB6CDE , 32'hFFFEF28E , 32'hFFFF56DA , 32'hFFF9B8AB , 32'h0006C4FB , 32'h000555ED , 32'hFFFEEF1F , 32'hFFFCAC56 , 32'h00052723 , 32'hFFF8E4E4 , 32'hFFFD3605 , 32'hFFFC8FBC , 32'hFFFE3AE4 , 32'h00026539 , 32'hFFF6ED78 , 32'hFFFEDE1B , 32'hFFFEC695 , 32'hFFFDE2B6 , 32'h00011613 , 32'h0005C55A , 32'h00042A3B , 32'h0003D100 , 32'hFFFC2C18 , 32'h0001923C , 32'hFFFC353B} , 
{32'hFFFEFE31 , 32'hFFFFB623 , 32'hFFFA599E , 32'hFFFADB66 , 32'h0002787C , 32'hFFFBD4E9 , 32'h0003914D , 32'hFFFF4F6A , 32'h0001470F , 32'hFFFCD98E , 32'hFFFDC823 , 32'h00022D9B , 32'hFFFFE74F , 32'h0000B4B1 , 32'h0001BDBA , 32'h0003BAA8 , 32'hFFF8834D , 32'h000356DE , 32'h00033837 , 32'h0001C0EA , 32'h00060414 , 32'h0000959A , 32'hFFF86069 , 32'hFFFCB57F , 32'hFFFD54CC , 32'hFFFB9674 , 32'hFFFA1557 , 32'hFFFB9EFE , 32'hFFFCD026 , 32'hFFFB3C04 , 32'h0001C758 , 32'h0002DF0D , 32'hFFFF3129 , 32'hFFFFBE11 , 32'h000258EB , 32'h00079185 , 32'hFFFF1C8F} , 
{32'hFFFE2361 , 32'hFFFBF633 , 32'hFFFFF264 , 32'hFFFB17FA , 32'hFFFEB8CE , 32'hFFFB9490 , 32'h000467A9 , 32'h00029A4E , 32'hFFFA5B0E , 32'h00059E4E , 32'hFFFF5365 , 32'h0002887F , 32'h00017A04 , 32'h000672BF , 32'hFFFE4910 , 32'hFFFEE36A , 32'h0002C4B9 , 32'h0006F95F , 32'h0001E542 , 32'hFFFEC762 , 32'hFFFFE8FA , 32'hFFFF7485 , 32'hFFFF07A4 , 32'h0005B222 , 32'h0001C061 , 32'h0003D60D , 32'hFFFF2744 , 32'h00016962 , 32'h000193ED , 32'h000101CA , 32'h000060EF , 32'h0003BB18 , 32'hFFFE070C , 32'h0001D6DE , 32'h0002868A , 32'hFFFDEF87 , 32'h00075516} , 
{32'hFFFEA6AF , 32'h00019697 , 32'h0001CD91 , 32'hFFFE1154 , 32'hFFFEC953 , 32'h0001B8B6 , 32'h00031C2E , 32'hFFFFF249 , 32'h000079E6 , 32'hFFFCD109 , 32'h00001155 , 32'hFFFBAF2E , 32'hFFFEFD5C , 32'hFFFFFC12 , 32'h000193AB , 32'hFFF8E441 , 32'hFFFCE811 , 32'h0006E7D6 , 32'hFFFE7C7B , 32'hFFFC58BC , 32'h0005F8CD , 32'h0000AB7D , 32'h000347F6 , 32'hFFFCB637 , 32'h00025145 , 32'hFFFD4939 , 32'h00030B75 , 32'h0000E996 , 32'hFFFED38E , 32'hFFF9F702 , 32'hFFFB8C91 , 32'h0002F528 , 32'h00034D16 , 32'h00006B2F , 32'hFFFEB5A5 , 32'h00022474 , 32'hFFFF7F7A} , 
{32'h041BF0E0 , 32'h00B32434 , 32'hFAF17150 , 32'hFE259E28 , 32'hFF2AB2A9 , 32'h038B7DD4 , 32'hFC4CD840 , 32'h01F8F94C , 32'hFB51B068 , 32'h0042BE85 , 32'hFA825930 , 32'h007D5F57 , 32'h01E64088 , 32'h03D6AF50 , 32'h00E8FA84 , 32'hFC9905E8 , 32'h04F0B028 , 32'h042F2658 , 32'h0123324C , 32'hFE46570C , 32'h01EA6F6C , 32'hFDD004F4 , 32'hFB556A48 , 32'hFFE27983 , 32'h021584E4 , 32'h03757E70 , 32'h08BBDA40 , 32'h01156700 , 32'h00DA7A8B , 32'hFEF3EA58 , 32'hFEAB8768 , 32'h0419CB80 , 32'h031A789C , 32'h0062FFEC , 32'h0126BB20 , 32'h028B246C , 32'h07C55580} , 
{32'hFFD4A753 , 32'hFFFCF917 , 32'hFFD9C8B3 , 32'h000EDED0 , 32'hFFE2856E , 32'hFFF1527D , 32'hFFF83B77 , 32'h0000B36A , 32'hFFED4BB0 , 32'h000BEE47 , 32'h0017C5BA , 32'hFFE91CFC , 32'h00090179 , 32'h000B15C2 , 32'h0006E53F , 32'hFFEBC045 , 32'h0006F088 , 32'hFFEBA0DC , 32'hFFEE453A , 32'h000F4CB9 , 32'hFFF247E5 , 32'h00201231 , 32'h0003DEFC , 32'h000B14BB , 32'hFFC51AFF , 32'h000541B5 , 32'hFFF3B8C1 , 32'h000249D2 , 32'hFFDE06A4 , 32'hFFFBEC18 , 32'h0005BEA2 , 32'hFFEDCE5D , 32'h000461D1 , 32'hFFFF5474 , 32'h0027B269 , 32'h000320A0 , 32'h00234C17} , 
{32'hFFBA7EAB , 32'h0695A8B0 , 32'h01F8CED0 , 32'h07DBD740 , 32'hED0E5A60 , 32'hF5F701B0 , 32'hF8198080 , 32'hFB6862F0 , 32'h055296C8 , 32'hFFC0213C , 32'h08F8BDC0 , 32'hEE4C3BC0 , 32'h00AB4D12 , 32'hF85FDFE0 , 32'h06FD8720 , 32'hED73D3A0 , 32'hE8E295A0 , 32'h0C9182F0 , 32'hF91E4DC0 , 32'h03F46A28 , 32'hFE1B8348 , 32'hF8C1F388 , 32'h00A9635E , 32'hFC68A8BC , 32'h13728B80 , 32'hFD812A00 , 32'h05AFC1E0 , 32'hF9E08FF8 , 32'hF6D85130 , 32'h082EB1E0 , 32'hF3F70F40 , 32'h0A629860 , 32'h00E9A160 , 32'h057A0A98 , 32'hFBD6B198 , 32'hF508F2A0 , 32'h02BBC790} , 
{32'hF93828D0 , 32'hF2CB1950 , 32'h0695ABB0 , 32'hF3813350 , 32'hEC0B82A0 , 32'hFCB8B188 , 32'h1B77E860 , 32'h03BB6D1C , 32'hFA876CD8 , 32'hF522CEA0 , 32'hF6328180 , 32'hF082E420 , 32'h101C9B00 , 32'hFFB963AF , 32'hFB04F0C0 , 32'hEAF0F540 , 32'hF5734770 , 32'h1B712000 , 32'hFD9EF78C , 32'h10508B20 , 32'h0A490310 , 32'hF9796690 , 32'hE05AF460 , 32'hEADDBA60 , 32'h062A54E0 , 32'hFC23A9D4 , 32'hF482F550 , 32'h08893090 , 32'hF98C6090 , 32'hF8FD4B78 , 32'hF5D64180 , 32'h06C559B8 , 32'hF582C7C0 , 32'h08E0F290 , 32'hDD9F4F80 , 32'h0DCC1880 , 32'hEE119620} , 
{32'hEEA79B80 , 32'h0BD79C20 , 32'hEAEF25E0 , 32'hF2362950 , 32'hE7BEA560 , 32'hE6AA6C80 , 32'h05EA91D8 , 32'hFB572698 , 32'hFFCA5B39 , 32'h06F2E2E8 , 32'h0C326000 , 32'h00FA04BA , 32'h04D32358 , 32'h004BA3CA , 32'hE8B228E0 , 32'hE989D5A0 , 32'hF6CA2C80 , 32'h11030F80 , 32'h011F2928 , 32'h1083C360 , 32'h01B66BAC , 32'hF5F47B60 , 32'hF2D68E00 , 32'hF635B8B0 , 32'h00FABFE9 , 32'h138CF480 , 32'hFF80E2AB , 32'hE72EE800 , 32'hED741120 , 32'h1475E360 , 32'hF7CDDD10 , 32'h1A84D3C0 , 32'hF240DFD0 , 32'h0E03B2E0 , 32'h014D77DC , 32'hFAEFC0F8 , 32'h013F2BD0} , 
{32'h0211C1D0 , 32'h08DCED20 , 32'hFA086628 , 32'hE77E6000 , 32'hFAD1D4D0 , 32'hF100D5E0 , 32'h11150B00 , 32'h050A6218 , 32'hF38CA230 , 32'hFE4255A8 , 32'hEFA5F8E0 , 32'hFC8371D4 , 32'h03C00390 , 32'hF77E5B10 , 32'hF55B7EC0 , 32'hF6A811C0 , 32'hEC5FFD20 , 32'h14466580 , 32'hFE1D39A0 , 32'h02598208 , 32'h0E6F2690 , 32'hFA318E90 , 32'h09DB5220 , 32'hFB8EACF0 , 32'hF558D870 , 32'h0B7A2110 , 32'h0F253EC0 , 32'hF9CE2B10 , 32'hF49CCB20 , 32'h0AB3F540 , 32'h0512DB48 , 32'h019F2F70 , 32'hF6A140C0 , 32'h17217220 , 32'h0950CE20 , 32'hF50BE7F0 , 32'hF8E7FC90} , 
{32'h07B1ABD8 , 32'h1927FFE0 , 32'h015D4DAC , 32'h03D565B0 , 32'hF1A01D20 , 32'hFCC13458 , 32'hF6953B70 , 32'h03CEC2A4 , 32'hFD65DA24 , 32'hF8875988 , 32'hF4AF9750 , 32'h0A677C30 , 32'hFCD49BE0 , 32'hF38FD8B0 , 32'hF2988830 , 32'hFEA3CE30 , 32'hE84E8D60 , 32'h040AA7D0 , 32'h08C3DA80 , 32'h0C3E7300 , 32'h01CC4DC4 , 32'hFE53CCDC , 32'hF88CD7B0 , 32'hFDACA408 , 32'h0AB27810 , 32'hFAEBE0A8 , 32'h0A1991D0 , 32'h05B36890 , 32'h0C83FAA0 , 32'h0208B3B0 , 32'hEFF719C0 , 32'h0C4E1770 , 32'hF72A6240 , 32'hFEAD02B8 , 32'hFDB480FC , 32'hF54E5350 , 32'hFEA5BC84} , 
{32'h0BF8E4B0 , 32'h127A4100 , 32'hFEEA9D5C , 32'hFCBA2B94 , 32'h0F82A2E0 , 32'hEADB0820 , 32'hECDABB00 , 32'h03D531A8 , 32'hF68CC290 , 32'hFE5D5390 , 32'hE9DDE320 , 32'h141A4C20 , 32'h02F48370 , 32'h0D0A11E0 , 32'hE3BAB440 , 32'hFF532183 , 32'hE5E8C440 , 32'h0726DB98 , 32'hF0E6C1B0 , 32'hFA8349D0 , 32'h0C459E80 , 32'h0362AE74 , 32'hF1F53180 , 32'hEA241EA0 , 32'h06130B30 , 32'h0B0B8E90 , 32'hF59E0F20 , 32'h06CDF2C8 , 32'h0149C1C4 , 32'h086AE580 , 32'h038B7118 , 32'h0F2ECF60 , 32'hF02CDDB0 , 32'h186A81C0 , 32'hF69E4400 , 32'h02B7EDF4 , 32'hF9587198} , 
{32'hF319A030 , 32'h12472F00 , 32'hFD7B0A08 , 32'h0385BD8C , 32'hF9F0D338 , 32'hF5557E30 , 32'h01DA4ADC , 32'h0B837E60 , 32'hFED16BE8 , 32'hF7E44470 , 32'h0729D000 , 32'h077A77D8 , 32'hFD4360FC , 32'hF536A920 , 32'hD9938380 , 32'hFE571EF8 , 32'hF3761920 , 32'h1A44D060 , 32'hFC5854D4 , 32'hF1CC89F0 , 32'h21F89CC0 , 32'h02FEBB38 , 32'h065D76C0 , 32'hF5478090 , 32'hE9B3DAC0 , 32'h13B2E200 , 32'h16310B60 , 32'h16674AA0 , 32'hFF1A20EA , 32'hFCAE2174 , 32'h0E8BC980 , 32'hE9B8A8C0 , 32'hE965EEC0 , 32'h066AFF58 , 32'hFBF9DD08 , 32'hF5102B10 , 32'hFBEB10A8} , 
{32'hF651F130 , 32'h11947B80 , 32'h09560360 , 32'hF8CCC9E0 , 32'hFB4331A0 , 32'hEC76ADC0 , 32'hE7827E40 , 32'h031C8C40 , 32'hFC31F1C0 , 32'hFC03B664 , 32'h00BF1529 , 32'h0017515D , 32'hF256D030 , 32'h1B25E140 , 32'hDE22D080 , 32'hF965C648 , 32'hF396A0F0 , 32'hFBC7FA40 , 32'h107F9300 , 32'hFEBB148C , 32'h18DF3F00 , 32'hFC9CA740 , 32'hF6B664A0 , 32'hFA537F68 , 32'hD6FEE540 , 32'h093A56B0 , 32'h09607CC0 , 32'hF679A010 , 32'hEF862D80 , 32'hF92CACB8 , 32'h0909FB60 , 32'hE18A8980 , 32'hF1B81CD0 , 32'h02B70B84 , 32'hFC274E3C , 32'hE5970220 , 32'hF8867F28} , 
{32'h0225C8B0 , 32'h36BCD540 , 32'hF7691370 , 32'hE65710A0 , 32'hF23C1F80 , 32'hECE761C0 , 32'h097F0930 , 32'h14000D60 , 32'hF50A1680 , 32'hFCF7FBB4 , 32'h02A1EE94 , 32'hF4CB4260 , 32'h084D4900 , 32'hF779F980 , 32'hC7211A00 , 32'h0D8C3A00 , 32'h04AE3C58 , 32'h004885F7 , 32'h04703038 , 32'hFF7EE11A , 32'h30E9F100 , 32'hFA4F4B88 , 32'hFC6D8ECC , 32'h13B27A40 , 32'hEDE55060 , 32'hFB4DEED0 , 32'h144D6D20 , 32'h0A162CC0 , 32'hEDFA5CC0 , 32'hFFF941E8 , 32'h01C0B708 , 32'hF4EEC100 , 32'hF5254DD0 , 32'hF3BB2550 , 32'h0C9B4C00 , 32'h002C7D2A , 32'h029D82FC} , 
{32'h0D46AC70 , 32'h1633DCA0 , 32'h068C6C30 , 32'hE9699440 , 32'h0C2AB280 , 32'hF11E13F0 , 32'h0C679ED0 , 32'h084A4270 , 32'hFBDE0EC0 , 32'h0062223D , 32'hFAB5E1C8 , 32'h03048FC0 , 32'hF6B50A50 , 32'h02C586D0 , 32'hE73E8A20 , 32'hFB9082F0 , 32'hFB3B98E0 , 32'h17BC05E0 , 32'hEEB90BC0 , 32'h054DAFC8 , 32'h03904984 , 32'hFBBDE9A0 , 32'hF2741E40 , 32'h06560328 , 32'h037492B0 , 32'hFE450EEC , 32'h0755BED0 , 32'h031BB584 , 32'h0B44CD90 , 32'h11B94980 , 32'h2340E1C0 , 32'h06E54F18 , 32'h00B03811 , 32'h067F8898 , 32'h0B442160 , 32'hFA464168 , 32'h09281960} , 
{32'hFABDA160 , 32'h0996A850 , 32'hF5998970 , 32'hF8484DE0 , 32'h0668E990 , 32'h0182C700 , 32'h032141C8 , 32'h08BB5E40 , 32'h00BC5462 , 32'h02150A10 , 32'h05CE5A90 , 32'hFBC91E20 , 32'hFAE7C1C8 , 32'h03F80EC4 , 32'hF0BD2B20 , 32'hF36E2810 , 32'h0F297AA0 , 32'h058CFB60 , 32'hFAB05458 , 32'hFC90C3EC , 32'hF456A580 , 32'hF12E6770 , 32'hF1C1CB40 , 32'h03AD6E54 , 32'h061876E0 , 32'h16678760 , 32'hFF33B093 , 32'hF0478370 , 32'hF6F765F0 , 32'hFB873940 , 32'h05B76700 , 32'h037AFBD8 , 32'h119BAD40 , 32'h095A1970 , 32'h05D493A8 , 32'h07A41288 , 32'h04644B78} , 
{32'hF63B66F0 , 32'h277CD940 , 32'hF79E9510 , 32'hF855A6B8 , 32'h116C53A0 , 32'h09E88D80 , 32'hFEF38270 , 32'h16208500 , 32'hF84BF258 , 32'h159B62C0 , 32'h1608DF60 , 32'hF2D8FCD0 , 32'hE9228B60 , 32'h104F9380 , 32'hDC4133C0 , 32'hEB80C7C0 , 32'h30F3DBC0 , 32'h05D1D2D0 , 32'hEE224D20 , 32'h07E81430 , 32'hD533DBC0 , 32'hE099E5E0 , 32'hE203C1C0 , 32'h09D31920 , 32'hFA387090 , 32'h16DCD6E0 , 32'h09891050 , 32'h02FC1FC0 , 32'h0AD74E30 , 32'h07AEA4C0 , 32'hF4819470 , 32'h05E826E8 , 32'h067DE678 , 32'h0B66E610 , 32'hFEF73EFC , 32'h0EE77340 , 32'hF9034BF0} , 
{32'h084AA9B0 , 32'h1AC2DA20 , 32'h06DF6128 , 32'hFFDAC30C , 32'h0AB88E10 , 32'h0EBEB4B0 , 32'h01C284FC , 32'h191405A0 , 32'h08EEE050 , 32'hEAEAC380 , 32'h0F8B02E0 , 32'hF6224890 , 32'hE692A440 , 32'h13E87200 , 32'h00BC78C5 , 32'h0C5EEB50 , 32'h1D0697A0 , 32'h0473E058 , 32'h03E3DFF4 , 32'hF5A15150 , 32'hF87ACB70 , 32'h0E715750 , 32'hF9B89DD0 , 32'hF5F936B0 , 32'hF50229A0 , 32'h0096F618 , 32'hFCA4DD6C , 32'h0AF4AF10 , 32'h000B9DBB , 32'h1915D7A0 , 32'hED19A540 , 32'h03D7916C , 32'hF26EFBF0 , 32'hFABD9CA8 , 32'h0277F644 , 32'hF5489320 , 32'h01E06298} , 
{32'h01C861EC , 32'h0F1332A0 , 32'hF63B5570 , 32'hF2D41580 , 32'h00D40D31 , 32'h0AF69850 , 32'h12DE12E0 , 32'h18867500 , 32'h05D89BE8 , 32'hEC779DE0 , 32'h0CAFD310 , 32'hF6A8BB10 , 32'hF735AA90 , 32'h07B43C48 , 32'h0BE957E0 , 32'h01558A3C , 32'h0C24F650 , 32'h11DC0600 , 32'hFB1564C0 , 32'h05C874B0 , 32'hF3EA08B0 , 32'hFF9D8552 , 32'h024F5EA8 , 32'hF3E61B50 , 32'hFF21D953 , 32'hFB392FE8 , 32'h03F8A044 , 32'h072F25A0 , 32'hFE10413C , 32'h08453DF0 , 32'hE9DCC0A0 , 32'h0EB9B600 , 32'hF0F73DB0 , 32'hF9FF72B0 , 32'h0159AD78 , 32'hFE3E769C , 32'h12FCF860} , 
{32'h029257A4 , 32'h116A2640 , 32'hF6D5EBD0 , 32'hF7A6DF70 , 32'hFFF0F358 , 32'hFB62EF40 , 32'h1FDC1460 , 32'h22C16180 , 32'h07859F98 , 32'hE2AA6EE0 , 32'h0CD43470 , 32'hFF161988 , 32'hCE1954C0 , 32'h32F06980 , 32'h238404C0 , 32'hF6BA0C50 , 32'hD64EE240 , 32'h00FDFA08 , 32'h1EC79260 , 32'hDBDC8D00 , 32'h0D1438D0 , 32'hDFA40A00 , 32'hE1849940 , 32'hF9FA5570 , 32'hDA84D440 , 32'hE0A57C20 , 32'hF63D0DD0 , 32'hF18AB870 , 32'hFC87C740 , 32'hE89DC760 , 32'h0570FF00 , 32'h2233DFC0 , 32'hFA41BC60 , 32'hE8580CA0 , 32'hE5D37120 , 32'h12B19060 , 32'h16FA6500} , 
{32'hFF68EA5E , 32'h022D39F0 , 32'hFEE23350 , 32'hFE3B24EC , 32'h01662500 , 32'hFCC8EF74 , 32'h08B8E2C0 , 32'h06E3F7C8 , 32'h00E68AA8 , 32'hFFF7B4B4 , 32'h028E19C0 , 32'hFFA61D11 , 32'hF6280260 , 32'h0E4F9B30 , 32'h0BDDDE90 , 32'hFD2611A0 , 32'hEFF53020 , 32'h07E2F9A8 , 32'h0E28F920 , 32'hF429BB00 , 32'h05AF8C20 , 32'hF089AB70 , 32'hF8B4DEB8 , 32'h0675C8C0 , 32'hF638AB10 , 32'hF8571C88 , 32'hFB1AEDE8 , 32'hFCF5DB1C , 32'hFC334554 , 32'hFDC9A740 , 32'h04077CA8 , 32'h082DE950 , 32'hFBA458B8 , 32'hF9FA0FB8 , 32'hF71EA840 , 32'h0935F530 , 32'h01152A98} , 
{32'hF730DEA0 , 32'hFF47FDE3 , 32'hFFBA578D , 32'hFC5FA660 , 32'hFCEE2AEC , 32'hF709F530 , 32'h099AC4C0 , 32'h055265A0 , 32'hF328BA40 , 32'hFE0C7938 , 32'h09137940 , 32'h0698F8F8 , 32'hEFDD1AC0 , 32'h1B4C9000 , 32'h0B4A4470 , 32'h0220464C , 32'hE51C9360 , 32'h08329470 , 32'h1FD28140 , 32'hEDE2E920 , 32'hF9860688 , 32'hEE452DC0 , 32'hF9AB8000 , 32'h143B6880 , 32'h192CD5A0 , 32'h019D26CC , 32'hF8F02698 , 32'h04B93E78 , 32'h0DAFFFE0 , 32'h05191C60 , 32'hF900DB08 , 32'hE289B720 , 32'hEF877560 , 32'h00702BED , 32'h13340020 , 32'h1EA24C80 , 32'h0553B2B8} , 
{32'h0009A1D5 , 32'hFFE6222B , 32'h0004D036 , 32'h0010DA1D , 32'hFFFF3D58 , 32'hFFF15D6B , 32'h00005B9A , 32'h00019E04 , 32'hFFEDE0D6 , 32'hFFE4AC3C , 32'hFFF4BA43 , 32'hFFEFB7B1 , 32'hFFEA3CAB , 32'hFFF603C1 , 32'h000E7A2F , 32'hFFF35788 , 32'h0014F5C1 , 32'hFFF668B1 , 32'h00060AE4 , 32'hFFE5E554 , 32'hFFF5C78C , 32'h0018052A , 32'hFFFD529B , 32'h00121B71 , 32'h002BC34F , 32'hFFD3FC6A , 32'hFFF30900 , 32'h0004ADEF , 32'h001EFE78 , 32'hFFEFEE32 , 32'h00167FA6 , 32'h0012BEE3 , 32'h0017B72C , 32'hFFFE2CC8 , 32'hFFF006CF , 32'hFFF3B5E6 , 32'hFFF5A761} , 
{32'hFFBFFA27 , 32'h00EF3FE2 , 32'h00874A09 , 32'h00220A80 , 32'h03D26920 , 32'hFFB56B6E , 32'h011407A0 , 32'h021CAFFC , 32'h005EC116 , 32'h0486C358 , 32'h02A253B0 , 32'h02000AD8 , 32'h0096A316 , 32'h059A4498 , 32'h079A1A98 , 32'hF7F3C6C0 , 32'hFD03406C , 32'h07A14C68 , 32'h08447720 , 32'hFF105634 , 32'h06C015B0 , 32'hF2993310 , 32'hFC74D5F4 , 32'h01C08FC8 , 32'hF5854DF0 , 32'hF9F0CA08 , 32'h000FC5DA , 32'hFCFC0B00 , 32'h007C76C2 , 32'h043CF9F8 , 32'h065855E0 , 32'h0A3E4130 , 32'h00992374 , 32'hFFE409C1 , 32'hFD593DE8 , 32'h01E24CDC , 32'hF8B93BB8} , 
{32'h00048B40 , 32'hFFFD2259 , 32'h000220C5 , 32'hFFFC9BA3 , 32'h000222BD , 32'h0002DBBF , 32'h000149DB , 32'hFFFF3D12 , 32'hFFFFA84F , 32'hFFFDE21C , 32'h000018FE , 32'h0002795D , 32'h0000971A , 32'h00022CB8 , 32'h00012298 , 32'h0004F36A , 32'h000308AE , 32'hFFFF6326 , 32'hFFFE6AD8 , 32'hFFFD4DED , 32'hFFFB65F1 , 32'h00006FBF , 32'hFFFEBAE4 , 32'h000543A9 , 32'hFFFC0736 , 32'hFFFCB241 , 32'h0003B8EC , 32'h0001FE03 , 32'h0000FFAF , 32'h0000A439 , 32'h00009F85 , 32'h0006CB7C , 32'hFFFE59D1 , 32'hFFFACB13 , 32'hFFFD0EC4 , 32'h00007994 , 32'h00010B50} , 
{32'h00024C75 , 32'h0002A1A2 , 32'h00024EAE , 32'hFFFD80ED , 32'hFFFC1E41 , 32'h00033695 , 32'h00030C28 , 32'hFFFA47A2 , 32'h00005D42 , 32'h00051D14 , 32'hFFFF9E89 , 32'h00049304 , 32'h00040265 , 32'hFFFC31FC , 32'h00021E28 , 32'h0004143A , 32'h00026CC2 , 32'h00015189 , 32'h0000516B , 32'h00037033 , 32'hFFFE9551 , 32'h0006895A , 32'hFFFB0991 , 32'hFFFE0D05 , 32'hFFFCEBBB , 32'hFFFECD32 , 32'hFFFB116E , 32'h0005567E , 32'h00021F1F , 32'hFFFE3C20 , 32'h000136F5 , 32'h0001693A , 32'hFFFA81CE , 32'hFFFC54D4 , 32'h00020D7A , 32'h000142AF , 32'hFFFD7620} , 
{32'hFFFE9B10 , 32'h000095AF , 32'hFFFE6CAC , 32'h0005134F , 32'h00042D79 , 32'h000172D4 , 32'hFFFAA629 , 32'h0004AA29 , 32'h00014310 , 32'hFFFD3A5B , 32'h0000B316 , 32'h00021093 , 32'hFFFBB64B , 32'hFFFDF71A , 32'hFFFE7C3B , 32'h0000E965 , 32'hFFFD7522 , 32'h0000493C , 32'hFFFC1385 , 32'hFFFCA356 , 32'h00003A12 , 32'h0000FB04 , 32'h0001A554 , 32'h00019E80 , 32'h00009583 , 32'h00054B0D , 32'hFFFBCBE5 , 32'hFFFF8424 , 32'hFFFEDE7E , 32'hFFF7FAE5 , 32'h00081CBC , 32'h00002988 , 32'h00034932 , 32'h00059C0B , 32'hFFFDBF7A , 32'hFFFC7A87 , 32'hFFFC8347} , 
{32'h0003F06C , 32'h00011407 , 32'h0004B9B4 , 32'h00005C43 , 32'hFFFF6891 , 32'hFFFDF325 , 32'hFFFB9A59 , 32'h00018481 , 32'hFFF844F1 , 32'hFFFC4248 , 32'hFFFF11E2 , 32'hFFFA0E74 , 32'h0002281F , 32'h0000F83E , 32'hFFFEEF4D , 32'hFFFE81A7 , 32'hFFFED056 , 32'hFFFA1BCB , 32'hFFFC2849 , 32'h000095EA , 32'hFFFD8324 , 32'h00075D2B , 32'h000065A9 , 32'h0003538D , 32'hFFF67A8B , 32'h00017AC3 , 32'h0001951C , 32'hFFFEC630 , 32'hFFFDB843 , 32'h0003C8C9 , 32'hFFFF272E , 32'h0000B888 , 32'h000094BF , 32'h0002996B , 32'h0003643D , 32'h000417B7 , 32'hFFFF4754} , 
{32'h00051F7A , 32'h0000854F , 32'h00019CB6 , 32'hFFFA4DF3 , 32'h0001F0AF , 32'hFFFD72BB , 32'h0002F9D8 , 32'h0000AA00 , 32'h0004C362 , 32'h00051967 , 32'hFFFF36B8 , 32'hFFFD1AA0 , 32'hFFFCDBEE , 32'hFFFDD40B , 32'h0000FAE6 , 32'hFFFC26D0 , 32'h00057FF3 , 32'hFFFD3E1E , 32'h000469D3 , 32'hFFFE8D9B , 32'hFFFFE487 , 32'hFFFCC466 , 32'h000291F8 , 32'h0000F433 , 32'hFFFD2586 , 32'hFFF52396 , 32'hFFFBAD19 , 32'hFFFFFC85 , 32'h0000B156 , 32'h0004A3AB , 32'hFFFAB460 , 32'h0001C25C , 32'hFFFF772B , 32'h0000FDC6 , 32'hFFFB46ED , 32'hFFFB74BC , 32'h0001C49F} , 
{32'h00085FE3 , 32'hFFFF5184 , 32'h00023D7D , 32'hFFFEBEBA , 32'h0005E349 , 32'hFFFF0EBE , 32'hFFFF8E60 , 32'hFFFD264F , 32'hFFFFACCC , 32'h00020CD7 , 32'hFFFED32C , 32'h0002ACA4 , 32'hFFFB2EDA , 32'h00031E8D , 32'h000037DE , 32'hFFFEE676 , 32'hFFFC6642 , 32'h0004275A , 32'hFFFCA83B , 32'hFFFEA6C3 , 32'h00020C5C , 32'hFFFE7164 , 32'hFFFFBA05 , 32'hFFFF8386 , 32'h0002A154 , 32'h00005CDF , 32'hFFFC249B , 32'hFFFF8141 , 32'hFFFBD751 , 32'h00037962 , 32'h0001C3A8 , 32'h00019916 , 32'h0003A94A , 32'h0005A673 , 32'h0001A530 , 32'h000014EE , 32'hFFFEEB01} , 
{32'hFFFBCF94 , 32'hFFFF9339 , 32'h00011B09 , 32'hFFFBD3A6 , 32'hFFFFAAAB , 32'hFFF9FAFF , 32'hFFFC8B15 , 32'hFFFD0965 , 32'hFFFD1750 , 32'h00011172 , 32'hFFFDBE29 , 32'h00020408 , 32'h00024686 , 32'hFFFD430F , 32'h0002D57A , 32'hFFFF0DD5 , 32'hFFFCF6C8 , 32'h0003EA58 , 32'hFFFD6019 , 32'h0000CA52 , 32'h000027FE , 32'hFFFEBE52 , 32'hFFFD2EEA , 32'h0001BDD2 , 32'h000128D4 , 32'h000110A4 , 32'hFFFD2A4C , 32'hFFFB6EEA , 32'hFFFC15AF , 32'hFFF9AB68 , 32'h000511E4 , 32'hFFFE0F3E , 32'h00014A6B , 32'hFFFAEC79 , 32'h00061A99 , 32'hFFFFDE8A , 32'hFFFBCE4E} , 
{32'h00068830 , 32'h00044089 , 32'hFFFAB777 , 32'h000294F3 , 32'hFFFDB18F , 32'hFFF8DED3 , 32'h0000552A , 32'hFFFE3F58 , 32'hFFF779C3 , 32'hFFF9BE65 , 32'h000C9AEA , 32'h0002BA54 , 32'h00001AC8 , 32'hFFFBD77E , 32'h000438DB , 32'h00080B48 , 32'hFFFEA45D , 32'h0004DFC4 , 32'hFFFAF7D6 , 32'hFFFA6640 , 32'h00065010 , 32'h00027FFF , 32'hFFFF1C66 , 32'hFFFB28E1 , 32'hFFFC964E , 32'h000B0269 , 32'hFFFA0FAB , 32'h0006208D , 32'h000025AC , 32'h000066CB , 32'h00032A61 , 32'h0004BFF0 , 32'hFFFF4622 , 32'hFFF9F916 , 32'h0009791A , 32'hFFFAF4A8 , 32'h0005E695} , 
{32'hFFCBBD52 , 32'h028986E0 , 32'hFA166EB0 , 32'hFAB97328 , 32'hF8622830 , 32'hFAEF9A58 , 32'h02F37750 , 32'h07625320 , 32'h030EF004 , 32'h0B8FE4F0 , 32'h006DD6D2 , 32'h031B1688 , 32'hF4B526F0 , 32'h065DD5B0 , 32'hFA1288A8 , 32'hFF151328 , 32'h07172528 , 32'h063B5BB8 , 32'hF7771810 , 32'h09309780 , 32'hFD52D6F8 , 32'hEA684800 , 32'hFE4ADD14 , 32'h03C16EA8 , 32'h03280BF8 , 32'h12526360 , 32'hF4092CA0 , 32'hFE14BDC4 , 32'h05C48BB8 , 32'h03B8A7FC , 32'h05023DC0 , 32'h041F4240 , 32'h09D42CF0 , 32'h0535B118 , 32'hFCC11608 , 32'hF9D970E0 , 32'hFD56C5F8} , 
{32'h033391B0 , 32'hFF000586 , 32'hFACAB860 , 32'h030838EC , 32'hFDA67F90 , 32'hFDA17020 , 32'h03AD342C , 32'h0266A5C8 , 32'hFA71F0F0 , 32'h08CC0380 , 32'hF0BD2ED0 , 32'hFD3FBD44 , 32'hFEEB4DF0 , 32'h039C0DE0 , 32'h07AFF480 , 32'hFD67FF44 , 32'hFE991E50 , 32'h0DB17D80 , 32'hFA505438 , 32'h0659F978 , 32'hFEA4AA80 , 32'hE9A4AEA0 , 32'h01F28B50 , 32'hF888B3D8 , 32'hFE963368 , 32'h02756FC0 , 32'h01DBC970 , 32'hFE8BBBCC , 32'h04BD4708 , 32'hF5178FD0 , 32'hFD46F9BC , 32'hFF585EBA , 32'hFDDF78E8 , 32'h10AC16A0 , 32'hFE3339C8 , 32'hF2B18240 , 32'hF8DB4210} , 
{32'hFCFBB548 , 32'hFF8F1DB0 , 32'h179E9020 , 32'hF5D36D80 , 32'hEEE2CDC0 , 32'h0741E028 , 32'h19B3B520 , 32'hF94A42C0 , 32'hE830F280 , 32'h0FF44100 , 32'hF12AA460 , 32'hF78C5750 , 32'h04A34FB0 , 32'hF9D84018 , 32'hFEC48874 , 32'h093A9860 , 32'hEDCCF240 , 32'h152DEAE0 , 32'h0179463C , 32'h0FB154C0 , 32'hF92B8D58 , 32'h01713584 , 32'hF8453088 , 32'hE2D4DB80 , 32'h02682520 , 32'hEFEE5540 , 32'hF0B886E0 , 32'hF2182600 , 32'hF1588AC0 , 32'h09983D80 , 32'hF7588530 , 32'h12E538A0 , 32'hFF812747 , 32'h08CD7CF0 , 32'h08DFA9B0 , 32'hF8B70840 , 32'h007D2D07} , 
{32'h03BC3D70 , 32'h095E9FB0 , 32'h07ADEFF0 , 32'hFDFAB288 , 32'h0C4930C0 , 32'hFC54BAEC , 32'hFBAFFD68 , 32'hF9F1B4A8 , 32'hFA3EAC68 , 32'h032490A4 , 32'hFE03404C , 32'h0C9BF220 , 32'h044929E0 , 32'h03754BBC , 32'hFDC4FDC4 , 32'h03C75470 , 32'hF629C4A0 , 32'h09A04D60 , 32'hFDD01A28 , 32'h090F29D0 , 32'hFE7A6B04 , 32'h0365C394 , 32'hF86A2848 , 32'h0A5C0390 , 32'h0E283940 , 32'hFB79CE08 , 32'h01DEC618 , 32'hF75EFB90 , 32'h09AB4D50 , 32'hFED318E8 , 32'hFF48068A , 32'h0B9BC610 , 32'hFB4FF5F0 , 32'hF894B6D0 , 32'h02C21624 , 32'h0A90A190 , 32'hF3B371E0} , 
{32'h07083BF0 , 32'hFF022D4F , 32'h055B2F20 , 32'h03B12C18 , 32'hFEAA18F4 , 32'hFD72C660 , 32'h0614FA70 , 32'h08D786E0 , 32'h054D6930 , 32'h01621F38 , 32'hFA8181B8 , 32'h0028658E , 32'hFEFC6D20 , 32'h00F56E6F , 32'hEB1677C0 , 32'h0B529B10 , 32'hF97E56F8 , 32'h10039EA0 , 32'h07C38270 , 32'h0080B645 , 32'h067467C8 , 32'h00547764 , 32'hFC4DC3B8 , 32'hFEBAA4C4 , 32'h0702D6A0 , 32'hF8F415E0 , 32'h046417C8 , 32'h09B45A90 , 32'hF937CD50 , 32'h056D63C0 , 32'h067ADB58 , 32'h00884844 , 32'hFDD8FEE4 , 32'h0404E5F8 , 32'hF92CE7A8 , 32'h00ECF0F2 , 32'hF7FCA6A0} , 
{32'h056F6BA8 , 32'h08F41800 , 32'h1A4D0D00 , 32'hF44E8BE0 , 32'hFACE0D60 , 32'hF6185D40 , 32'h07FDA8A8 , 32'hFE1278BC , 32'hF9A53300 , 32'hFC11DDE8 , 32'hF88FBD18 , 32'h05555D48 , 32'h0E5C3900 , 32'hFED180EC , 32'hE64211A0 , 32'hFC53E850 , 32'hEF2BBC00 , 32'h21AB9300 , 32'h0AC35D00 , 32'h049F23D0 , 32'h128A9E00 , 32'hF7F9D360 , 32'h02B18144 , 32'hF3587480 , 32'hE4C58020 , 32'h1603D9E0 , 32'h0A0261D0 , 32'h016D4310 , 32'h007C4085 , 32'hFF7C9933 , 32'hFC83D86C , 32'hF74DE110 , 32'hD7902300 , 32'h190F7560 , 32'h00C5E58B , 32'hE9FEC900 , 32'hF8823228} , 
{32'h0A5E9520 , 32'h101A2F80 , 32'h0EF97C30 , 32'h07199910 , 32'hE61E9900 , 32'hFF057754 , 32'hF813A418 , 32'hFD9E714C , 32'hFFBCB537 , 32'hFD885208 , 32'hFBBE47E8 , 32'h08E27DE0 , 32'h04305958 , 32'hFF977BB4 , 32'hECC5A7C0 , 32'h0829CE60 , 32'hFA68F7C0 , 32'h0D867150 , 32'hFB0C1AB8 , 32'hF83A7D60 , 32'h011D5558 , 32'h09912300 , 32'hF5C86B10 , 32'hF54C5C40 , 32'hF8D97768 , 32'hFCBD6228 , 32'h00AF8784 , 32'hFCF26BEC , 32'h0031ACF4 , 32'hF2DC6850 , 32'h0131E634 , 32'h0287F834 , 32'hF46CAA70 , 32'h15744E80 , 32'h05F9C6D0 , 32'h03DB19DC , 32'hF9F305C0} , 
{32'h0CAB91F0 , 32'h0F23B290 , 32'h0F5690F0 , 32'hF6FDEB10 , 32'hF1F3D820 , 32'hF3901A40 , 32'hFCA9CB24 , 32'hFE183FEC , 32'hFACA4A70 , 32'hEAA27820 , 32'h03D9DE00 , 32'h040D9E28 , 32'h08BE8710 , 32'hF7B0D340 , 32'hED212800 , 32'h074D0560 , 32'hF4D51AB0 , 32'h08EC1ED0 , 32'hF83BED38 , 32'hF8031788 , 32'h0C548440 , 32'h0118C52C , 32'h0E71C000 , 32'hF396B350 , 32'hE8E82F20 , 32'h0A8C12D0 , 32'h0CFD6DE0 , 32'hFE464B88 , 32'h0C65BE10 , 32'hED5FDEE0 , 32'h1278EF60 , 32'hF3A1A380 , 32'hEEDB4C80 , 32'h08C46310 , 32'h07C2C378 , 32'hFDE083FC , 32'hFAA921E0} , 
{32'h0AE04250 , 32'h128A20E0 , 32'h00C2A866 , 32'hF1A9E710 , 32'h048D64E0 , 32'hF38244F0 , 32'h05815D08 , 32'h07A3C550 , 32'hFBE50CB0 , 32'hF37DE130 , 32'hFB0DE000 , 32'h05634FB8 , 32'h000AD838 , 32'hF7CE3180 , 32'hEAAE16C0 , 32'h0B255D30 , 32'hFB9AC1A8 , 32'h0287CF60 , 32'hF7F23180 , 32'h0021F903 , 32'h0AC24690 , 32'h04B03BF0 , 32'hFDD597B4 , 32'hFEE2DFD8 , 32'h01A3A0CC , 32'h027EF714 , 32'hFE011CF8 , 32'h0B49E290 , 32'h189E7420 , 32'hFB4268A0 , 32'h09F7F840 , 32'hFD61AB9C , 32'h07C3A7A8 , 32'h0193F354 , 32'hFB9027C8 , 32'hFDBDE72C , 32'hFDB2A45C} , 
{32'h08172180 , 32'h1671DDA0 , 32'hFFC55297 , 32'hE92DA240 , 32'hF7D4A9D0 , 32'hFDAE5AEC , 32'h09AF2030 , 32'h067308C8 , 32'hFD7615B0 , 32'h0122F05C , 32'h03010144 , 32'hFE5AC2F8 , 32'h0750C3D8 , 32'h0A98F250 , 32'hF379AEA0 , 32'h1452CE80 , 32'h08D89880 , 32'hEC770440 , 32'hF953A8B8 , 32'hFF6A8D08 , 32'h05B2E9D8 , 32'hFFFF9655 , 32'h0170AC40 , 32'h0FFCA3E0 , 32'hFF01A1EF , 32'hF3424E50 , 32'hF539DFB0 , 32'h00A711CB , 32'hFE57DD14 , 32'hFE989D60 , 32'h065CCA78 , 32'h021F9EBC , 32'h00C3CC40 , 32'hF9FEC808 , 32'h035286A0 , 32'h0085014F , 32'h06677768} , 
{32'h0B305D60 , 32'h1039AC60 , 32'h01863AFC , 32'hEFDCAA40 , 32'h06022C18 , 32'h074F2AF0 , 32'h0033A044 , 32'hF914C830 , 32'h0537DAF8 , 32'h012666D0 , 32'h0F425590 , 32'hFB8EDC68 , 32'h0446ED88 , 32'h020DA298 , 32'hD7AD9D80 , 32'h0F578240 , 32'h035249B8 , 32'hFF1BAF13 , 32'hEE427AE0 , 32'hFFB37D4F , 32'hF7D82460 , 32'hF0882150 , 32'hE9947700 , 32'hFEDD4F5C , 32'hF1B08870 , 32'hF3532FA0 , 32'h013F3C8C , 32'hFAB1AD38 , 32'h035EB244 , 32'hEE7A2BA0 , 32'h07AD2240 , 32'hF6AA21F0 , 32'hF9238C78 , 32'hFDF4DC34 , 32'h034C3A2C , 32'hFBFBDF08 , 32'h0ED10560} , 
{32'hFEC7C330 , 32'h1A665640 , 32'h0406CDD8 , 32'hDD39DBC0 , 32'h07205758 , 32'hFFF6AE5C , 32'h0A146B70 , 32'h05F9B038 , 32'hF7A958B0 , 32'h01B8C1A0 , 32'h10F8DE20 , 32'hDEFE8500 , 32'h0C9CCB10 , 32'h05B49E10 , 32'hF1FF2E50 , 32'hFDB8C8D0 , 32'h0E976B60 , 32'hF28F83F0 , 32'hFDEAFFE8 , 32'hFD234420 , 32'hFFAA174E , 32'hF528C150 , 32'hFE254E08 , 32'hF0CAA6D0 , 32'hF5E9C240 , 32'hFF548D56 , 32'hF1B9E9D0 , 32'h04BA7950 , 32'hFFEFC87B , 32'h06705870 , 32'hFB141378 , 32'hF62B9250 , 32'hFE9B6ED4 , 32'hFD91851C , 32'hFB4D1F70 , 32'hF2144C90 , 32'hFE3B0080} , 
{32'h077607F0 , 32'h0E2729F0 , 32'h022FAC38 , 32'hE78878A0 , 32'h05A20808 , 32'h081885D0 , 32'h0B4BB690 , 32'h0046F546 , 32'h047FC788 , 32'h0424EAA0 , 32'h11B3B420 , 32'hF48590B0 , 32'hEFC42C40 , 32'h0153C444 , 32'h0E3E6EF0 , 32'hFDCA2A34 , 32'h143AA5C0 , 32'h119EAC60 , 32'hFA52EF68 , 32'h18ACBC80 , 32'hF80EDCF8 , 32'hFEA425B8 , 32'hFDD397E4 , 32'hF8B4F1C8 , 32'hFF8F157C , 32'hEBEDF6E0 , 32'h013CCBC0 , 32'h12A2FF80 , 32'h03822A40 , 32'hFE79AB3C , 32'hF82D8BA8 , 32'h049D2688 , 32'hF7954460 , 32'hF6981FA0 , 32'h0D3D60A0 , 32'hFF2C1C23 , 32'h0E07C620} , 
{32'h0DBE6D10 , 32'h2EE0D340 , 32'hEF2B4DE0 , 32'hDAC42500 , 32'hF231CCC0 , 32'h0DD18B40 , 32'h2F0CF780 , 32'h295E0AC0 , 32'h0AA408E0 , 32'hEDBFB960 , 32'h1DC328A0 , 32'hFC706EBC , 32'hEB513900 , 32'h008A1499 , 32'h041AC260 , 32'h097BD380 , 32'h1BAE2B00 , 32'h1B1ABDC0 , 32'h00903B08 , 32'h1F97E660 , 32'hDB4C4300 , 32'hFC93EE00 , 32'h1BCE0720 , 32'hED9558E0 , 32'hF78D0700 , 32'h0221976C , 32'h0D286790 , 32'h1789AB80 , 32'hFD8DC5F4 , 32'h09A4B590 , 32'hE9056A00 , 32'hFFC709B6 , 32'hFF1F700B , 32'h033A33F4 , 32'h085AA0A0 , 32'hEF543E40 , 32'h064B8690} , 
{32'hFAE02248 , 32'h1F0EAAA0 , 32'h02C3B448 , 32'h011DFC6C , 32'h09B35210 , 32'h051D77A0 , 32'hFACE0EE8 , 32'h0D19DFB0 , 32'hF9B405A8 , 32'h0143E6F4 , 32'hFFAC7125 , 32'hFFAE0E7C , 32'hFE1119F0 , 32'h1060D3E0 , 32'hF7AFBE80 , 32'h07879550 , 32'h0BE92D50 , 32'hFBC0F000 , 32'h15780D00 , 32'h120BA4A0 , 32'hF8A090F8 , 32'hF996E0A8 , 32'h105EEC80 , 32'hF75B8800 , 32'hF3A07A60 , 32'h0B68F970 , 32'h079F4E68 , 32'hF5189190 , 32'hEBA5C940 , 32'h02F4F20C , 32'hF427B7D0 , 32'hFDE9A2E0 , 32'h05663FC0 , 32'h04ECA1D0 , 32'h0AB01240 , 32'hF6FDD280 , 32'h1454AE00} , 
{32'hFE5F91F8 , 32'hFF3B9642 , 32'hFC6D9674 , 32'h0320CFFC , 32'h052FAFF8 , 32'hFDA998D4 , 32'h0955F4C0 , 32'h03BD7DEC , 32'hFBF31080 , 32'hFF9A7B5E , 32'h052CD958 , 32'hFD2507B0 , 32'h00FD90E9 , 32'h0A8C0C30 , 32'h03F8D938 , 32'hFA51D4A0 , 32'hF8ADA480 , 32'h0BA86E00 , 32'h0B8D7810 , 32'hFB51F140 , 32'h095138C0 , 32'hF45029B0 , 32'hF8F183A8 , 32'h0B783380 , 32'hFB8679A0 , 32'hF3A109F0 , 32'h040E1C60 , 32'h0059E077 , 32'h05128628 , 32'h05E6F788 , 32'hFE05F4CC , 32'h029A6768 , 32'h00423E4B , 32'hFDCFEFE8 , 32'hFEDB0694 , 32'h01EDCD0C , 32'hFA73A638} , 
{32'h004ECAD2 , 32'hFD45D458 , 32'h00DCE29E , 32'h015CA32C , 32'hFFDCE45E , 32'hFE92DF70 , 32'h01F0AF68 , 32'h0210E4AC , 32'h00E4628D , 32'hFFA20F09 , 32'h01FEDD04 , 32'h031BAEF0 , 32'hFEE473E8 , 32'h0237EE70 , 32'h019C097C , 32'hFE149E3C , 32'hFD3307FC , 32'h0268FDB8 , 32'hFC5A3A80 , 32'h0009C68C , 32'h014482E4 , 32'hFE6208D4 , 32'hFCC41660 , 32'h025E4644 , 32'hFF93B64B , 32'hFC8D0B04 , 32'hFF67E6AD , 32'hFEF63CAC , 32'h01FE0514 , 32'h001D051B , 32'h0094E529 , 32'h02BFA628 , 32'hFC826278 , 32'hFF4DC806 , 32'h028B53D0 , 32'hFED63C00 , 32'hFF800D5F} , 
{32'h0109EBE8 , 32'hFDA6C648 , 32'h033E76AC , 32'h00B2C6A7 , 32'h04A03538 , 32'hFEC07DCC , 32'h01A6F078 , 32'h03631EDC , 32'h01A1BF9C , 32'h04AFD5B8 , 32'h0519A290 , 32'h062DE2F8 , 32'h01837D1C , 32'h08057D40 , 32'h08B03700 , 32'hF4177BF0 , 32'hFCCBD380 , 32'h095FE5D0 , 32'h028B4180 , 32'h0061078E , 32'h0718A070 , 32'hF14ABE70 , 32'hF96E0320 , 32'h0233F014 , 32'hF47162F0 , 32'hF6900580 , 32'hFEAF8D4C , 32'hFD89FB8C , 32'h03C3A26C , 32'h03211FD0 , 32'h079AEDF8 , 32'h0D9A9610 , 32'hFD8CAF74 , 32'h009402DD , 32'h01AAD008 , 32'hFDFA80C8 , 32'hF67E2E50} , 
{32'h0063D5BC , 32'hFF7E2079 , 32'h0055C366 , 32'h00E458FE , 32'h0053DC36 , 32'h00153257 , 32'h0080BB6C , 32'h001A3300 , 32'h00266990 , 32'hFE9EFB4C , 32'h0043901E , 32'h00894139 , 32'h00D7D72F , 32'h0055AC4F , 32'hFFB9306D , 32'h006B3EB1 , 32'hFFE0774C , 32'h00548DFB , 32'hFF015E54 , 32'hFF58C231 , 32'h00025B04 , 32'hFE283E28 , 32'h00E408A6 , 32'hFF3E89F5 , 32'h00004B7A , 32'h0049DD14 , 32'hFFD5EBCB , 32'hFFED2D97 , 32'hFF704779 , 32'h0033FCAE , 32'h00AC2D41 , 32'h008D06C2 , 32'hFF8D8453 , 32'hFF7FD24A , 32'h0026D646 , 32'hFFC7FCEE , 32'h000AA210} , 
{32'hFFFF5150 , 32'h000098ED , 32'hFFFFF111 , 32'hFFFE7D16 , 32'hFFFF5F88 , 32'hFFFE0FE7 , 32'hFFFEDF5B , 32'hFFFF4773 , 32'hFFF6C491 , 32'hFFFDE8EF , 32'h00031026 , 32'hFFFCBD1C , 32'hFFFE90DD , 32'hFFFD654D , 32'h0000C69F , 32'h00012AB9 , 32'h00019FF7 , 32'h00042797 , 32'h00010DBC , 32'hFFFF9933 , 32'hFFFDF472 , 32'hFFFE2419 , 32'h0000A3F5 , 32'hFFFF2303 , 32'hFFFFF0D8 , 32'h0006EA19 , 32'hFFFF0DC2 , 32'h000067E1 , 32'h000050CB , 32'h0002F93B , 32'hFFFF7BCB , 32'h00003A67 , 32'hFFFDF676 , 32'hFFFDA39C , 32'h00012CAF , 32'h00021ACB , 32'hFFFFAF71} , 
{32'h0000FBAF , 32'hFFFFF52F , 32'hFFFE34AA , 32'h0001CECA , 32'hFFFBF127 , 32'h00008BFE , 32'h00015A28 , 32'hFFFFB9E4 , 32'hFFFDCF9D , 32'hFFFEA83A , 32'hFFFC91FD , 32'h00050F1B , 32'hFFFDAEB1 , 32'hFFFE4AB3 , 32'h00074CB0 , 32'hFFFFB08C , 32'hFFFCAA1D , 32'h00004D9C , 32'h00017503 , 32'hFFFAC975 , 32'h0000FDE7 , 32'h0003CB59 , 32'hFFFCD1E1 , 32'h000078A4 , 32'h0002D2B3 , 32'hFFFFE0F7 , 32'hFFFD1E2B , 32'h0004A7C8 , 32'hFFFB11AC , 32'hFFFA6A68 , 32'hFFFB4849 , 32'hFFFF5A78 , 32'h000131B9 , 32'h00003904 , 32'h00025AAA , 32'hFFFF0F6B , 32'h00035B36} , 
{32'h000119C9 , 32'h00014AAE , 32'h0001A14F , 32'h00047AD7 , 32'h000008CC , 32'h0000B9E4 , 32'hFFFA0B86 , 32'hFFFE9E1D , 32'hFFFB6750 , 32'hFFFBFF36 , 32'h0002A3F8 , 32'hFFFF5912 , 32'h0001E6EE , 32'hFFFE909F , 32'h00012D6B , 32'h00012916 , 32'h0002AF42 , 32'h0002F65E , 32'hFFFE943F , 32'hFFFD5B09 , 32'h000292D8 , 32'hFFF6BE78 , 32'hFFFEFD1B , 32'h00034D48 , 32'h0005D918 , 32'h0000CBDC , 32'h0003D3E0 , 32'h000437D8 , 32'h00031560 , 32'h00044616 , 32'h00033F60 , 32'h0000C139 , 32'hFFFCE18B , 32'hFFFEC57E , 32'hFFFDF492 , 32'hFFFC1CAE , 32'hFFFF39FA} , 
{32'hFFFA7DE6 , 32'h0000F3EA , 32'h000392F4 , 32'hFFFD5E82 , 32'hFFFEBD14 , 32'hFFFF5616 , 32'h00025E57 , 32'hFFFDE6C1 , 32'hFFFE3FAF , 32'h0001F762 , 32'h00022D28 , 32'hFFFE5477 , 32'h0000AE27 , 32'hFFFF12B2 , 32'h00021B64 , 32'h00003CDE , 32'hFFFFF052 , 32'h00047E5B , 32'h0000B71A , 32'hFFFDD91F , 32'hFFF9CAB3 , 32'hFFFFF68F , 32'h0000ABA6 , 32'hFFFF40F3 , 32'h0001FDC1 , 32'h0005704F , 32'hFFFF9CF3 , 32'hFFFEE774 , 32'h000132E1 , 32'hFFFEF3B5 , 32'hFFFDEEE0 , 32'h000225B9 , 32'h000274CA , 32'h00011B2C , 32'hFFFB7F44 , 32'h0002C612 , 32'h0003B5E5} , 
{32'hFFFFED73 , 32'hFFFE671F , 32'hFFFCE851 , 32'h0000DF97 , 32'hFFFEFDF6 , 32'h0000FE8A , 32'hFFFF8D5D , 32'hFFFC5C65 , 32'h0002A425 , 32'h00009C50 , 32'h00012439 , 32'hFFFE999F , 32'hFFFC4FE7 , 32'hFFFE0612 , 32'h00023263 , 32'h0004455B , 32'hFFFD5902 , 32'h0003447F , 32'h0003DFF9 , 32'h0003E0CB , 32'h0000D212 , 32'h0000500D , 32'h00014D17 , 32'h0003EA9C , 32'hFFFB617C , 32'hFFFF2A49 , 32'h00051812 , 32'hFFFE0485 , 32'h00008D7C , 32'h0001CD83 , 32'h00031D72 , 32'h00056002 , 32'h00024302 , 32'h0002AC80 , 32'hFFFD902B , 32'h0002EB53 , 32'hFFFF534E} , 
{32'hFFFBE992 , 32'h0002AB56 , 32'hFFFF357E , 32'hFFFDC22D , 32'h0000E1F6 , 32'hFFFDA790 , 32'hFFFF5239 , 32'h00044E93 , 32'h000048EC , 32'h00017E31 , 32'h00043D0A , 32'h0001425A , 32'h000559BF , 32'hFFFC58B1 , 32'hFFFDD642 , 32'hFFFF150D , 32'h0000500B , 32'h0000F407 , 32'hFFFDEB5E , 32'hFFFF4713 , 32'hFFFA3C33 , 32'h00028A18 , 32'hFFFEFAE8 , 32'hFFFC1A76 , 32'h00010CC8 , 32'h00011429 , 32'hFFFC636A , 32'h0002DD4C , 32'h000636B7 , 32'h00026826 , 32'hFFFDAA4E , 32'hFFFDCD26 , 32'hFFFEA2D6 , 32'h000380F9 , 32'h00018D2E , 32'hFFFE4BD4 , 32'hFFFA307B} , 
{32'h00005DD3 , 32'hFFFF8456 , 32'h00051BA9 , 32'h0005ECDB , 32'hFFFD8CC2 , 32'hFFFD733B , 32'hFFFD3294 , 32'h00004A02 , 32'hFFFCBFF4 , 32'h0005BCC1 , 32'hFFFE7CD5 , 32'h0000FBF2 , 32'h00013F54 , 32'hFFFEEB5A , 32'hFFFD0E29 , 32'h0006EF79 , 32'h0005BFE1 , 32'h0006161E , 32'hFFFB180E , 32'h00033447 , 32'h00043F36 , 32'hFFFF51C5 , 32'hFFFF0F3C , 32'h0002817F , 32'h0002E178 , 32'hFFFB8D6C , 32'h00017E57 , 32'hFFFF2187 , 32'h0000804C , 32'h0002947F , 32'h0001B9E6 , 32'hFFFEBC23 , 32'h0003F34C , 32'h00055F1F , 32'h0001137E , 32'hFFFBA3C3 , 32'h00016B94} , 
{32'hFFFF1969 , 32'hFFFFE291 , 32'hFFFCA030 , 32'hFFFD6C7E , 32'hFFFD0B93 , 32'hFFFBACC3 , 32'hFFFBBE98 , 32'hFFFC3AA6 , 32'hFFFFA9FE , 32'hFFFC8EDE , 32'h0004AD7F , 32'hFFFE4741 , 32'h00005802 , 32'hFFFC4278 , 32'h00019F38 , 32'h0000D3FC , 32'hFFFAE967 , 32'h0002B9A2 , 32'h00020155 , 32'hFFFF219A , 32'hFFFF20EC , 32'h00057721 , 32'hFFFA156E , 32'h0000131A , 32'h00049E2C , 32'h00021B38 , 32'h0000D480 , 32'h0003C797 , 32'h00043EEF , 32'hFFFD79E5 , 32'h0004D63E , 32'h00017AD0 , 32'hFFFB783E , 32'hFFFF628A , 32'hFFFF5D80 , 32'hFFFF3E4B , 32'h00069D5B} , 
{32'h0004E24F , 32'h000A39E1 , 32'hFFFB042E , 32'h0006C506 , 32'h0004A4FF , 32'hFFF8C088 , 32'h00016E5C , 32'h000501BF , 32'hFFF34CAD , 32'hFFFA28E2 , 32'h000DDF37 , 32'h0009836F , 32'hFFFFBC8E , 32'hFFFCAA9E , 32'h000928E4 , 32'h000A8DFA , 32'hFFFBBF79 , 32'h000472FE , 32'hFFF56005 , 32'hFFF995CF , 32'h0007DD22 , 32'h0000A01A , 32'hFFFB8C8D , 32'hFFF6FA7D , 32'hFFF8C945 , 32'h000E452E , 32'hFFF8B20A , 32'h0009C355 , 32'h00008DC0 , 32'h000008F1 , 32'h0002C981 , 32'h00093B62 , 32'hFFFD7A60 , 32'hFFFD87D9 , 32'h00092275 , 32'hFFFE94E1 , 32'h00041272} , 
{32'hFCF438D4 , 32'hFE1A0058 , 32'h01102238 , 32'hFAB67F88 , 32'hFD60C3D0 , 32'h01C98BFC , 32'hF8D0BA28 , 32'h01025620 , 32'hFFAAD1AC , 32'hFE36B5B4 , 32'hFEF6344C , 32'hFFE69E16 , 32'hFFAACA80 , 32'h029D076C , 32'hFE4B1E48 , 32'h006DA44F , 32'h00A8E5CC , 32'h026FA11C , 32'h00A4CFB3 , 32'h004F3196 , 32'hFF3C0ADA , 32'hFF5C537B , 32'h00F745B4 , 32'h00880CF8 , 32'h008BAB0D , 32'hFDC47450 , 32'h02129130 , 32'hFF80898A , 32'hFF74D8CF , 32'hFF69DB86 , 32'h009E5656 , 32'hFEA08DE4 , 32'h0274D4E8 , 32'hFE442184 , 32'hFED67ECC , 32'hFD68C074 , 32'hFE1D518C} , 
{32'h013700EC , 32'hF8684390 , 32'hFE016ADC , 32'hFB7A6F98 , 32'hF96AE728 , 32'hFC42C700 , 32'h0179857C , 32'hF734D370 , 32'h009CFB81 , 32'hFBF94F48 , 32'hF9E65E28 , 32'h08514150 , 32'h03C2D8DC , 32'hFE7CE590 , 32'h0206A7F8 , 32'hFD107174 , 32'hEF49C1E0 , 32'hF8ECBE90 , 32'h051A6B88 , 32'h052AFBA8 , 32'h0C6D4960 , 32'hFF9BE46D , 32'h044D6D70 , 32'hFF55F1DA , 32'hFE768D20 , 32'hFCA6E7D4 , 32'h0096DDD7 , 32'h00373596 , 32'h002FECE2 , 32'hECC2B020 , 32'h01ED1F48 , 32'h01B24C74 , 32'h0D947CA0 , 32'hF6A88FA0 , 32'h00305EEB , 32'h081ECE10 , 32'h05F39390} , 
{32'h08915B60 , 32'h0B72ADD0 , 32'h06CF7BB0 , 32'hFA6E8728 , 32'hF1DFE5B0 , 32'h02E89B3C , 32'h07C76588 , 32'h0E7CC100 , 32'h0C2B8D00 , 32'hF8FF64A8 , 32'h0AE58B40 , 32'h04578690 , 32'hFBB55450 , 32'hEBE66D60 , 32'h0CCF98B0 , 32'h0F17F980 , 32'h0CAD3310 , 32'h13857C20 , 32'hF2EB74A0 , 32'h13D800E0 , 32'h09389860 , 32'h085BB1C0 , 32'h0ECE9940 , 32'hF7F29DC0 , 32'hFD1824CC , 32'h0A4DA3B0 , 32'h0BBCE930 , 32'hF18CE9D0 , 32'hF208B550 , 32'hE8939AE0 , 32'h18F78980 , 32'hFA4ADE48 , 32'h0218EF38 , 32'h021EB530 , 32'h0537F3C8 , 32'hFF1752D9 , 32'hF857EFD0} , 
{32'h03B23F5C , 32'hEF582B40 , 32'h036A0A48 , 32'hF134A790 , 32'hE87DAA40 , 32'hE83A7C00 , 32'h06ECFE80 , 32'hF8075C60 , 32'hFF85A99D , 32'h0C324E80 , 32'hF7B5FB80 , 32'hF055C5B0 , 32'h0B9F47A0 , 32'h07516450 , 32'h130183E0 , 32'h0DDE9870 , 32'hF57DFE50 , 32'h1A2B9980 , 32'hF1C07B30 , 32'hF7401130 , 32'h0EC9C4E0 , 32'h0CE80700 , 32'h0D382A80 , 32'h023677B0 , 32'h082719D0 , 32'hEE148820 , 32'hE5F24DA0 , 32'hED0D9700 , 32'h0E0C7840 , 32'h0DE9D2D0 , 32'h0043EA80 , 32'hFC8364F0 , 32'hFEF22FF0 , 32'hF21E49F0 , 32'h02810328 , 32'hF101E5C0 , 32'hF40A16C0} , 
{32'h069AB008 , 32'h01DA6690 , 32'h00392605 , 32'h00F76491 , 32'hFE815B6C , 32'hF5E63300 , 32'h035202A0 , 32'hFCD991B4 , 32'hF8173508 , 32'hFBBB1C88 , 32'hFD65C8E0 , 32'h0EDE45D0 , 32'hF8F892D0 , 32'hFDDD8DC4 , 32'hF028BF80 , 32'h0699D6E8 , 32'hF33F1110 , 32'h13575420 , 32'hFA5FABD0 , 32'h07C2DD90 , 32'hFCDA1D28 , 32'h022F84BC , 32'hF8CCDFB0 , 32'hFB220DC0 , 32'hFFC95061 , 32'hFF26C821 , 32'h0B59BAF0 , 32'hF5E1CC20 , 32'hF769CE80 , 32'h0BAB5090 , 32'hFE622B54 , 32'h0040333C , 32'hF9A8CDA8 , 32'hFF32CD37 , 32'h065A22D8 , 32'hFFC97E5A , 32'hF928EB40} , 
{32'h031C8F14 , 32'h0FBE2D70 , 32'h0B0E1DF0 , 32'h04315220 , 32'hEE592BE0 , 32'hF750BCD0 , 32'hFAB64778 , 32'hFF10D741 , 32'h0065B3A1 , 32'hFAFB14B8 , 32'hFFD51617 , 32'hFF835A3A , 32'h01BBB600 , 32'hFF545174 , 32'hF84F4AE0 , 32'h015535F8 , 32'hFA8E6980 , 32'h08479A90 , 32'hFB61F148 , 32'hF9E59380 , 32'h0658CAC8 , 32'h00396F4C , 32'h0C11EF50 , 32'hF2A16610 , 32'hFE22831C , 32'hFFCACC88 , 32'h02946574 , 32'h061D0CD8 , 32'h0D04E340 , 32'hF4C2EB40 , 32'h08C564A0 , 32'hFA29D628 , 32'hF9AEEF70 , 32'h00F53411 , 32'h043EAD60 , 32'h0529BA30 , 32'h01C2C578} , 
{32'h0D12F5E0 , 32'h1EF08900 , 32'h1C2B90C0 , 32'hF4A23B70 , 32'hEE667CE0 , 32'hEFE2A0C0 , 32'hFF56FC63 , 32'h0422A958 , 32'hECF72480 , 32'hFAF61CC0 , 32'hFAE06838 , 32'hEC335180 , 32'h0F14F3F0 , 32'h02924B08 , 32'hEFAF6A20 , 32'h052333F8 , 32'hFAF088B0 , 32'h10D14680 , 32'h110202E0 , 32'h0114B530 , 32'h03166858 , 32'hFED8A53C , 32'h0AB371E0 , 32'hEDB93FE0 , 32'hFD6209EC , 32'hF672E840 , 32'hEDA398A0 , 32'hF93ED820 , 32'h0AACE880 , 32'hEE5342A0 , 32'h09C3A4D0 , 32'h02B70650 , 32'h0660FEC8 , 32'h08806610 , 32'h062842B8 , 32'h09A9DA90 , 32'h0E70B6E0} , 
{32'h05339400 , 32'h0A8CF530 , 32'h09DA9300 , 32'hF57FD190 , 32'hF0FFA4F0 , 32'hED3F5CC0 , 32'hFFE05C75 , 32'h0B8CB6C0 , 32'hF2575E80 , 32'h061C0FF8 , 32'h062BD4A0 , 32'hFA7D7088 , 32'h10D46500 , 32'h0D83BF60 , 32'hFBEF2698 , 32'h1647ED60 , 32'hEA98C0E0 , 32'h08F62160 , 32'hF7C1D610 , 32'h0194ECB4 , 32'h01B54A90 , 32'h023B9E94 , 32'h0201E414 , 32'hF0A89FA0 , 32'hF4D6FD10 , 32'h004740C4 , 32'hE0E62D20 , 32'hFF16D96B , 32'h10B5B260 , 32'hEFE46900 , 32'hFFF6013A , 32'hFB944B98 , 32'hFC91C324 , 32'hF76DD9A0 , 32'hFC2D4914 , 32'hF4A6DF20 , 32'hF8F58E90} , 
{32'h0114600C , 32'h09CCF440 , 32'h0636D3D0 , 32'hEE8F7140 , 32'hF9239540 , 32'hF4C381C0 , 32'h040DAEE8 , 32'hFB3C4910 , 32'hF5E885E0 , 32'hF7D67C30 , 32'h007AC14C , 32'hFEDDD7A4 , 32'h04C1CBE0 , 32'hF59C3B50 , 32'hFEB05AB8 , 32'h021850A0 , 32'h0753A690 , 32'hF4908CC0 , 32'hEFDEF040 , 32'hFF36E03D , 32'h02EEBF18 , 32'hF8844AA8 , 32'h07FEA8F0 , 32'hF6ADB960 , 32'hF4DD1110 , 32'h0D11E2B0 , 32'h052A5290 , 32'h04C7A4C8 , 32'h13F5A6A0 , 32'hF2D3D780 , 32'h05397EE8 , 32'hF4881130 , 32'hF893E060 , 32'hFE261BF8 , 32'h0EE75550 , 32'h03B88FE8 , 32'hFE4D41F0} , 
{32'h0994AA50 , 32'h10156400 , 32'h05529060 , 32'hF0779220 , 32'hFA8F6BE8 , 32'hFE11B5A4 , 32'h0A0C4430 , 32'hFC9DD00C , 32'hEF4A6080 , 32'hF0FD1BE0 , 32'hF7FD5960 , 32'hF5820960 , 32'hFE68211C , 32'h04821650 , 32'hFF3B3053 , 32'h1D334300 , 32'h0866EB20 , 32'hF2FC4E60 , 32'h0295A690 , 32'h02094050 , 32'hF68EB470 , 32'hF3E969C0 , 32'h0B8C40E0 , 32'hEF301C40 , 32'hF4D1B150 , 32'h0267513C , 32'hE48539E0 , 32'hF26AA260 , 32'h06340AE8 , 32'hFD62FD9C , 32'hFE31B810 , 32'hFF9CA8B7 , 32'h01B132D4 , 32'hEDE01180 , 32'h03E6B3AC , 32'h0F51DE70 , 32'h0E6FA180} , 
{32'h07BC1C00 , 32'h143B9520 , 32'h04C45060 , 32'hEC268E60 , 32'h079F0720 , 32'hFD7B5000 , 32'h07F40F58 , 32'h003DC411 , 32'hED64E3E0 , 32'hFA283F50 , 32'h011CBD60 , 32'hF7276DF0 , 32'h03A9CBD0 , 32'hFE73548C , 32'hEA988260 , 32'h16971C60 , 32'h08309460 , 32'h01BD2F0C , 32'h095AE430 , 32'h107F6420 , 32'hEA18CAE0 , 32'hF4D1CCF0 , 32'hF17BF460 , 32'hE6740200 , 32'hFE604FA8 , 32'hFF442407 , 32'hE06E59E0 , 32'hEED36EE0 , 32'hF9817060 , 32'hF7C22EA0 , 32'h0184AF7C , 32'h0324DE30 , 32'h08233350 , 32'hF8E870B8 , 32'hFF9474F5 , 32'h02E5E01C , 32'h13998940} , 
{32'h0D9FB1E0 , 32'h1C9507A0 , 32'hF9034920 , 32'hE383B640 , 32'hF68E2080 , 32'h0E8928D0 , 32'h1C6EB2E0 , 32'h19B59480 , 32'h0910B8D0 , 32'hED95DF60 , 32'h171C3980 , 32'hED103CA0 , 32'hFBB96570 , 32'h068BB000 , 32'hFA8ECE10 , 32'h22963400 , 32'h25E14740 , 32'h000D272B , 32'hE7AC7FC0 , 32'h12562180 , 32'hE40E26A0 , 32'h129F11C0 , 32'hF8EADB48 , 32'h1150F0A0 , 32'h1916CDA0 , 32'hFF1ED586 , 32'h0EAB50B0 , 32'h0D30CEA0 , 32'hFBF9CF58 , 32'hEB185140 , 32'h04F945B0 , 32'hE5963120 , 32'hF69FFD80 , 32'h004CF667 , 32'h17F82960 , 32'hF84C4688 , 32'h2295CB00} , 
{32'h180C5D40 , 32'h239EFC40 , 32'hFF6DC907 , 32'hE7CEC320 , 32'h03A30834 , 32'hF468EA70 , 32'h1A1AC420 , 32'h016E8568 , 32'hE99B9440 , 32'h0A510D00 , 32'hFD209424 , 32'hD83F0B00 , 32'h0531D198 , 32'h13C6FFA0 , 32'hF68DCBC0 , 32'h1703B420 , 32'h04163AB8 , 32'hED971D60 , 32'hFECD1B04 , 32'h1CD52D60 , 32'hEF6FDE80 , 32'hEE95C300 , 32'hFE414B64 , 32'hE6E8FCE0 , 32'h0D5AAFC0 , 32'hFB2AE4D0 , 32'hEFF3EDE0 , 32'h0B668630 , 32'h0682D090 , 32'h12F9C120 , 32'h058919D0 , 32'h019BEBA4 , 32'h05D61DF0 , 32'hFEC85554 , 32'h12C2CEC0 , 32'hE4FF5200 , 32'hFB284F08} , 
{32'hFF09AD37 , 32'h14FD4AA0 , 32'hEFE29BC0 , 32'hEBDE8C60 , 32'hEE6BFF40 , 32'h010AEEAC , 32'h0AA44C10 , 32'h0BC7B070 , 32'hFD7B1888 , 32'hFA001760 , 32'hF93C40C0 , 32'hFE9A8AE4 , 32'hF7A5E8E0 , 32'h0505F330 , 32'hFD910EEC , 32'h024B67A4 , 32'h0189A494 , 32'hF19D3BF0 , 32'hFA9769C0 , 32'hF9C96518 , 32'h104F4B00 , 32'hEDC2FE00 , 32'hFE332934 , 32'h01F41D18 , 32'h15040340 , 32'h1B08D900 , 32'hFCD44C00 , 32'hF33584E0 , 32'hF4FF3300 , 32'h06005B18 , 32'hFDEB9670 , 32'h03567408 , 32'h11730880 , 32'h06D5F7F0 , 32'h0180659C , 32'h00DEA6A6 , 32'hFB9819A8} , 
{32'hF8D6BC70 , 32'h03CDDE68 , 32'hFB5E5028 , 32'h0D0BAF70 , 32'hFDB496EC , 32'h05253750 , 32'hFE0BC78C , 32'h105F3800 , 32'h0052365B , 32'hF6E97E80 , 32'hFE97A044 , 32'h06434710 , 32'hF9D00AF0 , 32'h0B3F3300 , 32'h036CBDA8 , 32'h07DB3230 , 32'h00B408D2 , 32'hFB8955B8 , 32'h197F3DE0 , 32'hFB8A58B8 , 32'h0A641030 , 32'hF8F71AC0 , 32'h091E0860 , 32'hFCA91070 , 32'h1020F840 , 32'h0EE03C00 , 32'hFBCE54D8 , 32'hF30E7830 , 32'hFCDF79C0 , 32'h0A7F5130 , 32'hF91C07C0 , 32'hEBAD6640 , 32'h066EBF10 , 32'h0FC70E90 , 32'hFF55ECD1 , 32'hFC58BE10 , 32'h096B2020} , 
{32'h0366CA24 , 32'h0ADBD230 , 32'h032BDDE8 , 32'hF62B6AA0 , 32'hFF0C538D , 32'h00E22D17 , 32'h037C1C24 , 32'h00360B06 , 32'hF5C90450 , 32'h01E672D4 , 32'hFCDD80B0 , 32'hF4764DE0 , 32'h05D4B9B8 , 32'h037A49DC , 32'hFD8C0570 , 32'h0A30FF00 , 32'hFCF38A88 , 32'hF9DC3F70 , 32'h021BB2A0 , 32'h08656730 , 32'hFBDFD3D8 , 32'hFA26D998 , 32'hFDA99A84 , 32'hF93A4FC0 , 32'h007F2AF5 , 32'hF6B31DF0 , 32'hF5FA9370 , 32'hFC0816D0 , 32'hF9948358 , 32'hFD54A918 , 32'hFE5B452C , 32'h03C8DEDC , 32'h01E3562C , 32'hF9856EE8 , 32'h042490D8 , 32'hF97918D8 , 32'h03BC8888} , 
{32'hFC09427C , 32'hFCB7D560 , 32'h013F3454 , 32'hFF9D4344 , 32'h01D6C0B8 , 32'h003ACCF5 , 32'h0598E0D8 , 32'h02202A64 , 32'hF581DBB0 , 32'hFCDF11AC , 32'h0A925330 , 32'h0B6F4640 , 32'h01C96A9C , 32'h0EB971D0 , 32'h01AAB794 , 32'hFA0B0B08 , 32'hF5772F60 , 32'h029E629C , 32'h176B4A20 , 32'hFB6F03D0 , 32'hFC42D940 , 32'hF41B3A90 , 32'hFE7BF894 , 32'h11798020 , 32'h16755A20 , 32'h04A1FDD8 , 32'h0145C3F0 , 32'hFEBFCEF0 , 32'h0CF93070 , 32'h07D29990 , 32'hF7B725B0 , 32'hED27D840 , 32'hF0BB1FA0 , 32'h0058E760 , 32'h1E086CE0 , 32'h0BC61FA0 , 32'hFEA1595C} , 
{32'h00CD76E1 , 32'hFEF40624 , 32'hFFBFED59 , 32'h0075708E , 32'hFFF7B9DE , 32'hFFD5E8F6 , 32'h004EFB10 , 32'h003BB36B , 32'hFF2AC300 , 32'hFDEE5150 , 32'h00A2AB24 , 32'h0152A1B8 , 32'h0190CECC , 32'h001D919E , 32'h00C24254 , 32'h00C1170D , 32'hFFE1D286 , 32'h0075AAE7 , 32'hFE5B7DD4 , 32'hFF71B630 , 32'hFFE03D6C , 32'hFE60BAC4 , 32'hFFF8C38C , 32'hFF124278 , 32'hFF8638CC , 32'h00EC9E08 , 32'hFF85D129 , 32'hFFC52979 , 32'hFF9B06C4 , 32'h0047A1D9 , 32'hFFE8E1CB , 32'h00A607AD , 32'hFFB40FF4 , 32'hFF8C530C , 32'hFF83BFE2 , 32'hFF4F20D0 , 32'h009DEC74} , 
{32'hFCCF74FC , 32'hFE27ABE0 , 32'h01B6D57C , 32'hFF0DF115 , 32'h0185559C , 32'h0040645D , 32'h039229FC , 32'h00C553E5 , 32'hF8580D30 , 32'hFEAEC450 , 32'h0806D970 , 32'h07F4A8E8 , 32'h00D86705 , 32'h0ACC6DE0 , 32'h010276E4 , 32'hFB7487E0 , 32'hF90919B0 , 32'h0175A2C8 , 32'h124B14A0 , 32'hFCFC20B8 , 32'hFD6406C0 , 32'hF913C7F8 , 32'hFEE29F9C , 32'h0D478960 , 32'h11AD9920 , 32'h03524B98 , 32'h0170CC90 , 32'hFF98B06E , 32'h09D60AF0 , 32'h055B4EA8 , 32'hF9E38950 , 32'hF1BAC600 , 32'hF56CB510 , 32'h00B7AE91 , 32'h16268B20 , 32'h09A3E970 , 32'hFE1B30A0} , 
{32'hFFFFA895 , 32'hFFFC7631 , 32'h0000D93C , 32'hFFFDE2D7 , 32'hFFFC92B7 , 32'hFFFEE1C9 , 32'hFFFDB019 , 32'h00010C81 , 32'h0003136B , 32'h0001E8CF , 32'h0000E095 , 32'h00042EA1 , 32'hFFFBC2DC , 32'hFFFB763D , 32'hFFFB856B , 32'hFFFDD2C5 , 32'h0000E4A4 , 32'hFFFFF84F , 32'h00020A26 , 32'h000283E7 , 32'h000365C7 , 32'hFFFFDC22 , 32'hFFFEBFDA , 32'hFFFD6E9D , 32'hFFFD090A , 32'hFFF778AD , 32'h00026C6A , 32'hFFFC0412 , 32'hFFFC6E2B , 32'hFFFEE5A8 , 32'hFFF9740D , 32'h00001062 , 32'h00001C22 , 32'h0001D04A , 32'h0000928D , 32'h0001B51F , 32'h00046CB2} , 
{32'h00063ED7 , 32'h0002C715 , 32'hFFFFE71B , 32'h000478E3 , 32'h000197E7 , 32'hFFFB2F1D , 32'hFFFF9433 , 32'h00014ACA , 32'h00031991 , 32'hFFFD5DE4 , 32'h00008ADF , 32'h00023B7B , 32'h0001E487 , 32'hFFFF2077 , 32'h000339B1 , 32'hFFF90715 , 32'hFFFFF636 , 32'hFFFEBC08 , 32'hFFFE59CD , 32'hFFFE1F90 , 32'hFFFA51DB , 32'h0004AE68 , 32'hFFFFFFCD , 32'h0003E07B , 32'hFFFF5FF8 , 32'h00037E92 , 32'hFFFB0D3F , 32'hFFFE40E3 , 32'hFFFCBB4F , 32'h000278EC , 32'hFFFBDAE3 , 32'hFFFC6E7A , 32'h00001E6A , 32'hFFFEDA85 , 32'h000048F9 , 32'h00013950 , 32'h0001BD8E} , 
{32'h0001176A , 32'h0001E2EB , 32'h00015E5E , 32'hFFFF2021 , 32'h0001EE87 , 32'h00020B46 , 32'hFFFE0510 , 32'hFFFC7BDE , 32'h00019F42 , 32'hFFFD1D10 , 32'h0005BE69 , 32'h000422E6 , 32'h00006549 , 32'h000736B9 , 32'hFFFE582A , 32'hFFFC4C00 , 32'hFFF920DF , 32'h000483A5 , 32'hFFFDB2E2 , 32'h00000F82 , 32'hFFFB8D20 , 32'h0001AE01 , 32'hFFFC9112 , 32'hFFF621B2 , 32'h0003923D , 32'h0001FA04 , 32'h000A78AE , 32'h000109F2 , 32'h0001D7F2 , 32'hFFFE68F0 , 32'h00000431 , 32'h00024F7B , 32'h00045E28 , 32'hFFFEF4A8 , 32'hFFFF6D38 , 32'h00037DCE , 32'hFFFCFACA} , 
{32'h0001C33C , 32'h00022C42 , 32'h0002B83C , 32'h00054B8C , 32'hFFFF7EB5 , 32'h00023615 , 32'hFFFF74AE , 32'hFFFA75FE , 32'hFFFDD1C6 , 32'h0000DE5C , 32'h00008E3E , 32'hFFFF0AAE , 32'h0000BEF3 , 32'h0001B237 , 32'hFFFF436F , 32'hFFFE1091 , 32'hFFFDFAA3 , 32'hFFFD09FB , 32'h00024894 , 32'h00013D93 , 32'hFFFFC54C , 32'h0000AC80 , 32'h00000F41 , 32'hFFFD40BE , 32'hFFFE316E , 32'h00030675 , 32'h0001B515 , 32'h00016A6F , 32'h000896FB , 32'hFFFF3660 , 32'h0003BEF1 , 32'hFFFEB62C , 32'hFFFE1175 , 32'hFFFFAC5E , 32'h0001AD75 , 32'hFFFA14E0 , 32'hFFFA49AE} , 
{32'h0002F7F2 , 32'h00000A82 , 32'hFFFF7921 , 32'h000300C7 , 32'hFFFA3216 , 32'hFFFF5537 , 32'hFFFBA241 , 32'h00008304 , 32'h0001450A , 32'h0002906D , 32'h00018514 , 32'h000221CB , 32'h0001EE66 , 32'hFFFA8409 , 32'hFFFF8E6D , 32'h000346BB , 32'hFFFEAA2B , 32'hFFFFCEBC , 32'hFFF9981F , 32'hFFFFA1E4 , 32'h00004240 , 32'h00045063 , 32'h0000F4DF , 32'h0001580E , 32'hFFFA807D , 32'h00007BEE , 32'h00049E95 , 32'h00020AB8 , 32'h0000262D , 32'h000164DF , 32'h0001A8D6 , 32'hFFFEAEF4 , 32'hFFFD9883 , 32'h00077EC2 , 32'hFFFF5F31 , 32'h0006B2E1 , 32'hFFFD1A01} , 
{32'h0002245E , 32'hFFFD9163 , 32'hFFFD3DF9 , 32'hFFFBD381 , 32'h0002B014 , 32'h00029B5F , 32'h0004BFBC , 32'h0002BC2A , 32'hFFFE2119 , 32'hFFFABC96 , 32'hFFF70862 , 32'hFFFFEF8D , 32'hFFFD801B , 32'hFFFC5835 , 32'hFFFF23AB , 32'h00018215 , 32'h00024546 , 32'hFFF95B18 , 32'hFFFEA747 , 32'h00002D26 , 32'h0001A8A7 , 32'hFFFF1B65 , 32'hFFFEA802 , 32'hFFFCCDBF , 32'hFFFE62D2 , 32'hFFFFD133 , 32'h00009BC8 , 32'h00006863 , 32'hFFFD3E1B , 32'hFFFE991E , 32'h0004102C , 32'hFFFE2367 , 32'hFFFD7340 , 32'hFFFF9A99 , 32'h000003AE , 32'hFFFF2799 , 32'hFFFC98C0} , 
{32'hFFFE9DAC , 32'hFFFCAA23 , 32'hFFFC14C6 , 32'h0000E06D , 32'hFFFE744B , 32'h00034CB3 , 32'hFFFFD21F , 32'h00027AE0 , 32'h000085D6 , 32'hFFFC3AB5 , 32'hFFFF9EB4 , 32'h00000B0E , 32'hFFFC0B64 , 32'hFFFFCBBE , 32'hFFFD820F , 32'hFFFEC01F , 32'hFFFDAA7C , 32'h0008BDBE , 32'h00020071 , 32'hFFFD22FB , 32'h0002636E , 32'hFFFFA4F1 , 32'hFFFEB15E , 32'hFFFEB588 , 32'h00021395 , 32'h00002D33 , 32'hFFFBE841 , 32'h00004DCA , 32'hFFFF7C17 , 32'hFFFFBEA8 , 32'hFFFAE006 , 32'h000205E5 , 32'h00038548 , 32'hFFFE5B3E , 32'hFFFDA3FA , 32'hFFFE9FCB , 32'h00046C28} , 
{32'hFFF71A2A , 32'hFFFF9527 , 32'h0000BF76 , 32'h000104AC , 32'h0001DC97 , 32'h000164F0 , 32'hFFFF07EA , 32'hFFFDD8D6 , 32'hFFFCC790 , 32'h0000259D , 32'h000335C7 , 32'hFFFFF778 , 32'hFFFF0A4C , 32'h00026734 , 32'h0001A3C9 , 32'h0001101C , 32'h0000CDF2 , 32'hFFFE832E , 32'hFFFF5077 , 32'h00042080 , 32'h0006E4A9 , 32'hFFFD7D07 , 32'hFFFFD448 , 32'hFFFCC4FD , 32'hFFFF91BF , 32'hFFFC6ECA , 32'hFFFDF355 , 32'hFFFC8AD0 , 32'hFFFF223E , 32'hFFFFF96E , 32'hFFFF1302 , 32'h00021CBC , 32'h0005B61B , 32'hFFFD6118 , 32'hFFFED31A , 32'h00008779 , 32'hFFFD5B1D} , 
{32'h019F7284 , 32'hFF786997 , 32'h00ADCC2E , 32'hFF3AB458 , 32'hFFBE21CC , 32'h00F0FF49 , 32'hFF4E607F , 32'h0019E206 , 32'h01A7F670 , 32'h015F6400 , 32'hFFBED2B1 , 32'hFDE636D0 , 32'h02F87CDC , 32'h0083CBE6 , 32'hFFDD0BBE , 32'hFF0E2B38 , 32'h0047F424 , 32'hFED78994 , 32'hFEC085CC , 32'h012341B4 , 32'h039832A4 , 32'h02E2DC28 , 32'hFD3148A4 , 32'h033F8138 , 32'hFC570F9C , 32'h014DFDA8 , 32'hFFA1BA8E , 32'hFAAA1938 , 32'hFD883F58 , 32'hFD4309D0 , 32'hFDF730CC , 32'h06558A78 , 32'hFE3ABCD4 , 32'hFF15F695 , 32'h04118670 , 32'hFEFBA9E4 , 32'hFDCA73A4} , 
{32'h00743074 , 32'hFD83290C , 32'hFF8EAFBE , 32'hFC67BB60 , 32'hFC9FE8C0 , 32'hFFE9BC80 , 32'h0127F6D8 , 32'hFD396710 , 32'h00C9A379 , 32'hFBEB3910 , 32'hFD0CAC10 , 32'hFF8E44FA , 32'h0099F887 , 32'hFF107B6B , 32'hFFF97982 , 32'h00A90C1B , 32'hFD42C2CC , 32'hF9BDE560 , 32'h029D34EC , 32'h006E6B20 , 32'h03A7B784 , 32'h00FADD9F , 32'h05AA3AD0 , 32'hFBDC1120 , 32'h01885D3C , 32'h033F1874 , 32'hFEAF5C60 , 32'h038F96AC , 32'h0206A57C , 32'hFA5DBB50 , 32'hFCB6F230 , 32'hFFB49EF5 , 32'h0238020C , 32'hFD21AD1C , 32'h02A73BE8 , 32'h02FE495C , 32'hFC10B1B4} , 
{32'h06CDDB18 , 32'hFDCBFF64 , 32'h02EF2EE8 , 32'hFCACEF00 , 32'hFED34928 , 32'h03E939A0 , 32'hFD193980 , 32'h005FBA67 , 32'h06F32998 , 32'h058DD1A0 , 32'hFEB9EBE0 , 32'hF72D8BF0 , 32'h0C7D2B60 , 32'h02219E44 , 32'hFF7F4232 , 32'hFC002000 , 32'h00FD7D69 , 32'hFB7039C8 , 32'hFADDFD68 , 32'h04D277A0 , 32'h0F07B410 , 32'h0BC6B0E0 , 32'hF430A160 , 32'h0D62A6C0 , 32'hF0EC3E90 , 32'h0599E9F8 , 32'hFE68BA04 , 32'hE9BD8BC0 , 32'hF5DDD880 , 32'hF47BC800 , 32'hF79B7B60 , 32'h1A4AE940 , 32'hF8BE1278 , 32'hFC447F68 , 32'h10DDFF20 , 32'hFBBF1F28 , 32'hF6C9C3D0} , 
{32'h0DC1E760 , 32'h143BA120 , 32'h20CB2180 , 32'hFE8C88BC , 32'hD912D280 , 32'h0A0E4920 , 32'h07522310 , 32'h0768AF98 , 32'h0031FE5B , 32'h0B1B1170 , 32'hF4C777B0 , 32'hF0C49060 , 32'h17F0A7A0 , 32'h0221874C , 32'hFB38A9F8 , 32'h04D78CF0 , 32'h0B7ADBF0 , 32'h008C690D , 32'hF93A1DB8 , 32'hF6530E30 , 32'h133C4F20 , 32'h0358B218 , 32'hEFDAD7A0 , 32'h18649DC0 , 32'hF5CF61F0 , 32'hFDC8E0A4 , 32'hF6600970 , 32'hFE469894 , 32'hF042F710 , 32'hEF404E60 , 32'hF6431BD0 , 32'h10AA7760 , 32'hE9600FC0 , 32'h02765770 , 32'h03DBEDF4 , 32'h05C3D5C8 , 32'hEE332680} , 
{32'h022C5CEC , 32'h199EF880 , 32'h21E09800 , 32'hFE9E21B4 , 32'hF201AC60 , 32'hF7CDA170 , 32'h0B254420 , 32'hF959C728 , 32'h08906A20 , 32'h063823D8 , 32'hE5882BC0 , 32'h0E22B750 , 32'h0AEE44C0 , 32'h02C7CA80 , 32'h077BFAE0 , 32'h098132A0 , 32'hF74826C0 , 32'h0F5BED30 , 32'hFF875AD9 , 32'hF53DBA30 , 32'h0AE8F7B0 , 32'hFC72AF38 , 32'hF7838450 , 32'h039EB088 , 32'h00AF46FE , 32'hF4E848E0 , 32'hF95DEDA8 , 32'hFB580C50 , 32'h0BA77750 , 32'hF0D0C580 , 32'hF9FCF108 , 32'h06C54DC8 , 32'h07EBC9F0 , 32'hFFEC2AE0 , 32'hFA5BAE18 , 32'h0C1C2340 , 32'hFF5FC5C9} , 
{32'h05232F98 , 32'h0CFD28B0 , 32'h1817EA60 , 32'hF735E800 , 32'hF333CBE0 , 32'hFFA78D9F , 32'h0F3BE3B0 , 32'h05A26698 , 32'hF79E6F50 , 32'h05A7D650 , 32'hE9F7F1A0 , 32'hFAFAEBF0 , 32'h010EA948 , 32'h03C0A6B0 , 32'h0A35DF30 , 32'h0136D3A4 , 32'hF44F6900 , 32'h08DC4E20 , 32'hF7739300 , 32'hFD485068 , 32'h000BFBB0 , 32'hF4AE3590 , 32'h01ABC9A0 , 32'hFC28BF90 , 32'h0A086CF0 , 32'hFAFDAAD8 , 32'hF8155A18 , 32'h049D5758 , 32'h0CFE6EF0 , 32'hF7894F90 , 32'hF4329140 , 32'h05FBA568 , 32'hF4E46B20 , 32'h11571A40 , 32'hF24C9380 , 32'h002BC349 , 32'hF315ED20} , 
{32'h0BD5E3B0 , 32'h0260DB28 , 32'h0FE92820 , 32'hF4E617A0 , 32'hF15728E0 , 32'h0DD2BEB0 , 32'h1F713F20 , 32'h06BAC690 , 32'h08530780 , 32'hFF85C728 , 32'h0A2377A0 , 32'hFD4583A4 , 32'h0F69C590 , 32'hEF3AE820 , 32'h0C3BC6B0 , 32'h0EC26350 , 32'h09487D80 , 32'h20CAF240 , 32'h02D56C8C , 32'h07AD2CD8 , 32'hF13D22B0 , 32'hFEF8DFBC , 32'h09F32F60 , 32'h0F27D3C0 , 32'h0248E220 , 32'hF93BEC70 , 32'h0B280D90 , 32'h09ABE8B0 , 32'hF9F45600 , 32'hF65CCC30 , 32'h024EA758 , 32'h028361C8 , 32'hFF5AA338 , 32'h07BDAE58 , 32'hFEDE6564 , 32'h04BBE378 , 32'hE5DFE1A0} , 
{32'h09B9FB50 , 32'h10514900 , 32'h046713B0 , 32'h029AC2E4 , 32'hE86486E0 , 32'hEFBBBFE0 , 32'h085CED40 , 32'h0E0CC490 , 32'hFA2B0B80 , 32'hF49E2810 , 32'h15315220 , 32'h0B99B2B0 , 32'h01217790 , 32'hF9C354F0 , 32'hFB23E538 , 32'h06C26090 , 32'h02795AF0 , 32'h164AD800 , 32'h00C66EAA , 32'h08DA4900 , 32'h024F5F74 , 32'h0F1954A0 , 32'h0683E258 , 32'h03550514 , 32'hFC60F61C , 32'h07B8DDB0 , 32'h0EEC42B0 , 32'hF808C8A8 , 32'hFECF1F10 , 32'hDCF50300 , 32'h0D8FD620 , 32'hF00FC2F0 , 32'hF9016100 , 32'hFFA9F5B3 , 32'h00A406CF , 32'hFE385500 , 32'hED4231A0} , 
{32'h0235950C , 32'h1D3CAA80 , 32'h08843CC0 , 32'hDC730580 , 32'hF08AC240 , 32'h01863934 , 32'h09C7AF50 , 32'hFBC5A350 , 32'hECEF3AC0 , 32'h030BD23C , 32'h10CF8A40 , 32'hF2F313B0 , 32'h18E98D40 , 32'h116EFCC0 , 32'h089D04C0 , 32'h0A5A4370 , 32'h0C538E40 , 32'hE19AE940 , 32'hDB853F80 , 32'hEBC30380 , 32'h1FA04360 , 32'hEF061820 , 32'hF9751960 , 32'h12EC0180 , 32'h086681E0 , 32'hF4388AF0 , 32'hF9049E58 , 32'hF816FC00 , 32'hF7501490 , 32'hF0E7F0A0 , 32'hFD24F744 , 32'hF87AE890 , 32'hEE79CFC0 , 32'h00F56E3B , 32'h05367F80 , 32'hF88D75B0 , 32'h01C3B2D8} , 
{32'h0AD97790 , 32'h164C2880 , 32'h02245118 , 32'hDB3FC900 , 32'hFAAFBBC8 , 32'h051AE6B0 , 32'h0C9AD2D0 , 32'hFDCA5120 , 32'hEF4B49A0 , 32'h2127F8C0 , 32'h06444B70 , 32'hE84C6800 , 32'h1A7CC4E0 , 32'hF646BB00 , 32'hF5D06870 , 32'h3081E180 , 32'hF35ECEE0 , 32'hEF747180 , 32'hF9D4F8A0 , 32'h0CC38A80 , 32'hF5717200 , 32'hEBCE0500 , 32'h05E3AC78 , 32'hF72F87C0 , 32'h16008B60 , 32'hEFA4C520 , 32'hF65BE280 , 32'hF3231980 , 32'h014CBC90 , 32'hEAF7D040 , 32'h00F70905 , 32'h08DC6220 , 32'hFBADDB78 , 32'hFEEE7D70 , 32'h06D0E968 , 32'h0157D520 , 32'hFE0F5710} , 
{32'hFDE505B4 , 32'h11913280 , 32'h0B19A250 , 32'hF3BDA820 , 32'hEEB41AE0 , 32'hFCB8FB20 , 32'h1AEDAEE0 , 32'h06EC0C40 , 32'h0C90EC30 , 32'hFAD488E8 , 32'h02F7620C , 32'hF5DFC510 , 32'h092C8B00 , 32'h00EE8894 , 32'h0F208F50 , 32'h1831DCE0 , 32'h04195930 , 32'h08275CA0 , 32'h00E533EB , 32'h05A00400 , 32'hFDDC2798 , 32'hFC6286F0 , 32'h031FDA84 , 32'h02E646F0 , 32'h019E4208 , 32'hEEC21C00 , 32'h15EF6AA0 , 32'h05BABB10 , 32'h15949780 , 32'hEA104020 , 32'hF8336458 , 32'hF2E9C5F0 , 32'h0BE45910 , 32'h04AD5898 , 32'h075BBE48 , 32'hFEFD5AE8 , 32'hF991D6E8} , 
{32'h063DD598 , 32'h09CC4570 , 32'hFCB1C0BC , 32'hF582C460 , 32'h00FDBF95 , 32'h01D11E40 , 32'h088505B0 , 32'h093A1BD0 , 32'h07A71B80 , 32'hF5258E20 , 32'h07F46E18 , 32'hFFA1FA34 , 32'hFCED2724 , 32'hFBDFA400 , 32'hF7D30350 , 32'h0A212090 , 32'h064AFA50 , 32'h05E54F50 , 32'hF79D6110 , 32'h027BBF40 , 32'hF54DB330 , 32'h03ACD764 , 32'h032BA0E0 , 32'hF5E71640 , 32'h04A28230 , 32'hEDB58520 , 32'h063790B0 , 32'h060655B8 , 32'h0C80AED0 , 32'h05038720 , 32'hF51D6730 , 32'hF9C265C8 , 32'h00CECDD1 , 32'h0A62DFA0 , 32'h06C943A0 , 32'hFCF37FB4 , 32'h1B9B3FE0} , 
{32'h0AAE6060 , 32'h1A60E420 , 32'hF28D62F0 , 32'hDA07A140 , 32'h0FB69C00 , 32'h1199F860 , 32'hFEA0C4FC , 32'h1DA4FC00 , 32'h0F2DAA30 , 32'h2D6EB380 , 32'h2B611780 , 32'hD056A380 , 32'hF1D409D0 , 32'hF991B750 , 32'hE9596980 , 32'h00944C32 , 32'h248EE7C0 , 32'hFF24EB55 , 32'h00046DA7 , 32'hF05A33C0 , 32'h004973DC , 32'hFB2F8850 , 32'hCEAD4540 , 32'h0002D8D2 , 32'h1AC506C0 , 32'h1CCC09A0 , 32'hFA536138 , 32'h017BF694 , 32'h02E30A88 , 32'h071F9870 , 32'hF59E7920 , 32'hFF4F2834 , 32'hF2179420 , 32'h0AE9E260 , 32'hF8B75C08 , 32'hF64E8D30 , 32'hF5D56D00} , 
{32'h082D5250 , 32'h0F518FF0 , 32'hF12A92A0 , 32'hFA772718 , 32'h115D65C0 , 32'h1122BDC0 , 32'h0AC5E1D0 , 32'h13C692E0 , 32'h04ECFF00 , 32'hF7436B00 , 32'h0C348F10 , 32'hE4F60D20 , 32'hF8AECE88 , 32'h0DC03F40 , 32'hD86F2400 , 32'hF3B4B230 , 32'h1E674960 , 32'h1AAC2E00 , 32'hF20440D0 , 32'hF6CBA9D0 , 32'hFB07EF50 , 32'hEFE4B6E0 , 32'hEB6C15A0 , 32'h01A8A440 , 32'h16F2DF00 , 32'h26BEDE00 , 32'hF7D38BB0 , 32'hE85BAAE0 , 32'h011CA8F4 , 32'h128DA200 , 32'hFE60CD88 , 32'hFF2531E7 , 32'h0896D650 , 32'h0D33BBD0 , 32'h01DD284C , 32'h088B8390 , 32'h01A928F8} , 
{32'h045E55E0 , 32'h075E97A0 , 32'hFB6AE418 , 32'h0648D7D8 , 32'h07292DB8 , 32'h01C6E0B0 , 32'h0E103260 , 32'h08DE5280 , 32'h02009558 , 32'hFF899B42 , 32'h05474E38 , 32'hF33BAF70 , 32'hFC226D14 , 32'hFD8E351C , 32'h01302988 , 32'h0058439B , 32'h0B5A8260 , 32'hFE4761DC , 32'hFE0E35C4 , 32'hF9442F08 , 32'hF9F44C68 , 32'hFF97CF72 , 32'hFD629FAC , 32'hFACE4BD8 , 32'h011C1720 , 32'h06FD4420 , 32'hFB35DA58 , 32'h0398D380 , 32'h06E38EB0 , 32'h0DA241A0 , 32'hF8033580 , 32'h051C50A0 , 32'hF3C715A0 , 32'h049189B8 , 32'h0046D4EB , 32'hFE226720 , 32'hF8007A28} , 
{32'hFFC6DD00 , 32'h03F1781C , 32'h0091A5E8 , 32'hFA86B250 , 32'h042D49B0 , 32'h01591DFC , 32'h0653EB70 , 32'h09E989D0 , 32'hF764F7D0 , 32'hF93099C0 , 32'h04932CC0 , 32'hFB360D48 , 32'hFE180A0C , 32'h0B7E3500 , 32'h0170C370 , 32'h02A8C354 , 32'h011CC764 , 32'hFC2F8DD4 , 32'h0D2F9F20 , 32'hFA97F4B8 , 32'hF218BD10 , 32'hF6DA70F0 , 32'hFE7CB558 , 32'h0AD6F120 , 32'h15A02C60 , 32'h08B70680 , 32'hFF84DC68 , 32'h09C6EA10 , 32'h167AFB40 , 32'h0C0C7310 , 32'hF253EA80 , 32'hF11DA8C0 , 32'hF0626F30 , 32'h05A54158 , 32'h187165E0 , 32'h03CA58D0 , 32'hF37B7970} , 
{32'hFF56265F , 32'h0075FAA7 , 32'hFEE876A8 , 32'h00FE8B27 , 32'hFFA2A531 , 32'h000EAFB3 , 32'h00A14D2E , 32'h00D193E9 , 32'h005D98FF , 32'hFFB08373 , 32'hFEEAAD18 , 32'hFF616CDE , 32'hFF129415 , 32'h007DA40E , 32'h0097BD85 , 32'h0084F88B , 32'hFE6262D4 , 32'h01187DB4 , 32'h00085AEF , 32'hFEF1F83C , 32'hFF12C621 , 32'hFEB9F500 , 32'hFF906B31 , 32'h0008188A , 32'hFEC0F66C , 32'hFF0A9CD5 , 32'hFF232CD6 , 32'hFF782062 , 32'h0096328F , 32'h0065D6EB , 32'h000A84D1 , 32'h00736F8D , 32'h00106A3B , 32'h00564879 , 32'hFF7D879D , 32'hFEDF8CB0 , 32'h003707C6} , 
{32'hFC6E9930 , 32'hFD6AFA3C , 32'h013E6B6C , 32'hFE2AD700 , 32'hFFF44981 , 32'hFD11D0E4 , 32'h02CD88F0 , 32'h04883600 , 32'hF7DAF820 , 32'hFB537C18 , 32'h048B0FC8 , 32'h0AC79570 , 32'hFFD44CC7 , 32'h0952AC20 , 32'h0353DEE4 , 32'hF94F25F8 , 32'hF6CEB690 , 32'h01A26784 , 32'h13956880 , 32'hFC72269C , 32'hFCA07D40 , 32'hF9C1AE08 , 32'hFA85E8B0 , 32'h0B5CC540 , 32'h117C40A0 , 32'h004D562E , 32'hFF2F1390 , 32'h024A9DAC , 32'h0E2589F0 , 32'h04894B98 , 32'hF34EAB80 , 32'hF0303100 , 32'hF1364280 , 32'h02995B48 , 32'h1811A380 , 32'h092791C0 , 32'hFC3AEC5C} , 
{32'hFE2FC948 , 32'hFE68B648 , 32'hFFA683AC , 32'hFEFC9D20 , 32'hFF63FE05 , 32'hFFDBE1A2 , 32'h01C83BD4 , 32'h00A0303B , 32'hFA0443C0 , 32'hFE3BE72C , 32'h03D1E948 , 32'h04A16908 , 32'h0071C5CE , 32'h0585C958 , 32'h02C9C0B8 , 32'hFE0B79B0 , 32'hFC1766A4 , 32'h00F79ACA , 32'h090CA440 , 32'hFE6B6160 , 32'hFE6C1E4C , 32'hFD212BFC , 32'hFD3D6F00 , 32'h07844960 , 32'h08E3C820 , 32'h01C85AB8 , 32'hFFA8E7C2 , 32'hFF22786F , 32'h0601A0C8 , 32'h0313AF7C , 32'hFB50C630 , 32'hF8D577C0 , 32'hFB22CFE0 , 32'h00DE05FA , 32'h0AD1A100 , 32'h04536160 , 32'hFF390D5E} , 
{32'h00662015 , 32'hFEF23F00 , 32'hFF29B7A1 , 32'hFF016CDA , 32'hFEA052D4 , 32'hFF62BBA8 , 32'hFF782E10 , 32'hFFC9DD13 , 32'hFDBD3658 , 32'hFEA6C9A4 , 32'h002E7CF1 , 32'h00B24C18 , 32'h00AD33E3 , 32'hFFE6AD69 , 32'h023E4004 , 32'h00884201 , 32'h006CAA20 , 32'h002811AF , 32'hFF816EB4 , 32'h00594F97 , 32'h000A95AB , 32'h0110DD0C , 32'hFDE470E8 , 32'h00595FBD , 32'h000E2429 , 32'h007AD6C6 , 32'hFF172C95 , 32'hFFA21DD9 , 32'h009F161C , 32'hFFF6A7F5 , 32'hFE655FB0 , 32'h0086D7FC , 32'h00B16F77 , 32'h006EC2FB , 32'hFEF58470 , 32'hFFB6F4F0 , 32'h00080F46} , 
{32'h00019B55 , 32'h00041A0E , 32'h00011CDF , 32'h0004E44B , 32'hFFFDB020 , 32'hFFFECF41 , 32'hFFFB9D8A , 32'hFFFACED8 , 32'h000020E6 , 32'hFFFDF4A3 , 32'h0006346C , 32'h0002DF3D , 32'h0001A0E3 , 32'h0001CA57 , 32'h0005D8B3 , 32'hFFFEC966 , 32'h0001F33B , 32'hFFFFDDA4 , 32'hFFFDCE73 , 32'h00028DF7 , 32'hFFFBAB0F , 32'hFFFF1376 , 32'hFFFCFC81 , 32'h000405E3 , 32'h0000381B , 32'h0003F48B , 32'h0006F10A , 32'h0003A6BB , 32'hFFFF63B3 , 32'h00024D58 , 32'h00005D29 , 32'h00018CC8 , 32'h00020998 , 32'hFFFCB562 , 32'h00018B83 , 32'hFFFE402A , 32'hFFFF4F2E} , 
{32'h0002FB7D , 32'h0000430A , 32'hFFFD730D , 32'hFFFE588F , 32'hFFF73369 , 32'h000335BD , 32'hFFFA74D7 , 32'h0002A744 , 32'h0009603B , 32'h00031F9E , 32'hFFFDD0F1 , 32'h00000BEC , 32'h00025158 , 32'hFFF9F9E5 , 32'hFFFFDAE9 , 32'h0004E55A , 32'h0003B078 , 32'h0001C486 , 32'hFFFD5693 , 32'hFFF9CDEA , 32'h0000824A , 32'hFFFE7280 , 32'hFFFCEAA5 , 32'h00035098 , 32'hFFFCE0FD , 32'h00021705 , 32'h0000D716 , 32'h00039A55 , 32'h00008D37 , 32'h0003AD6D , 32'h00015EB7 , 32'h0001E61F , 32'h00033B2C , 32'hFFFF629F , 32'hFFFFD6A7 , 32'hFFFE6C57 , 32'h0002F5BD} , 
{32'hFFFEE715 , 32'h00015B8D , 32'h00002C54 , 32'hFFFBC3A3 , 32'hFFFB486F , 32'h000017D8 , 32'hFFFD0C7E , 32'hFFFF6A3B , 32'h00085602 , 32'h0004A5B5 , 32'h000072C4 , 32'h000594FF , 32'hFFFCB5E4 , 32'h000569D5 , 32'hFFFD2AA6 , 32'h00023045 , 32'h00019022 , 32'h00007CAA , 32'h0000710B , 32'hFFFDE26C , 32'hFFFD78A0 , 32'hFFFC417F , 32'hFFFC6558 , 32'hFFFFE3A0 , 32'h00033045 , 32'h00019008 , 32'hFFFD6523 , 32'h000B4423 , 32'h0002DBA8 , 32'hFFFEF7DB , 32'hFFFE3783 , 32'hFFF5F11B , 32'h00015160 , 32'hFFFF37BA , 32'h00028E56 , 32'hFFFE6D0C , 32'h0002D3F5} , 
{32'hFFFE6C97 , 32'hFFFA5BC5 , 32'hFFFEF568 , 32'hFFFD695C , 32'h000459CB , 32'h00017A8A , 32'hFFFF38D5 , 32'hFFFE0235 , 32'h0007986F , 32'hFFFF8FAE , 32'hFFFF2174 , 32'h0001B2A7 , 32'h00060073 , 32'hFFFE15F1 , 32'hFFFDC2DF , 32'h00037E89 , 32'hFFFD500D , 32'h0003B71B , 32'h0000EFA8 , 32'h0000D682 , 32'hFFFB08E5 , 32'hFFFC568D , 32'h00036B0F , 32'h00050AEA , 32'h00021552 , 32'h00004D2D , 32'hFFFEE74E , 32'hFFFF8D93 , 32'h0001A63C , 32'h00028724 , 32'hFFFC4E96 , 32'hFFFC575B , 32'hFFFF9964 , 32'h000074C2 , 32'hFFFE7A32 , 32'hFFFA501E , 32'h0005BADE} , 
{32'h00035910 , 32'h000217A9 , 32'h0002854E , 32'h0003047C , 32'h00005FA0 , 32'hFFFF0075 , 32'hFFFAFA21 , 32'hFFFE6223 , 32'hFFFA6AB4 , 32'h00048384 , 32'hFFF9795D , 32'hFFFC8C3C , 32'hFFFD033E , 32'h00025448 , 32'hFFFDA5CE , 32'h000167A0 , 32'hFFFDB5DA , 32'h00009E83 , 32'h0002A6A6 , 32'h00000A8A , 32'hFFFC6CC6 , 32'h00025005 , 32'hFFFBF89F , 32'h0001AFC3 , 32'hFFF7144E , 32'hFFFCAAEA , 32'hFFF9859B , 32'hFFFB0458 , 32'hFFFE4046 , 32'h00061B55 , 32'hFFF7E6B5 , 32'h00013F59 , 32'hFFFF8425 , 32'hFFFB7C62 , 32'h0001F2EF , 32'hFFFF9916 , 32'hFFFE6AE5} , 
{32'hFFFEF473 , 32'hFFFFF279 , 32'hFFFBAD26 , 32'hFFFF3EBD , 32'hFFFEA845 , 32'hFFFF3E0F , 32'h00000727 , 32'h00005CC2 , 32'hFFFF85F6 , 32'hFFFFE128 , 32'h00018F31 , 32'h00036621 , 32'h00004DBC , 32'hFFFFAE13 , 32'h0000B7B2 , 32'h00020D76 , 32'h00024B4D , 32'h000104D8 , 32'h00023265 , 32'hFFFC1938 , 32'h00054616 , 32'hFFFE8C97 , 32'hFFFE9C34 , 32'hFFFEBF4F , 32'h00022BB8 , 32'h0004D8D2 , 32'hFFFDDF4C , 32'hFFF99BA0 , 32'h0000986E , 32'hFFFD8ADD , 32'hFFFD0C4E , 32'h00046545 , 32'hFFFDAF30 , 32'h00009E94 , 32'h00016C29 , 32'hFFFE1FF7 , 32'h000178DB} , 
{32'h00028601 , 32'h0000AF64 , 32'hFFFA13C7 , 32'hFFFDD724 , 32'hFFFC02C4 , 32'h00062E68 , 32'hFFFA692E , 32'h00021972 , 32'h0000A2EA , 32'h0000181B , 32'h0002020F , 32'hFFFF5BDD , 32'h00074250 , 32'hFFF88AA7 , 32'hFFFE27B5 , 32'hFFFB2E7C , 32'hFFFA4803 , 32'h0000371F , 32'h00075D04 , 32'hFFFE138B , 32'h0003AB31 , 32'hFFFF35D6 , 32'h00020112 , 32'hFFFD8E46 , 32'hFFFDCAE9 , 32'h00040FF9 , 32'hFFFC3657 , 32'h00023135 , 32'hFFFD36AD , 32'h00049176 , 32'h00036F49 , 32'h0004AB44 , 32'h00018DB9 , 32'h0004B5ED , 32'h00006425 , 32'hFFFB5F20 , 32'hFFFF7913} , 
{32'h00005B39 , 32'h0001EAFC , 32'hFFFD4059 , 32'hFFFE9A64 , 32'h00056DDE , 32'hFFFF71AF , 32'h00012B67 , 32'hFFFD2BFB , 32'hFFFC45FD , 32'h0000E688 , 32'hFFFE62AD , 32'hFFFE708E , 32'h00001C5F , 32'h000106AC , 32'h0003363C , 32'h00019357 , 32'h0002A697 , 32'h0005D898 , 32'h0003ED67 , 32'hFFFFFEB2 , 32'h0008025C , 32'hFFFDCC53 , 32'h0004D46B , 32'h00002B3B , 32'h0006F081 , 32'h00015C3B , 32'h000217D9 , 32'hFFFC6845 , 32'h0003AE11 , 32'hFFFE9CED , 32'h00051059 , 32'h0000B8DF , 32'h0005133F , 32'hFFFDF09B , 32'hFFFBADFA , 32'hFFFD1C8F , 32'h0000FC15} , 
{32'hFFFFD411 , 32'h00047670 , 32'hFFFEC2D0 , 32'hFFFEEA37 , 32'hFFFF86FB , 32'h00030056 , 32'h00013276 , 32'h00012CD5 , 32'h0002D922 , 32'hFFFCB800 , 32'hFFFE8EB3 , 32'h00049662 , 32'hFFFFF8ED , 32'hFFFDFFF4 , 32'h0006C19D , 32'h00028B3C , 32'h0001D524 , 32'h00019677 , 32'h0005F866 , 32'hFFFC6962 , 32'hFFFEC20D , 32'hFFF978E3 , 32'h00007588 , 32'hFFFE40BE , 32'h0002D34A , 32'hFFFF96BD , 32'hFFFB7DF9 , 32'hFFFC95C3 , 32'h0002EC0D , 32'h000380D5 , 32'h0001BC4E , 32'h00053FC6 , 32'hFFFBC614 , 32'hFFFF145A , 32'h0003DE08 , 32'hFFFF7509 , 32'hFFFD6AB0} , 
{32'hFD095750 , 32'hFF27A722 , 32'h026CDD40 , 32'h00C64CC6 , 32'h02C2DEEC , 32'h02CFD5F4 , 32'hFD3F4270 , 32'h011C0224 , 32'h015E68B0 , 32'h01190194 , 32'hFBC686E8 , 32'hFA533E90 , 32'hFFA402BC , 32'h00D2FDCC , 32'h0280A670 , 32'h02175594 , 32'h03EDBF18 , 32'hFD384E08 , 32'h00EE81C9 , 32'hFE346D18 , 32'h089AB9B0 , 32'hFFEFE4E4 , 32'h019F1CD8 , 32'h0125F57C , 32'h02EFF4A0 , 32'hFF3EC37D , 32'hFB0A9320 , 32'h01008834 , 32'hFE81471C , 32'hFD19B6FC , 32'h02BDEC90 , 32'h035190F4 , 32'h00A3422A , 32'h07545080 , 32'h0191C550 , 32'hFFDE5D0D , 32'h0547D920} , 
{32'h0412F9D0 , 32'hFEA56E78 , 32'h01ADF528 , 32'hFE02A2B8 , 32'hFF5A8814 , 32'h02576DE4 , 32'hFE407258 , 32'h004FD25A , 32'h042EB890 , 32'h037117B0 , 32'hFF5BD7E3 , 32'hFABBA530 , 32'h077D6580 , 32'h014E449C , 32'hFFAA548F , 32'hFDAA59FC , 32'h00ACA7B4 , 32'hFD2575A8 , 32'hFCDE8A10 , 32'h02DEE2B4 , 32'h090B7530 , 32'h07437CC0 , 32'hF8E64830 , 32'h081D7090 , 32'hF6DAEFF0 , 32'h033EE638 , 32'hFF1AF9A8 , 32'hF29FEB70 , 32'hF9DDAE28 , 32'hF9211900 , 32'hFAE94050 , 32'h0FDE9A00 , 32'hFB8C3870 , 32'hFDB906B0 , 32'h0A345140 , 32'hFD83E35C , 32'hFA6E84F0} , 
{32'h030D3B78 , 32'h0111BAE0 , 32'h00BCE2A7 , 32'hFE884D98 , 32'hFF7FCF45 , 32'h0A51F5D0 , 32'hFFF599FB , 32'hFDF2C238 , 32'h0AD87300 , 32'hFDF6CA28 , 32'hFB5C6260 , 32'hF8EF4518 , 32'h09F50870 , 32'h039E0FE8 , 32'hFE36CFD8 , 32'hFA4F1278 , 32'hFDACB5C0 , 32'hFF9D118E , 32'hFC9011F0 , 32'h057D78E0 , 32'h0A67A420 , 32'h0B470450 , 32'hF6B26510 , 32'h0C9D8370 , 32'hF7D541A0 , 32'h06A668E8 , 32'hFB2E67B8 , 32'hF4FD2910 , 32'hFCB14EB4 , 32'hFB0D4660 , 32'hFD738918 , 32'h0E6C77C0 , 32'hFDEA6E60 , 32'hFC7A9E98 , 32'h095911B0 , 32'hFB6B4750 , 32'hFA7389B8} , 
{32'h06C692C0 , 32'h0CC2BB60 , 32'h05A83F88 , 32'hF03D2E00 , 32'hFC243684 , 32'h07A342E8 , 32'hFF612AA7 , 32'h0CC86300 , 32'h0168FF00 , 32'h0A294CD0 , 32'hF7D0D0B0 , 32'hE5BA4580 , 32'h155EA0C0 , 32'h08BA9460 , 32'hFAF46DB8 , 32'h0A4E6B50 , 32'h09F78440 , 32'hE2552EC0 , 32'hED7016E0 , 32'hFFB8D880 , 32'h27A5C580 , 32'hF8597708 , 32'hF0F72390 , 32'h1F24ADA0 , 32'h05DD9960 , 32'hF5ED26D0 , 32'hF8F34B18 , 32'hF5395A20 , 32'hE9F6E980 , 32'hEE077180 , 32'hFBA0D3B0 , 32'h0DAEA930 , 32'hEBA60F20 , 32'hFED87894 , 32'h0A60CB10 , 32'hF1353F30 , 32'h01095A60} , 
{32'h0A7E0D00 , 32'h045DBD80 , 32'h04030AA8 , 32'hEBCA2640 , 32'hFC99BA38 , 32'hFD6599F0 , 32'h058F13C0 , 32'hF98AB820 , 32'hFA419120 , 32'h10791700 , 32'hFE2E1C48 , 32'hF7828280 , 32'h0BF1AFE0 , 32'hF8029398 , 32'hF3E5C3F0 , 32'h00A04949 , 32'h0959EE10 , 32'hF2E62980 , 32'hE191C600 , 32'h079F06E8 , 32'hFFFA95E9 , 32'hEEA4A100 , 32'hF47B0A60 , 32'h1976EFC0 , 32'h074A45F8 , 32'hEEFAF460 , 32'h05C19638 , 32'h12FA0580 , 32'h04609BE0 , 32'hF4266760 , 32'h02C5B114 , 32'hFEE14600 , 32'hF1618CA0 , 32'hEFDA6120 , 32'h058BFC70 , 32'hFEE3EA80 , 32'hFDBF0C44} , 
{32'h0B73D7E0 , 32'h0E90A390 , 32'h0E431630 , 32'h04D0FF38 , 32'hE5EF3CE0 , 32'hFE2BAC38 , 32'hF68CBDD0 , 32'h018F69D0 , 32'h0301E2E8 , 32'h0081E96F , 32'hFC1B1078 , 32'hF4AD9160 , 32'h0EF5D8D0 , 32'hFC4B2028 , 32'h0147FE74 , 32'hF9182258 , 32'h0088EF62 , 32'h06D17568 , 32'hFCBA37A0 , 32'hFE373C68 , 32'h0D593CE0 , 32'h0ACE2370 , 32'hFA3B4CB8 , 32'h0A6A2670 , 32'hF80E8990 , 32'h0E671540 , 32'hFDED4CB4 , 32'hEE857560 , 32'hFB2D03D8 , 32'hE81AA380 , 32'hFBBAC588 , 32'h1655CA40 , 32'hF6964A30 , 32'hFA784428 , 32'h1302D620 , 32'h09549140 , 32'hF5C44AD0} , 
{32'h0C5759C0 , 32'hFCBEBB5C , 32'hFE73B318 , 32'hFD9C3E48 , 32'hFA104AE0 , 32'h01BAE7DC , 32'hFBFC9928 , 32'h075EF0D8 , 32'hF47F2330 , 32'hF9F16EE0 , 32'h00537F14 , 32'hFF0D34E0 , 32'hFBEF8348 , 32'hF38A2EF0 , 32'h0C860A90 , 32'h0285C240 , 32'hFDD42584 , 32'hFB6523F0 , 32'h04415470 , 32'h04E5FCE0 , 32'hFFC431B1 , 32'h07186450 , 32'hFAB5CAC0 , 32'h18DB4200 , 32'hF606D700 , 32'h0BEBADD0 , 32'h0026DCDC , 32'hF179FF80 , 32'hFBFE8268 , 32'hF91D6030 , 32'hF194A8B0 , 32'h0666B4D8 , 32'hFF8B9D3B , 32'h07210D68 , 32'hFDD7784C , 32'h033880A0 , 32'hF138E030} , 
{32'h0CFDA460 , 32'hFC7326C0 , 32'h077A3A68 , 32'hF58E7800 , 32'hF2B5ECE0 , 32'h07C050E0 , 32'h00A9D086 , 32'hE8F8DA20 , 32'hF88BE678 , 32'h182B50E0 , 32'hF4966CD0 , 32'h09050050 , 32'h05F17E40 , 32'hEDE6D540 , 32'h089BDA30 , 32'hFB410AE0 , 32'h10F6BA40 , 32'h095653F0 , 32'hE976C1E0 , 32'h07B334F8 , 32'hEED9F900 , 32'hF0404410 , 32'hF156ABF0 , 32'h0E6C9D50 , 32'h059D0FF8 , 32'h03676AFC , 32'h0761B770 , 32'h229289C0 , 32'h045B9D80 , 32'h04B6DAC8 , 32'h05E0B558 , 32'h0608F8D0 , 32'hFA4F94F8 , 32'hF2E76C10 , 32'h008436AA , 32'h0FBAE4D0 , 32'h0F44D5E0} , 
{32'h068F1BB8 , 32'h016A3BF4 , 32'h0FF26180 , 32'h02619374 , 32'hF8080D68 , 32'h0BF9C160 , 32'hFEBE001C , 32'h08B67780 , 32'hFBE87C48 , 32'h099E04A0 , 32'hFAF43978 , 32'hFE5511A4 , 32'h16D978A0 , 32'h00C71F37 , 32'h0AF8D360 , 32'hF9677FB0 , 32'h05B772C0 , 32'h0610AF88 , 32'h0F335910 , 32'hFACDFA08 , 32'hFA54AC90 , 32'hF76D4B10 , 32'hFEBFC654 , 32'h05523D20 , 32'hFB62EEF8 , 32'h005F5226 , 32'hF66A5EB0 , 32'h10D42580 , 32'h020FFFF0 , 32'h033463CC , 32'hFE3ED8E4 , 32'h03A7E2D8 , 32'h008A6ECF , 32'h042D3BF8 , 32'h02CC1448 , 32'h0074F3BA , 32'h0E68A9E0} , 
{32'h098A77F0 , 32'h050F8628 , 32'hFFA6BA2A , 32'h00EB611A , 32'hFB5F0BB8 , 32'h058D9B78 , 32'h05B01FA0 , 32'hFF831ABF , 32'hFAD53748 , 32'h01AB7594 , 32'hF9EB3738 , 32'hF6F811D0 , 32'h094CFF90 , 32'h0A2886F0 , 32'hFA4066C0 , 32'h09932220 , 32'h018A4BF4 , 32'hF4911480 , 32'hF79539B0 , 32'hFF99D170 , 32'h0E827950 , 32'hFBA1B900 , 32'h05CBDC70 , 32'h0F117FE0 , 32'h00CE3310 , 32'hEE5E04A0 , 32'h02E7CA64 , 32'h034B34F0 , 32'hF5A04280 , 32'hF747C0B0 , 32'hF613C9C0 , 32'hF8C0E8D8 , 32'hF5040A00 , 32'hFC7446F0 , 32'hFEAA6850 , 32'hF8823560 , 32'hFF152B67} , 
{32'h08C611E0 , 32'h0FAE8890 , 32'hFF5AD729 , 32'hF752FD40 , 32'h02876500 , 32'hFE3F77A4 , 32'h023A3580 , 32'h080F3B10 , 32'hFFB3D95E , 32'h00EF901D , 32'hFF2D085E , 32'hFDB2E5DC , 32'h05A83A70 , 32'h006A5B3A , 32'hF85264B8 , 32'h0853CF00 , 32'h01C0903C , 32'hF14CB690 , 32'hF526DB90 , 32'h022867CC , 32'h10201FE0 , 32'hF9BBA568 , 32'hFC732C38 , 32'h0EB07270 , 32'h08A02010 , 32'hFA2C19A8 , 32'hFE5E609C , 32'h06E460C8 , 32'hFAB51828 , 32'hF7EC93A0 , 32'hF96FD640 , 32'h000A5ED0 , 32'hF9AC1540 , 32'hFC04FDA4 , 32'h003AC1F5 , 32'hF2C9FBA0 , 32'hFC7ED144} , 
{32'hFB455808 , 32'h00629298 , 32'hF76C4F70 , 32'hEB358860 , 32'hFEC00604 , 32'h0C134AA0 , 32'hE96007A0 , 32'h098B90F0 , 32'hF2CAA2F0 , 32'h0D0BC2C0 , 32'h0053506C , 32'hF5CA0620 , 32'hEF6EC660 , 32'hF13EB420 , 32'hFC000540 , 32'hFFCD0385 , 32'hFED4AAA4 , 32'h031C7B28 , 32'h0A350310 , 32'h05A68650 , 32'hF85EC018 , 32'h00A95EF3 , 32'hE6B4BC80 , 32'h07777148 , 32'hF4C21A60 , 32'hEBF7AC60 , 32'h02F8AF04 , 32'hFA4F9548 , 32'h0169F1A4 , 32'h18922680 , 32'hE42A6BA0 , 32'hF0D26F40 , 32'h28C83140 , 32'h16425BA0 , 32'h0846C3B0 , 32'h0E974680 , 32'hEAA12BE0} , 
{32'hFA045300 , 32'h09B3FD00 , 32'hF4F2F620 , 32'h004287E3 , 32'h041DECA8 , 32'h02705854 , 32'hFEAA5320 , 32'h07BD2300 , 32'hF891E1B8 , 32'hFE09DD58 , 32'h08062310 , 32'hFBDD5430 , 32'h03122E6C , 32'hFB025A38 , 32'h01273AE0 , 32'hFCE84610 , 32'hFEF5B868 , 32'hFBD6A5C0 , 32'hFBFC1638 , 32'hFDF9C1FC , 32'hFCBB49BC , 32'hFF723558 , 32'h013494A8 , 32'h058D4110 , 32'h03EFEF50 , 32'hFB314618 , 32'hFE6076C4 , 32'h05E55F68 , 32'h05CCEF68 , 32'hFD8C2484 , 32'h04B05578 , 32'hF96316F8 , 32'h0DEE9220 , 32'h00BCC93B , 32'hFCDF7EDC , 32'hFFD00D59 , 32'h01FEF340} , 
{32'h005A9D71 , 32'hFFC06008 , 32'hFF6B03E2 , 32'hFFCCF6CF , 32'hFF9FC287 , 32'hFF3BF805 , 32'h002A4C3A , 32'h01C1E988 , 32'hFDEDFE8C , 32'h0079A9D5 , 32'hFF2EDF6E , 32'hFFECA15D , 32'h00A262A1 , 32'h00193ADC , 32'h007FCF77 , 32'hFFB836E1 , 32'hFFA57212 , 32'hFEDE1E6C , 32'hFF9B24D3 , 32'h00782264 , 32'hFF188A8C , 32'h01DE8C90 , 32'hFF36EAB3 , 32'h02505938 , 32'hFF8E3D13 , 32'hFEAA40C8 , 32'h00F5FAA6 , 32'h00262522 , 32'h0137ACC4 , 32'h002B7EA1 , 32'hFF83D8D2 , 32'hFF614936 , 32'h00DE1D6D , 32'h00BB53A7 , 32'hFF33C785 , 32'hFF6506CD , 32'h003F8938} , 
{32'h0D373000 , 32'hFC7A9DBC , 32'hFE2DEC28 , 32'hF28AE130 , 32'h00375F28 , 32'h00F73B7D , 32'hFBB1CD78 , 32'h05C95968 , 32'hEFBFAE40 , 32'hF3F36190 , 32'hFB2B26F8 , 32'hFE1262DC , 32'hFB36E8D8 , 32'hE5EC5FC0 , 32'h09855BE0 , 32'hFE5366C8 , 32'hFCFD5D44 , 32'hF3AF65A0 , 32'h05050B78 , 32'h0B80C950 , 32'hF68F56F0 , 32'h04A747E0 , 32'hF42072E0 , 32'h1C4C9100 , 32'hEC094780 , 32'h01C8993C , 32'hF9650E30 , 32'hEEECABC0 , 32'h0D6686A0 , 32'hFE57E790 , 32'hE2ECF240 , 32'hFED69FC8 , 32'h028E221C , 32'h0F352FF0 , 32'h04AE6D68 , 32'hFA4BE0F8 , 32'hFDCFA300} , 
{32'h0C13F300 , 32'hFC82C2CC , 32'h02C14300 , 32'hFDF21A64 , 32'hFE71EC54 , 32'hEFC63940 , 32'hFD998ED8 , 32'h0BB533A0 , 32'hE1E94D60 , 32'hF3588020 , 32'hFDE6157C , 32'hF862F7E8 , 32'hF804F500 , 32'hEFC81EE0 , 32'h07A15978 , 32'hF4D5C7A0 , 32'h0A8C3B70 , 32'hF9DFC900 , 32'h0E857C80 , 32'h030D47C8 , 32'hF8E0CD78 , 32'h11905B80 , 32'hF9DFBE40 , 32'h1B916BE0 , 32'hFCEDC154 , 32'hFDF8321C , 32'hFFD2A8A2 , 32'hF6C9D120 , 32'h0508E898 , 32'hFB73E5A8 , 32'hF41D5CD0 , 32'h0138D7E8 , 32'h09823940 , 32'h100C6E00 , 32'hEF933440 , 32'hFC422E44 , 32'hF75430A0} , 
{32'h000BA4D0 , 32'hFFEBC28D , 32'h000B1ED3 , 32'h000362DE , 32'h0005002A , 32'hFFEFC896 , 32'h00004612 , 32'hFFF636A8 , 32'hFFE5F1C1 , 32'hFFE88D34 , 32'h0018B145 , 32'hFFFF09E3 , 32'hFFFE2C0D , 32'hFFFBB810 , 32'h001DB651 , 32'hFFF7222A , 32'h000DCC35 , 32'hFFF3ACA8 , 32'hFFFDB450 , 32'hFFD42706 , 32'hFFFEDAC1 , 32'h001B9B50 , 32'hFFFFC2AB , 32'h000CD7E1 , 32'h002D3A9D , 32'hFFD88AA7 , 32'hFFE9C364 , 32'h0004BA13 , 32'h001ECD1D , 32'hFFF0688A , 32'h000DE82D , 32'h001085FD , 32'h001BFC69 , 32'h00094198 , 32'hFFF311C5 , 32'hFFF1FB78 , 32'hFFF8B5D3} , 
{32'h002F12E2 , 32'hFFAC3F8A , 32'h0035D757 , 32'hFFD83C36 , 32'hFFE6536A , 32'hFFC70E5C , 32'hFFC54190 , 32'h00120C3D , 32'hFF54B423 , 32'hFF5BA442 , 32'h00621514 , 32'h00246054 , 32'h0042FC5C , 32'h000F1F22 , 32'h0088A58F , 32'hFFF53A5E , 32'h004C00D1 , 32'hFFF6849B , 32'hFFD02069 , 32'hFFF473E4 , 32'h0015F543 , 32'h00863492 , 32'hFF800D7E , 32'hFFE0348E , 32'h0061E562 , 32'hFFE5C674 , 32'hFF984539 , 32'h0042CF0F , 32'h004C62DE , 32'hFFAFEE54 , 32'h00170EC7 , 32'h0021603D , 32'h0060D281 , 32'h001EB4C0 , 32'hFF719078 , 32'h005A34EE , 32'hFF9FE5B5} , 
{32'h002B42A8 , 32'hFFA8F830 , 32'h0034C6D2 , 32'hFFD2DC60 , 32'hFFD5B234 , 32'hFFB73A7A , 32'hFFBC3B06 , 32'h000E5CBD , 32'hFF3AF9DC , 32'hFF4C10A2 , 32'h006DCD98 , 32'h003C6788 , 32'h0055FEAC , 32'h00276CDD , 32'h00A04DF9 , 32'hFFFB4BA1 , 32'h004EF400 , 32'h0002D1F1 , 32'hFFC05DEE , 32'hFFF96758 , 32'h00222623 , 32'h009C66DC , 32'hFF6E6B40 , 32'hFFC4D8FD , 32'h006CF487 , 32'hFFEAC100 , 32'hFF8F9015 , 32'h00576A0E , 32'h004A1B36 , 32'hFFAE7403 , 32'h001441CC , 32'h003017F7 , 32'h005E6D5D , 32'h00292AEE , 32'hFF6C9A5F , 32'h005E9AC0 , 32'hFF9A9FF6} , 
{32'hFFFEC95C , 32'hFFFDB335 , 32'hFFFA9060 , 32'hFFFF88BB , 32'h00011907 , 32'h0001EE2A , 32'hFFFF9E79 , 32'h0000249A , 32'hFFFFCF95 , 32'h000077E4 , 32'hFFFF2BE7 , 32'h00000D01 , 32'hFFFCF477 , 32'h0001A385 , 32'h000047E6 , 32'hFFFDF1F8 , 32'h00022C1D , 32'hFFFF0416 , 32'h0004E6CB , 32'h0001153A , 32'hFFFFA062 , 32'hFFFBF73B , 32'h00051378 , 32'h0008868E , 32'hFFFEE487 , 32'h00045BBE , 32'hFFFF8A03 , 32'hFFFCBFD3 , 32'h0002AFFB , 32'hFFFE9C77 , 32'h0002DB0C , 32'hFFFBC03F , 32'hFFFC4700 , 32'hFFFF7498 , 32'hFFFDDD56 , 32'hFFFE2138 , 32'hFFF9CDFD} , 
{32'hFFFF95A9 , 32'h000202E5 , 32'hFFFDD844 , 32'h0003230A , 32'h0000F55F , 32'hFFFF481C , 32'hFFFBD4F1 , 32'hFFFE5F8B , 32'h000326FC , 32'h0004EE51 , 32'hFFF9A75D , 32'hFFFCA092 , 32'hFFFCCA0B , 32'h0000854B , 32'h00040351 , 32'h000004E2 , 32'hFFFC26C4 , 32'h0007104F , 32'h00007DCF , 32'h0005E69A , 32'hFFFF1626 , 32'h00028200 , 32'hFFFA3674 , 32'hFFFF3999 , 32'h00009899 , 32'h000026AA , 32'hFFF9046E , 32'hFFFECD78 , 32'hFFFD4A6D , 32'hFFFD1812 , 32'h0001612B , 32'hFFFCB31E , 32'hFFFF8E52 , 32'h0001370E , 32'hFFF78632 , 32'hFFFDCA7E , 32'hFFFC1CD1} , 
{32'h0004E691 , 32'h0001F6CD , 32'hFFFE116B , 32'h0000B92B , 32'hFFFED608 , 32'hFFFF6996 , 32'h00054FF9 , 32'h0001D9C2 , 32'hFFFE2779 , 32'hFFFFF18E , 32'hFFFF7181 , 32'h00053991 , 32'hFFFF6D03 , 32'hFFFFE1C9 , 32'hFFFE5C64 , 32'hFFFCF6C0 , 32'h00024DAC , 32'hFFFAD456 , 32'hFFFBC32B , 32'h0001B23C , 32'h00010C87 , 32'h00007DC7 , 32'h000137C4 , 32'h00003822 , 32'h00017D20 , 32'h00031855 , 32'h0003E2B1 , 32'hFFFF78C4 , 32'hFFFED4F2 , 32'hFFFF051F , 32'h00065BBF , 32'hFFFC7754 , 32'h00014069 , 32'h0000C5D7 , 32'hFFFF0176 , 32'h000808E0 , 32'h0006ED46} , 
{32'h000018E2 , 32'hFFFE35BC , 32'h0001689C , 32'hFFFF711E , 32'h0000B2B5 , 32'hFFFFAE77 , 32'hFFFE9887 , 32'hFFFCB211 , 32'hFFFC0663 , 32'h0004A19C , 32'hFFFBA373 , 32'h00047B48 , 32'hFFFE08D4 , 32'hFFFCBEC4 , 32'h00001BE6 , 32'h00057162 , 32'h000480D5 , 32'hFFFC089E , 32'h0002A8C1 , 32'hFFFEE7AF , 32'hFFFC67AD , 32'h0009187A , 32'hFFF79DEB , 32'hFFFF8F24 , 32'hFFFE3E22 , 32'h00004F17 , 32'hFFFD208F , 32'h00001C82 , 32'h000113BE , 32'h0001577A , 32'h00051EF6 , 32'hFFFE69DF , 32'hFFFB6B75 , 32'h0001840C , 32'hFFFC9E88 , 32'h000457AC , 32'h0001CC28} , 
{32'h00036C4A , 32'h00024F93 , 32'hFFFD7678 , 32'hFFFB9C92 , 32'hFFFFFCF1 , 32'hFFFEC2A4 , 32'hFFFBC215 , 32'hFFFAE019 , 32'hFFF57BDE , 32'h00020C47 , 32'h0005C787 , 32'h0002AEEC , 32'h0001ACA2 , 32'h0001B254 , 32'hFFFE3087 , 32'hFFFEC7B6 , 32'h00008EA0 , 32'hFFFE0024 , 32'h0002A2F6 , 32'h000457EE , 32'hFFFDC4A9 , 32'hFFFE062B , 32'h00020521 , 32'hFFFF5ECB , 32'hFFFF047B , 32'hFFFBA063 , 32'h000CEC02 , 32'hFFFD1973 , 32'h00012884 , 32'hFFFFCD81 , 32'hFFFCD12C , 32'hFFFCE189 , 32'h000114B8 , 32'hFFFDB1EC , 32'h0002FBDA , 32'h0000E852 , 32'hFFFA870C} , 
{32'h00007300 , 32'h0000357C , 32'h00012905 , 32'hFFFE0160 , 32'hFFFFC7E1 , 32'h00043159 , 32'hFFFA1C9F , 32'h0000D3B2 , 32'h0009D81D , 32'hFFFD8AAB , 32'hFFFA4BBB , 32'h00007CF6 , 32'h0002D8C5 , 32'h00029A69 , 32'h0000C8EC , 32'h0001C1C8 , 32'h00011FBC , 32'hFFFF5FAA , 32'h00015A1A , 32'hFFFDC288 , 32'h00041AFE , 32'h00009300 , 32'hFFFF1E96 , 32'h00069FB3 , 32'h00025121 , 32'hFFFC109C , 32'hFFFE1F01 , 32'h00003FCF , 32'h0002AE22 , 32'h0004B898 , 32'h0007BDBF , 32'hFFFF7D63 , 32'h0000D53F , 32'h00053B86 , 32'h0002D6F9 , 32'h0005C78A , 32'h000244F0} , 
{32'h00039CB3 , 32'h00068611 , 32'hFFFF848B , 32'h00048839 , 32'h000166F0 , 32'h0000EAAD , 32'h0000B211 , 32'h000445EA , 32'hFFFCD8BF , 32'h0007D73C , 32'h0003DC17 , 32'hFFFF4D3A , 32'hFFFE14C0 , 32'h00013FDA , 32'hFFFDBFA1 , 32'hFFFD1F7C , 32'h0002ED95 , 32'hFFFEDF4E , 32'hFFFF135F , 32'h00036721 , 32'h00031A13 , 32'hFFFBAD1D , 32'h00013973 , 32'h00016FCD , 32'h000647CC , 32'hFFFFCC0A , 32'hFFFFC491 , 32'h000083C3 , 32'hFFFC4B7B , 32'hFFFE6BF9 , 32'h000203F1 , 32'h00022816 , 32'h0001DAC5 , 32'hFFFF07AF , 32'hFFFE549B , 32'hFFFE5300 , 32'h00039969} , 
{32'h0000E09C , 32'hFFFE57D9 , 32'hFFFCDAE7 , 32'hFFFDB0BC , 32'h0001706C , 32'hFFFBD83B , 32'hFFFD32AF , 32'h00020DBD , 32'hFFFFE7C6 , 32'hFFFF75EC , 32'h0002D8FD , 32'hFFFDD81E , 32'hFFFBB9B7 , 32'h000563FA , 32'hFFFB2B84 , 32'h0000FCD5 , 32'hFFFC8CD1 , 32'hFFF98975 , 32'h00008F02 , 32'hFFFF7C1F , 32'hFFFAF326 , 32'hFFF9ADCD , 32'h000487C1 , 32'hFFF9F40C , 32'hFFFF79D6 , 32'h000328E6 , 32'hFFF94E38 , 32'hFFFBCB47 , 32'h00014F3C , 32'hFFFC5C91 , 32'h0001FB2A , 32'h000818E1 , 32'hFFFD9735 , 32'h0005B12F , 32'h00001B05 , 32'hFFFD1090 , 32'h0002E6FB} , 
{32'h0005BEBC , 32'hFFFC97BB , 32'h00033AE7 , 32'h00018CB7 , 32'hFFFBF26E , 32'h0001451E , 32'hFFFFD887 , 32'hFFFE3061 , 32'h0002C05F , 32'h0000B8DF , 32'h0003047C , 32'hFFFE3AB8 , 32'h0002E267 , 32'h00000118 , 32'h00013FBF , 32'h000116FD , 32'h00008CD1 , 32'h00003EC1 , 32'h00035B18 , 32'h00026C43 , 32'h0000DD4D , 32'h00025E58 , 32'hFFFE8356 , 32'hFFF9633E , 32'h0003984A , 32'hFFFE83E3 , 32'h0003692E , 32'hFFFFA119 , 32'h0000AD85 , 32'h00032541 , 32'h00046F33 , 32'hFFFE4C21 , 32'hFFFDFC59 , 32'h0000E091 , 32'hFFFEF830 , 32'hFFFE6B5E , 32'hFFFFE900} , 
{32'h000F9A6F , 32'hFFEBC3B3 , 32'hFFE3A05F , 32'h002F79C7 , 32'hFFF2787A , 32'hFFECA83F , 32'h0000B89A , 32'h005228F3 , 32'h0031A8A8 , 32'h0016646B , 32'hFFA4D83B , 32'hFFD8A1A7 , 32'hFFD54DFC , 32'hFFDF508C , 32'hFFE0DA14 , 32'hFFFAC43B , 32'hFFF2277C , 32'hFFFE64D0 , 32'h001E4C35 , 32'h00252178 , 32'hFFEBA360 , 32'hFFEC8401 , 32'hFFFC9A7E , 32'h00079DA7 , 32'hFFF86CDB , 32'hFFFC68A5 , 32'h000778B5 , 32'hFFFA9C17 , 32'h00153250 , 32'hFFFB8C07 , 32'h000F1491 , 32'h000266EC , 32'hFFF8214C , 32'hFFE98AED , 32'h00136845 , 32'h0005C04B , 32'h000FDDE4} , 
{32'h000D23B2 , 32'hFFEB8FBE , 32'hFFE76EDC , 32'h00326BA5 , 32'hFFEC6F5B , 32'hFFEF5392 , 32'h0007B3E5 , 32'h00507147 , 32'h0035A1D1 , 32'h001BBACA , 32'hFFA80591 , 32'hFFDE939D , 32'hFFD92F18 , 32'hFFDED814 , 32'hFFE21E19 , 32'h0000D466 , 32'hFFF0A5AE , 32'hFFFE806A , 32'h001AE3D7 , 32'h0020E3BF , 32'hFFE85F18 , 32'hFFF102E1 , 32'hFFF6FD85 , 32'h000EAC5B , 32'hFFFA536E , 32'hFFFDB310 , 32'h0001D632 , 32'hFFFBBAF7 , 32'h00114911 , 32'hFFFE2DA9 , 32'h001115C7 , 32'h00021FC5 , 32'hFFF6FFA6 , 32'hFFE8A6B0 , 32'h00107241 , 32'h0006D548 , 32'h001671BD} , 
{32'hFFFD4F90 , 32'hFFFD7D36 , 32'h00045089 , 32'hFFFF1CFA , 32'h00018E00 , 32'hFFFCEAA2 , 32'hFFFF11E0 , 32'hFFFC10AF , 32'h00048164 , 32'hFFFEC63D , 32'h000182BA , 32'h00026D9C , 32'hFFFF1B4F , 32'hFFFD64D4 , 32'h000000D7 , 32'hFFFFC34C , 32'h0001B00D , 32'h0005798C , 32'h000214ED , 32'hFFFD9949 , 32'hFFFD2F12 , 32'hFFFB3969 , 32'h0002F5FA , 32'hFFFFE5B9 , 32'hFFFE3036 , 32'hFFF7C2B2 , 32'hFFFEA8A3 , 32'hFFFCDACB , 32'hFFFC023A , 32'h00025AD3 , 32'hFFFB8786 , 32'h0005ABAB , 32'h000618FB , 32'h0001B168 , 32'hFFFF4258 , 32'h0002CC4A , 32'hFFFDA0CC} , 
{32'hFFF9D137 , 32'hFFFC940B , 32'hFFFE314D , 32'hFFF9F5C6 , 32'hFFFEABA8 , 32'hFFFFD294 , 32'h00093355 , 32'hFFFEACD8 , 32'hFFFA121D , 32'hFFFDA4DA , 32'h00027D0A , 32'h00042A7A , 32'hFFFCE074 , 32'hFFFBD56F , 32'h0000BBF1 , 32'h00031986 , 32'h0002C81D , 32'h0002A6C1 , 32'hFFF99E10 , 32'h00052BB7 , 32'hFFFC9C67 , 32'h000664E8 , 32'hFFF829D1 , 32'hFFF85FF8 , 32'h00034659 , 32'hFFF7E2F1 , 32'h0006E633 , 32'hFFFBFEC3 , 32'hFFFB7822 , 32'hFFFB558E , 32'h00016738 , 32'h000190EE , 32'h00023D1C , 32'h0000E633 , 32'hFFFE82CE , 32'h00025C77 , 32'h00010CEC} , 
{32'h0006EC4C , 32'h00098657 , 32'h0009DB07 , 32'hFFFA50B8 , 32'h000A5771 , 32'hFFF30C2A , 32'h000842BB , 32'h000496D5 , 32'hFFFBC356 , 32'h000781CB , 32'hFFFE6290 , 32'h00033E4F , 32'hFFF68FA8 , 32'h0003DF09 , 32'h0007F9F0 , 32'h000C3684 , 32'hFFF7DE70 , 32'h0012A811 , 32'h0003F9C5 , 32'hFFF9B4B7 , 32'h00091DA9 , 32'hFFF9226F , 32'hFFF83E76 , 32'h000287CD , 32'h0007CE46 , 32'hFFFE8BA3 , 32'hFFF84029 , 32'h0006A4C7 , 32'hFFF5B43F , 32'hFFFBDDF1 , 32'hFFFEB2AF , 32'hFFFAA84C , 32'hFFFDBDD6 , 32'hFFFBC2D4 , 32'hFFF49B53 , 32'h000A36F2 , 32'h0001930A} , 
{32'h0DCE1B00 , 32'hFBA3E3F8 , 32'hFD971B38 , 32'hFA83F240 , 32'hFEFAE714 , 32'h0463F458 , 32'hFA6FD618 , 32'h04F437B0 , 32'hF5895CE0 , 32'hF7028880 , 32'h01BA3A4C , 32'hFA200118 , 32'hF9304E90 , 32'hF0186670 , 32'h072264F0 , 32'h01D4D9AC , 32'hFDA63F40 , 32'hF8A11FF8 , 32'h05CC6C78 , 32'h03B41144 , 32'hF8ACEA70 , 32'h03736734 , 32'hF748FD90 , 32'h18E02540 , 32'hF1D36770 , 32'h02EACC6C , 32'h000B9766 , 32'hEED0EDC0 , 32'h04EA5E68 , 32'hFF7B4282 , 32'hEF3B45A0 , 32'h00CDF258 , 32'h0594E740 , 32'h0EF203C0 , 32'hFB0E3E70 , 32'h005168A3 , 32'hF71D79E0} , 
{32'hFF69CD04 , 32'hFFE3A669 , 32'hFF0A3D3B , 32'h0018FA7F , 32'hFF0C925B , 32'hFF45FC1B , 32'h0005FE55 , 32'hFF6497D0 , 32'h00309BCE , 32'hFF31275A , 32'h00023B75 , 32'hFF75A666 , 32'h00115D99 , 32'h0045CFBC , 32'h009B3752 , 32'hFFA54690 , 32'h006F4D63 , 32'h000C6BFE , 32'h006BD198 , 32'h0053273C , 32'hFFBCFD54 , 32'h003ED099 , 32'hFF985A2C , 32'h00F1B035 , 32'h0036AB89 , 32'hFFE32215 , 32'hFEB96968 , 32'h000A1D4D , 32'h00777789 , 32'hFFFF8891 , 32'h00D5AAAD , 32'h0040CF94 , 32'hFFD2779A , 32'h00586E94 , 32'hFF601F6D , 32'hFF909DA9 , 32'h00259410} , 
{32'hFFC92443 , 32'hFFC1A1C4 , 32'hFFC6FA87 , 32'h0005EC80 , 32'hFFB2F854 , 32'hFFF1D3E7 , 32'h0044A85A , 32'hFFECEA02 , 32'h00037922 , 32'hFFC10AF6 , 32'hFFEDBE91 , 32'hFFE7C288 , 32'h002A992E , 32'h00173C80 , 32'hFFE6DA41 , 32'hFFC2505D , 32'h00166446 , 32'hFFF5068E , 32'h002B1DB8 , 32'h00091312 , 32'hFFFA420F , 32'h00554961 , 32'hFFD8F1D0 , 32'h0033631F , 32'h00296AC0 , 32'h0003097E , 32'hFFC5F9DD , 32'h000C30C8 , 32'h0048E63A , 32'h00050AB6 , 32'h0025FC0F , 32'h00096140 , 32'h00127950 , 32'h001AA72B , 32'hFFD9EA50 , 32'hFFE7A653 , 32'h0011EB56} , 
{32'h0B05AD90 , 32'hFD15D63C , 32'hFF324731 , 32'hFC7261D4 , 32'hFF71319D , 32'h04ACABC0 , 32'hFBE1BC60 , 32'h040BA5B0 , 32'hF8526438 , 32'hFA2675C0 , 32'h020129A8 , 32'hFC31B2A8 , 32'hFB2D95E8 , 32'hF3F24880 , 32'h058BB290 , 32'h012B42E4 , 32'hFEF66E04 , 32'hFA57F648 , 32'h04444178 , 32'h02FC9E68 , 32'hFA396EB8 , 32'h018A7AC4 , 32'hF9C97D58 , 32'h11AEFF00 , 32'hF47B6E30 , 32'h0204CCB4 , 32'h00CB777F , 32'hF2C15E20 , 32'h0348738C , 32'hFEA2D928 , 32'hF2F56C60 , 32'h00EB3FFF , 32'h04935978 , 32'h0AE9B9C0 , 32'hFBF9B460 , 32'h007BFBB6 , 32'hFA005BA8} , 
{32'h035F880C , 32'hFF128C57 , 32'h008392D5 , 32'h023114F8 , 32'h02CAB458 , 32'h07B60020 , 32'hFB548BD8 , 32'hFCE6128C , 32'hFFEE2AD1 , 32'hFE96FE54 , 32'hFEF91548 , 32'h05AC3958 , 32'h0C19D700 , 32'hEF6F2FA0 , 32'hFA7A2D88 , 32'hF8D1ED60 , 32'h0FB8C090 , 32'hFA222F18 , 32'hFA02C3D0 , 32'h0F38C5C0 , 32'hFFCF8EBC , 32'h052F4DD8 , 32'h05382D70 , 32'hFE4F71A0 , 32'hFC5EBBA8 , 32'h02231AAC , 32'h05FAB6D0 , 32'hFD29621C , 32'h0148F568 , 32'h04218DD8 , 32'hFE1B3E00 , 32'h076E7908 , 32'h03F67AB8 , 32'hFF99CD19 , 32'h03C9E464 , 32'hEF1F4AC0 , 32'hFF5C03AA} , 
{32'h0056B65D , 32'h0000EE0F , 32'h003BF0DB , 32'h003331B9 , 32'h017AACF0 , 32'h01619638 , 32'hFF4207FA , 32'hFE7F3524 , 32'h0066B908 , 32'h005E2AB8 , 32'h00B630F2 , 32'h00DA9C55 , 32'h01123BEC , 32'hFE7D04B4 , 32'hFF703E3A , 32'h00382C20 , 32'hFFAB2D8A , 32'hFF8DEE35 , 32'h0076CD5C , 32'h00A84AF2 , 32'h00FABA08 , 32'h0000450C , 32'h002A0D9C , 32'hFEDB3188 , 32'hFF7C5B2C , 32'hFF8357B7 , 32'h019B1CB0 , 32'hFE6537EC , 32'hFFDF29FE , 32'hFF9F9ACE , 32'hFED0E3D8 , 32'h0045DFC1 , 32'h01801998 , 32'hFFBDACBE , 32'h01F2CC30 , 32'hFEC84DE0 , 32'h01323424} , 
{32'hFF4E4C19 , 32'h00BC50DB , 32'hFFF5B902 , 32'hFCA79428 , 32'hFFCE3BC8 , 32'h0082D799 , 32'hFEABA6FC , 32'hFEECD188 , 32'hFB3AA300 , 32'hFE2BB770 , 32'h00241940 , 32'h002AC1F8 , 32'hFFDDADFB , 32'hF65A1D60 , 32'h01F061B4 , 32'hFC559FE8 , 32'h0021B003 , 32'hFBDF8930 , 32'h024523B8 , 32'h088F9D80 , 32'hFE9FC178 , 32'h001383F0 , 32'hFEE6D600 , 32'h084A0750 , 32'hF52FF310 , 32'h02398584 , 32'hFAD0FFB0 , 32'hF7561F40 , 32'h0260EBA8 , 32'h01487938 , 32'hF8722C20 , 32'h00394560 , 32'hFEC07BC4 , 32'hFFD54661 , 32'h059DC578 , 32'hFE9C87C8 , 32'h070D0E48} , 
{32'h0B2F6FC0 , 32'hFCA35240 , 32'hFEAB9FA0 , 32'hFB9FDC20 , 32'hFFA22C9E , 32'h03E77F50 , 32'hFBA1B000 , 32'h04357608 , 32'hF7A56610 , 32'hF9717DA0 , 32'h0177E228 , 32'hFBB5D768 , 32'hFA5127B0 , 32'hF34DB500 , 32'h0588B808 , 32'h01C16078 , 32'hFDD9054C , 32'hFA347F88 , 32'h044BF610 , 32'h02DA6010 , 32'hFA5A40E8 , 32'h025D7048 , 32'hF94473B8 , 32'h13448140 , 32'hF4818E70 , 32'h026B9CF8 , 32'h009A0C06 , 32'hF2515D60 , 32'h03A05D68 , 32'hFFAE6FA8 , 32'hF267B050 , 32'h00A102E3 , 32'h0482F750 , 32'h0BA30B30 , 32'hFC715578 , 32'h004C1638 , 32'hF8FC2D38} , 
{32'h0F93F3C0 , 32'hFB4BB3C8 , 32'hFE257788 , 32'hF9D36C88 , 32'hFF710B6F , 32'h04CCFA88 , 32'hFA01F7C0 , 32'h05E19DD0 , 32'hF41A3730 , 32'hF7B24040 , 32'h01B95678 , 32'hFA3AD1D8 , 32'hF868AB98 , 32'hEEE1D740 , 32'h07CE1310 , 32'h01865FAC , 32'hFD3D3A7C , 32'hF8549EA0 , 32'h058442E0 , 32'h03FB446C , 32'hF805A928 , 32'h040A22E8 , 32'hF65BBBC0 , 32'h1AB8B920 , 32'hF1082460 , 32'h01E18F18 , 32'h01A9D4C8 , 32'hEE822460 , 32'h060CA2E0 , 32'hFFE0AA1F , 32'hEE134220 , 32'h01137AFC , 32'h0650C248 , 32'h0F4C1C10 , 32'hFA5360F0 , 32'hFFAD047A , 32'hF749B1A0} , 
{32'h0172B258 , 32'h000C83FC , 32'hFFD08D40 , 32'hFF9D06BF , 32'h003BC9F4 , 32'hFF874ADD , 32'hFFAC8F39 , 32'h0037AF4C , 32'hFEC3FB84 , 32'h003B53DC , 32'hFF70D05E , 32'h0022A3D9 , 32'hFFB712D6 , 32'hFF2452BE , 32'h00905B5D , 32'hFEF4C058 , 32'h0059C96F , 32'h003113BB , 32'h000161E4 , 32'h004F4916 , 32'hFF4A3B7A , 32'h0145CD14 , 32'hFEEA697C , 32'h01E0EFB4 , 32'h00289894 , 32'hFE95AD90 , 32'h00B515DE , 32'h002D1B58 , 32'h01750A58 , 32'h000520E4 , 32'hFF65C78A , 32'h00B5AF1F , 32'h00AD8424 , 32'hFFBFEC5B , 32'hFEA17978 , 32'hFEECD1C0 , 32'h0052E7F1} , 
{32'h00B4B0BA , 32'h00198A61 , 32'h0019CF21 , 32'hFFB415FE , 32'h0025C8EC , 32'hFFBE338B , 32'hFFD3ABE5 , 32'h001B6F37 , 32'hFF763FA1 , 32'h002B721E , 32'hFFE246F2 , 32'h002DDC34 , 32'hFFAE158C , 32'hFF9A461A , 32'h00633DA0 , 32'hFF75B288 , 32'hFFF7EC2B , 32'h00033459 , 32'h00294525 , 32'h0001AC3F , 32'hFFA97074 , 32'h0062AE4E , 32'hFF7435D3 , 32'h0100AC74 , 32'h00281664 , 32'hFF72968B , 32'h00335E86 , 32'h0004E469 , 32'h00FDB28C , 32'hFFDE9687 , 32'hFF967718 , 32'h002BAF4B , 32'h0012A84F , 32'hFFF6343A , 32'hFF90B032 , 32'hFFBCA56C , 32'hFFEEAD6C} , 
{32'hFFFFC2D6 , 32'h00009C68 , 32'hFFFB3E0C , 32'h00015561 , 32'hFFFFEE50 , 32'hFFFE4466 , 32'h000164C7 , 32'h0000A37A , 32'h0000CA24 , 32'h0003AE9F , 32'hFFFAC8D2 , 32'h00013D86 , 32'h000030F6 , 32'hFFFF97BC , 32'hFFFC6A3A , 32'h0003573B , 32'hFFFCF19E , 32'h000296D7 , 32'h0002D831 , 32'hFFFF125E , 32'hFFFA7EB2 , 32'hFFFDCE53 , 32'h000374AB , 32'hFFFF8B0C , 32'h00035336 , 32'hFFFF8B6D , 32'hFFFD4DDE , 32'h00022E32 , 32'h0000F08F , 32'h00003222 , 32'hFFFD7B5B , 32'h00034541 , 32'hFFFE9279 , 32'h000128A6 , 32'hFFFFB923 , 32'h000559C7 , 32'h00025046} , 
{32'h00022113 , 32'hFFFF6E5D , 32'h00034393 , 32'hFFF954D7 , 32'h00016603 , 32'hFFFFA2FB , 32'hFFFEF4E7 , 32'hFFFB2362 , 32'h0004CEE7 , 32'hFFFD68D5 , 32'hFFFDAAC6 , 32'hFFFD0FB6 , 32'h00001F78 , 32'h00004C7C , 32'h0002F185 , 32'h0002571A , 32'hFFFD669D , 32'hFFFE8723 , 32'h000338A8 , 32'h00030FB4 , 32'hFFFBA0AE , 32'h0005C170 , 32'h0001C4F3 , 32'h00036FA5 , 32'h00037232 , 32'hFFFD4219 , 32'h00040DC7 , 32'hFFF7B9A9 , 32'h0005C7A4 , 32'h0001FE4A , 32'h0000FFBE , 32'h000486E2 , 32'hFFFAFFAA , 32'h0004BD00 , 32'hFFFFBEC2 , 32'hFFF8DB60 , 32'h0002086A} , 
{32'h0003247A , 32'hFFFE3405 , 32'hFFFF7659 , 32'hFFFFBA94 , 32'h0006B81C , 32'h0001AB7D , 32'h00014F83 , 32'h00013C27 , 32'hFFFE073E , 32'h00096DB2 , 32'h00009938 , 32'h0000E0A6 , 32'h000196E6 , 32'hFFFFAD7F , 32'h0000EDE3 , 32'hFFFE0DED , 32'h0005DB14 , 32'hFFFDA29C , 32'h000227DE , 32'hFFFDE849 , 32'hFFFF91B5 , 32'hFFFEFD90 , 32'h000607C5 , 32'h00001280 , 32'hFFFEDD23 , 32'h0000369A , 32'hFFFE6439 , 32'h0000488F , 32'hFFFFDDC5 , 32'h0003A533 , 32'h00012A96 , 32'hFFFDB4DE , 32'h0001B5F7 , 32'h00039A8C , 32'h0005DC48 , 32'hFFFE7577 , 32'h0000281F} , 
{32'h0002D7A6 , 32'h000009C5 , 32'h00011CEF , 32'h00002451 , 32'hFFFDE608 , 32'hFFFFD61B , 32'hFFFACE33 , 32'hFFF868A3 , 32'h000310FC , 32'hFFFB100E , 32'hFFFF48FC , 32'h0001EFA2 , 32'h000943C8 , 32'h00007FFF , 32'h0000D37A , 32'h0003748B , 32'hFFFE8FE6 , 32'hFFFCF1FD , 32'h000324ED , 32'h00008279 , 32'hFFFF6327 , 32'h0003DA00 , 32'h00022BF2 , 32'hFFFD0E30 , 32'h00011C20 , 32'hFFFCBADF , 32'hFFFC9D6B , 32'h0001BD97 , 32'hFFFF4938 , 32'h00028AE7 , 32'h00023C8E , 32'h000222B0 , 32'hFFFB2A2B , 32'h000372B7 , 32'h0008B470 , 32'h00046F3E , 32'h0000FA6F} , 
{32'hFFFF0D4D , 32'hFFFED588 , 32'h0001323E , 32'hFFF953EA , 32'hFFF69353 , 32'h00008FFD , 32'h00014E5B , 32'hFFFFF040 , 32'h00062D75 , 32'hFFFF112F , 32'h00027F7A , 32'h0002CDE2 , 32'h0002B9B3 , 32'h0002899F , 32'h0002534B , 32'h00040A6D , 32'h0006F1AF , 32'h000380AC , 32'hFFFF20C1 , 32'h00041270 , 32'hFFFDCB82 , 32'h000268D3 , 32'hFFFF469D , 32'h0006A32A , 32'h0000E4DE , 32'h0005CB87 , 32'hFFFC8FC5 , 32'h00009AE8 , 32'h00032377 , 32'h00009D44 , 32'hFFFE9CAC , 32'hFFFBDDB8 , 32'hFFFCF10B , 32'hFFFA8443 , 32'h00030F35 , 32'h00034AF6 , 32'hFFFEC479} , 
{32'hFFF975C7 , 32'h00022CC4 , 32'hFFFFB946 , 32'hFFF88274 , 32'hFFFFFF84 , 32'hFFFEDBEB , 32'hFFFED1E7 , 32'hFFFDE0BD , 32'h0000D29C , 32'h0001C533 , 32'h00057F0D , 32'hFFFD7A8E , 32'hFFFF3641 , 32'hFFFA1A77 , 32'hFFFC014C , 32'h00017531 , 32'hFFFED8FC , 32'h000169C4 , 32'h00004223 , 32'hFFFFCD82 , 32'hFFFFBAEB , 32'hFFFB492E , 32'h00065ECF , 32'hFFFB809F , 32'h0001E151 , 32'hFFFF21C6 , 32'h000212D5 , 32'h0001FE41 , 32'hFFFC0741 , 32'hFFFDD133 , 32'h00012D88 , 32'h0001854B , 32'hFFFC0308 , 32'h00041764 , 32'hFFFB5FD6 , 32'h0002E3B0 , 32'h000367B4} , 
{32'hFFFCF2B8 , 32'hFFF9F6F9 , 32'hFFFB80F7 , 32'hFFFCE930 , 32'h0000D6FC , 32'h0006D231 , 32'hFFFF1F46 , 32'hFFFDFA70 , 32'h00037090 , 32'hFFFEB526 , 32'hFFFEAF24 , 32'h00013E08 , 32'hFFFABC1D , 32'h0001BF22 , 32'h00016D3B , 32'hFFFC295A , 32'hFFFEE148 , 32'h0001C4CF , 32'h00001832 , 32'h00026882 , 32'h00053E3C , 32'hFFFF896D , 32'hFFFB9C55 , 32'h0001144F , 32'hFFFA1742 , 32'h000A7EAB , 32'hFFFD5E28 , 32'hFFFEEB16 , 32'hFFFD92DF , 32'hFFF98687 , 32'hFFF9E22E , 32'h00012466 , 32'h0002B0FB , 32'hFFFF541A , 32'h0001E584 , 32'hFFFC8C9C , 32'hFFF92BBA} , 
{32'hFFFCECB8 , 32'hFFFAA25D , 32'h0001B806 , 32'hFFFFC571 , 32'h00043B24 , 32'hFFFCDE04 , 32'hFFFC634B , 32'hFFFDC6B6 , 32'h000386D4 , 32'h00042F6D , 32'h0000592C , 32'hFFFA1CFD , 32'hFFFD9055 , 32'h00009154 , 32'h0001E243 , 32'hFFFCA333 , 32'h00029C4B , 32'h00008E36 , 32'h0001C06F , 32'h000324FE , 32'h0002BA13 , 32'h00039AC4 , 32'hFFFC639A , 32'hFFFF5858 , 32'hFFFFCBBF , 32'hFFFEF07D , 32'hFFFFD113 , 32'h00044962 , 32'h0002CE0A , 32'hFFFE4BE6 , 32'h000580C6 , 32'h00056D66 , 32'h000199F6 , 32'h0003CD48 , 32'hFFFA4489 , 32'hFFFE0079 , 32'h0008D06E} , 
{32'hFFFF34BD , 32'hFFFB3C2E , 32'h000431A2 , 32'h0004BC4B , 32'hFFFFAAD2 , 32'hFFFFF41A , 32'h000649EB , 32'h0007F05A , 32'hFFFEDE68 , 32'hFFFE1CEB , 32'h000413D0 , 32'hFFFC0410 , 32'h0001C186 , 32'h00029D56 , 32'h000B2E3E , 32'hFFFD1454 , 32'h000008E8 , 32'hFFFB93EB , 32'hFFF767CF , 32'h000289E2 , 32'hFFFE6AB6 , 32'h000146F1 , 32'h00044E54 , 32'h0000FE88 , 32'hFFFB6CFF , 32'h00016083 , 32'h00000650 , 32'hFFFDFE08 , 32'hFFFB7BC9 , 32'h0000C135 , 32'hFFFDF646 , 32'h00065CE4 , 32'h0002966A , 32'h0002835D , 32'hFFF88F39 , 32'hFFF783BF , 32'h00015994} , 
{32'h0004A3F2 , 32'h000B360F , 32'hFFFE3E22 , 32'hFFFEE411 , 32'hFFFF5A98 , 32'hFFFEB125 , 32'hFFFD6B88 , 32'hFFF9181F , 32'hFFFF7345 , 32'hFFFFDB6F , 32'hFFFBD894 , 32'hFFFC6ED9 , 32'hFFFA357D , 32'h00039AF1 , 32'hFFFE97A8 , 32'h0001E311 , 32'hFFF9BCFA , 32'hFFF7F7B9 , 32'h0000AF4D , 32'hFFFCAE34 , 32'h000015D1 , 32'h000209FC , 32'hFFFA2D42 , 32'hFFFF9FC8 , 32'h0001A753 , 32'h00034D6F , 32'hFFFC7A94 , 32'hFFFBDF8F , 32'h00005609 , 32'h0004DC51 , 32'hFFFF65B0 , 32'hFFFD77D8 , 32'hFFFB2F7D , 32'hFFFD4ABF , 32'hFFFECC96 , 32'h00004A15 , 32'hFFFADEAB} , 
{32'h00045B93 , 32'h0000E1D1 , 32'hFFFEE2CB , 32'hFFFBEA4F , 32'h00031E8A , 32'h000003F5 , 32'h00027436 , 32'hFFFECD7A , 32'h00057ED8 , 32'h000036F4 , 32'h00013042 , 32'hFFFC2672 , 32'hFFFB9756 , 32'h0002B47A , 32'hFFFDC6DD , 32'h00010C02 , 32'h00049D4D , 32'hFFFBCE9E , 32'h00008FC8 , 32'h0002D43C , 32'h00010191 , 32'hFFFFE698 , 32'hFFF68A39 , 32'hFFFBC02A , 32'h0000F5F0 , 32'h0001F731 , 32'h00033447 , 32'h0000A997 , 32'h0002F7AB , 32'hFFFE3DBB , 32'h00015F92 , 32'hFFFAC1A0 , 32'h0001A65A , 32'hFFFD37E0 , 32'hFFFBF75F , 32'hFFFC2678 , 32'h00076A0B} , 
{32'h00002DFD , 32'h000000E5 , 32'hFFFE34BB , 32'h0001C7D1 , 32'h0002F5DA , 32'hFFFD34C7 , 32'hFFFF68EA , 32'h0000B0A9 , 32'hFFFF9C6D , 32'hFFFD70B7 , 32'h0004C05F , 32'hFFFB054A , 32'hFFFE2DE4 , 32'h00093BA6 , 32'hFFFDC931 , 32'hFFFFF494 , 32'hFFF8C1EF , 32'hFFFE0DF9 , 32'hFFFA3D14 , 32'h00054847 , 32'h00010F83 , 32'hFFFA9F1B , 32'h0001B3AE , 32'h000334CD , 32'hFFFFAFF5 , 32'hFFFE1B4E , 32'hFFFF8C93 , 32'h0002A1FE , 32'h000243E8 , 32'hFFF9729B , 32'h00055570 , 32'hFFFFE040 , 32'h0001830D , 32'hFFFEC2D2 , 32'hFFFC033F , 32'h000939A4 , 32'h0007BA6D} , 
{32'h0003BE30 , 32'h00013A00 , 32'h00018543 , 32'hFFFB4313 , 32'hFFFEF79B , 32'hFFFAB971 , 32'hFFFF70FA , 32'hFFFA8992 , 32'hFFFB346A , 32'hFFFF610B , 32'hFFFCF045 , 32'hFFFB236B , 32'h0000F9BC , 32'hFFFF44E5 , 32'hFFF9AF50 , 32'hFFFE0A37 , 32'h0003CD3A , 32'h00021EDF , 32'hFFFE2D54 , 32'hFFFD5F77 , 32'h0005369A , 32'h0002C84F , 32'h00042954 , 32'h000329D2 , 32'h00040925 , 32'h000609D8 , 32'h000A64A2 , 32'hFFFD71AD , 32'hFFFCF6DC , 32'h0001968F , 32'hFFFB4E28 , 32'h00007921 , 32'hFFFC90FA , 32'hFFFCA9E2 , 32'hFFFFC389 , 32'hFFFE64BC , 32'hFFFD8AA3} , 
{32'h00074BEE , 32'h0000AC98 , 32'h00063B2C , 32'hFFFE72DC , 32'h00099BAC , 32'hFFFEF21C , 32'h0005BEBC , 32'hFFF94C47 , 32'h0004A805 , 32'hFFFF4A90 , 32'hFFFD4985 , 32'h0003B3C7 , 32'hFFF99A3C , 32'h0000DC9F , 32'hFFFE5264 , 32'hFFFFA942 , 32'h0002D0DD , 32'hFFFE0954 , 32'h0001713C , 32'h000818EB , 32'hFFFF97CD , 32'h0000A0A9 , 32'hFFFE805C , 32'hFFFCB34A , 32'hFFFA76E9 , 32'h0000676C , 32'hFFFF3EA8 , 32'hFFFBB2AB , 32'hFFFDCC4C , 32'h0000E297 , 32'hFFFFD25B , 32'h0000C1C7 , 32'h0001B9B8 , 32'h0003494B , 32'hFFFBF46D , 32'hFFFDA382 , 32'hFFFDE506} , 
{32'h00047F73 , 32'hFFFA23CA , 32'hFFFAA705 , 32'h0000AAD6 , 32'h0003E1CA , 32'hFFFCBCD4 , 32'hFFF96441 , 32'h0000BCA8 , 32'hFFFEC9A8 , 32'h00014ADB , 32'hFFFF8414 , 32'hFFFAC647 , 32'hFFFB0EE6 , 32'h0002CDCD , 32'h0002E040 , 32'h00079E93 , 32'h00002306 , 32'hFFFF7CAB , 32'hFFFBBEBF , 32'h00019C69 , 32'h0003247A , 32'h00019B5F , 32'hFFFC59B7 , 32'h0004C045 , 32'h0002E436 , 32'hFFFAB101 , 32'h00021A51 , 32'hFFFFCDC0 , 32'h0003A42D , 32'h00025A1F , 32'h00006B70 , 32'hFFFDAED3 , 32'hFFFE2FEA , 32'h00034531 , 32'hFFF90279 , 32'h0000AAC8 , 32'hFFFD067E} , 
{32'h000286C0 , 32'hFFFED975 , 32'h0004896A , 32'hFFFE2E43 , 32'h000621E5 , 32'h0001812D , 32'h0003EFAE , 32'h00000FAF , 32'hFFFE66EC , 32'h00080FE4 , 32'hFFFD1483 , 32'hFFFD33E5 , 32'h0004D1CF , 32'hFFFB8B21 , 32'hFFF948F8 , 32'h00002225 , 32'h0000B0B1 , 32'h00025298 , 32'h000726AB , 32'hFFFD81BD , 32'hFFFF9F1D , 32'h0000D4DB , 32'hFFFF0C09 , 32'h0001AC9E , 32'hFFFFC868 , 32'h0000333A , 32'hFFFD3FCB , 32'h00002856 , 32'h00061856 , 32'hFFFD2317 , 32'h00052C16 , 32'hFFFBE820 , 32'hFFFD8125 , 32'h0002FA08 , 32'hFFFEB27E , 32'h000058E0 , 32'h00017D8C} , 
{32'h0000DFDE , 32'h0004B591 , 32'h00013D7C , 32'h00038168 , 32'h0006B29D , 32'h0008DD5C , 32'h0002AE74 , 32'hFFFF9111 , 32'hFFFE1B22 , 32'h000176E0 , 32'hFFFE1377 , 32'hFFFDBAF3 , 32'hFFFFD55F , 32'h00013A1D , 32'hFFFE68F6 , 32'hFFFC06F6 , 32'h00030FA9 , 32'h00039D74 , 32'hFFFD88BF , 32'hFFFEC662 , 32'hFFFCB92F , 32'h0004A076 , 32'hFFFFA85E , 32'h0003E68F , 32'h0000BB4A , 32'hFFFB995C , 32'hFFFF6E5F , 32'hFFFE968D , 32'hFFFF8F35 , 32'h0001CBEC , 32'hFFFE4E8C , 32'hFFFC9999 , 32'h0001702D , 32'h00051DF5 , 32'hFFF9ACE4 , 32'h00022B4D , 32'h00039146} , 
{32'h00002E26 , 32'h000107DD , 32'hFFFBA558 , 32'h000350BC , 32'hFFFEE7DF , 32'h00024496 , 32'h00060DF4 , 32'h00033FF8 , 32'hFFFAA17A , 32'hFFFEA504 , 32'h0000ED0F , 32'hFFFF68A2 , 32'hFFFE2059 , 32'h0002F064 , 32'h00050C78 , 32'h0005E9D0 , 32'hFFFFF0F7 , 32'h000318A2 , 32'hFFFD7AEF , 32'h00031C6F , 32'hFFFF9C58 , 32'hFFFD4D12 , 32'hFFF7F6B9 , 32'hFFFA6489 , 32'h00055DD4 , 32'h00083CBC , 32'hFFFBFDEF , 32'h00055707 , 32'h0000D045 , 32'hFFFFCF26 , 32'h00040D8E , 32'hFFF95555 , 32'h0001F23C , 32'hFFFC37FA , 32'hFFFD7AFD , 32'hFFFC0F11 , 32'hFFFE2DF2} , 
{32'h000295DB , 32'h00006438 , 32'h00007D92 , 32'hFFFF1E8E , 32'hFFFEAD15 , 32'hFFFEF88F , 32'hFFFAB358 , 32'h00053E24 , 32'h0003BE5E , 32'h000096E2 , 32'hFFFE6A39 , 32'hFFF91454 , 32'hFFFEFEAD , 32'h00060482 , 32'hFFFC4017 , 32'hFFFF7555 , 32'hFFFF5AFF , 32'hFFFDBDD6 , 32'hFFFD16C3 , 32'hFFFD3047 , 32'hFFFCCFCB , 32'h0001365D , 32'hFFFEBC71 , 32'h0000FE34 , 32'hFFFF00B3 , 32'hFFFDD4D2 , 32'h0001DC34 , 32'h0001DAC1 , 32'hFFFCB1B1 , 32'hFFF6C15A , 32'h0007CC18 , 32'hFFFF6C6E , 32'h00034B95 , 32'hFFFEA97B , 32'h00037A34 , 32'h00056B94 , 32'hFFFE44C2} , 
{32'h0004D686 , 32'hFFFDF838 , 32'h00047A1B , 32'h0002558C , 32'h000293BE , 32'hFFFBA045 , 32'hFFFE6A02 , 32'hFFFD75EF , 32'hFFFC442F , 32'hFFFFE755 , 32'h0005D4CE , 32'h0003525B , 32'h00031E1D , 32'h0003ED95 , 32'hFFF9552C , 32'h000234FB , 32'hFFFC0B99 , 32'hFFFEAE2F , 32'hFFFF362B , 32'hFFFF569A , 32'h00030B13 , 32'h00039525 , 32'hFFFEFC82 , 32'hFFFE7C32 , 32'hFFFC9BE7 , 32'h0001929F , 32'h000341F4 , 32'hFFFD9AB6 , 32'hFFFD7D14 , 32'h0004171A , 32'h00003B7D , 32'h000491D8 , 32'hFFFEA409 , 32'h00026ABA , 32'hFFFF76AD , 32'hFFFD6338 , 32'h0003404D} , 
{32'hFFFEAEC9 , 32'h00025CBF , 32'hFFFAE6A9 , 32'hFFFD6348 , 32'h0000A985 , 32'hFFFC465E , 32'h00035C10 , 32'h00030FCC , 32'h00044C11 , 32'h0000B545 , 32'h0004F419 , 32'hFFFFDEDB , 32'hFFFF2B1C , 32'hFFF9F155 , 32'hFFFC65A8 , 32'h00064802 , 32'h00041CC4 , 32'h0001F978 , 32'hFFFF2AD1 , 32'hFFFF4353 , 32'hFFFFB2F4 , 32'h00002BB4 , 32'h0000557B , 32'hFFFE5DA5 , 32'h00006A94 , 32'h00020B17 , 32'h00004ED6 , 32'hFFF7A9E0 , 32'hFFFCC2EB , 32'h00032E1F , 32'hFFFEA22D , 32'hFFFBBB9D , 32'h00053FF7 , 32'hFFFED2DE , 32'h0000FFF0 , 32'hFFFBE8DE , 32'hFFFD4321} , 
{32'hFFFCAB3C , 32'hFFF6D960 , 32'h00050816 , 32'h00099382 , 32'hFFFB7E0F , 32'h00010832 , 32'h00026B4E , 32'hFFFE72B6 , 32'hFFFF9DDE , 32'h0003C117 , 32'hFFFBF951 , 32'hFFF8A614 , 32'hFFFE5B16 , 32'hFFFED681 , 32'h00035844 , 32'h00086F66 , 32'h00036D94 , 32'h0000A0BE , 32'h0000735F , 32'h00012AA7 , 32'h00056DB7 , 32'hFFFF2CE8 , 32'h0001ECA5 , 32'hFFF9C5D7 , 32'h00051F58 , 32'h0001C89F , 32'h00046B0C , 32'hFFF6D2A3 , 32'h00042A4D , 32'h00017D6A , 32'hFFFDAFBD , 32'hFFFA21EA , 32'hFFF992A6 , 32'hFFFDFCF6 , 32'hFFF63E2A , 32'hFFF9CD48 , 32'h0003F49A} , 
{32'h0002E5BE , 32'h00061A68 , 32'hFFFE324C , 32'hFFFDC8F1 , 32'hFFFB6271 , 32'h0001E0C6 , 32'hFFFEE050 , 32'hFFFEA99D , 32'h000077EF , 32'h0006D065 , 32'h00007994 , 32'hFFFBF959 , 32'hFFFF32FD , 32'hFFFD8926 , 32'hFFFF485F , 32'hFFFC8130 , 32'hFFFD12BF , 32'hFFFF5114 , 32'h0000D061 , 32'h000063C0 , 32'hFFF8E045 , 32'hFFFE757C , 32'hFFFDF386 , 32'hFFFC21BD , 32'hFFFEB447 , 32'hFFFEE40A , 32'hFFFEEB93 , 32'h0001A28B , 32'h0001A866 , 32'h00014F8B , 32'hFFFE0CED , 32'hFFFE02A6 , 32'h000069D7 , 32'h00013801 , 32'hFFFC906C , 32'hFFFB3DA1 , 32'hFFFD13CE} , 
{32'h0000B043 , 32'hFFFA474D , 32'h0001D53C , 32'h00029212 , 32'hFFFD5874 , 32'hFFFD0474 , 32'hFFFCDD9D , 32'hFFFE32B9 , 32'hFFFEA590 , 32'h0003CBDE , 32'hFFFF9FCE , 32'h00032D3A , 32'hFFFEC067 , 32'hFFFFACA6 , 32'hFFFF1D11 , 32'hFFFEE7C7 , 32'h0000F422 , 32'h000162C7 , 32'hFFFEDF3A , 32'hFFFC7F97 , 32'h00041911 , 32'h00012EE8 , 32'hFFFCADE5 , 32'h00032B8D , 32'h00009591 , 32'hFFFD2ED0 , 32'hFFFD49D1 , 32'hFFFFEA5B , 32'h0002025F , 32'h0003692C , 32'hFFFDDA99 , 32'h00005607 , 32'h00008CEF , 32'hFFF94712 , 32'hFFFCED37 , 32'hFFFC7719 , 32'h000226DB} , 
{32'h00042E3D , 32'hFFFBDCD4 , 32'h00011DA7 , 32'h00057DCC , 32'h0003FE73 , 32'h00007D97 , 32'h000088CD , 32'h0003804E , 32'h00031A1A , 32'hFFFFC79D , 32'h000321D9 , 32'hFFFEC029 , 32'h0002BF16 , 32'hFFFE4839 , 32'hFFFF2932 , 32'hFFFFB239 , 32'hFFFF5245 , 32'h00007808 , 32'h0001538B , 32'hFFFF5AB0 , 32'h0002D8EB , 32'h00004643 , 32'hFFFFB859 , 32'h00067748 , 32'hFFFA7D08 , 32'h0000E478 , 32'hFFF9B1EE , 32'h0005F173 , 32'h00010454 , 32'h0003CD5A , 32'h00025582 , 32'h00069E41 , 32'hFFFBD585 , 32'h00017B08 , 32'hFFF932FC , 32'h00042BFF , 32'h0002B1DA} , 
{32'h0001EF02 , 32'hFFFF75A2 , 32'h0000166F , 32'h0000F68F , 32'h0000CAD2 , 32'hFFFF6283 , 32'hFFFE1C07 , 32'hFFFB33A6 , 32'hFFFE5444 , 32'hFFFB0852 , 32'hFFF85561 , 32'h0002CEFD , 32'hFFFC5C3E , 32'h0004A2F9 , 32'hFFFF618F , 32'h00036C99 , 32'h0001714C , 32'hFFFF7190 , 32'h0003207F , 32'h00009C37 , 32'h00011363 , 32'hFFF8B389 , 32'h00029CD0 , 32'hFFFF5C4C , 32'hFFFD9E8B , 32'h0001D89E , 32'hFFF92EF7 , 32'hFFFE907E , 32'hFFFC8291 , 32'h0002191B , 32'hFFFFE665 , 32'h0002A8C4 , 32'h00028B89 , 32'hFFFB43F7 , 32'hFFFD69C8 , 32'hFFFE92B9 , 32'hFFFEC00F} , 
{32'h0009CB95 , 32'hFFFDDF6F , 32'h0000F55B , 32'hFFFDEA3E , 32'h0000F428 , 32'hFFF8C3E6 , 32'h0003D510 , 32'h00023E41 , 32'h0003CE79 , 32'h00046382 , 32'h000284A9 , 32'hFFFFCB99 , 32'h00032ACB , 32'h00056B86 , 32'h000069DF , 32'hFFFEF029 , 32'h00004A94 , 32'hFFFF9250 , 32'hFFFCEBBA , 32'h0006368D , 32'hFFFFB27A , 32'h00026425 , 32'hFFFEC859 , 32'h00034C3A , 32'hFFFFC9D1 , 32'hFFFE7DDA , 32'h0002189F , 32'hFFFE5F27 , 32'hFFFFAAAB , 32'hFFFD86A9 , 32'hFFFD2CB2 , 32'h000139AF , 32'hFFFA366D , 32'hFFFDE81B , 32'h0004E3D0 , 32'hFFFE7F56 , 32'hFFFDACA5} , 
{32'hFFFC41DE , 32'h0002F0B4 , 32'h0001B4E6 , 32'h000647BD , 32'hFFFEC07B , 32'hFFFC76CE , 32'hFFFACB9E , 32'h0000D744 , 32'hFFFF416C , 32'h0003ABDA , 32'hFFFD9109 , 32'hFFFD5EE8 , 32'h0000ED93 , 32'hFFF9093B , 32'h00018BDE , 32'hFFFCA217 , 32'h0001C4E7 , 32'hFFFC0346 , 32'hFFFF499B , 32'hFFFBF6FA , 32'hFFFF1E43 , 32'hFFFC4654 , 32'h0003A479 , 32'hFFFF065A , 32'hFFFAF392 , 32'hFFFE6559 , 32'hFFFF6C83 , 32'hFFFDD2BF , 32'h00039E86 , 32'hFFFEE16B , 32'hFFFD8D73 , 32'h0003C5F1 , 32'hFFFE19A4 , 32'h00031F85 , 32'h0003EC7B , 32'hFFFEA761 , 32'hFFFFD7E0} , 
{32'hFFFC3D81 , 32'h00011154 , 32'h0006C9CA , 32'hFFFD8125 , 32'h00019A30 , 32'hFFFFEE39 , 32'hFFFE118A , 32'hFFFFE19C , 32'hFFFAC77F , 32'hFFFD575A , 32'hFFFE1A89 , 32'hFFFE6D36 , 32'h00019C83 , 32'h00000FC6 , 32'h000509FD , 32'hFFF7A15A , 32'hFFFF1E8A , 32'hFFF8F4DB , 32'h0001CD82 , 32'h0005A701 , 32'hFFFE358E , 32'h00021585 , 32'h0003FAB4 , 32'hFFFC1245 , 32'h0003CE5D , 32'h00021434 , 32'hFFFAA344 , 32'h0004F426 , 32'hFFFDC6EF , 32'h000041A1 , 32'hFFFD08B5 , 32'hFFFEB0CE , 32'h0003CA55 , 32'h000489B8 , 32'hFFFCC466 , 32'h0002A2EA , 32'hFFFE279E} , 
{32'h0004AE0B , 32'h00055A9C , 32'hFFFBFDF7 , 32'h0002209D , 32'h00028267 , 32'h00026F5D , 32'hFFFD2364 , 32'h0001AD08 , 32'h0006A680 , 32'hFFFE4E25 , 32'hFFFF8616 , 32'h00040CE0 , 32'hFFFB2A37 , 32'hFFFC25F6 , 32'h0000C7CF , 32'hFFFB65A6 , 32'hFFFF0799 , 32'hFFFF89C2 , 32'h0001AB70 , 32'hFFFEC108 , 32'hFFFF6F07 , 32'h0001FAD4 , 32'h0002D8F7 , 32'h00037ACE , 32'h000512FD , 32'h000190E4 , 32'hFFFC46D4 , 32'hFFFD894B , 32'hFFFAFADF , 32'hFFFE6BC4 , 32'hFFFD52EF , 32'h0005D6F1 , 32'hFFFF3B60 , 32'hFFFDE77B , 32'hFFFDF42C , 32'h0001CBCE , 32'h00019739} , 
{32'hFFFBD3E0 , 32'h0000A3DD , 32'h00060198 , 32'h00027E76 , 32'hFFFBD361 , 32'hFFFEFCAE , 32'hFFFCFCDC , 32'h00004675 , 32'h00016D6D , 32'hFFFB2B5A , 32'h0000FC95 , 32'h0003F142 , 32'hFFFFEDEF , 32'hFFFA62BC , 32'hFFFE443D , 32'hFFFEF102 , 32'hFFFEF035 , 32'hFFFD0A8B , 32'hFFFF7C9A , 32'hFFFC1371 , 32'h00018680 , 32'hFFF8754B , 32'h0009853C , 32'hFFFB41DE , 32'hFFFBE642 , 32'hFFF9FC08 , 32'hFFFC5E91 , 32'h0001F513 , 32'hFFFFAE92 , 32'hFFFC9069 , 32'hFFFCD10A , 32'hFFFE648A , 32'h0003E74B , 32'h0001B6B7 , 32'h0005D508 , 32'hFFFFF259 , 32'h0002A951} , 
{32'hFFFC6BA9 , 32'h000016DD , 32'h000616FE , 32'hFFFFEC87 , 32'hFFFFAC3F , 32'hFFFF1612 , 32'h00022106 , 32'hFFFFB749 , 32'h0001D559 , 32'h0001645A , 32'hFFFE48C4 , 32'hFFFFDC80 , 32'h0001967A , 32'h000008E7 , 32'h0001E59C , 32'h000095A3 , 32'h0005936E , 32'hFFF75539 , 32'h000434AE , 32'h0004ADA3 , 32'h0001113D , 32'hFFFDE2F6 , 32'hFFF9B907 , 32'hFFFC87CE , 32'hFFFD3CE9 , 32'hFFFE6BDB , 32'h0003626D , 32'h00024214 , 32'hFFFEAB6D , 32'h0003D472 , 32'h0000DE6A , 32'h00025408 , 32'hFFFEAFAE , 32'hFFFEB798 , 32'hFFFF5C67 , 32'hFFFCAC54 , 32'hFFFF0F2A} , 
{32'hFFFF8AF2 , 32'h0004B457 , 32'hFFFE1EE7 , 32'h00072DB9 , 32'h00022B8A , 32'hFFFE1617 , 32'h00008030 , 32'h000096F4 , 32'hFFFFD5BB , 32'h0001B011 , 32'hFFFD62A2 , 32'h00027FEC , 32'h00001AB0 , 32'h00037717 , 32'hFFFB37EE , 32'h0006B602 , 32'hFFF9ED7E , 32'h0002B05C , 32'h0004566A , 32'hFFFD97B8 , 32'h0000B391 , 32'h0000C1C6 , 32'h00023D2C , 32'h0002E62E , 32'h000539E6 , 32'hFFFE78C2 , 32'hFFFFFE6C , 32'h00000B71 , 32'hFFFF0818 , 32'h00026405 , 32'h0000BB02 , 32'hFFFDF9A2 , 32'h00013439 , 32'h00046901 , 32'h0003D6CC , 32'h00026373 , 32'hFFFFF102} , 
{32'h00010AB9 , 32'h00020D0A , 32'hFFFBAC48 , 32'h0005B8B7 , 32'hFFF79DCA , 32'hFFFE9481 , 32'h00061A7D , 32'h00008C1A , 32'h00019DF6 , 32'hFFFEB88F , 32'h0000E40C , 32'hFFFE96BB , 32'h00054993 , 32'hFFFED6EC , 32'h0000C9A3 , 32'h0000EAF1 , 32'h0006E0A3 , 32'h0001E21E , 32'hFFFBF7DC , 32'hFFFBCE1B , 32'hFFF8D313 , 32'h00017845 , 32'h00067EBA , 32'hFFFCD3A8 , 32'h000029A7 , 32'hFFFE8A94 , 32'hFFFB2BAD , 32'hFFFF9283 , 32'hFFF8FBC5 , 32'hFFFD178A , 32'h00005473 , 32'hFFFB04D0 , 32'h0001FE7C , 32'h00003500 , 32'hFFFE087B , 32'h0004C999 , 32'hFFFCC9B4} , 
{32'hFFFEAEB6 , 32'hFFFE1594 , 32'h0003D353 , 32'hFFFE0DD7 , 32'hFFFD189B , 32'h0002FC9B , 32'hFFFF1CE8 , 32'h0003AB3A , 32'h00001866 , 32'hFFFB0E79 , 32'hFFFE6D36 , 32'hFFFD62A2 , 32'h0004A4B6 , 32'hFFF6DCE7 , 32'h0007A7B1 , 32'hFFFAF786 , 32'hFFFD4D85 , 32'h0004FB4A , 32'h00047D87 , 32'hFFFD973D , 32'h00038984 , 32'h00041214 , 32'hFFFDC618 , 32'hFFF75CA8 , 32'h000081B7 , 32'h00015DEF , 32'hFFFFCC84 , 32'hFFF88460 , 32'hFFFCDAE4 , 32'h00016946 , 32'hFFFC9943 , 32'hFFFE38FD , 32'h00050A84 , 32'h0000CD11 , 32'hFFFB3477 , 32'h0001AAD5 , 32'hFFFD9986}
};

logic signed [31:0] US_1 [37][37] ='{
{32'hE943E960 , 32'h0E147B70 , 32'hD8748240 , 32'h1211A7E0 , 32'hF0B520C0 , 32'hBACA6100 , 32'h12FC2F00 , 32'h0F07FF40 , 32'h13D552E0 , 32'hBDEE6580 , 32'h12A75080 , 32'h12129220 , 32'h043A21B0 , 32'h1CCD3020 , 32'hD66F65C0 , 32'hDC06EC80 , 32'h27C16A40 , 32'h0CC65700 , 32'h2395B7C0 , 32'h1DCF0260 , 32'hB9326380 , 32'hE7CF4B40 , 32'h10960F60 , 32'h043D0808 , 32'h01FC7D2C , 32'h09E70DB0 , 32'h33D32BC0 , 32'hDFBF5480 , 32'h30AE0480 , 32'h0E681840 , 32'hE491F8A0 , 32'hFFAA14FD , 32'hF783BBE0 , 32'h1159E620 , 32'hCAC66A80 , 32'h0380F86C , 32'hA9579E00} , 
{32'hE809C760 , 32'h0D74F6D0 , 32'hB49BB200 , 32'hF0B86510 , 32'h22C00340 , 32'h1F5A4700 , 32'h299C2240 , 32'hEBA4B760 , 32'hFA13DFE0 , 32'hF1719B20 , 32'hF8E1AC20 , 32'h21C4A280 , 32'hED9C3D40 , 32'hEA32B5C0 , 32'hD5BA3B80 , 32'h0BD018E0 , 32'hFC2096EC , 32'hA5557400 , 32'h15F9BE20 , 32'h02D0BBC0 , 32'hCE56A7C0 , 32'h0F712B90 , 32'h05A070F8 , 32'h30FBC7C0 , 32'hEA775080 , 32'hE040AD80 , 32'hC0B7B500 , 32'h2D636380 , 32'h0A7B9DC0 , 32'hC2A28640 , 32'h1C179F60 , 32'hEEC33320 , 32'h25C69F80 , 32'h0BCFA930 , 32'hE04202C0 , 32'hE38A3420 , 32'h102F9480} , 
{32'hC82854C0 , 32'hC2857A40 , 32'hE043AA20 , 32'hDF6A51C0 , 32'h2D306F00 , 32'h071B9EE0 , 32'h2CE7A300 , 32'hFA579CB0 , 32'h2C7E4080 , 32'h10167A20 , 32'h255C0440 , 32'hCDD97640 , 32'hD4B03D80 , 32'h0E3B9860 , 32'h1AD62060 , 32'h38505080 , 32'h045DCA78 , 32'h39E3C080 , 32'h37A31640 , 32'hEFD86900 , 32'h3237E100 , 32'h0B54D590 , 32'h1B0F4100 , 32'h0647AF48 , 32'hFD1C7528 , 32'h15039360 , 32'hDF22CA80 , 32'h0C48AF50 , 32'hDB853340 , 32'hF8CC9238 , 32'hE4767220 , 32'h1F772860 , 32'h10D576E0 , 32'hF7692DE0 , 32'hDEB8D1C0 , 32'h070E1980 , 32'hC4E9FA80} , 
{32'hF8FD3E48 , 32'h12BE66E0 , 32'h13FB6260 , 32'hBC70AF00 , 32'h1497BCE0 , 32'hCEF37600 , 32'h01E86C38 , 32'hF96B7DB8 , 32'hF6790ED0 , 32'hEF4EA060 , 32'h50AF4380 , 32'h015B1B00 , 32'hCA7D5340 , 32'h0DD45E40 , 32'hE1562020 , 32'hF12B08F0 , 32'hEAEC6AC0 , 32'hFE2CC5F8 , 32'h0838C3C0 , 32'hF75A05A0 , 32'hFCA9DEA0 , 32'hE1F23720 , 32'h2511DD00 , 32'h145D0F00 , 32'h0DEC8730 , 32'hCE844A40 , 32'h12456CC0 , 32'h09709180 , 32'h034DDC20 , 32'h140911E0 , 32'h209D8380 , 32'h4142B600 , 32'hED128BC0 , 32'h1AA36640 , 32'h03394ABC , 32'h4CF7F100 , 32'h52385C00} , 
{32'h33AACB80 , 32'h069BDDE0 , 32'h20E952C0 , 32'h31E16400 , 32'hF01448D0 , 32'hD014CC00 , 32'hF10A4590 , 32'h0646A9D0 , 32'hF480E1F0 , 32'hB9651800 , 32'hCBB38400 , 32'hEFBBBF60 , 32'h174D3620 , 32'h1DFA9D00 , 32'hE71F7E40 , 32'h25DCEE40 , 32'hF9E9CC50 , 32'h2AC66440 , 32'h2431EEC0 , 32'hF863C5F8 , 32'h1899A5C0 , 32'hE4571A40 , 32'h2680D080 , 32'h0F111380 , 32'hEEE2AC80 , 32'hDF4BD700 , 32'hB02CA580 , 32'h1F61F880 , 32'h138D5360 , 32'hF0DE8B30 , 32'hD0E9D680 , 32'h023A8A40 , 32'h36DACC00 , 32'hDCE46AC0 , 32'hEF0BEA80 , 32'h1C04F0E0 , 32'h241A3480} , 
{32'hFC4C85D0 , 32'h1927F9E0 , 32'h2EA80680 , 32'hF42CA700 , 32'hF288FF30 , 32'hEC32A6C0 , 32'h00DA47E7 , 32'hD5AE0640 , 32'hEEFA5B20 , 32'h0A8DDE00 , 32'hDAA47940 , 32'h3AB39B80 , 32'h0492FDD8 , 32'hFD5E12BC , 32'h00869973 , 32'h0CD17DE0 , 32'hF9D386D8 , 32'hDA4FA680 , 32'hF138AFC0 , 32'h12F29320 , 32'h55441F80 , 32'h260EA180 , 32'hED1E3AC0 , 32'h0AA59630 , 32'hF8B39510 , 32'h0D8F1AC0 , 32'h00DFECBB , 32'hE41D4A20 , 32'hFE57CB34 , 32'hDC20E5C0 , 32'hF766BA00 , 32'h17370AC0 , 32'h1E477E20 , 32'h5C5C1F80 , 32'hCCD33C40 , 32'h480AEE80 , 32'hC8F19580} , 
{32'hF26D22F0 , 32'h3DA58280 , 32'hED984360 , 32'hF07F4F50 , 32'h1E5421A0 , 32'hEAACE7E0 , 32'hD9488CC0 , 32'hEB93D9C0 , 32'hF70F40A0 , 32'h1D876AE0 , 32'h49A10380 , 32'h11B20C20 , 32'h181BF2A0 , 32'h39F59CC0 , 32'hD2FCE800 , 32'hF54990B0 , 32'hF198D700 , 32'h09A138F0 , 32'h0A38FDB0 , 32'hD7DBFBC0 , 32'h16D13C00 , 32'h1BCE65C0 , 32'hF629CDA0 , 32'hDC3D5B40 , 32'h31D3BC40 , 32'h32D84DC0 , 32'hCD87BAC0 , 32'hE3E32F40 , 32'h0B5E42D0 , 32'hF9F44140 , 32'h04CC1508 , 32'hA176F380 , 32'h181C0E40 , 32'hDB725240 , 32'hFC950464 , 32'h14A127C0 , 32'hFFBC0694} , 
{32'h0E3549A0 , 32'h1BAE7B80 , 32'hF1970A00 , 32'hEC292B00 , 32'h365A12C0 , 32'hEFD4C680 , 32'hE5D11780 , 32'hEBAF88E0 , 32'hEA13BC80 , 32'hFA3E0940 , 32'hD4F18280 , 32'hFC0F9DC4 , 32'hE04D1600 , 32'h0176708C , 32'hEC661160 , 32'h0351467C , 32'hAF9BE100 , 32'hE829B480 , 32'h25B3B980 , 32'h24458500 , 32'h2EC55A00 , 32'hCB6D5940 , 32'h09EA3C40 , 32'hECDF9840 , 32'hCB74EBC0 , 32'h4BF06C00 , 32'h322AF7C0 , 32'h028C86E4 , 32'h16DA2DE0 , 32'h25B933C0 , 32'h26243F80 , 32'h19F35960 , 32'h1DC8B0E0 , 32'hD9A2F6C0 , 32'hF44193C0 , 32'hCBF72240 , 32'hFC7ACE60} , 
{32'hC639EE00 , 32'hC4A2F700 , 32'h28214440 , 32'hD0CC8880 , 32'hD78C3300 , 32'hE73F5840 , 32'hFCD6BD20 , 32'hF1EDE8E0 , 32'hD7494180 , 32'h15DE1E20 , 32'hD7FEFB00 , 32'h3ABABF40 , 32'hFB7A6738 , 32'h1F269720 , 32'hF79B8C60 , 32'hD8466F40 , 32'hEBB11F80 , 32'hEAB8E580 , 32'h260A0700 , 32'hDB66E7C0 , 32'hF32008F0 , 32'hCC3F1A80 , 32'hF72ECFD0 , 32'hFE5F2818 , 32'h097C3F70 , 32'hEC4BA760 , 32'hCC71BAC0 , 32'hB87F3B00 , 32'hE5586120 , 32'hE7C9B9C0 , 32'hED8FBEC0 , 32'h1BE5DD80 , 32'hE1590E40 , 32'hD2A0B780 , 32'h071774F0 , 32'hD4FB3A80 , 32'hF7801C00} , 
{32'h1299B740 , 32'h06713D58 , 32'hF2B76160 , 32'hF813F1A0 , 32'h0C944A10 , 32'h4ED67000 , 32'h263A1040 , 32'hEB6433E0 , 32'h1A4037E0 , 32'h03C6B2C0 , 32'hE88D1A00 , 32'h10346F40 , 32'hFC9C1930 , 32'h34578E40 , 32'hB3DA9300 , 32'h0021EA2D , 32'h09624950 , 32'h3166F2C0 , 32'h088CB1B0 , 32'hEDD54B40 , 32'h204A1200 , 32'hC2565500 , 32'hB5898A00 , 32'hBBE41300 , 32'hF4D1C980 , 32'hB1D94480 , 32'h13303020 , 32'h0E3EAEC0 , 32'h0D0F2FB0 , 32'h08DBB3B0 , 32'h0B27F680 , 32'hF8EB1FF8 , 32'hF7489D30 , 32'h1CCDB8A0 , 32'hF6D24C30 , 32'hFFC85C3D , 32'hF7FDE4F0} , 
{32'hD088DF80 , 32'hAD3B3500 , 32'h06B231A8 , 32'h010CA0FC , 32'hFE35449C , 32'hEE812840 , 32'h102A3B40 , 32'h20813700 , 32'h072B66D0 , 32'hE400D220 , 32'hD3833E80 , 32'hF8699CA0 , 32'h0504A660 , 32'hF381A7E0 , 32'h04515408 , 32'h05889910 , 32'hDAD04440 , 32'h15F77140 , 32'hDFA00C80 , 32'h242D9880 , 32'hEDE4AE20 , 32'hED87BAE0 , 32'hE532C820 , 32'hD8477480 , 32'h2FD2DB00 , 32'h286716C0 , 32'hF9202EE8 , 32'h13CB0580 , 32'h16EEC6A0 , 32'hE2D64160 , 32'h54D79D00 , 32'hD0D6F780 , 32'hF5046510 , 32'hF82B9270 , 32'hC2B646C0 , 32'h3CC2A640 , 32'h24992140} , 
{32'h1B192840 , 32'hDA902040 , 32'hF7220970 , 32'h1FC122C0 , 32'hFA6CE6F0 , 32'hB8EBDF00 , 32'hDF4DA680 , 32'h0537E300 , 32'hF58ADF60 , 32'h22154280 , 32'h1B1F6EC0 , 32'hF7E85BD0 , 32'hE48FB1C0 , 32'h03FA8044 , 32'hF65F3130 , 32'h306A2280 , 32'h15CA6C80 , 32'hEADF6F80 , 32'hEF877560 , 32'h23A1B000 , 32'h254B3240 , 32'hCA3ADB80 , 32'h0ED698A0 , 32'h18EA07A0 , 32'hFAB4E668 , 32'hC4BC0040 , 32'hDDE38E80 , 32'hFA750C88 , 32'hEADBBCC0 , 32'h1C746D40 , 32'h4FEE4B80 , 32'hC2403D00 , 32'hEDF72820 , 32'h24B91840 , 32'h1B77C0C0 , 32'hDE55F8C0 , 32'hC7AAC180} , 
{32'hFC1DEA00 , 32'hEE96B080 , 32'h1F2D6D40 , 32'h1ED66640 , 32'hF181D220 , 32'hFFE6216E , 32'h210D2200 , 32'hFF1EB3E2 , 32'h1277DE60 , 32'h2DDEBBC0 , 32'h40E15400 , 32'h49558A80 , 32'h176AA420 , 32'hE7EBFC80 , 32'h02D571FC , 32'hDA09C840 , 32'hE9A057C0 , 32'h44906200 , 32'h04DB9690 , 32'h3F9544C0 , 32'hF06BB940 , 32'h1DA88200 , 32'hE04A86A0 , 32'h0F787D20 , 32'hC9B073C0 , 32'hFB108CF0 , 32'hCF727C80 , 32'hFFB37020 , 32'h23655340 , 32'h2984C480 , 32'h257F5340 , 32'h23A23FC0 , 32'h3D501140 , 32'hEC495100 , 32'hFCD6E008 , 32'hF06D69C0 , 32'h046CC810} , 
{32'hBE73C380 , 32'h269A7000 , 32'hA579B100 , 32'h4DF4EB80 , 32'hD819F900 , 32'hC3D63F00 , 32'h22C6B5C0 , 32'h02BC4158 , 32'hCE45A800 , 32'h22C9AF80 , 32'hF4C952B0 , 32'hE7D7F1E0 , 32'h0B941EF0 , 32'h1B726520 , 32'h0DA1EE90 , 32'h1224D9E0 , 32'hE8802BA0 , 32'hFDBB29F8 , 32'hF1A30C90 , 32'hF19F3520 , 32'h168EE080 , 32'h195346C0 , 32'hD9ED6C40 , 32'hE99A8200 , 32'hE1CB92E0 , 32'hD9345880 , 32'h1E9510C0 , 32'hF2F31E10 , 32'hDC572E80 , 32'hFE646604 , 32'h09C21E60 , 32'h25A9E840 , 32'h02AC91C8 , 32'hDF673D00 , 32'hFBAB2A30 , 32'h17524220 , 32'h1DF01580} , 
{32'h05FDF658 , 32'h0786E698 , 32'h03928AF0 , 32'hD7A64A40 , 32'hC07E8CC0 , 32'h0175EEBC , 32'hFE0CBB60 , 32'hC2106540 , 32'h21CAFBC0 , 32'h044529C8 , 32'h07E50FD0 , 32'hE0F93F00 , 32'hCE96E140 , 32'h22562440 , 32'hFB8F41A8 , 32'hFDDCBF18 , 32'h298BB480 , 32'hEEC65F20 , 32'h94CA2C80 , 32'h1EC68B80 , 32'hE1D67A80 , 32'hE9311860 , 32'h2394C580 , 32'hC84F9800 , 32'hCDCC3C80 , 32'h0FA95960 , 32'hEEDB6300 , 32'hFCEBAF08 , 32'hE63904A0 , 32'hEF606040 , 32'hFC66A8F0 , 32'h0634AAD8 , 32'h36211A80 , 32'hD38251C0 , 32'hEB1E71A0 , 32'h05BA4FB8 , 32'hF8A298A0} , 
{32'h14A8A500 , 32'hEF648560 , 32'h0CCFAC80 , 32'hDBFDD300 , 32'h0FD52740 , 32'hDD50E3C0 , 32'h2EA23AC0 , 32'h0B753A70 , 32'hDB962C40 , 32'hFAB50978 , 32'hFC66C604 , 32'h03E9F2B0 , 32'h17F9AF40 , 32'h32858100 , 32'hEB9ABF00 , 32'hF5540030 , 32'hB0DBC400 , 32'hF6ADB530 , 32'hD93ABD80 , 32'h31128C40 , 32'hF1628CD0 , 32'h38E475C0 , 32'h11A4D7E0 , 32'hD815D900 , 32'h318FAC80 , 32'hE249CE80 , 32'h00B7687A , 32'h553C8E00 , 32'hEAF62D80 , 32'h026D0B34 , 32'hDDA2FA00 , 32'h0DA81290 , 32'hF98DBE00 , 32'hFDD7E18C , 32'h2DF13900 , 32'hE7F8DFE0 , 32'hC52E9A00} , 
{32'h08BDC460 , 32'hFAEDCEC8 , 32'hE7B57EE0 , 32'h12BD29E0 , 32'h0BC19700 , 32'hFFE33ADC , 32'hC2B86840 , 32'hD8664400 , 32'hFBDFEB10 , 32'hEB0E9A80 , 32'hF1D631F0 , 32'h0FF65400 , 32'hC7E7F940 , 32'hF5DB5560 , 32'hC4175D80 , 32'hFFD7EEF4 , 32'h223DCDC0 , 32'h3B7C5880 , 32'hF9669CD8 , 32'h4B19E100 , 32'h0FC7FB50 , 32'h2C4273C0 , 32'hDD5BA340 , 32'h27D5F940 , 32'h4E103A00 , 32'hFFCE3009 , 32'h136589A0 , 32'hEDEBF780 , 32'hD2576500 , 32'hCEAD0B80 , 32'hFEF58738 , 32'h25386F00 , 32'hFC2CB2D0 , 32'hE3B79DE0 , 32'h00DEF34D , 32'hDA0BD700 , 32'h18561800} , 
{32'h13FB6C20 , 32'h2D9C1400 , 32'h0A061130 , 32'hF9DDB360 , 32'h3866BD40 , 32'hDB4AF080 , 32'h11B189A0 , 32'h4079A100 , 32'h1FED4840 , 32'h1B0FEDC0 , 32'h09BF4B50 , 32'h2F515F40 , 32'hF0B28FC0 , 32'hEBF210C0 , 32'h3937D1C0 , 32'hEC1D3FA0 , 32'h0FEFA4C0 , 32'hF6E976A0 , 32'h139AB5C0 , 32'h3E7C1C40 , 32'h0021A659 , 32'hC41E33C0 , 32'hE5847C00 , 32'hDCB1ED40 , 32'hF3F14970 , 32'hEFA50720 , 32'h082C84D0 , 32'h09AAFAD0 , 32'hB4452F00 , 32'hCA87B8C0 , 32'hC8A11C00 , 32'hDAD40CC0 , 32'h01430AA8 , 32'hECD35D60 , 32'hEC334860 , 32'h0C905320 , 32'h16327BE0} , 
{32'hC63169C0 , 32'h2FD8A4C0 , 32'hF0750460 , 32'hEA48FCC0 , 32'hD5472E40 , 32'h1D63C6A0 , 32'h0F4D0320 , 32'hFFBAFA35 , 32'h1BF9DE40 , 32'h3AD90080 , 32'hBF78BE00 , 32'hF993C950 , 32'h0CBC8A40 , 32'hD108E040 , 32'hD3A11F00 , 32'hF734FBF0 , 32'hF8701CE0 , 32'h126EEF60 , 32'h1E8FA420 , 32'h42C90380 , 32'h0E173FE0 , 32'hFC10CADC , 32'h5DFCCC00 , 32'h04658E18 , 32'h1EF45660 , 32'hE8826840 , 32'hF77E65F0 , 32'hF5F09710 , 32'hF9712CA0 , 32'h3809B740 , 32'hEDDF0020 , 32'hD728DC00 , 32'hF7DAD2D0 , 32'hFF6A706B , 32'h0F3003F0 , 32'h1DC850C0 , 32'h0C74C740} , 
{32'h07B18A80 , 32'h25DCF300 , 32'hE3E348A0 , 32'hED986500 , 32'h2CBCC300 , 32'h1E3F8700 , 32'hF53761E0 , 32'h2CF34600 , 32'hEC61D420 , 32'h022D2AFC , 32'hFA51C668 , 32'h13076240 , 32'h41910C00 , 32'hF138CA60 , 32'h04BF0790 , 32'hEB482340 , 32'h1808D180 , 32'h11BE5780 , 32'hB0C94480 , 32'hEBF2E880 , 32'h2441F900 , 32'hD561CA80 , 32'h22F88F00 , 32'h2B8FA100 , 32'h18C91420 , 32'hEDB04880 , 32'hEA6710A0 , 32'h046D19D8 , 32'h0436F018 , 32'hFA832BC0 , 32'h28BF8580 , 32'h3CE95F00 , 32'hE8CFF9E0 , 32'hBA390680 , 32'hD45E7EC0 , 32'h11820560 , 32'hC510A000} , 
{32'hFD078390 , 32'h0F13E860 , 32'h0A915B90 , 32'h363D2E80 , 32'h11B70020 , 32'h16588F00 , 32'hE314C4E0 , 32'hFDDC841C , 32'h01FCD238 , 32'hF6D24180 , 32'hFD6C5C10 , 32'hEDB61BC0 , 32'hAA768480 , 32'hE40A62E0 , 32'hE8B29A40 , 32'hDEBA4140 , 32'hDD6F4AC0 , 32'hE69FDE00 , 32'hFA352E78 , 32'h0AA4BC20 , 32'hF1AF01E0 , 32'h0F870010 , 32'hD78FFBC0 , 32'hF70113C0 , 32'hDA4AE2C0 , 32'h07203998 , 32'hB6DBF600 , 32'h0EA40A40 , 32'h07834448 , 32'h200D1100 , 32'hE1BCBE20 , 32'h06953F38 , 32'hA3EC0E00 , 32'hDE077B40 , 32'h0364C2AC , 32'h44C4C480 , 32'hCE48D8C0} , 
{32'h58F6E100 , 32'hEB2A1D40 , 32'hD7D46740 , 32'h0B905B10 , 32'hE4FC9320 , 32'h01F92374 , 32'h1A00E660 , 32'hD1995740 , 32'h401B7100 , 32'h0F3DE6D0 , 32'h0688E080 , 32'hE7D64400 , 32'h2C67AC40 , 32'h1E29B860 , 32'hFC7DEA48 , 32'hCB3A14C0 , 32'hAF015100 , 32'h099928E0 , 32'h0B530020 , 32'h0053F328 , 32'hFDE87ED4 , 32'hFCA5B2D0 , 32'h14C0F7C0 , 32'h37DBC780 , 32'hED2D1F20 , 32'h0E2C2140 , 32'h03741A04 , 32'hDC567700 , 32'hC737CDC0 , 32'hDD2497C0 , 32'h0EA1E300 , 32'hF2BD03C0 , 32'hCE19E440 , 32'h09CF7620 , 32'hE0FDED40 , 32'h0F768650 , 32'h09335290} , 
{32'h45849E00 , 32'h166EBAE0 , 32'hDFA3B540 , 32'hC0DDE380 , 32'hB2B0B800 , 32'hE8F0B580 , 32'h4F236300 , 32'h347152C0 , 32'hD39C7D40 , 32'hFBA645E8 , 32'hFA0615A8 , 32'h1C134F00 , 32'hCD0545C0 , 32'hCF4D5940 , 32'hDFD83040 , 32'h2336BC40 , 32'h0C12E5F0 , 32'h24680440 , 32'hFBC73678 , 32'hDF466F80 , 32'h0D9BCD30 , 32'h03076BE4 , 32'hDC66C780 , 32'h15C5D5E0 , 32'h0084E2DF , 32'h3A849C00 , 32'hF32CBEF0 , 32'h02A0024C , 32'hF586B170 , 32'h0FE062A0 , 32'h00CE1A80 , 32'hED6E99C0 , 32'hF0E44430 , 32'hF2F96420 , 32'h057602D8 , 32'h0030EEDF , 32'hFBB73DE8} , 
{32'h08DE0C40 , 32'hE9B2FEC0 , 32'hCE4B7800 , 32'hD0EAF200 , 32'h1114D6E0 , 32'h12728C40 , 32'hF7036090 , 32'hCDE5FA00 , 32'hC9C7E1C0 , 32'hD78E8100 , 32'hF36DD180 , 32'h047FD630 , 32'h2794E200 , 32'h28E277C0 , 32'h3A2A1D00 , 32'hFCE8AD94 , 32'h27533640 , 32'hF5059B50 , 32'h096C8D20 , 32'h35879100 , 32'hF545D840 , 32'hF5C91210 , 32'hCD756B80 , 32'h1D09F860 , 32'h0394F070 , 32'h08563130 , 32'hE05DD340 , 32'h02A36B74 , 32'hD803CA80 , 32'h6C7FFA80 , 32'hEA4407E0 , 32'hEF3CC460 , 32'h00ADA6D7 , 32'h07054B70 , 32'hEF440340 , 32'h20010680 , 32'h16B49CA0} , 
{32'h0209B240 , 32'hFD3C71D4 , 32'hE1DEE1A0 , 32'h084018F0 , 32'hCBF693C0 , 32'h1AA8C020 , 32'hE445FA40 , 32'h1EA259C0 , 32'h5CF06400 , 32'hC349A980 , 32'h10053840 , 32'h475FA800 , 32'hE4313800 , 32'h07135110 , 32'h2583A880 , 32'h2B2053C0 , 32'hC55FEFC0 , 32'hCC2D3180 , 32'hFCBD96F8 , 32'hEF6B13C0 , 32'h19132BA0 , 32'h059A72B8 , 32'hF6977A00 , 32'hFE3A7220 , 32'h37511100 , 32'hDEF90D00 , 32'h0EAEC0F0 , 32'hEE544DE0 , 32'hF9633330 , 32'h2F620580 , 32'hFF1FF02B , 32'h076268F0 , 32'h24B22DC0 , 32'hD8E50140 , 32'h083CF380 , 32'h06ED06E8 , 32'hF426C680} , 
{32'hD0347940 , 32'hF2DFA740 , 32'h059C27D8 , 32'h10DF3DC0 , 32'h2E777140 , 32'hFE2238E8 , 32'hF9C658F8 , 32'h0033B002 , 32'h0075EDAE , 32'hD08D2480 , 32'hE16E1CA0 , 32'h4C2FF480 , 32'hEC825980 , 32'h0AA2D5F0 , 32'hE871A9A0 , 32'hF541D670 , 32'hF4642770 , 32'h3A1CBB00 , 32'hCB165480 , 32'hC79FAB40 , 32'hF1CE5280 , 32'h0F149A60 , 32'h29234980 , 32'h231655C0 , 32'hBC023580 , 32'h0CE00170 , 32'h20147400 , 32'h0D721DD0 , 32'hB1CA7900 , 32'h164EE320 , 32'h055BB570 , 32'hCAED5600 , 32'h083F3320 , 32'h1220F480 , 32'h232C94C0 , 32'h0B6CD310 , 32'h006A06A6} , 
{32'h170F7D80 , 32'h0E413EC0 , 32'hF22C5120 , 32'hFF0CF0CA , 32'h39CC2C80 , 32'hB2483D80 , 32'h31F36680 , 32'hA0991180 , 32'h33E6E300 , 32'hED751700 , 32'hD7AF8080 , 32'h15062860 , 32'h0916DB60 , 32'hB54AED00 , 32'h1DCBAEA0 , 32'hFD37A41C , 32'h14D76A00 , 32'h0B4CBF70 , 32'hF256D140 , 32'hD6D2AC00 , 32'hFD9F8658 , 32'h1141C1E0 , 32'h02ED2BE0 , 32'hC5DBF080 , 32'h205C9100 , 32'hEE8B6DA0 , 32'hE3B7D7A0 , 32'hEAE990A0 , 32'h1305A0A0 , 32'h1A627B60 , 32'h0FF7F990 , 32'h0CAD0180 , 32'hE78B8FC0 , 32'hF6DEF910 , 32'h121441C0 , 32'hED32B7C0 , 32'h077D84F0} , 
{32'h0D6974D0 , 32'h04944DF8 , 32'h04C4E258 , 32'hC5280C00 , 32'hFB4AA608 , 32'hF8CA4038 , 32'hED6B1E60 , 32'hFF517F8F , 32'h043F1218 , 32'h01AD6F50 , 32'hE6C5F7C0 , 32'h1A2B8660 , 32'hECA6E7A0 , 32'h2DE1F8C0 , 32'h30DE0F40 , 32'h11F9EFA0 , 32'h16D06FA0 , 32'h1377EE60 , 32'h1B2F7960 , 32'h12B3C060 , 32'h14525A20 , 32'h5680FE00 , 32'h112F29E0 , 32'h07C94370 , 32'hC1C36540 , 32'hC57697C0 , 32'h223F2C80 , 32'h03D7C690 , 32'h3DFF5440 , 32'hE7118120 , 32'h1BC463C0 , 32'hD317F140 , 32'hC04E4BC0 , 32'hC260BBC0 , 32'hE5B2D680 , 32'hFF06CAD0 , 32'h052BF850} , 
{32'h0DA94440 , 32'h1C0403C0 , 32'h35B1E100 , 32'h19EB0F80 , 32'hE96EC780 , 32'h0DFDFBF0 , 32'h07480B30 , 32'h0E2E88B0 , 32'h02BE8414 , 32'hEABA56C0 , 32'h01963A10 , 32'h06C0E8B0 , 32'h1166ACA0 , 32'h0EC29D10 , 32'hEA537A20 , 32'hFC13AFFC , 32'h33A29E40 , 32'hE06A66E0 , 32'h47581780 , 32'hF325A3C0 , 32'hF4E64600 , 32'h2D40B540 , 32'h1A6FB140 , 32'hC867DD40 , 32'h04266E90 , 32'h13267EA0 , 32'hF8212C88 , 32'h21BFE500 , 32'h9ED5B980 , 32'h1F1F4840 , 32'h56370C80 , 32'h20331440 , 32'hECE921C0 , 32'hF3847400 , 32'hD1FDA9C0 , 32'hF3293350 , 32'hF91861B0} , 
{32'hF9AB8730 , 32'hE6E40780 , 32'hF681CEF0 , 32'hCB8BA7C0 , 32'h0208BD4C , 32'h02DF6634 , 32'hECF33460 , 32'h12972A60 , 32'hF3164BC0 , 32'hB4289F00 , 32'h20D2B8C0 , 32'hCEDA9940 , 32'h3A691BC0 , 32'hAE14F800 , 32'hD4BAB400 , 32'hF421F1A0 , 32'hF4498130 , 32'hF56BF460 , 32'h1123A020 , 32'h17540520 , 32'h19A54D00 , 32'h1B8A4480 , 32'hE9982860 , 32'hD9BEE900 , 32'hC8D18A40 , 32'hD7129680 , 32'h05AFF3B0 , 32'hC29CA280 , 32'hDEA28000 , 32'hE61A11A0 , 32'h09756370 , 32'hF14507A0 , 32'h1B51C1A0 , 32'hE8C4E240 , 32'h2A94CB00 , 32'h193A1580 , 32'hE78D16E0} , 
{32'h19453380 , 32'hEA4386C0 , 32'h1AC12A00 , 32'h0944E8E0 , 32'h173CC040 , 32'h04F874D8 , 32'h039E1C64 , 32'h0C3D96E0 , 32'hD2534B00 , 32'h126DB7E0 , 32'h088F64A0 , 32'hE27929A0 , 32'hD8B46380 , 32'hD89F4FC0 , 32'hF50E0F30 , 32'hE97127A0 , 32'hDE0E5100 , 32'hFDC88750 , 32'hE4036AC0 , 32'hDF4D2440 , 32'hF98B6330 , 32'h20D0E180 , 32'h0BBFF910 , 32'hFC679400 , 32'h137010C0 , 32'hC126E240 , 32'h167AD360 , 32'hD9C5FE40 , 32'hF16CABC0 , 32'h36912F00 , 32'hDAA80F80 , 32'hDA0E3580 , 32'h2461A9C0 , 32'hFBAB4570 , 32'h82118580 , 32'hD8788100 , 32'h09D9EC60} , 
{32'h1448D6A0 , 32'hD0D9CDC0 , 32'hE6E728C0 , 32'hEEFC3D60 , 32'h2410CE80 , 32'hD5F7B740 , 32'hFC259F0C , 32'h5176AA00 , 32'h401A1080 , 32'h25D76C00 , 32'hC834DB80 , 32'hEB42EDC0 , 32'hF7CC2980 , 32'h2B4DE640 , 32'hCFC6EB00 , 32'hBFBAF080 , 32'h3353C080 , 32'hD24AC740 , 32'hF08681E0 , 32'hF31955B0 , 32'h20186340 , 32'h303B7F40 , 32'hECE2EA80 , 32'h09BE80F0 , 32'hF36A76D0 , 32'h0DD22C40 , 32'hEE56D060 , 32'hEED0FAC0 , 32'h0B6033E0 , 32'h240FBAC0 , 32'hFB94E5B8 , 32'h18599EA0 , 32'h21952840 , 32'h07E75BC8 , 32'h13DAF9A0 , 32'h07EA26C8 , 32'h1D14E240} , 
{32'hDB6B0100 , 32'h095AA0F0 , 32'hF8C7A920 , 32'hFD5F8290 , 32'hF8F02A88 , 32'hFBA32FB8 , 32'hFE990CD0 , 32'h1DB9FDE0 , 32'h1896E840 , 32'hD54C71C0 , 32'h24BECBC0 , 32'h0F084570 , 32'h23ED0000 , 32'h0702AEE8 , 32'hE4F0EE80 , 32'h27FA7B80 , 32'hF75748E0 , 32'hFA8D1968 , 32'hCD78D400 , 32'h1F3C28C0 , 32'h2F6369C0 , 32'h0841EE40 , 32'h0EE63C80 , 32'hE3B7C640 , 32'hDEB97A80 , 32'h1A9BCD80 , 32'hD1E9DF40 , 32'hF0925360 , 32'h07A2EAC0 , 32'h0C125240 , 32'hD66C5AC0 , 32'h0F54DBB0 , 32'hAA1A2A80 , 32'h31E5C280 , 32'hD5403840 , 32'hAF9D9F00 , 32'h3C10FDC0} , 
{32'hFAE3B118 , 32'hF79572A0 , 32'hD4E07380 , 32'h151997E0 , 32'hDBDB7700 , 32'h1353CE40 , 32'h0B257990 , 32'hFF786282 , 32'hDC98B100 , 32'hCC4C08C0 , 32'h125421C0 , 32'h03A30FB0 , 32'hD1BD0380 , 32'hFB82C9E8 , 32'h3615BB80 , 32'h80000880 , 32'h0F756D60 , 32'h0BDE67B0 , 32'h0BF53EA0 , 32'hFD6898C0 , 32'h55A6D180 , 32'hF978FE50 , 32'h2B0DE200 , 32'hE13A4880 , 32'h0ED59340 , 32'hFDC20FDC , 32'hED89C500 , 32'h1FB6B980 , 32'h11B5EC60 , 32'hEBF19460 , 32'h0C42A660 , 32'hEC8559A0 , 32'h0B98B780 , 32'h1C3C6580 , 32'h0BE5DA70 , 32'hE70F8460 , 32'h047F04A8} , 
{32'hC5353BC0 , 32'h36AB0040 , 32'h26843940 , 32'hD1CB6D00 , 32'hD7F53A80 , 32'hD0CAFEC0 , 32'hE379DC40 , 32'hF190A1D0 , 32'h37C3B2C0 , 32'hF2BA6210 , 32'hF4279310 , 32'hC99E5640 , 32'h0F5D6F00 , 32'hED0025E0 , 32'h05D0C9D8 , 32'hD7290300 , 32'hF0E1E2A0 , 32'h0E44CF80 , 32'hFCA31454 , 32'hE5841DA0 , 32'h0ED7C9B0 , 32'hF5B7CD50 , 32'hB0B73780 , 32'h3E66F2C0 , 32'hFEB58850 , 32'hF0737890 , 32'hFE9436A8 , 32'h4F5D5B00 , 32'hF0D42740 , 32'h0A6C4800 , 32'h07A1D4F8 , 32'hEC62EDC0 , 32'h063D44E8 , 32'h023814B4 , 32'hE79D0CC0 , 32'hD5DBC700 , 32'hF1C7EE80} , 
{32'h02799658 , 32'hB1BD4180 , 32'hFA173DE8 , 32'h14666DC0 , 32'hEACC0740 , 32'hEDEFC700 , 32'hF7208210 , 32'hD090E400 , 32'h0121E1DC , 32'h1E8A3C00 , 32'h28C53800 , 32'h2BB82980 , 32'h25D53180 , 32'hD4CA2D80 , 32'hCBD1DF40 , 32'hFDEDB94C , 32'h24E85380 , 32'hD27FA880 , 32'h081E3070 , 32'hF12C91A0 , 32'h312AD100 , 32'hED53D5A0 , 32'h05E77130 , 32'h01EEA3EC , 32'hF6A0B0C0 , 32'h0EF7AF20 , 32'h39034E80 , 32'h54240D80 , 32'h07250BE0 , 32'h07AFA5A0 , 32'hCC4EFC80 , 32'hF1285FB0 , 32'hEB1B4060 , 32'hC6C53080 , 32'hED7972A0 , 32'h17DFCA60 , 32'h0D766E60} , 
{32'hE7693160 , 32'h0ECAC270 , 32'h4AE7D400 , 32'h25602C40 , 32'h18BA4EA0 , 32'h11422100 , 32'h7657F700 , 32'hF00218F0 , 32'h0296970C , 32'hD588AB40 , 32'h10485760 , 32'hE2683DC0 , 32'hF58E6D00 , 32'h21677740 , 32'hF55D1F30 , 32'hFE2FE638 , 32'h156C75E0 , 32'hD3C3D800 , 32'hED96BEE0 , 32'h1EFEB7A0 , 32'h2EED8FC0 , 32'hF9B1DDF0 , 32'hF4F936B0 , 32'h3DBB8BC0 , 32'h12944FE0 , 32'h06A25DD0 , 32'h15C03AE0 , 32'hD5377D00 , 32'h0810EA40 , 32'h05F60C68 , 32'h07549EF8 , 32'hDDCEDA40 , 32'hFB597400 , 32'hC8887E00 , 32'h1B1ADCE0 , 32'hF970EE00 , 32'h0AD795F0}
};

logic signed [31:0] US_2 [300][100] ='{
{32'hF8CA1178 , 32'h9FEF0C80 , 32'h292E3B00 , 32'h1CFEDC40 , 32'h0B9A2400 , 32'hF2AFD410 , 32'h15E70060 , 32'h011A89B8 , 32'hE3DC0BC0 , 32'hE5A73820 , 32'hEA952040 , 32'h0EB115A0 , 32'h07DFB280 , 32'hEAA8FCE0 , 32'h0D0215C0 , 32'hF9CF1E90 , 32'hEEC07EA0 , 32'h0949EB50 , 32'h04CE1DE0 , 32'hF804F980 , 32'h024051B8 , 32'hEE6CA200 , 32'h16917B60 , 32'hF5E5F6C0 , 32'hE74C0340 , 32'hF2F3BA20 , 32'hF73AED50 , 32'hF503A0F0 , 32'h05248D80 , 32'hFA065470 , 32'hFFA1B4CD , 32'hFFAF49D3 , 32'hEE939120 , 32'hFFB3DF10 , 32'h034BA19C , 32'h02BE4060 , 32'hFE739A30 , 32'hF1E37310 , 32'hFC523F60 , 32'hFFF3EBF1 , 32'hFA470E70 , 32'hFC3868C8 , 32'h017B58EC , 32'h15742C80 , 32'hF0C7A220 , 32'hF62E6850 , 32'hFE77D4A0 , 32'hFB9C1250 , 32'h03A79F48 , 32'h06B50DE8 , 32'hFFFA362F , 32'h028B5294 , 32'hFF1CBA36 , 32'h015CB9D8 , 32'hF8543F78 , 32'h0235D3F4 , 32'hFA222BB8 , 32'h04725E48 , 32'h077A4F68 , 32'h0A189D30 , 32'hFEFA6464 , 32'h033A16B0 , 32'h02E43754 , 32'h02ECB610 , 32'h02763F88 , 32'hFFFAE524 , 32'hFCBF77C8 , 32'hFADB1740 , 32'h03AF1548 , 32'h004B7711 , 32'h03EBC950 , 32'h0183AA08 , 32'h004BCD97 , 32'h07F928C8 , 32'hFDCFDEDC , 32'h029911EC , 32'hFB65D230 , 32'h015CD588 , 32'h06539848 , 32'hFD0DFA70 , 32'h031A516C , 32'h01460270 , 32'hFD966AF4 , 32'hFB26E0C8 , 32'hFACE8EF0 , 32'hFEED91DC , 32'h02732150 , 32'hFE8C8C24 , 32'hFD2212E8 , 32'h0033952D , 32'h0000BDBD , 32'h0000E9D2 , 32'hFFFFB3F5 , 32'hFFFE2D27 , 32'h0001E0EB , 32'h000019BB , 32'hFFFFB21A , 32'hFFFF0744 , 32'h000005A2 , 32'hFFFF0353} , 
{32'h22A88DC0 , 32'hB68CCC00 , 32'h1EE64C20 , 32'h3EA41180 , 32'hFFE817E8 , 32'hCD93AF00 , 32'hF51487E0 , 32'h36C9F600 , 32'h194C7060 , 32'h2F4B3BC0 , 32'h047757D8 , 32'h04F386A0 , 32'h0D9B47B0 , 32'hF18E1350 , 32'hEFA48C60 , 32'hF1A6C290 , 32'h04F2DFE0 , 32'h1BB83700 , 32'h2DCB5A00 , 32'h08052EB0 , 32'hF7BB9970 , 32'hEF12FFC0 , 32'hDCAC4740 , 32'hF610DF60 , 32'h03CFC348 , 32'h0264C31C , 32'hE7A085A0 , 32'h0189711C , 32'h0085D048 , 32'h125E84E0 , 32'h1138A5C0 , 32'h0232CEAC , 32'h01F531C0 , 32'h087452B0 , 32'h0462F960 , 32'h08162500 , 32'hFDF72DB8 , 32'hF4B45A90 , 32'h1145E0E0 , 32'hF2595EB0 , 32'h06817F88 , 32'hF9D82EE0 , 32'h12224300 , 32'hFB73CB58 , 32'hFFBC959C , 32'h04E0DC88 , 32'h0AFE23C0 , 32'h01C0CA08 , 32'hFA56A308 , 32'hFE5FDA00 , 32'h025E05F0 , 32'h0AB11180 , 32'hF64B15E0 , 32'hF9B0B4E8 , 32'hFBBFF7C0 , 32'h011233AC , 32'hF9CA7BA0 , 32'hFFFFC687 , 32'h03E8710C , 32'h069DA168 , 32'h010116E0 , 32'hFCB350CC , 32'h0B1A7730 , 32'hFE520A50 , 32'h026E9A54 , 32'h01FE7694 , 32'h01D59030 , 32'hFCD6A5A8 , 32'hFD347EA8 , 32'hFB0E3068 , 32'hF9442B38 , 32'hFE5C89A8 , 32'h046A5850 , 32'h007AAFEB , 32'hFF20C3A4 , 32'hFA5C0D70 , 32'h029CCB70 , 32'hFDD2DC8C , 32'h02C20CE0 , 32'h023FABC4 , 32'h04991528 , 32'h025676EC , 32'h01BE5808 , 32'h016246F8 , 32'h0069C01E , 32'h03482894 , 32'h00F8F99A , 32'hFF80C4A6 , 32'hFDDEEB38 , 32'h00734180 , 32'hFFFFD533 , 32'h00001CFE , 32'hFFFF25DA , 32'hFFFDB92C , 32'hFFFEEEFC , 32'h0000D06A , 32'hFFFFC59A , 32'h000200FD , 32'hFFFFB727 , 32'hFFFF616A} , 
{32'h00035320 , 32'hFFFA742D , 32'h00014447 , 32'hFFFDB5D6 , 32'h00004DF1 , 32'hFFFEBDC1 , 32'h0000E063 , 32'h00032CAC , 32'h0003FD2F , 32'hFFFD6AC4 , 32'hFFFAA477 , 32'h0000A2D7 , 32'h00014EED , 32'hFFFC4857 , 32'h0003D142 , 32'hFFFDDE1B , 32'hFFF9D753 , 32'h0001418E , 32'hFFFF3789 , 32'hFFFD1E69 , 32'hFFFD93A7 , 32'h000130F7 , 32'hFFFD08DE , 32'h000584FA , 32'h00026BB0 , 32'hFFFEFA93 , 32'h00038F48 , 32'hFFFFDA2E , 32'hFFFF1191 , 32'h0001BC2A , 32'h000046EE , 32'h0000F3D6 , 32'h00009FBA , 32'h00009AC2 , 32'h000246B4 , 32'h000270DB , 32'hFFFD3D8B , 32'h000412ED , 32'hFFFE4A8D , 32'h0003F857 , 32'hFFFAF0AC , 32'hFFFBE76D , 32'hFFFF152B , 32'h0001C36D , 32'h00023C78 , 32'h00034411 , 32'hFFFFEBCF , 32'hFFFCF663 , 32'hFFFCC06B , 32'h0001C34B , 32'h0001F9FC , 32'h00031DFA , 32'h00023B83 , 32'h000349B4 , 32'hFFFDC8DC , 32'hFFFF9F35 , 32'h0003E9B2 , 32'h000416D2 , 32'hFFFF7411 , 32'hFFFC0BB0 , 32'hFFFC26CC , 32'hFFFF7F60 , 32'hFFFEABB2 , 32'h0003493E , 32'h00019F96 , 32'hFFFFE944 , 32'h000234AE , 32'h00022AC2 , 32'hFFFE4257 , 32'hFFFC9FA5 , 32'hFFFE1A4C , 32'hFFFFD7C9 , 32'hFFFDBFD4 , 32'h0004A073 , 32'hFFFC7CE5 , 32'hFFFC777C , 32'h0000F77F , 32'h0000291F , 32'h000067CB , 32'hFFFE7162 , 32'hFFFDF454 , 32'hFFF833C1 , 32'h0000BDC3 , 32'hFFFD4449 , 32'h0000BB1E , 32'hFFFEF936 , 32'h000464FB , 32'h00009A65 , 32'h0004633C , 32'hFFFFB3BB , 32'h0000714A , 32'hFFFAF120 , 32'hFFFCB607 , 32'h00017FE6 , 32'hFFFF43EF , 32'hFFFD1412 , 32'h00014ECD , 32'hFFFF6274 , 32'hFFFC72DD , 32'hFFFDDF66} , 
{32'hE5345920 , 32'h0A138C60 , 32'hFD2968DC , 32'h28CF9780 , 32'h034BE738 , 32'h01377C90 , 32'hEBB0F620 , 32'hE9B90460 , 32'hEE3E8840 , 32'h1917CE60 , 32'hFAE28650 , 32'hF4D36CE0 , 32'hDE7B0640 , 32'h12AE13C0 , 32'h005343B2 , 32'h0472DDF8 , 32'h05CEFD10 , 32'h1D691300 , 32'hFC4FF65C , 32'hF09274B0 , 32'hF5EA7890 , 32'h18870E40 , 32'hE24E9820 , 32'hFE075FF8 , 32'hFA7B3BE0 , 32'h0CCD2B90 , 32'h06ADD000 , 32'hF757C0E0 , 32'hEF8B7760 , 32'hEC65B140 , 32'hFF1B4BFD , 32'hF6A88630 , 32'h19811180 , 32'h0A315BC0 , 32'hF92E77C8 , 32'h09BFE980 , 32'h03D0F40C , 32'hF9170218 , 32'h10B46820 , 32'hFD7E8548 , 32'hF5E2E3B0 , 32'hF55E0550 , 32'hEC8D73C0 , 32'hFF881B17 , 32'hFD37E04C , 32'h0E1C1BC0 , 32'hFB18FB70 , 32'hF603D6C0 , 32'hFEAB524C , 32'hFF3EB3A8 , 32'hFB69D510 , 32'hFCD169F4 , 32'h0806AD80 , 32'hFA3A3BA0 , 32'h0669F130 , 32'h0031D324 , 32'hFDAAEBA0 , 32'hFD8B82BC , 32'h0353AB00 , 32'h01168BD8 , 32'hFD801E58 , 32'h01437BB4 , 32'h00A4B678 , 32'h00C3AFC3 , 32'h03F36BC8 , 32'hF574EC50 , 32'hF9DFE670 , 32'hFEBA3054 , 32'hFCF5CD08 , 32'hFF6FE76E , 32'h00266777 , 32'h0860C5E0 , 32'h00004FB9 , 32'h010A8E78 , 32'h08A25FD0 , 32'hFFE6C608 , 32'hFA9EA600 , 32'h00E71A60 , 32'h061D0B20 , 32'h028435C8 , 32'hFF91F675 , 32'hFF68F0E8 , 32'hFF961AE9 , 32'hFE4896A4 , 32'h02BC92BC , 32'hFB8D6CF0 , 32'h0149AFD4 , 32'h0100EA1C , 32'hFEBA8970 , 32'hFF996877 , 32'h0000994F , 32'hFFFF6F5C , 32'h0000B091 , 32'hFFFE2D44 , 32'h0001D170 , 32'h000151B8 , 32'h0000E704 , 32'h0000E225 , 32'hFFFDA883 , 32'hFFFF679B} , 
{32'h0002C7F0 , 32'hFFFD64FF , 32'hFFFEE15A , 32'hFFFFE1E7 , 32'hFFFEA28E , 32'hFFFE51AC , 32'h0001694B , 32'hFFFF3619 , 32'h00016D44 , 32'h00011468 , 32'h00015552 , 32'hFFFEEFB8 , 32'hFFFF4291 , 32'h0002F854 , 32'h0000A85A , 32'h0002631F , 32'hFFFBD5C6 , 32'h000429E3 , 32'hFFFD116A , 32'h0002D35A , 32'h00005F87 , 32'h0001D8B1 , 32'hFFFF5B65 , 32'h0001209F , 32'h00001AA7 , 32'h00031BA2 , 32'hFFFF37B6 , 32'h000117D8 , 32'hFFFA9B8F , 32'h0001D89A , 32'hFFFB294F , 32'hFFFE9FBE , 32'h00058806 , 32'h000315D9 , 32'hFFFDF02F , 32'hFFFFB665 , 32'h00016396 , 32'h000160D8 , 32'hFFFF6EC7 , 32'h0002848A , 32'hFFFE3F01 , 32'h0002A3DD , 32'hFFFD2CE7 , 32'h00013E3D , 32'h0003E1DB , 32'h00033DB3 , 32'hFFF9CA6D , 32'h0004B9D8 , 32'hFFFDEB21 , 32'hFFFAD79B , 32'h00023AE9 , 32'hFFFE84E2 , 32'hFFFEDD14 , 32'hFFFF2D23 , 32'hFFFD4CD2 , 32'h000155A8 , 32'h0004EFA6 , 32'hFFFD404C , 32'h000222A8 , 32'hFFFC7431 , 32'h0002184B , 32'h00005AD9 , 32'hFFFBFBBE , 32'hFFFC60E8 , 32'hFFFCF84F , 32'hFFF9A5CA , 32'h000091F0 , 32'h00007947 , 32'h000121DD , 32'hFFFF2227 , 32'hFFFD153C , 32'hFFFD37DD , 32'hFFFD12AA , 32'hFFFBA429 , 32'hFFFF76C4 , 32'hFFFC4EFD , 32'hFFFF6DC6 , 32'hFFFCC84C , 32'h000055EB , 32'hFFFD1200 , 32'h00009C73 , 32'hFFFB5065 , 32'hFFFD7B32 , 32'hFFFF485C , 32'hFFFD7E8E , 32'hFFFE4249 , 32'hFFFE8DFA , 32'hFFFE2FD3 , 32'h00015F63 , 32'hFFFB35EE , 32'hFFFB5921 , 32'h000026ED , 32'h00015B0F , 32'h000063F6 , 32'hFFFE8C4F , 32'hFFFB0D54 , 32'hFFFFD42F , 32'hFFFD345B , 32'hFFFE66ED , 32'hFFFECF23} , 
{32'hFBF3E878 , 32'hF52599C0 , 32'h04CEDF90 , 32'hF73423F0 , 32'hF03050C0 , 32'h002B58C6 , 32'h090B6480 , 32'hEA941500 , 32'hFC174D4C , 32'hF9820128 , 32'h072E4268 , 32'hFF6E28D6 , 32'hFD4DC05C , 32'h0011A610 , 32'hFC7F05B4 , 32'hFB7E1CF0 , 32'hFFDDF82F , 32'h02E1A194 , 32'hFC0E4DE4 , 32'h12ACFDE0 , 32'h127985A0 , 32'h04FA77A8 , 32'hFD96431C , 32'hE8F4A940 , 32'hFE4F4000 , 32'h0A6BB3C0 , 32'h0ABDB0E0 , 32'h05F48D30 , 32'hFF2C8E74 , 32'hF45862C0 , 32'hFF2DA647 , 32'h075D51A0 , 32'h02EE2BDC , 32'hFB1B76F0 , 32'h116E9120 , 32'h07A6FEB8 , 32'h00440C32 , 32'hFBC67810 , 32'hFD427F60 , 32'hF3FD7D90 , 32'h033D0CF4 , 32'hFD28B31C , 32'hFAE0B800 , 32'hFAC849B0 , 32'h02E55BF4 , 32'h0E5025A0 , 32'h0BD81C50 , 32'hF709DFB0 , 32'h046518D0 , 32'hFF5E20D6 , 32'hF9BD5368 , 32'hFC274E00 , 32'h0988E3A0 , 32'hFCCA9FD4 , 32'hFDDDBFC0 , 32'h01ED7464 , 32'hF8DBD7C8 , 32'h0249454C , 32'h013379A8 , 32'hFE6FDAA0 , 32'h070ACC60 , 32'hFE28E4B8 , 32'h053C4390 , 32'h0364A838 , 32'hFC41F584 , 32'hFB1C2798 , 32'hFFB8155D , 32'hFEFD89B8 , 32'hFD15F1F4 , 32'hF93D9E40 , 32'h0080B4A9 , 32'hF9950388 , 32'hFE7CA968 , 32'h0382B198 , 32'hFE7CB244 , 32'h024958F0 , 32'h01C4D510 , 32'h02EB6B20 , 32'hFF91211F , 32'hFD8DDF48 , 32'h00923238 , 32'hFC993240 , 32'hFB7F0410 , 32'h00895AE6 , 32'hFFBD8697 , 32'hFE22D800 , 32'hFF300B20 , 32'hFCC0CEC0 , 32'h032AACC0 , 32'h00D88E13 , 32'h0001A81D , 32'h000166D3 , 32'hFFFFB94B , 32'h000096AB , 32'hFFFFB08A , 32'h00008E6E , 32'h00017E60 , 32'hFFFE053D , 32'hFFFE7065 , 32'hFFFE45D7} , 
{32'h00051947 , 32'h00009114 , 32'hFFFFDF0B , 32'h0002DCF6 , 32'h00011693 , 32'hFFFE3922 , 32'h00008067 , 32'h0000846B , 32'h00067A05 , 32'h00008CED , 32'hFFFF79FF , 32'hFFFC85E0 , 32'h0003475D , 32'h000260CB , 32'hFFFB8CC1 , 32'h0000A6B1 , 32'hFFFA7BAD , 32'h00018939 , 32'hFFFEF190 , 32'hFFFAC9C4 , 32'h00009888 , 32'h00005DE7 , 32'hFFFFF705 , 32'h000147FB , 32'h000034EF , 32'h00000046 , 32'hFFFFAF49 , 32'hFFFD623D , 32'hFFF83013 , 32'h0007B301 , 32'hFFFD0B62 , 32'h0000C69D , 32'hFFFE9392 , 32'hFFFDE8AB , 32'hFFFBE9FF , 32'hFFFE8FD9 , 32'h000251BB , 32'h0003ECCE , 32'hFFFB821B , 32'h000082F6 , 32'hFFFB4D65 , 32'hFFFF1027 , 32'hFFFC1F03 , 32'h00016099 , 32'hFFFFFABF , 32'hFFFE1A50 , 32'hFFFF6449 , 32'h0001AACE , 32'h00007939 , 32'h0000EB41 , 32'hFFFE74F2 , 32'hFFFFB513 , 32'h00064743 , 32'hFFF9B3DC , 32'h00008594 , 32'hFFFB575F , 32'h0001CBC1 , 32'h00010F81 , 32'h0000FEC8 , 32'hFFFF5CD1 , 32'hFFFF5438 , 32'hFFFD8AD5 , 32'hFFFEE9C5 , 32'hFFFCCCEA , 32'hFFFF7DB2 , 32'h0006A841 , 32'hFFFFF63C , 32'h0002AF05 , 32'h00018F3B , 32'hFFFF14FA , 32'h0000A445 , 32'hFFFD4983 , 32'hFFFFAB1A , 32'hFFFF830A , 32'hFFFEA180 , 32'hFFFFC3C1 , 32'h00024A4C , 32'h00049F7B , 32'h0002B5C3 , 32'hFFFEB6AE , 32'hFFFC7CC1 , 32'h00000CE8 , 32'h0000D74D , 32'hFFFEF994 , 32'h00023A97 , 32'h000277A6 , 32'h0001680D , 32'h00010777 , 32'hFFFF7DC7 , 32'h0000D1F5 , 32'hFFFFDA8F , 32'hFFF9B7A2 , 32'hFFFEBD26 , 32'hFFF853EA , 32'hFFFC41AA , 32'h0001D2FD , 32'h00005B56 , 32'hFFFB2B8A , 32'h00075680 , 32'hFFFD22EE} , 
{32'hFFFFE56F , 32'hFFFDFC28 , 32'h0003233E , 32'h000491D1 , 32'hFFFF4558 , 32'hFFFD71A2 , 32'h0002E302 , 32'h00017202 , 32'hFFFFF373 , 32'h0002C856 , 32'h0003637D , 32'h0002EBB4 , 32'h00027AAD , 32'hFFFE225B , 32'hFFFFEF63 , 32'hFFFF5033 , 32'h0001286A , 32'h0002F0B7 , 32'hFFFDAD90 , 32'hFFFE1D4A , 32'h0000CEB1 , 32'hFFFF5A3F , 32'h00038AE0 , 32'hFFFD4B3B , 32'hFFFFE758 , 32'h0002A51A , 32'h0003928E , 32'hFFFFD619 , 32'hFFFC3CE6 , 32'h00020771 , 32'h00027126 , 32'hFFFDB6DC , 32'h000029C0 , 32'hFFFEE7AD , 32'h00003F7B , 32'h00023B79 , 32'h0001DE4C , 32'h00028472 , 32'h0000DC20 , 32'h0002A5B2 , 32'h000367F7 , 32'h00023C7C , 32'h00018A1A , 32'h00019FD3 , 32'h0000C41F , 32'hFFFB9B25 , 32'hFFFFEF36 , 32'h00010DE5 , 32'hFFFDE438 , 32'hFFFF1986 , 32'h00047647 , 32'hFFFFF43E , 32'hFFFD1C7F , 32'hFFFCB1FF , 32'h00015D20 , 32'hFFFB62F5 , 32'hFFFF6603 , 32'h00006124 , 32'hFFFB9380 , 32'hFFFF799F , 32'h0001DB95 , 32'hFFFFC6A3 , 32'hFFFE3199 , 32'h0003B1EA , 32'hFFFE2FCE , 32'hFFFF990B , 32'hFFFFAC8C , 32'h00009B8B , 32'hFFFED8C3 , 32'hFFFE8C41 , 32'hFFFF81D8 , 32'hFFFF6FFA , 32'h0003707B , 32'h000217A9 , 32'h0001701D , 32'hFFFE307B , 32'h00014517 , 32'hFFFDF089 , 32'hFFFD7CF8 , 32'hFFFF8921 , 32'h000259B2 , 32'h00015447 , 32'hFFFCD407 , 32'hFFFF3334 , 32'hFFFEFE86 , 32'hFFFA6D28 , 32'h0002D809 , 32'h00025F7F , 32'h00009F22 , 32'hFFFECFAB , 32'h0000F911 , 32'hFFFC89B9 , 32'hFFFD6D0A , 32'hFFFFAD1A , 32'h00036321 , 32'hFFFEC504 , 32'hFFFAFA2E , 32'hFFFE59B5 , 32'h0002F50E , 32'hFFFEE586} , 
{32'h000284DC , 32'hFFFC9FC6 , 32'h00016EBA , 32'h00016A24 , 32'hFFFEDDA4 , 32'h00036ABD , 32'h00033288 , 32'h00014B52 , 32'hFFFBB953 , 32'h0002E057 , 32'h00041210 , 32'h000417E8 , 32'h00059651 , 32'h00007011 , 32'h00040B00 , 32'hFFFDFAC0 , 32'h00000204 , 32'hFFFC3B30 , 32'h00011E85 , 32'hFFFAA499 , 32'hFFFE67CC , 32'h000535B3 , 32'hFFFFD549 , 32'hFFFDCDC6 , 32'h00014EFD , 32'hFFFEA3A4 , 32'hFFFF3A0C , 32'hFFFEA327 , 32'hFFFAD5CB , 32'hFFFE4565 , 32'hFFFC1920 , 32'hFFFF79CE , 32'h0000110E , 32'hFFFCB0A3 , 32'h00035F87 , 32'h00009828 , 32'h0000F4A7 , 32'hFFFAED1E , 32'h000190E9 , 32'hFFFE5016 , 32'hFFFF5193 , 32'h0000906B , 32'hFFFCAC06 , 32'h00053BE0 , 32'hFFFE0803 , 32'hFFFF8EA6 , 32'h000242F3 , 32'h000433B2 , 32'hFFFF9C1C , 32'hFFFA59C0 , 32'h0005288A , 32'hFFFFC974 , 32'hFFFF81B2 , 32'hFFFBBE6E , 32'hFFFDED2F , 32'h0002464A , 32'h00022815 , 32'h00004C8D , 32'hFFFE32E6 , 32'h00016410 , 32'h000296FF , 32'h000556A2 , 32'h00015227 , 32'hFFFD86F5 , 32'hFFFF1F0D , 32'hFFFBB234 , 32'h0003DFC5 , 32'h00002375 , 32'hFFFA819C , 32'h0002B2D5 , 32'hFFFFBC80 , 32'hFFFDB172 , 32'h00029917 , 32'h0002ED35 , 32'h0004BAB5 , 32'h00018C55 , 32'hFFFC07CB , 32'hFFFEFAD1 , 32'h00033B38 , 32'hFFFF558C , 32'h00068D2B , 32'h00010F66 , 32'h00027CBE , 32'hFFFD1C6F , 32'hFFFE16B6 , 32'hFFFD8598 , 32'h00031171 , 32'h0004A06D , 32'hFFFFBB4D , 32'h000119FB , 32'hFFFD9889 , 32'h0000869E , 32'h0000FB09 , 32'hFFFCA0AF , 32'h0005CBC6 , 32'hFFFE9402 , 32'hFFFFBA53 , 32'hFFFCDC23 , 32'h00013B01 , 32'h0000BC8C} , 
{32'h00031CA0 , 32'hFFFD3622 , 32'h00033F89 , 32'h000443E9 , 32'hFFFD7627 , 32'hFFFEA864 , 32'hFFFB2433 , 32'hFFFEF1F7 , 32'h00005BBB , 32'hFFFDC19B , 32'hFFFD53BC , 32'h0001C7AF , 32'hFFFF40BE , 32'hFFFE66C4 , 32'hFFFD68BC , 32'h00080C50 , 32'hFFFDB8EE , 32'hFFFEA856 , 32'h0002A783 , 32'hFFFD93F1 , 32'h00035A92 , 32'hFFFDD32F , 32'h00020F0F , 32'h000050AB , 32'hFFFE0314 , 32'hFFFFA9FE , 32'h0002D7E4 , 32'h00031355 , 32'h0001FCB6 , 32'hFFFB786D , 32'hFFFFD402 , 32'hFFFE6062 , 32'h0003B593 , 32'h00042089 , 32'h00015C25 , 32'h0000CCC2 , 32'h00059AD1 , 32'h00000CF1 , 32'h000250E2 , 32'h00046BC2 , 32'h0002683E , 32'hFFFD2FE0 , 32'hFFFECBE2 , 32'h0004CE63 , 32'hFFFFAA6F , 32'hFFF9743B , 32'hFFFC021F , 32'hFFFD43B9 , 32'h00005358 , 32'hFFFE3911 , 32'h0000C85E , 32'h00049FBB , 32'hFFFD3BC3 , 32'hFFFFE6E9 , 32'hFFFD8B22 , 32'h00036771 , 32'hFFFA8524 , 32'h00021EBE , 32'h00041EE3 , 32'hFFFDD89F , 32'hFFFB68D1 , 32'h00027F77 , 32'hFFFE44D3 , 32'h00032C35 , 32'hFFFA5935 , 32'h000206D1 , 32'hFFFF0959 , 32'h00022B65 , 32'h000175CA , 32'hFFFB076F , 32'h0001BCFC , 32'hFFFDFD03 , 32'h00034E83 , 32'hFFFE574B , 32'h0004A03E , 32'h0004021B , 32'hFFFC23E4 , 32'h00060518 , 32'h00009083 , 32'hFFFB4A3C , 32'h000468F0 , 32'h00038465 , 32'h00033EE4 , 32'hFFFD9C77 , 32'hFFF9B2CC , 32'hFFFCEFC2 , 32'h0002E3B8 , 32'h0002C88B , 32'h00046BFD , 32'h000448C2 , 32'h000416CA , 32'hFFFFE2E6 , 32'h0002F372 , 32'hFFFCAEA4 , 32'hFFFBC2E5 , 32'h00018F84 , 32'h0002C95C , 32'hFFFE46ED , 32'h00014212 , 32'h00008EA8} , 
{32'h22A86500 , 32'hEDA07A00 , 32'h08B7DA20 , 32'hFA786AF8 , 32'hF4F20FA0 , 32'h105C0E20 , 32'h23E57340 , 32'h09535300 , 32'hE75F4480 , 32'h0F944290 , 32'h0AF04FB0 , 32'hF64BD000 , 32'hFCD6C720 , 32'hFC2EAF04 , 32'hFD63DB58 , 32'h18B3BB80 , 32'hF6DA9920 , 32'h11A00C00 , 32'hF4DF5770 , 32'h08EF8D80 , 32'hF037AB70 , 32'hFA7C6B30 , 32'h09897170 , 32'h0CD33D30 , 32'hF9A4C838 , 32'h09F9F880 , 32'h06E0FF88 , 32'h0319BE8C , 32'h08AB6220 , 32'hFD672B80 , 32'h0B61F040 , 32'h06814358 , 32'hEF3AD640 , 32'hE84A68A0 , 32'h0539F918 , 32'h06255378 , 32'hF59C2430 , 32'h0A5064F0 , 32'h0708B0C0 , 32'hF99851A0 , 32'hF8F1DE08 , 32'h01B5291C , 32'hE9FB3EC0 , 32'h0A5C0490 , 32'h01A4BE68 , 32'h0A241B50 , 32'hFE7539F8 , 32'hFD62A228 , 32'hFD488B8C , 32'hFFAF1CD3 , 32'hF9530180 , 32'h065A4510 , 32'hF141E360 , 32'h0B96F810 , 32'h0620D6E0 , 32'h051341C8 , 32'h04D2D2C8 , 32'hFF866E37 , 32'hF6762330 , 32'h00316B9B , 32'hFEF4322C , 32'hFF16C3B4 , 32'hFDF4E424 , 32'h01562754 , 32'h03F1C04C , 32'hFF280548 , 32'h0486D520 , 32'hFB5BD680 , 32'hFAAEE1E8 , 32'h017B41D4 , 32'hFD4D6CD0 , 32'hFEBACD70 , 32'h08DF6940 , 32'h00D61A69 , 32'h0383D368 , 32'h01663CE0 , 32'hFE145780 , 32'h094E22D0 , 32'h00EEE17E , 32'h027000F4 , 32'h00C7E1C1 , 32'h00EDFC0E , 32'hFB05F608 , 32'hFCED207C , 32'h01EBE0A4 , 32'hFEAE9CF0 , 32'hFE48ECCC , 32'hFF12006A , 32'h015C0360 , 32'h00842198 , 32'h00006B44 , 32'h000162E2 , 32'h00005B8B , 32'hFFFD2DD4 , 32'hFFFEEC95 , 32'hFFFF1026 , 32'hFFFB0D22 , 32'hFFFF9BAD , 32'hFFFE56C5 , 32'hFFFED423} , 
{32'h2805D3C0 , 32'hF4553090 , 32'hC4565BC0 , 32'hE934BC20 , 32'h2789E800 , 32'hFA878FC8 , 32'hE132CFE0 , 32'h06B779F8 , 32'hF6382970 , 32'hFD5CC610 , 32'hBC334180 , 32'h0E491210 , 32'hF5EBA6E0 , 32'h07B47B80 , 32'h12A91D00 , 32'hF4003040 , 32'h0391DCE8 , 32'h055DD5D8 , 32'h0BC01670 , 32'h05D98350 , 32'h040C9FC8 , 32'h1DFF2920 , 32'h15BF8AE0 , 32'h14412320 , 32'hF1A63970 , 32'hF6814400 , 32'hF7FFE7B0 , 32'hEEEE67A0 , 32'h080882F0 , 32'hFF343200 , 32'h00DF389A , 32'h0A8EC1F0 , 32'h05744100 , 32'hF923D5C8 , 32'h02B5440C , 32'h0A1D3C30 , 32'hF362D450 , 32'hF4DF5060 , 32'h034E6E3C , 32'hEDE42900 , 32'hFE400564 , 32'h07CF2760 , 32'hEFF0EBA0 , 32'hFA6987B8 , 32'hFF10ECAB , 32'hF5866C50 , 32'h0CB09EA0 , 32'h0058AD73 , 32'h02457EC8 , 32'hFE387AD4 , 32'h092C0A20 , 32'h00E51114 , 32'hFC897CDC , 32'hFEF8C888 , 32'hFCEFEEF0 , 32'hFD2745AC , 32'h0320B1E8 , 32'h02623BF8 , 32'hFF67115F , 32'hF8D2FA10 , 32'hF837A768 , 32'h028C9E48 , 32'hFCFBCE74 , 32'hFBF4C408 , 32'hFE39D244 , 32'h0423B220 , 32'h031FC4A4 , 32'h01D56D68 , 32'h045B40A8 , 32'hFF12CA3F , 32'hFEC3D994 , 32'h01EAB9D0 , 32'hFFE0F93A , 32'h018B4868 , 32'h01CE0C40 , 32'hFF18B7ED , 32'h03541CF8 , 32'hF8FBAFB8 , 32'hFF059DAD , 32'h0358C65C , 32'h05683BC0 , 32'h05A394D8 , 32'h02B2286C , 32'hFD5C60C4 , 32'h00EB4128 , 32'hFFC8E0F5 , 32'hFE987B34 , 32'hFFFE5EB3 , 32'h02099338 , 32'hFEE197B4 , 32'hFFFEBA4D , 32'h00018A65 , 32'hFFFCC062 , 32'h000060A5 , 32'hFFFDE8AF , 32'hFFFEF610 , 32'hFFFFEEAA , 32'hFFFF531B , 32'h00005FFE , 32'hFFFE0A4D} , 
{32'h0BA0E730 , 32'h25CF1100 , 32'hF5D409D0 , 32'h05DCE0F0 , 32'hF5813290 , 32'h07FB1AC0 , 32'hE2E57340 , 32'h07E6E7C0 , 32'hF46A5150 , 32'h0E363B00 , 32'h01DDFA64 , 32'h02212434 , 32'hF74DCCC0 , 32'hEE8EF780 , 32'hEE70DBA0 , 32'h0128DD08 , 32'h05B57E18 , 32'hFFD510C3 , 32'h10DD3E20 , 32'hFF860264 , 32'hFEEBA818 , 32'hF20AA170 , 32'hFAB6D128 , 32'hFAD5CC20 , 32'h017A3014 , 32'h0573CD90 , 32'h03EDD8A0 , 32'hFD8E05D0 , 32'h0ABC0950 , 32'h083D9750 , 32'hFD7F9F10 , 32'hF8010170 , 32'h0D506520 , 32'hFA41F768 , 32'h0EE4A080 , 32'h079579D0 , 32'h015D1B1C , 32'h06978A98 , 32'hFED55F8C , 32'hF2AC40F0 , 32'hFF15CDD2 , 32'h0BA40540 , 32'h11AAF220 , 32'h0308ABD0 , 32'hFAB48330 , 32'hEA0E7280 , 32'hF5B2C930 , 32'hF51AB0B0 , 32'h03D1BA78 , 32'h0874B310 , 32'hF600CDF0 , 32'h00DA8DDA , 32'hFD21B70C , 32'h11BFD5E0 , 32'hF5DBA520 , 32'h05B3A258 , 32'hFF8AE18D , 32'hFD0EE58C , 32'h04B89D18 , 32'hFDB960E4 , 32'hFAB45388 , 32'h01F61C7C , 32'hF56DDA40 , 32'hF6FA7570 , 32'h08B698D0 , 32'hFF406ABC , 32'hFA69CE90 , 32'h00EC01B5 , 32'hFD7C40F0 , 32'h036F3628 , 32'h027529AC , 32'hFD56DB7C , 32'hFA0B4780 , 32'h06943880 , 32'h02E64970 , 32'h02EE4578 , 32'hF818E308 , 32'hFCF790E0 , 32'hFF030E3B , 32'hFDB0FF18 , 32'hFE61792C , 32'hFE7D8A1C , 32'hFE8A213C , 32'hFF581D4F , 32'h037E8130 , 32'h00E2FBA0 , 32'h01D764E0 , 32'h0178CD28 , 32'h01657C64 , 32'hFFEA1522 , 32'hFFFC5E61 , 32'h00004A37 , 32'h0001576F , 32'hFFFD9602 , 32'hFFFD81DE , 32'h000101B2 , 32'h000124F3 , 32'hFFFF4BB4 , 32'h00006511 , 32'h00000C95} , 
{32'h0000B1B1 , 32'h0000091A , 32'h0001C092 , 32'hFFFC892E , 32'hFFFCB0E1 , 32'hFFFF93D9 , 32'h0003033F , 32'hFFFC0489 , 32'hFFFF4793 , 32'hFFFC3BFA , 32'h000453FB , 32'h000068FB , 32'h00005FA6 , 32'h00023BA1 , 32'h000446F7 , 32'h00027635 , 32'h0001A53D , 32'h00007E41 , 32'h0003F1D6 , 32'h00013A05 , 32'h0000C026 , 32'hFFFEF8BC , 32'hFFFD3CC4 , 32'h00024ABB , 32'hFFFD4229 , 32'hFFFBE5D4 , 32'hFFFF796A , 32'h000030E9 , 32'h000271C6 , 32'hFFFF640F , 32'h0000DF1F , 32'h0002BFB8 , 32'hFFFC6A9A , 32'h0000DEDB , 32'hFFFE5D67 , 32'hFFFE77E6 , 32'h000022F6 , 32'h00032B80 , 32'hFFFC8605 , 32'h0001DA54 , 32'hFFFCE198 , 32'hFFFBA09D , 32'hFFFF98CC , 32'h00004677 , 32'hFFFEE7F0 , 32'hFFFB3043 , 32'hFFFBE632 , 32'h00008297 , 32'h0002E312 , 32'hFFFDE5A4 , 32'hFFFD4439 , 32'hFFFE9EAE , 32'h00058B33 , 32'hFFFDD9B2 , 32'h00006A0E , 32'h00008797 , 32'hFFFE3947 , 32'h0000BECE , 32'hFFFEB19C , 32'h0000B7BB , 32'h0001B99D , 32'hFFFC70D2 , 32'h00002130 , 32'h0000E02B , 32'hFFFE3F32 , 32'h0001AB27 , 32'h0001C236 , 32'hFFFE0CFD , 32'hFFFEFF69 , 32'h0003F47F , 32'h0002E6E4 , 32'hFFFE919F , 32'hFFFD0D8F , 32'hFFFFA418 , 32'h0002766A , 32'h000048DF , 32'h00008737 , 32'hFFFD7DDA , 32'h00004832 , 32'h000161F6 , 32'h0001676E , 32'hFFFFA4CC , 32'h000106F1 , 32'hFFFF607D , 32'h00033264 , 32'hFFFF045E , 32'hFFFEE036 , 32'hFFFE063F , 32'hFFFFDBE7 , 32'h00017EA6 , 32'h0001FB71 , 32'hFFFD788B , 32'hFFFF129A , 32'h0004BFA2 , 32'h00022D93 , 32'h000269F9 , 32'h0001DE4C , 32'hFFFD96AE , 32'h00004525 , 32'hFFFD9730} , 
{32'h000403D2 , 32'hFFFE9ED7 , 32'h0004D2E2 , 32'hFFFFF8C2 , 32'h00014505 , 32'hFFFE1DA6 , 32'h0000BAD8 , 32'h00002DFE , 32'hFFFF5D45 , 32'hFFFF04A0 , 32'hFFFC09C6 , 32'hFFFDA6C8 , 32'hFFFF37B5 , 32'hFFFE375D , 32'h00007CC9 , 32'hFFFCEE15 , 32'h0001A51E , 32'hFFFFC6CA , 32'hFFFC753B , 32'h0001F55D , 32'hFFFE2EED , 32'h00009E8B , 32'h000173C5 , 32'hFFFE21D2 , 32'h000072EF , 32'h0002CD5D , 32'hFFFCBEF2 , 32'hFFFA7A16 , 32'h0000B37B , 32'h00004C44 , 32'hFFFF5583 , 32'h000159F9 , 32'hFFFD7D2E , 32'hFFFEC427 , 32'hFFFD58EE , 32'h000035AF , 32'h0000B784 , 32'h00072712 , 32'hFFFEE8F7 , 32'hFFFEDD7B , 32'h00009F4E , 32'h0004C878 , 32'h0000E45C , 32'h00047961 , 32'h00023FAE , 32'h00013035 , 32'hFFFC5EF7 , 32'h00019475 , 32'h0004555D , 32'h0000C37E , 32'hFFFD21CD , 32'h0000631C , 32'h000169A6 , 32'hFFFD012F , 32'hFFFFB6A7 , 32'h00021EF6 , 32'hFFFC2C72 , 32'hFFFB9A13 , 32'h00009FD3 , 32'hFFFFE483 , 32'hFFFE93A9 , 32'hFFFF6EE3 , 32'h00033757 , 32'hFFFEA72C , 32'hFFFE7FDE , 32'hFFFE1901 , 32'h0000C4FF , 32'h000076E5 , 32'h00003E3E , 32'hFFFF5E3A , 32'hFFFE8AE3 , 32'h0004C9F7 , 32'hFFF7E827 , 32'h00041C40 , 32'hFFFFBCF5 , 32'hFFFD9EA9 , 32'h00024734 , 32'hFFFDC46C , 32'h0002B6ED , 32'hFFFD96EB , 32'hFFFF551C , 32'h0006C61B , 32'hFFFBA390 , 32'hFFFD63F1 , 32'h000000A8 , 32'h00016A0F , 32'h00025B43 , 32'hFFFE2D53 , 32'hFFFDF894 , 32'hFFFFA90C , 32'h0002A333 , 32'hFFFFD06E , 32'h00022854 , 32'hFFFD92C9 , 32'hFFFC7CF2 , 32'hFFFFE375 , 32'hFFFE5C4E , 32'h00006064 , 32'h000100B8 , 32'hFFFD1C77} , 
{32'hB3D42880 , 32'h174CCDA0 , 32'h30A34DC0 , 32'hEDE4F340 , 32'hEAB94C60 , 32'h02EAA9BC , 32'h05D83D08 , 32'h03E24680 , 32'hE541F3C0 , 32'hF01F3030 , 32'hD6317BC0 , 32'h101CA060 , 32'h01AE1274 , 32'h026F7E44 , 32'hF4683030 , 32'hF2474B80 , 32'h14EC1D20 , 32'hF57A7EB0 , 32'h130C2B00 , 32'h0FE64180 , 32'hF5AFC2D0 , 32'hF9F3AB20 , 32'hED8FB8E0 , 32'hFC18E3AC , 32'hFEC8220C , 32'h0ABEAFA0 , 32'h007BD2C3 , 32'h06BC3C28 , 32'h12637960 , 32'h09D15E50 , 32'hFBD95280 , 32'h069F70B8 , 32'h03BCD544 , 32'h04382FC8 , 32'h0614A640 , 32'hF132BF10 , 32'h09E33550 , 32'hFF251090 , 32'h043A6840 , 32'hFF22372B , 32'h06C9BD30 , 32'hFD8BC16C , 32'h02FFA448 , 32'hFAA86548 , 32'hF44AD1C0 , 32'hF3C826F0 , 32'hFD86BAB8 , 32'hFF82265B , 32'hFBBDA998 , 32'h0139659C , 32'hF8767DE8 , 32'hFC401338 , 32'h10307B20 , 32'hFF386EFB , 32'h037D6F6C , 32'h058916A0 , 32'hF5493F80 , 32'h05467300 , 32'hFABF4AB8 , 32'h00A84010 , 32'h0592ECD0 , 32'hFC2AD7A4 , 32'hFB270DC0 , 32'h06B01C10 , 32'hFBF9B628 , 32'hFB082BF8 , 32'h01F904CC , 32'h000B344B , 32'h0F22A770 , 32'hFFC0D70B , 32'hFDD55A68 , 32'hFE43314C , 32'hFF64A942 , 32'h070E82A8 , 32'h054BA7A0 , 32'hFEA37D98 , 32'h02249A54 , 32'h0711D018 , 32'h022F5F2C , 32'hFF8474BF , 32'hF5C70AA0 , 32'h00F8E57E , 32'h05BA9540 , 32'hFFFF4E6D , 32'h01DAEFB4 , 32'h02CB4950 , 32'h00C25642 , 32'hFCCD11F0 , 32'h03855BF8 , 32'h00ADC4FB , 32'hFFFEF42A , 32'h00009A9D , 32'hFFFC13A8 , 32'h0001D66C , 32'hFFFFA8DA , 32'hFFFEEBF0 , 32'hFFFE6DFF , 32'h000084A7 , 32'hFFFF7D53 , 32'h0000F38F} , 
{32'h0003479C , 32'hFFFFD4B4 , 32'hFFFA1C40 , 32'h00061993 , 32'hFFFFC8FB , 32'h0000B1B2 , 32'hFFFB156F , 32'h0001042A , 32'hFFFD326A , 32'hFFFEF069 , 32'hFFFB3B4A , 32'h0001FD8C , 32'h0000A6BB , 32'hFFFD5B0C , 32'hFFFD11EE , 32'h00006CF1 , 32'hFFFCA82C , 32'hFFFC7DAF , 32'h00027ABC , 32'h0000F719 , 32'hFFFF7142 , 32'hFFFC75BC , 32'h0001362B , 32'h0001DBAF , 32'h00019797 , 32'hFFFD9658 , 32'hFFFF975B , 32'h0001F24A , 32'hFFFFDE64 , 32'hFFFD5BCB , 32'h0000925E , 32'hFFFF7286 , 32'hFFFFF6B3 , 32'hFFFCC5E4 , 32'hFFFD0806 , 32'h00015498 , 32'h0000DFE5 , 32'hFFFECA84 , 32'h000229A1 , 32'hFFFF9A92 , 32'hFFFEA1BB , 32'h0001800A , 32'h00024F87 , 32'hFFFEA3DF , 32'hFFFDAFF9 , 32'hFFFDF43C , 32'h00025F0F , 32'hFFFBF29D , 32'h0000AD58 , 32'h00013F5A , 32'hFFFF740D , 32'hFFFCCC43 , 32'h00050F1D , 32'hFFFD6D45 , 32'hFFFE7A60 , 32'h00039842 , 32'h00030C05 , 32'h00024E64 , 32'h0001FF06 , 32'h00009208 , 32'h00004D9B , 32'h0001AEB7 , 32'hFFFF84EE , 32'hFFFB7F9B , 32'h0004CD3D , 32'h0000BCAB , 32'hFFFFC837 , 32'hFFFCC4EF , 32'hFFFF02AA , 32'hFFFF132F , 32'hFFFE5A77 , 32'h00014729 , 32'hFFFDFF68 , 32'hFFFFF4B5 , 32'h0001E68D , 32'h0004CC8E , 32'hFFF9F96D , 32'hFFFCA5E4 , 32'h000189DC , 32'hFFFFD2FB , 32'h00009F2E , 32'hFFFA9CB0 , 32'hFFFE77E9 , 32'h00008D53 , 32'hFFFCBE6F , 32'hFFFD0536 , 32'h000089DD , 32'hFFFCBE9B , 32'hFFFFA3CD , 32'hFFFDB417 , 32'h00050865 , 32'hFFFD5350 , 32'hFFFBD4D8 , 32'h0002C98A , 32'hFFFD17FF , 32'hFFFF02F8 , 32'h00036320 , 32'hFFFF5B33 , 32'h00006BFF , 32'hFFFBEC48} , 
{32'hD7EB14C0 , 32'h1E2A3120 , 32'h10E3B380 , 32'h314F8640 , 32'hFC4F27C8 , 32'hDDE5A380 , 32'h23712A40 , 32'hFAC23608 , 32'hD2C94380 , 32'h047138F8 , 32'hF804FF18 , 32'h0125A5DC , 32'h155ED340 , 32'hF09BC230 , 32'hFE8DE368 , 32'h13C98A00 , 32'h0182EB5C , 32'hF458E990 , 32'h0471EE38 , 32'h0BFC2C30 , 32'h18A3CBE0 , 32'h00BFB3AD , 32'h0511C100 , 32'h05236B98 , 32'hFF36C056 , 32'h0B7257C0 , 32'h06D20AC8 , 32'hF8ABBB10 , 32'hFEFF41CC , 32'hEA6ADB00 , 32'h10C84240 , 32'h04B04710 , 32'h09B9AB20 , 32'h01ABCF84 , 32'hF8471520 , 32'h0C341430 , 32'h0945FB30 , 32'hFE396830 , 32'h05CCB058 , 32'hF907A878 , 32'hFFD0CE2F , 32'h02C86B44 , 32'h05AB58F0 , 32'h085C0EF0 , 32'h03B67A60 , 32'h0407A930 , 32'h028F1E70 , 32'hFEA9C8DC , 32'h13E71180 , 32'h0688F100 , 32'h07233528 , 32'hFDF2DD20 , 32'hF264A2A0 , 32'hF361B190 , 32'hF8E0CC80 , 32'h08459000 , 32'hFC991D0C , 32'hF5752300 , 32'hF8869BB0 , 32'hFED127A0 , 32'h016BF248 , 32'hFD9D9B4C , 32'h0816CDB0 , 32'hFD6B90EC , 32'hFBC3DDA8 , 32'hFB9DE730 , 32'hFB0DA440 , 32'hF94FAF98 , 32'h04919B38 , 32'hFF50970A , 32'h01E49E00 , 32'h06631488 , 32'hFBFF3CA0 , 32'h00F85B8E , 32'h03B68B28 , 32'h038290C0 , 32'hFE931708 , 32'h018308D8 , 32'hFB3B4240 , 32'hFE7B91F0 , 32'hFC81C254 , 32'h019DE524 , 32'hFF2FC087 , 32'h00ECFCC0 , 32'h0296AAAC , 32'h01D4D7D8 , 32'hFA9488F0 , 32'h01F0ABB0 , 32'hFFDB8626 , 32'h00A1FEDB , 32'hFFFFDE9D , 32'hFFFCE077 , 32'hFFFF49EF , 32'h0001A36E , 32'hFFFECDF2 , 32'h00005852 , 32'h0000DAD3 , 32'h0000BC7A , 32'h000183FE , 32'hFFFF4580} , 
{32'h04A4BDD8 , 32'h0A063CE0 , 32'hF24A95F0 , 32'h041B8768 , 32'h05173370 , 32'h1D5E4980 , 32'h037BBA34 , 32'hFE8A2C98 , 32'hFC0BA4FC , 32'hF8447928 , 32'h0A18C0B0 , 32'hF6DFC580 , 32'h075D5DB8 , 32'h049263F8 , 32'hFDB9D150 , 32'h0135824C , 32'h06D1BC70 , 32'h06B82800 , 32'h024D0FBC , 32'h0CE1DA20 , 32'hF7BA2620 , 32'hFF189DA5 , 32'h15480BC0 , 32'hF646FC20 , 32'hF8D4CD28 , 32'hFD426580 , 32'h0BFB8330 , 32'h0A1B67A0 , 32'hF86FD598 , 32'hFDF1FA74 , 32'h0A2F6630 , 32'hF82E8010 , 32'h10731FA0 , 32'hEB595620 , 32'hEFF25AA0 , 32'hEDF14A20 , 32'h0045ACB1 , 32'hFEB78C04 , 32'h09CF9370 , 32'h077F22F0 , 32'hF0D1AE60 , 32'h0C010480 , 32'hFB03A460 , 32'hFAE59418 , 32'h00CE5EAF , 32'hF16D94F0 , 32'h0EC21B00 , 32'h04EA8EB0 , 32'h087D8C70 , 32'h02247370 , 32'hF3F7AAA0 , 32'hFFA32BBA , 32'hFB60B858 , 32'h02DBDDFC , 32'hFCC61768 , 32'hFD74E3BC , 32'hFD6CC550 , 32'h0082933C , 32'h036047EC , 32'h00789D53 , 32'hFD16C04C , 32'h083D14B0 , 32'h004CCFE7 , 32'h0163FAB0 , 32'h07EB6198 , 32'h01F1A100 , 32'hFE9CC118 , 32'h04A1E640 , 32'hFCE2E134 , 32'hFDCE9D24 , 32'h073AFE38 , 32'hFA9C61F0 , 32'hFC9FC7CC , 32'h02E5E3A0 , 32'hFE231C54 , 32'hFB14EB80 , 32'h0DDA0980 , 32'h012FD2F4 , 32'h03D665D0 , 32'h04F16F70 , 32'hFE3D347C , 32'h0468F050 , 32'hFE534850 , 32'hF9732198 , 32'h008B3920 , 32'h02F8B45C , 32'h02D6FFE4 , 32'hFF11B942 , 32'hFFE1CEC7 , 32'h005405F4 , 32'hFFFECA36 , 32'hFFFF2CEA , 32'h00017121 , 32'h00002B2C , 32'hFFFC887A , 32'hFFFF1C89 , 32'h00001AC6 , 32'h00008095 , 32'hFFFE0B9D , 32'hFFFF9391} , 
{32'hFFFF1A52 , 32'hFFFFF80B , 32'h0003EE66 , 32'h0000D640 , 32'h000409DA , 32'h000305F0 , 32'hFFFD5033 , 32'h0001557A , 32'h0000CA50 , 32'hFFFEBF33 , 32'h000541C2 , 32'hFFFFC7D7 , 32'h0000726E , 32'h00007DED , 32'h000519CA , 32'hFFFAD4DA , 32'hFFFE6194 , 32'hFFFEC595 , 32'h0001D810 , 32'hFFFDBF1F , 32'hFFFF967F , 32'hFFFEAA8B , 32'hFFFCE187 , 32'h00035644 , 32'hFFFD2DB8 , 32'h0002C924 , 32'h000121E1 , 32'h0000709C , 32'h0000BF80 , 32'h00026C6E , 32'h00021270 , 32'hFFFE3755 , 32'hFFFEC542 , 32'hFFFB7744 , 32'hFFFFDC3D , 32'hFFFD05B2 , 32'h00018795 , 32'h000166DC , 32'h000237BB , 32'hFFFCC0CF , 32'h00023AA0 , 32'hFFFA0751 , 32'hFFFCDAF6 , 32'hFFFF70B9 , 32'hFFFAB1EC , 32'hFFFA76A5 , 32'hFFFC6E11 , 32'h00020FCF , 32'hFFFC914D , 32'hFFFD4CC2 , 32'h00010DB2 , 32'h00002180 , 32'h00022913 , 32'hFFFEFD43 , 32'h0001A8C7 , 32'h000288AD , 32'hFFFF560C , 32'h0001C4CE , 32'h00039829 , 32'h00029015 , 32'h0000DAD9 , 32'hFFFE78A6 , 32'h0001FDA0 , 32'hFFFF1C96 , 32'h000162ED , 32'h0002627C , 32'hFFFCD1AB , 32'hFFFADFC3 , 32'hFFFE8BA7 , 32'h0003EEA7 , 32'hFFFF0F1B , 32'h0003AD3E , 32'h00013C43 , 32'hFFFD3770 , 32'h00047079 , 32'hFFFFB897 , 32'h0003BB75 , 32'hFFFF1424 , 32'hFFFB595F , 32'h00022BED , 32'hFFFF5398 , 32'hFFFEF384 , 32'h0002FBED , 32'hFFFE260A , 32'h0004A369 , 32'hFFFEE893 , 32'hFFFE84B7 , 32'hFFFE0461 , 32'hFFFE3040 , 32'hFFFC7A63 , 32'hFFFE75CF , 32'hFFFDD591 , 32'h0002CC3F , 32'h00018A77 , 32'h0000A767 , 32'hFFFB7E36 , 32'hFFFFD18C , 32'h00005635 , 32'hFFFFBFB6 , 32'h00048799} , 
{32'h0001C1F1 , 32'h0001A685 , 32'hFFFB744F , 32'hFFFC22EF , 32'hFFFF8F31 , 32'hFFFFAC15 , 32'hFFFEDF76 , 32'h000052AA , 32'hFFFCCDFF , 32'h0004EFF4 , 32'hFFFDEFE9 , 32'hFFFDC046 , 32'hFFFCCFB9 , 32'h00005554 , 32'hFFFF3F61 , 32'hFFFBE7EB , 32'hFFFCBF79 , 32'h0003855D , 32'hFFFE01B3 , 32'hFFFF507D , 32'hFFFFD893 , 32'h00029A89 , 32'h00006695 , 32'hFFFDDC6E , 32'h000184C0 , 32'hFFFF179E , 32'h00056E11 , 32'h0002429D , 32'h00011DC7 , 32'hFFFF13E1 , 32'hFFFC9681 , 32'h0003BD75 , 32'hFFFF8025 , 32'h00026096 , 32'hFFFF5E12 , 32'h000045CA , 32'hFFFFD8F7 , 32'hFFFDEFE8 , 32'hFFFD1ACF , 32'hFFFFD2EE , 32'h000089E6 , 32'hFFFD540F , 32'h0001BA53 , 32'h0004D08B , 32'h0001D396 , 32'hFFFF1C74 , 32'hFFFC4B0C , 32'h0003B82D , 32'h00051DD9 , 32'hFFFBA4A9 , 32'hFFFEB443 , 32'hFFFF05B7 , 32'hFFFF57B7 , 32'h0004EEE9 , 32'hFFFE8064 , 32'h0006DB44 , 32'h0002C2DD , 32'h000130BC , 32'h00009262 , 32'h00012B33 , 32'hFFFD2286 , 32'h0000B4F4 , 32'h0008BA45 , 32'hFFFF1F97 , 32'h00002233 , 32'h000024B2 , 32'h0001CD9D , 32'hFFFD8128 , 32'h0002E2F5 , 32'hFFFFE7E9 , 32'h0004F825 , 32'hFFFF4CF6 , 32'hFFFFB3AE , 32'h0000511C , 32'h000314E1 , 32'hFFFF9030 , 32'h00036CB1 , 32'h00040AB7 , 32'h00000386 , 32'h0001A976 , 32'hFFFF912C , 32'hFFFAA131 , 32'hFFFCDDC3 , 32'h0004CCF3 , 32'hFFFE10AF , 32'hFFFFA612 , 32'hFFFEF942 , 32'h0005C035 , 32'hFFFC3312 , 32'hFFFE5EFF , 32'h0001A8BC , 32'hFFFB6AD2 , 32'hFFFE4E49 , 32'hFFFFCE9B , 32'hFFFE10A5 , 32'h00007471 , 32'h0000A3F6 , 32'hFFFC8E9E , 32'hFFFE81AB , 32'hFFFFAC6F} , 
{32'hFC98BA04 , 32'h00ABF813 , 32'h07C12448 , 32'h06D63FC8 , 32'hFFCAE336 , 32'hF7DAFB80 , 32'hF9959BC0 , 32'hFDDB7804 , 32'hFFB2498A , 32'h0084E3B5 , 32'h073A6960 , 32'hFD71E258 , 32'h07588718 , 32'h014157E8 , 32'h06641280 , 32'h011492FC , 32'h06777498 , 32'hFB143DF0 , 32'h068E7A90 , 32'h017AE78C , 32'hFB418518 , 32'hFBBD4DC8 , 32'hFD5F71C8 , 32'hFEE66070 , 32'h03626D78 , 32'h081FB990 , 32'hFE84C3EC , 32'hF66A35B0 , 32'hFCEEC718 , 32'hF74184F0 , 32'hFADA51F0 , 32'h0824D520 , 32'h02802E18 , 32'h0068B9BA , 32'hFF9DCFDD , 32'hF9072C00 , 32'hFFA90CED , 32'h0185C4C8 , 32'h0017BED8 , 32'hFC06C6B4 , 32'hFF6F2085 , 32'hFFBF5BD4 , 32'h01A7D450 , 32'hFE0B193C , 32'hFE09B39C , 32'hFC81D2D0 , 32'hF9D78880 , 32'hF7A7C7A0 , 32'hFB87D508 , 32'h023BE5CC , 32'hFCE73AE8 , 32'h01E10270 , 32'h00FE001F , 32'h032DB3B0 , 32'h02E4FD10 , 32'h01488C08 , 32'hFF603CA0 , 32'hFFF2F4E4 , 32'h013ADDB0 , 32'h013E9EE0 , 32'hFEC55FEC , 32'h04ABADC0 , 32'h001A9B5A , 32'hFB8B7498 , 32'h032AD7D8 , 32'hF68911F0 , 32'hFFD48684 , 32'h01C0295C , 32'hFD96ADD0 , 32'hFEA62884 , 32'h040E4308 , 32'hFDF7CF78 , 32'hFDBC1BDC , 32'hFE3411B8 , 32'h008500E0 , 32'h0029A739 , 32'hFD1614F0 , 32'hFEA4460C , 32'h0138612C , 32'h02052C94 , 32'h01572A04 , 32'hFF8E79C5 , 32'hFFED4476 , 32'h002D9D23 , 32'h00863E6D , 32'h02BF60B4 , 32'h014C0120 , 32'h01B13C7C , 32'h02AAC58C , 32'hFF93C6D4 , 32'h00023934 , 32'hFFFE3517 , 32'hFFFE10F4 , 32'hFFFDE579 , 32'h0000E21C , 32'h000050CF , 32'h000133FB , 32'hFFFE7D3C , 32'h0003E956 , 32'h00001A3E} , 
{32'h0A23E830 , 32'hFB39CE08 , 32'h27A8A400 , 32'hF4A95990 , 32'hEAF99580 , 32'h087B3980 , 32'hF8F34208 , 32'hE426C4E0 , 32'h0BB22370 , 32'hFB63F730 , 32'hFA23D3A8 , 32'hFBAEB860 , 32'hFDCECDD8 , 32'hF42E07F0 , 32'h0061EA19 , 32'hF5435E80 , 32'hF6AF9A60 , 32'hF8ECAC68 , 32'h0D1701F0 , 32'h043F1748 , 32'hF88BA5F8 , 32'hFC85A790 , 32'hF35E7B90 , 32'hFB5DA600 , 32'hF4857F80 , 32'h021CA028 , 32'hF2D53EC0 , 32'h024BA350 , 32'hF9FEFD10 , 32'hF8F893B8 , 32'hEAB1B520 , 32'h01D71844 , 32'h088FA440 , 32'hF4A17E70 , 32'hFEBA6930 , 32'hF96F1378 , 32'h0F031CF0 , 32'hF9E4C3B0 , 32'hFB868C68 , 32'h0BFA84A0 , 32'h04F8AB30 , 32'h09798140 , 32'hF6941890 , 32'hFDC88704 , 32'hF46F4BE0 , 32'hF61A9C30 , 32'hFDDC8A08 , 32'hFD1E4A40 , 32'h09855A00 , 32'hFD135E34 , 32'h079C2F80 , 32'hF7232110 , 32'hFD8821D8 , 32'hF67ADD50 , 32'hF61C40D0 , 32'hF83D4CB0 , 32'hF6AA85D0 , 32'hF790AF90 , 32'hFAD412F8 , 32'h0820ADA0 , 32'hFD0354AC , 32'hFF934707 , 32'h00381978 , 32'hFE689654 , 32'hF5581430 , 32'h02A0C444 , 32'h0644B118 , 32'h019F9BDC , 32'hFF8DC74C , 32'h05F1E720 , 32'h02AFA36C , 32'h081B57C0 , 32'hFD9C9C50 , 32'hFA001488 , 32'h030801C8 , 32'h0518CC90 , 32'hFE5D0A98 , 32'h0327DAE0 , 32'h076A19F8 , 32'h04DBFF48 , 32'h043CF0C0 , 32'hFF0DD98F , 32'hFE0194E0 , 32'h02AE89F8 , 32'h00812B73 , 32'h043DEA30 , 32'hFE6990C4 , 32'h00E8AD9A , 32'hFFC47288 , 32'hFFFBA7D4 , 32'hFFFEBAA8 , 32'hFFFD4399 , 32'hFFFF61B1 , 32'hFFFEB004 , 32'h0000C6B1 , 32'h0000BDBF , 32'hFFFCBF8D , 32'hFFFF8E4D , 32'h00034FA0 , 32'hFFFF2320} , 
{32'hE5198AA0 , 32'h050BB4C0 , 32'h14BDEE60 , 32'hE1A1AE80 , 32'hF33ABDE0 , 32'hEF8569A0 , 32'h06615F20 , 32'hEF89A6E0 , 32'h098E7AF0 , 32'hE4E25240 , 32'hFB6560E8 , 32'h145D75E0 , 32'h0DBEA620 , 32'hFE6885CC , 32'hF947C700 , 32'hEFB38100 , 32'hF5829C40 , 32'hF5468B40 , 32'hF096E670 , 32'h156912C0 , 32'hF40BA350 , 32'hF613BC50 , 32'hFBFA9B50 , 32'hF508A8A0 , 32'hF501A290 , 32'h166E03C0 , 32'h037C6B80 , 32'h098236E0 , 32'hF7E899D0 , 32'hE97721C0 , 32'h0C59A720 , 32'h00C0E39E , 32'hECC51EA0 , 32'hF19521C0 , 32'hFB727FB0 , 32'h01E3B12C , 32'hF5E6B9F0 , 32'h00E790FA , 32'h003B622E , 32'h050E2C38 , 32'h04DDF490 , 32'h0A296570 , 32'h0505D7A0 , 32'h030CBE40 , 32'hFD58B7DC , 32'hFD4BBCE4 , 32'h056E04B0 , 32'h027B6138 , 32'h02BFBECC , 32'h00D5F235 , 32'hFBC87E08 , 32'h02226BDC , 32'hFDDA5180 , 32'hFBB72BB8 , 32'hFA971350 , 32'h06703968 , 32'h0B440FF0 , 32'h00ECE20E , 32'h087B8270 , 32'hF5650C70 , 32'h08300E60 , 32'hFE2BA4A4 , 32'h08D30DB0 , 32'hF2F65540 , 32'h05817E80 , 32'h02CB8CE0 , 32'hFB5CC8C0 , 32'h01C5F14C , 32'h008577D7 , 32'hFEBB3E48 , 32'h036346A0 , 32'h06A96518 , 32'h031FEAB0 , 32'h053A1020 , 32'h00A56C80 , 32'hF97C9C60 , 32'hFF5E4B97 , 32'h016778E0 , 32'hFDF1D8DC , 32'hFE928774 , 32'hFE845EC4 , 32'hFFBD29D8 , 32'h04377158 , 32'h01C72E1C , 32'h00AC4518 , 32'hFC68A7A0 , 32'hFFEBD68A , 32'h00A20BF9 , 32'hFDB28258 , 32'hFFD0D7B7 , 32'hFFFF3E7B , 32'hFFFE0DCF , 32'h000072FE , 32'h00015FFC , 32'h00002BAD , 32'h000274E9 , 32'hFFFC06C8 , 32'h0000F1F8 , 32'h0002CF88 , 32'hFFFF95C1} , 
{32'hD3A65F00 , 32'h163760E0 , 32'h22ECAA40 , 32'hFE359D1C , 32'hFF459953 , 32'h0BBFDA00 , 32'h0EBFC200 , 32'hF5676DD0 , 32'hF2791110 , 32'h166335A0 , 32'hEAFD9D20 , 32'h08E19FE0 , 32'hFD6CA718 , 32'hFCC0FFCC , 32'hED53C0C0 , 32'hE645BD80 , 32'h138079A0 , 32'h0218CEC0 , 32'h08ED8480 , 32'hF39DE070 , 32'h007FEEC3 , 32'hF2855010 , 32'h008467C6 , 32'h014991F4 , 32'h140C5D40 , 32'hF174D540 , 32'hFE0B40A4 , 32'hF64C7A40 , 32'hFC7FE1EC , 32'hE9B4B140 , 32'h062A4070 , 32'h0CE00160 , 32'hFF69CA5E , 32'h0561B1B0 , 32'hF7D759E0 , 32'h0298ADB4 , 32'hFAB4D7F8 , 32'hFA19FC38 , 32'hFB7AEE78 , 32'h0BAE2990 , 32'h01E350E4 , 32'h056C3C68 , 32'hF4858DC0 , 32'hFD150C28 , 32'hFF8F6874 , 32'hFB23F918 , 32'hF2C1ECF0 , 32'h0238C4E8 , 32'hF18A8630 , 32'hFF15B3F6 , 32'h02D59C88 , 32'hF85B9360 , 32'hFF34537B , 32'h0B1850D0 , 32'h09ECA8C0 , 32'h074145D0 , 32'h03E73A28 , 32'hEFFD4060 , 32'h08380E90 , 32'hFF788360 , 32'hFF074D54 , 32'hF7985DA0 , 32'h0C281600 , 32'hF492A9C0 , 32'h0D723D50 , 32'h024F4764 , 32'h03CDD610 , 32'hFE5B3508 , 32'hFEAE94CC , 32'hFCFCD754 , 32'hFE3EA6D0 , 32'h004734BF , 32'h0652D210 , 32'hF7E9ED50 , 32'hF99C5AA0 , 32'h07DD3708 , 32'h001B41E1 , 32'hFFB98820 , 32'hFFD7B932 , 32'hFB1BA7A0 , 32'h008D575E , 32'h029DA4D8 , 32'h013CE4DC , 32'hFAFD2D50 , 32'h0200BEC8 , 32'hFF740708 , 32'h00B9B46F , 32'hFEBCC880 , 32'hFE52B278 , 32'hFF84AC8B , 32'h0001714F , 32'h0001B2C4 , 32'hFFFDAFE1 , 32'h0000D799 , 32'hFFFE8AEF , 32'hFFFDAEAF , 32'h000097E7 , 32'h000054D4 , 32'hFFFF5321 , 32'h00015642} , 
{32'h00011F00 , 32'hFFFDBAF1 , 32'h0002FEE5 , 32'hFFFDF089 , 32'h0001C186 , 32'h00063E30 , 32'hFFFB2202 , 32'h0001226E , 32'h00036460 , 32'h00003D7A , 32'hFFFA5771 , 32'hFFFF71F2 , 32'hFFFEE25E , 32'h0005D35B , 32'h0003524F , 32'hFFFEF3A6 , 32'h000325EF , 32'hFFFF3032 , 32'h00028519 , 32'h000206A5 , 32'h00022244 , 32'h00002F8F , 32'h00014814 , 32'h0000AF88 , 32'hFFFB388B , 32'h0000CE7F , 32'hFFFD6648 , 32'h00068F97 , 32'hFFFE1FF3 , 32'h00016B5D , 32'hFFFDFD20 , 32'h00023CE2 , 32'h00031667 , 32'hFFFE50DA , 32'h00018598 , 32'h00023B8A , 32'hFFFF4230 , 32'hFFFFCDFC , 32'hFFFBF857 , 32'h00010098 , 32'hFFFEAD0E , 32'h00024457 , 32'h0002473F , 32'h00030DED , 32'hFFFF1D7C , 32'h000462DA , 32'hFFFAFC34 , 32'h000289EF , 32'hFFFE1387 , 32'hFFFF3A11 , 32'h0000E063 , 32'hFFFFBDD0 , 32'hFFFEBA0B , 32'h00021FB5 , 32'hFFFDBD11 , 32'h0000F969 , 32'hFFFFF307 , 32'h0001221C , 32'h0004DDE2 , 32'h0005572B , 32'h00035327 , 32'h0001D769 , 32'h0003CF05 , 32'hFFFB5798 , 32'h0000F610 , 32'hFFFDA528 , 32'hFFFE6646 , 32'h0003775C , 32'h00021E07 , 32'h00058F75 , 32'hFFFE6CDC , 32'h00007934 , 32'h000009AF , 32'hFFFEB2F0 , 32'h00019433 , 32'h0000B503 , 32'hFFFEAD2C , 32'h0002D5B0 , 32'h00021748 , 32'h0004DE83 , 32'h00002911 , 32'h0001896C , 32'h00026036 , 32'hFFFCCBA8 , 32'h00060B69 , 32'h00019501 , 32'hFFFF57C5 , 32'hFFFBCEE4 , 32'h00003867 , 32'hFFFF3F24 , 32'hFFFBA96D , 32'h00029AD9 , 32'hFFFCED4A , 32'hFFFCDDE4 , 32'h0002615C , 32'hFFFFED5B , 32'h00024407 , 32'h0000584E , 32'hFFFBE297 , 32'h000040F1} , 
{32'h00087438 , 32'hFFD72676 , 32'h00CE60E6 , 32'hFDD84ED8 , 32'hF3781A30 , 32'h021988D4 , 32'h031429F8 , 32'hFFD0B014 , 32'h04B365E0 , 32'h0857A6E0 , 32'h014AB8D0 , 32'h02EE6E50 , 32'hFAF9DA60 , 32'h07955838 , 32'h040F06F0 , 32'hFABE64A0 , 32'h070EF170 , 32'hFEB830CC , 32'hFF6B2072 , 32'h02E0E498 , 32'h00E97627 , 32'h089509F0 , 32'h05AF1158 , 32'hF86419A0 , 32'h006A4D4E , 32'h0D456660 , 32'hF677CCA0 , 32'hFAB51408 , 32'h0820C480 , 32'hFF0CB772 , 32'h00F12F3A , 32'hFD5896A0 , 32'h06C355F0 , 32'hF9774420 , 32'h05D61518 , 32'hFDF24D70 , 32'hF7E23120 , 32'hFAFBF408 , 32'h09F012F0 , 32'hFEE4F65C , 32'h013F5704 , 32'hFCE3B608 , 32'h08620C30 , 32'hF40CDDF0 , 32'h070BF100 , 32'hFF72C417 , 32'hFDC60DD8 , 32'hF7098C10 , 32'hFB3809A8 , 32'hF9CEC518 , 32'h00B41509 , 32'hFEEFD69C , 32'hFFD722EB , 32'hFB26A778 , 32'hFD355BB0 , 32'hFF4D2357 , 32'h04646DB0 , 32'h05D23518 , 32'h0271A8AC , 32'h0242B250 , 32'h005AAF60 , 32'hFCD1AD0C , 32'hFBE8FAA8 , 32'hFBEA3490 , 32'h03352A70 , 32'hFDC7BFA0 , 32'hFB594810 , 32'hFB4878D0 , 32'h0092FC59 , 32'h026C8F10 , 32'h067C6C68 , 32'h01612F58 , 32'h043DB4E0 , 32'hFE54432C , 32'hFFD488AF , 32'hFD706414 , 32'h00482012 , 32'hFF9C70AB , 32'h049B5A40 , 32'hFB357198 , 32'hFD410784 , 32'hFF2C7359 , 32'hFEA1C53C , 32'hFEE6DCE4 , 32'h01C1D198 , 32'hFB401390 , 32'hFD95B680 , 32'hFD999664 , 32'hFD680890 , 32'hFFD39413 , 32'h00005D56 , 32'hFFFEE37E , 32'hFFFCC152 , 32'hFFFE42E4 , 32'hFFFF1275 , 32'hFFFF1CE6 , 32'hFFFDC6F9 , 32'hFFFF2140 , 32'h0000D83A , 32'h00004489} , 
{32'hF8573CB0 , 32'h07B14098 , 32'h00BEE9D8 , 32'h06345288 , 32'h024D743C , 32'h01CF4828 , 32'hFC250AC0 , 32'h0004A711 , 32'h07064498 , 32'hF60B7550 , 32'hFF6297C2 , 32'h01172388 , 32'h02005660 , 32'h0C606440 , 32'h01E29E60 , 32'hF6C36DA0 , 32'hFD8F2F8C , 32'hFB616608 , 32'h08A3A6B0 , 32'hFD35A710 , 32'h0B3ACA70 , 32'hFFD69A98 , 32'h023F3DCC , 32'hFC62436C , 32'hFFE0D3BE , 32'hFD685D7C , 32'h01DC509C , 32'h007E0406 , 32'h04D4F170 , 32'hFC1B0558 , 32'h00B85E55 , 32'hFDEABC48 , 32'h03605CCC , 32'h0371D180 , 32'hFDCC8414 , 32'hFF38FC9D , 32'hFFBDA7A7 , 32'h01530504 , 32'hFF291D32 , 32'h01ADEA7C , 32'h00DE9B18 , 32'h047412B0 , 32'h012573FC , 32'hFEA1F6E0 , 32'h05791D58 , 32'hFE017690 , 32'hFD55DFAC , 32'hFFA00A10 , 32'h010C3158 , 32'hFA409AC8 , 32'h00DACB0D , 32'hFB2A8D38 , 32'hFE07FD2C , 32'h00F2C8D9 , 32'h04E958E8 , 32'hFE124B00 , 32'hFCF88FEC , 32'hF97A3130 , 32'h01B8D93C , 32'hFB707D88 , 32'h05B849A8 , 32'h00B67189 , 32'hFFE29F22 , 32'hFF8B1203 , 32'hFC351718 , 32'h037398CC , 32'hFDA7D028 , 32'hFF40567A , 32'hFBFE9060 , 32'h053C3988 , 32'h047E6B60 , 32'h02C9C8FC , 32'hFEABAC78 , 32'h0228D694 , 32'h00D54F54 , 32'h046DCFC0 , 32'h01340A58 , 32'h00C743D1 , 32'hFFAC222E , 32'hFAD8EEE8 , 32'h005C7297 , 32'h02DAB764 , 32'hFE57E3E8 , 32'h01445FF8 , 32'h01A1A75C , 32'h00A2EECB , 32'hFD04D250 , 32'hFDD109B4 , 32'h0012F81B , 32'h0044DF1E , 32'h0001AAA1 , 32'hFFFC7603 , 32'hFFFED5F5 , 32'hFFFFCEC5 , 32'h00043DEC , 32'h000187CE , 32'h00027D7E , 32'hFFFCF4B1 , 32'hFFFEF3BE , 32'h00010DFF} , 
{32'hFFFFA691 , 32'hFFFC7266 , 32'hFFFFF626 , 32'hFFFCBB54 , 32'hFFFE8D86 , 32'hFFFBF7D4 , 32'hFFFE4C28 , 32'h00028DB4 , 32'hFFFC5EC2 , 32'hFFFFDA5F , 32'hFFFDB4A2 , 32'hFFFF778F , 32'hFFFEE7BC , 32'h0004451A , 32'hFFFC56B5 , 32'h00018E90 , 32'hFFFD809D , 32'hFFFECDE3 , 32'hFFFF954D , 32'hFFFE7E07 , 32'hFFFAEFA4 , 32'h00001300 , 32'hFFFCEF1C , 32'h0000CE47 , 32'h0003CCE2 , 32'h000574E3 , 32'h00024A8F , 32'hFFFF6AB9 , 32'hFFFEA08A , 32'h0000B595 , 32'h00039959 , 32'hFFFC39F8 , 32'hFFFA4223 , 32'h000057E2 , 32'hFFFFA8D2 , 32'h000139CA , 32'hFFFEF60A , 32'hFFFF79AA , 32'h0003DE27 , 32'h0000E426 , 32'h00014F2B , 32'h00029EC2 , 32'hFFFEC3AC , 32'hFFFE47B0 , 32'hFFFAC2C9 , 32'hFFFF211D , 32'hFFFFDDDB , 32'hFFFCA6D5 , 32'hFFF768A0 , 32'hFFFBE005 , 32'hFFFFEA04 , 32'h0002C5CF , 32'h00009953 , 32'hFFFF0E86 , 32'hFFFF3060 , 32'hFFFE2BD5 , 32'h0004D915 , 32'h00021E49 , 32'h0002F78F , 32'h000121E1 , 32'h0000AD8F , 32'hFFFE2BED , 32'hFFFFED00 , 32'h0001F151 , 32'hFFFDB676 , 32'h0003A241 , 32'hFFFE6881 , 32'h00018D51 , 32'h0000875C , 32'hFFFF1C7C , 32'hFFFEE289 , 32'h000238AD , 32'hFFFC38AA , 32'h0001A5A3 , 32'h000031D1 , 32'hFFFFBE3F , 32'hFFFCFE15 , 32'hFFFEB05C , 32'hFFFF9356 , 32'h00020EC4 , 32'h000131D0 , 32'h000145F5 , 32'h00004F65 , 32'h0001ED91 , 32'h0003BF19 , 32'hFFFBACFD , 32'h00005039 , 32'hFFFBC260 , 32'h000219C9 , 32'hFFFFF1C6 , 32'h000214B8 , 32'hFFFD7D27 , 32'h0003FA68 , 32'h00003480 , 32'h00028441 , 32'hFFFBD4AE , 32'h0001934A , 32'hFFFAACEE , 32'hFFFFFE60 , 32'hFFFC2EEB} , 
{32'hDDF09C80 , 32'hF3C554B0 , 32'h33A25F00 , 32'hDBB99DC0 , 32'h0FDB4B10 , 32'h1379EEC0 , 32'hD850D500 , 32'hD8051540 , 32'hEC8BD5E0 , 32'h027276BC , 32'h0A289950 , 32'h1BB8B320 , 32'hF9772C68 , 32'hEC8633C0 , 32'hFB835EF0 , 32'h0A322A30 , 32'h2128EF00 , 32'h03E11140 , 32'h0536F5A8 , 32'hD7DD8D40 , 32'h1B0C3AC0 , 32'hF97543C8 , 32'hDC6D2700 , 32'hF40117E0 , 32'h04072ED0 , 32'hFDD44DE8 , 32'h024563B0 , 32'hFBF43878 , 32'hF0341D40 , 32'h091EE450 , 32'hFDD39CA8 , 32'h005FFB89 , 32'h0EC792B0 , 32'hEF4AAEC0 , 32'hF4EC8A70 , 32'h12391A60 , 32'h0234D5AC , 32'h1730AEC0 , 32'h11CCF1E0 , 32'h07657988 , 32'hF46AC0F0 , 32'h01A7D034 , 32'hF949E870 , 32'h0C59ED80 , 32'h04A0D6A8 , 32'h011FEA30 , 32'h0B12E7F0 , 32'hF73F8C70 , 32'h0720C660 , 32'h0C561B70 , 32'hF8CEF990 , 32'hFC55E500 , 32'hFAF45650 , 32'h0304BD64 , 32'hFDAE843C , 32'h01633ADC , 32'h121EE960 , 32'h00FC73B8 , 32'hFB922BE0 , 32'h0003E34A , 32'hF31E5230 , 32'h048161B8 , 32'h036C6F58 , 32'h039C1EDC , 32'hFB52CF98 , 32'h0609FAB8 , 32'h09894AC0 , 32'hFE7EDB90 , 32'h024FD550 , 32'hFDC03B38 , 32'h03F6A534 , 32'h010EE798 , 32'hFDF51FE0 , 32'hFABF6F60 , 32'hFC977C04 , 32'h01B6E328 , 32'hFFE87934 , 32'h01EA566C , 32'h02D1611C , 32'hFE8B7444 , 32'hFEA4117C , 32'hFE9F8C64 , 32'h01E65448 , 32'hFFE04F76 , 32'hFBCEEEB8 , 32'hFFFAC24E , 32'hFD770C58 , 32'h0054FA17 , 32'h007D9AE9 , 32'h0010BC11 , 32'hFFFFBAC5 , 32'h0001624E , 32'h00007E35 , 32'hFFFCBC0E , 32'hFFFD6EEE , 32'hFFFF8E31 , 32'h000117FC , 32'hFFFF70B0 , 32'hFFFFFCDE , 32'h00009129} , 
{32'hFFFCA07F , 32'h0004B9DF , 32'hFFFE5DDD , 32'hFFFF4A5D , 32'hFFFF9FA8 , 32'hFFFE265C , 32'hFFFD7BB9 , 32'h0004D7F9 , 32'h0001D23B , 32'h0007FAE2 , 32'h00026EB8 , 32'h0000D4E6 , 32'h000228F8 , 32'hFFFF7D6E , 32'hFFFF058C , 32'hFFFE0146 , 32'h0000D541 , 32'hFFFDE861 , 32'h00011166 , 32'hFFFFAD0C , 32'hFFFFED77 , 32'hFFFE4F43 , 32'hFFFB1208 , 32'h00045DEB , 32'h00013A48 , 32'hFFFE2E0F , 32'hFFFB5D8F , 32'h000083D5 , 32'h000021E7 , 32'hFFFE9C64 , 32'h0002048B , 32'hFFFE102F , 32'h0000C578 , 32'hFFFF44C5 , 32'h00030FB2 , 32'h000805EB , 32'hFFFE2641 , 32'hFFFD91FB , 32'h00030775 , 32'hFFFAAEB8 , 32'hFFFE271B , 32'h0005AAFF , 32'hFFFE01B1 , 32'hFFFEF0F6 , 32'h00029E60 , 32'hFFFE1814 , 32'hFFFCEC2A , 32'h000021A8 , 32'hFFFC643D , 32'hFFFACD17 , 32'hFFFD3ECB , 32'h000563E8 , 32'hFFFFC026 , 32'h0002BB55 , 32'hFFFC8173 , 32'h0002C641 , 32'hFFFE97A1 , 32'hFFFCAD8C , 32'hFFFEB75D , 32'hFFFF5F2A , 32'hFFFE96C8 , 32'h00013F12 , 32'h00012ED0 , 32'hFFFE4AEE , 32'h000033E5 , 32'hFFFEDFA5 , 32'h0004CE3C , 32'hFFFEE201 , 32'hFFFD71E7 , 32'h0000610F , 32'h0001E80F , 32'hFFFFF076 , 32'h000138C6 , 32'h00065D2A , 32'hFFFEC0DA , 32'h00054D88 , 32'h0002DEE7 , 32'hFFFD69C1 , 32'h0001AE23 , 32'h000052AE , 32'h00013211 , 32'hFFFE3F80 , 32'h000398CE , 32'hFFFB0ECE , 32'h000043BE , 32'h0001677A , 32'hFFFEDFAC , 32'h0000B4BB , 32'hFFFF5514 , 32'h000031DE , 32'h00025587 , 32'h0001A889 , 32'h00024631 , 32'h000283FC , 32'hFFFB92CB , 32'hFFFA7CC4 , 32'h00000F1A , 32'h000368EE , 32'h00038B29 , 32'h00000132} , 
{32'h0DC59420 , 32'h22D2A580 , 32'hF8ED5088 , 32'h0379EFA8 , 32'h02658CD0 , 32'h13317520 , 32'hF2C0AD10 , 32'hFD0514D8 , 32'h0CD31730 , 32'hFBBD3930 , 32'hFE92F1BC , 32'hF30EA610 , 32'hF7851B30 , 32'hF089E4D0 , 32'hF5669030 , 32'h16CB8F80 , 32'h01D0A21C , 32'hFEB8C8B4 , 32'h0D3F0690 , 32'h1B440D20 , 32'h0A685020 , 32'hFF54AE20 , 32'hF6442430 , 32'hF9FEEE58 , 32'h0A76CDE0 , 32'h04BE8F20 , 32'h0A6345B0 , 32'hF89782B0 , 32'hFE215614 , 32'h0288A7BC , 32'hFEE7E480 , 32'hFF827398 , 32'h02DCAA18 , 32'hF0515480 , 32'h0AE5E190 , 32'hFECF1648 , 32'h06737550 , 32'h05A940F8 , 32'hF7697F00 , 32'hF3982920 , 32'hFE81B92C , 32'hF8562D48 , 32'h0361D294 , 32'h0213E394 , 32'h01A2D28C , 32'hFEC4D560 , 32'hFD2BF29C , 32'hFD59D8B0 , 32'h0690AB50 , 32'hFD6155A8 , 32'h0945E6E0 , 32'h0CFD27C0 , 32'h012C04E4 , 32'hFB41A878 , 32'h05768C30 , 32'h030019F8 , 32'h069346F8 , 32'h00B519E1 , 32'h0003A8EB , 32'hFD44BAEC , 32'hF8CA5748 , 32'hF31CCC40 , 32'h02A4CE84 , 32'hFE3C7FBC , 32'hF87A10F0 , 32'hFE1DB38C , 32'hFF231B62 , 32'h00783C17 , 32'hFE4E19A4 , 32'h02A5BE70 , 32'h07C95FC8 , 32'hFB229CC0 , 32'h037FC81C , 32'h027E422C , 32'hFACA0DF8 , 32'h00FA2713 , 32'h05F75728 , 32'h00DA9F10 , 32'h00DCA6C0 , 32'hFCC1D424 , 32'h01E8B630 , 32'h033251C8 , 32'hFE7888E4 , 32'h005546BF , 32'h00FC6596 , 32'hFCB0C42C , 32'h00193125 , 32'hFFBECBEE , 32'h01D94640 , 32'h002DAB80 , 32'hFFFE3949 , 32'h00000E75 , 32'h0000CCAD , 32'h00033990 , 32'h0003515F , 32'hFFFE90BD , 32'h00015922 , 32'h00063125 , 32'h00021B33 , 32'hFFFEC7E1} , 
{32'hFFFFC0C4 , 32'hFFFFB1EF , 32'h0002C6B6 , 32'h00013C64 , 32'hFFFE80AA , 32'h00020891 , 32'hFFFEE6A1 , 32'h00003716 , 32'hFFFD4EDB , 32'hFFFAB8A5 , 32'h0000C8C3 , 32'hFFFD3727 , 32'hFFFE6D56 , 32'h0003B942 , 32'hFFFF7EC3 , 32'h00037663 , 32'h0000EBF2 , 32'hFFFE22D3 , 32'h0002D20E , 32'h0001EE4C , 32'h0001DD04 , 32'hFFFC56E7 , 32'hFFFF074E , 32'h0000E84E , 32'h0000F3B6 , 32'h000058FC , 32'h00002899 , 32'hFFFEDAC2 , 32'hFFFF5866 , 32'h00018AA0 , 32'hFFFCAB7D , 32'hFFFCD4EB , 32'hFFFC3FF4 , 32'hFFFD4A6E , 32'hFFFD5E07 , 32'hFFFB6B42 , 32'hFFFF5E73 , 32'hFFFE95E0 , 32'hFFFFDAE1 , 32'hFFFD0665 , 32'hFFFF8A5F , 32'hFFFFDD4A , 32'hFFFA516C , 32'hFFFF55DA , 32'hFFFECB54 , 32'hFFFDA2EE , 32'hFFFC8574 , 32'h00021264 , 32'h000397C4 , 32'hFFFD3DBA , 32'hFFFE73AE , 32'hFFFFABEB , 32'h00030050 , 32'hFFFD3E6D , 32'hFFFBBE67 , 32'h0002DEB8 , 32'hFFFF3C91 , 32'h0001CB8D , 32'hFFFF93EF , 32'h00054C5B , 32'h0000D049 , 32'hFFFF1CD0 , 32'h000409A2 , 32'h00012E0D , 32'h0002311D , 32'h00010C55 , 32'hFFFD4BA8 , 32'hFFFE481F , 32'hFFFE8288 , 32'h0006D4FB , 32'h00066B31 , 32'hFFFF3993 , 32'hFFFC3BC5 , 32'h0000BEA8 , 32'hFFFCCD52 , 32'hFFFD861B , 32'h0001DCCA , 32'hFFFE4EDE , 32'h00021C3E , 32'h0002F8D8 , 32'h0003D944 , 32'hFFFE6B01 , 32'hFFFF34A0 , 32'hFFFC7B50 , 32'hFFFDB186 , 32'hFFFF2893 , 32'h0000C007 , 32'hFFFD6EA6 , 32'hFFFE978D , 32'h0002FDD6 , 32'h000472EE , 32'hFFFF4040 , 32'h00059B56 , 32'h0006FE80 , 32'hFFFF3E6D , 32'hFFFE5F58 , 32'h0000BBDF , 32'hFFFE46CE , 32'hFFFE5095 , 32'h00003FEF} , 
{32'hFFFF4BF4 , 32'hFFFAC5B2 , 32'h00017945 , 32'h00016A47 , 32'h0001D39B , 32'hFFFD928F , 32'h00037C5A , 32'h00019D4A , 32'hFFFEB6D1 , 32'hFFFDD8BC , 32'hFFFEEB0F , 32'hFFFFE81E , 32'hFFFF1261 , 32'h000248D9 , 32'hFFFDEC0F , 32'h00032A0E , 32'h0000C536 , 32'hFFFD9A7B , 32'h00051997 , 32'hFFFD1CCB , 32'h0001C0CD , 32'hFFFFA82F , 32'h00034BA6 , 32'hFFFEFA9A , 32'hFFFF7341 , 32'hFFFCEFAD , 32'h00006DD3 , 32'hFFFF0EBB , 32'h0003E8B0 , 32'h000079C7 , 32'hFFFC7890 , 32'hFFFF7019 , 32'h0001E927 , 32'h0003DF73 , 32'h0003601B , 32'hFFFF9273 , 32'h000075F1 , 32'hFFFB179C , 32'hFFFF23DD , 32'h0001FDBE , 32'h00010934 , 32'h00022286 , 32'h0000E68A , 32'h00019062 , 32'hFFFFA4D3 , 32'h000283EC , 32'h000040F2 , 32'h0002E877 , 32'h00009750 , 32'hFFFD3994 , 32'hFFFE176C , 32'h000003D0 , 32'hFFFFD649 , 32'hFFFB9262 , 32'h00044D27 , 32'h00028908 , 32'h0000D8BD , 32'h00041D7B , 32'h0001AC33 , 32'hFFFBDEF4 , 32'hFFFC8C7F , 32'h000249DD , 32'hFFFE36F9 , 32'hFFFF72BE , 32'h0000ED43 , 32'hFFFFB606 , 32'h0003EE03 , 32'hFFFE1B47 , 32'hFFFAC1C4 , 32'hFFFF8758 , 32'hFFFED25E , 32'hFFFD5581 , 32'hFFFC38CC , 32'h000372F1 , 32'hFFFD5007 , 32'h0000484D , 32'hFFFE8064 , 32'h0000835B , 32'h0000B183 , 32'hFFFCB129 , 32'h00047BC8 , 32'h0001AF61 , 32'h000438B2 , 32'h0000E6CF , 32'h0000C8AC , 32'h00029690 , 32'hFFFDC7B6 , 32'h000305C2 , 32'hFFFFCEC0 , 32'hFFFDF0C0 , 32'hFFF74D60 , 32'hFFFC0134 , 32'hFFFD032D , 32'h0000FBAC , 32'hFFFFC365 , 32'h0002684F , 32'h0003D667 , 32'h00033B6C , 32'h000224E3 , 32'h0003ABAD} , 
{32'hFFFFC33F , 32'hFFFF3907 , 32'hFFFB923D , 32'h00010A71 , 32'hFFF78F05 , 32'hFFFF1EC8 , 32'h0001034D , 32'h00015212 , 32'h000073E3 , 32'h000577BE , 32'hFFFA1757 , 32'h0001ED5A , 32'hFFFAEF83 , 32'h000166F4 , 32'h000352C6 , 32'hFFFDE55F , 32'h00062AAE , 32'h0003C047 , 32'h0007C382 , 32'h0004EF32 , 32'hFFFDBC58 , 32'hFFFE6529 , 32'h0001F914 , 32'hFFFEC205 , 32'h0004E21F , 32'hFFFEB66D , 32'hFFFF6DFE , 32'hFFFD0EEF , 32'h0005F469 , 32'hFFFF9F5D , 32'hFFFF0F0E , 32'h000029E4 , 32'h0001CEF4 , 32'h00018A5D , 32'hFFFFF315 , 32'hFFFE1AB9 , 32'hFFFAFAE8 , 32'hFFFC8BC7 , 32'h0003B104 , 32'h00027D50 , 32'hFFFF244F , 32'hFFFEC2A5 , 32'hFFFF9E3E , 32'hFFFC7A98 , 32'hFFFB7853 , 32'hFFFDB21D , 32'h0004152A , 32'hFFFF20C3 , 32'hFFFF03F7 , 32'h000083D8 , 32'h00033317 , 32'hFFFFE1EE , 32'h00020A22 , 32'h00018662 , 32'h00005231 , 32'hFFFF4BB8 , 32'hFFFEC4DF , 32'hFFFFE283 , 32'hFFFF4F28 , 32'h00013426 , 32'hFFFFEE63 , 32'hFFFF3297 , 32'hFFF7260E , 32'h00044FA1 , 32'hFFFC9434 , 32'hFFFFCF7A , 32'hFFF80532 , 32'hFFFDF9A1 , 32'hFFF9B513 , 32'h0000AF37 , 32'h0000E306 , 32'h0000F2FE , 32'hFFFA0024 , 32'hFFFE8E9C , 32'hFFFDF672 , 32'hFFFA4845 , 32'hFFFB5D4B , 32'h00021A9F , 32'h0002A002 , 32'h00056FDD , 32'h0000AC00 , 32'h00030AB2 , 32'h00004255 , 32'h0006A287 , 32'h00034D48 , 32'hFFFEFAAE , 32'h0001023B , 32'hFFFFA08A , 32'h0001B5CD , 32'h00041171 , 32'hFFFC5FD7 , 32'h00008BC1 , 32'hFFFDAF4E , 32'h0000A209 , 32'hFFFF02C5 , 32'h00015BD9 , 32'h00049B55 , 32'h00004ADE , 32'hFFFF8C12 , 32'h00022B70} , 
{32'hCF5629C0 , 32'hE1AF7980 , 32'hBAFB1980 , 32'h175E1D60 , 32'h3354A440 , 32'hDB294380 , 32'hFCCAFC54 , 32'h03E4D58C , 32'hFD348400 , 32'hDE5BEFC0 , 32'h05E90478 , 32'hEB3CBA40 , 32'h1204A8C0 , 32'h05F1A108 , 32'hE11AB4A0 , 32'h08F087B0 , 32'hEA1D1AE0 , 32'hE79FD3C0 , 32'hF9D3FC38 , 32'h10086600 , 32'h169F4300 , 32'hF7BAC120 , 32'hEFAA0540 , 32'h064A92D0 , 32'h0366DEC4 , 32'h1314FFC0 , 32'hDFF4CFC0 , 32'h021DF2BC , 32'hFCACAAF4 , 32'h0FCCD190 , 32'hFC0FA924 , 32'hF8CA3778 , 32'hFD5320E8 , 32'h14F74B60 , 32'hF4831220 , 32'hF270D070 , 32'hF3492AE0 , 32'h0AC846F0 , 32'hFFB726E5 , 32'h03BF2B48 , 32'hF0593580 , 32'h0DE7DBD0 , 32'hEF967160 , 32'hFEF30BF0 , 32'h03AEF95C , 32'hF9CDF088 , 32'hFD64A3AC , 32'h0F320B90 , 32'h075326E0 , 32'h065BEA18 , 32'h031556D0 , 32'hF8982358 , 32'hF59A1C20 , 32'hF83EB3E8 , 32'hFD558CF8 , 32'h091EC230 , 32'hFD9B7E50 , 32'hF8E05300 , 32'h04810CC0 , 32'h050B26D0 , 32'h02007D6C , 32'hF6FB4F50 , 32'hFC7C01D8 , 32'h05925180 , 32'h098C8430 , 32'hFD2A08B4 , 32'h045AA320 , 32'hF6BC72E0 , 32'h033EE9A0 , 32'h090EB100 , 32'h05E3D3F8 , 32'h00CBD009 , 32'hFEC56B80 , 32'hFDADE154 , 32'hFFA16CE4 , 32'h0109AAE4 , 32'hF876BF30 , 32'hFEDDA51C , 32'hFED19E50 , 32'h0551ECC8 , 32'h00EB7D7A , 32'hFD22CEA8 , 32'h019F5E8C , 32'hFD7BDB94 , 32'h0311110C , 32'hFEF19EF0 , 32'hFE95D750 , 32'hFFD2E589 , 32'h012FDC08 , 32'hFFD60B06 , 32'hFFFF914C , 32'h000068B8 , 32'h0001D4C5 , 32'hFFFEFA5C , 32'hFFFFD0F4 , 32'h00000684 , 32'hFFFF925E , 32'hFFFF8691 , 32'hFFFEE086 , 32'h00015E52} , 
{32'h0E0D8110 , 32'h13A36D20 , 32'h290D2DC0 , 32'hD63B3440 , 32'h31948600 , 32'hEDACE540 , 32'hE76CC840 , 32'h0196F46C , 32'h27668940 , 32'hFE11C398 , 32'hE13C3B00 , 32'h0555F090 , 32'h02DF61B8 , 32'h139E6A60 , 32'h0315335C , 32'hFBCC5AE0 , 32'hF8940A60 , 32'h0F5D8C90 , 32'hF30DC6B0 , 32'hF120B070 , 32'hFAD64058 , 32'h092C82A0 , 32'hEDAF83E0 , 32'h0DA55B80 , 32'h03777E30 , 32'h08BC55A0 , 32'hE77C02E0 , 32'h0FFD2AF0 , 32'h173C9380 , 32'hE493A220 , 32'hFDADAD14 , 32'hEE192A20 , 32'hF4EEDD60 , 32'h09710B60 , 32'hF96C8808 , 32'h0A675C20 , 32'hFCEAE12C , 32'h0E1DD780 , 32'hFE9FE3FC , 32'h0B7B54D0 , 32'hFA5816D8 , 32'h01C3C338 , 32'h051CCCF8 , 32'hFA047C68 , 32'hFA450E20 , 32'hF7790090 , 32'hF69C7210 , 32'hFBF83DC8 , 32'hF9A87BF0 , 32'hF55F5B40 , 32'hFD5EB100 , 32'hFAB33B30 , 32'hF6B06440 , 32'h06065F90 , 32'hEFEEA0C0 , 32'h03CC4C6C , 32'h01701F54 , 32'h02F4DF90 , 32'hFA2BA970 , 32'hFDF1BACC , 32'h01249A3C , 32'h069067C8 , 32'hFE541FC8 , 32'h06E62D38 , 32'h00FC91AB , 32'hF1071EA0 , 32'hFAA81B88 , 32'h020BA77C , 32'hFBA582E8 , 32'h003D8256 , 32'hFAC26488 , 32'hFEFC6770 , 32'hFF6D5E42 , 32'h01D37B50 , 32'hFAC47AA8 , 32'hFB4F9380 , 32'h0163DAE4 , 32'h00E1C349 , 32'h0145BF2C , 32'hFDC88A14 , 32'hFED645F4 , 32'h00A14A52 , 32'hFDF2C95C , 32'h01BFF85C , 32'hFD623E58 , 32'h00FC5EBD , 32'h012C864C , 32'hFE5163A0 , 32'h005D2691 , 32'h008C0204 , 32'hFFFF81B8 , 32'h00013CA0 , 32'h00013AE1 , 32'hFFFFC26D , 32'h00000F73 , 32'h000242BB , 32'h00017A68 , 32'hFFFE7259 , 32'h00007E16 , 32'hFFFDC7BA} , 
{32'h11DF7EE0 , 32'hE1FBAF00 , 32'hD32AB8C0 , 32'h2438D480 , 32'h0D2A8A90 , 32'hCEBB6180 , 32'hED6A6660 , 32'h19C642E0 , 32'hF630A610 , 32'h0F6B0A30 , 32'hE16BC0E0 , 32'h1973F520 , 32'h093F5AD0 , 32'h1E50ECA0 , 32'hF2221740 , 32'h0AB05BD0 , 32'hFF2DBE38 , 32'hFF0D13B4 , 32'hEC0BE040 , 32'h010EB7F8 , 32'h209AE340 , 32'hFB51BDA8 , 32'hFC17A0B4 , 32'h086DF660 , 32'h0860F730 , 32'h08409D00 , 32'hFB2CBEF0 , 32'h03D08B88 , 32'hFBEBB440 , 32'h0A710D40 , 32'hEB1061A0 , 32'h04835D70 , 32'hF698A440 , 32'hDF8DF3C0 , 32'h0A0995F0 , 32'hF89D7ED0 , 32'h12618E00 , 32'hFBEA2E18 , 32'hFC2E403C , 32'h08F11FD0 , 32'h0382B2B8 , 32'h0243FD80 , 32'hF5AE8410 , 32'hFE04FF48 , 32'h02EE2FA4 , 32'h06A74EF8 , 32'hFE1E12F4 , 32'hFEA346CC , 32'hF3CD86A0 , 32'hEE213AA0 , 32'h01484338 , 32'hFC01912C , 32'h052E2D20 , 32'h007D698A , 32'h0AB76970 , 32'hFAA14F58 , 32'hFED74994 , 32'h054DBD58 , 32'hFBC9A280 , 32'h0E9F6550 , 32'h09471F30 , 32'h07FF16C8 , 32'hFCE035B0 , 32'hF4AC45E0 , 32'h0706A9E0 , 32'h025C2B68 , 32'hFC011818 , 32'hFFD20FD7 , 32'hF91BE698 , 32'h01FAC2BC , 32'h05636C48 , 32'h009761CA , 32'h03113614 , 32'h05098BB0 , 32'h0249A50C , 32'h00DD6695 , 32'hFD1AF33C , 32'hFEA3FEE4 , 32'h0100CAF0 , 32'h01034C7C , 32'h0036E837 , 32'h00A8300B , 32'hFCEBBBA8 , 32'hFBA3C098 , 32'hFDCDE72C , 32'h03ACB0C8 , 32'h0053FA96 , 32'h0266A1C0 , 32'hFFDD6D9F , 32'h00C8A1D0 , 32'h000270EB , 32'hFFFFC671 , 32'hFFFEB7AB , 32'hFFFE61A4 , 32'hFFFF3857 , 32'h0000CD6E , 32'h0000AD46 , 32'hFFFFF735 , 32'h0000A278 , 32'h0001267C} , 
{32'hFFFE0950 , 32'hFFFD8D0A , 32'hFFFEAB7E , 32'hFFFE9763 , 32'hFFFE2C31 , 32'h0002A3B8 , 32'hFFFFA7F5 , 32'hFFFCB913 , 32'hFFFF503E , 32'h0007DA43 , 32'h0000812E , 32'hFFFF2B89 , 32'hFFF9FED5 , 32'hFFFFF113 , 32'hFFFE60B6 , 32'hFFFEAF5F , 32'hFFFFB360 , 32'hFFFE16E9 , 32'hFFFE3B23 , 32'hFFFCC32F , 32'h0001820F , 32'h0003EEB0 , 32'h0006C774 , 32'hFFFFD918 , 32'h00011E38 , 32'h000432AA , 32'hFFFDB407 , 32'h000161EC , 32'hFFFF3EF6 , 32'hFFFF90CF , 32'hFFFBFEFD , 32'hFFFEC026 , 32'hFFFE4006 , 32'hFFFA4219 , 32'hFFFFD404 , 32'hFFFDF177 , 32'hFFFDF2B7 , 32'hFFFA9F1B , 32'h000064C3 , 32'h00025A27 , 32'h0000C45D , 32'hFFFF11DA , 32'h0001FF67 , 32'hFFFE2212 , 32'hFFFDBFE2 , 32'h00027A2A , 32'hFFFE33D2 , 32'hFFFFACA3 , 32'hFFFCCA7B , 32'hFFFE0F8A , 32'h0002A888 , 32'hFFFCDB48 , 32'h0000BBD3 , 32'hFFFA35B8 , 32'hFFFFC937 , 32'hFFFBA09A , 32'h0000B8FD , 32'h00003AE5 , 32'hFFFE63B3 , 32'h00033891 , 32'h000298A8 , 32'hFFFD97E9 , 32'hFFFCE464 , 32'hFFF8FEE1 , 32'hFFFB9473 , 32'hFFFDB1E3 , 32'hFFFA438B , 32'h00015717 , 32'hFFFFC948 , 32'hFFFF51C2 , 32'h0000F5CF , 32'h00043F3A , 32'h00012B40 , 32'hFFFF48C4 , 32'hFFFF01EC , 32'hFFFE1B57 , 32'h000119DA , 32'h000123CF , 32'hFFFE3CA7 , 32'h00018799 , 32'h0000FD82 , 32'h00035BC4 , 32'h00017F8E , 32'h0001F551 , 32'h00001E0E , 32'h000249D3 , 32'hFFFBD931 , 32'hFFFEC88E , 32'hFFFFE505 , 32'hFFFFF4AC , 32'hFFFD5860 , 32'hFFFDB98C , 32'h00016390 , 32'hFFFE31DA , 32'h00008B17 , 32'h00016DF4 , 32'h00046A66 , 32'hFFFF94EB , 32'h0002E9AB , 32'h0000CF58} , 
{32'h21D39700 , 32'h20CB0080 , 32'h07118720 , 32'h0B25EA90 , 32'hFCC9CAE4 , 32'hDF4CBA80 , 32'hECACA240 , 32'hFC8557BC , 32'h467B8800 , 32'h1F960C00 , 32'h00729907 , 32'hFCEF4D30 , 32'h0B4472C0 , 32'h088C2B90 , 32'hDEF3CBC0 , 32'hF0BEA870 , 32'hFB4917E8 , 32'hE8BE4A40 , 32'hF7CD3DF0 , 32'hE877FC80 , 32'h092A1180 , 32'h01AD5AFC , 32'h1A67B7A0 , 32'h0201D424 , 32'h06D4D0C8 , 32'hF9E05F80 , 32'hF3C28EF0 , 32'h03D11DE0 , 32'hF3554D50 , 32'h1140F420 , 32'h0037E6E4 , 32'h02AA46CC , 32'h015CA6D4 , 32'hF86BB120 , 32'hF6FEEB70 , 32'hF926CBC0 , 32'h05C14750 , 32'h07220638 , 32'hF210C9A0 , 32'hFBDBE0C0 , 32'h069554E0 , 32'h0344C1DC , 32'hF26EEEE0 , 32'h0A0C0170 , 32'h039FA514 , 32'h03EDEC04 , 32'hFDA2C6B4 , 32'hF2268AF0 , 32'hFD5BCB40 , 32'hFD59AE40 , 32'hF5050D00 , 32'hFD2DFE64 , 32'hFBD98CF0 , 32'hFB5DF3D8 , 32'hFB9352B0 , 32'h09156410 , 32'hF8E8BD10 , 32'hFA416D08 , 32'hFB12EF80 , 32'hF6E891A0 , 32'hFD387358 , 32'hF993C830 , 32'hFE3E2EB8 , 32'h0778C6E8 , 32'hF6E41BF0 , 32'hF02FAF40 , 32'h024A6474 , 32'hFE41D0F4 , 32'h07D58420 , 32'hFE9F536C , 32'h014203AC , 32'h03620DD8 , 32'hFF8D24A7 , 32'h0AAC10F0 , 32'hFC860B1C , 32'h017EC70C , 32'h04064750 , 32'hFE3F4828 , 32'h001D5577 , 32'hFF8C4FA1 , 32'h02F74DE0 , 32'h03B56540 , 32'hFFDAFF04 , 32'hFD5B72C0 , 32'h01E0A518 , 32'hFB59EA08 , 32'hFF4C7CD6 , 32'hFD10BAA8 , 32'hFC7985A0 , 32'h00E1CCD0 , 32'h000339EB , 32'hFFFFA0C8 , 32'hFFFE534D , 32'hFFFF7F71 , 32'hFFFFB968 , 32'hFFFEBCE5 , 32'hFFFF62EC , 32'h000215BE , 32'hFFFEF5EF , 32'h00000BEF} , 
{32'h133E05E0 , 32'hFD104B48 , 32'h342552C0 , 32'h15657680 , 32'h1296F080 , 32'h18F15520 , 32'h08936420 , 32'hFEDB0F94 , 32'h1A3990E0 , 32'h0720BD20 , 32'hED4D9760 , 32'hF1AB0BE0 , 32'hE1045C40 , 32'hDAF41BC0 , 32'hF7D2FCA0 , 32'h0314A4F0 , 32'hE36153E0 , 32'h055EDB28 , 32'h11DD5300 , 32'h0B9A8AD0 , 32'h16A3F4E0 , 32'hE90F9780 , 32'h10F4D5A0 , 32'hFE9EA4FC , 32'hFDDAA104 , 32'h09CFC4C0 , 32'h1179E7C0 , 32'hF8CECC18 , 32'h022A5FE4 , 32'h02A26934 , 32'hF3376430 , 32'hFCF0CF00 , 32'h0D5E9590 , 32'h0BC449C0 , 32'hF254FE50 , 32'h00A95699 , 32'hF56CE430 , 32'h01C921F8 , 32'hF8A07268 , 32'hFB58D630 , 32'h007D968C , 32'hFE8B1AC0 , 32'hF46B41E0 , 32'h0543EE38 , 32'h034D3C74 , 32'h043269D8 , 32'hF2AA7DE0 , 32'hF36FD9D0 , 32'h08AF9D60 , 32'hF9C93C58 , 32'hF98DBD68 , 32'hF5964A90 , 32'hFBE49630 , 32'h02DB90A8 , 32'hFE0C7498 , 32'h00937127 , 32'hF9770D88 , 32'h0F13C250 , 32'hF9E8D368 , 32'hFACFFF08 , 32'h0BCE4F00 , 32'h024F8160 , 32'h02B5C918 , 32'h02645598 , 32'hFD6CD818 , 32'hFD88F634 , 32'hF45B6B90 , 32'h045DDDF0 , 32'hF5F1CFB0 , 32'hFB24FB20 , 32'hFF19EDB6 , 32'h02E69064 , 32'hFDF3E018 , 32'hF3D266B0 , 32'hFED0B9B0 , 32'hFE46B120 , 32'hFD9D0800 , 32'hFB867820 , 32'h0375CC9C , 32'h001411DD , 32'hFFD446E3 , 32'h00B988E2 , 32'hFD65DAA4 , 32'h00B49242 , 32'h015CA3AC , 32'h002DA32E , 32'h00444F15 , 32'hFEB69FC8 , 32'h005EE015 , 32'hFFFABA54 , 32'h0000B376 , 32'h00005ECF , 32'hFFFD8D8F , 32'h000225CC , 32'hFFFD43C0 , 32'hFFFEE8A0 , 32'h0000C775 , 32'h0001F662 , 32'hFFFFBE75 , 32'h0000CE86} , 
{32'h000058BB , 32'h000592CF , 32'h000125A4 , 32'h000268AD , 32'hFFFF08D0 , 32'h0000D27B , 32'hFFFF91FF , 32'h0003BBB4 , 32'h0000E41A , 32'h0003A9B5 , 32'h00011D84 , 32'hFFFD055E , 32'h0003D5C5 , 32'hFFF8D352 , 32'hFFFD0802 , 32'h00028237 , 32'h0001167C , 32'h0002CE43 , 32'hFFFDE538 , 32'hFFFE88CA , 32'h0001326D , 32'hFFFE44CA , 32'h00027260 , 32'hFFFF9A8A , 32'h00011E74 , 32'h00018A1F , 32'h0002D191 , 32'hFFFDC2BC , 32'h000093CF , 32'hFFFC72BB , 32'hFFFC81CB , 32'hFFFF44E7 , 32'h00002BF7 , 32'h0002FB8A , 32'h00036947 , 32'hFFFBE399 , 32'hFFFDBFF9 , 32'hFFFEBAB7 , 32'hFFFC9F22 , 32'hFFFC7C28 , 32'h000132AB , 32'hFFFE5E19 , 32'h0001CB25 , 32'hFFFCEC17 , 32'h0003544E , 32'hFFFD4392 , 32'h00026AB8 , 32'hFFFB459A , 32'h00007F4D , 32'hFFFE3B4C , 32'h00024544 , 32'h0002FE17 , 32'hFFFF8957 , 32'h0000C106 , 32'h00010EA4 , 32'hFFFFB538 , 32'hFFFBA31B , 32'h000061FE , 32'h00031B70 , 32'h00024D78 , 32'hFFFF93C1 , 32'h000163CF , 32'h00032DBE , 32'h000191F6 , 32'hFFFE9528 , 32'hFFFC0B1A , 32'h00000CC2 , 32'h00022BD7 , 32'h0002CB3C , 32'h00013203 , 32'h0001CA6F , 32'h00046571 , 32'h00012D58 , 32'h00056C04 , 32'h000352BC , 32'h0000E9FE , 32'hFFFDB608 , 32'hFFFA94EE , 32'h00001313 , 32'hFFF8EA03 , 32'h00002ADF , 32'hFFFF88A9 , 32'hFFFED195 , 32'h00007446 , 32'hFFFEF98F , 32'h0003420F , 32'hFFFF6810 , 32'hFFFE6AD8 , 32'h000106AC , 32'hFFFFC8AA , 32'h000464F5 , 32'hFFFDF59F , 32'hFFFFC6B7 , 32'hFFFEDB23 , 32'h00028CD3 , 32'hFFFBF313 , 32'hFFFFF4F8 , 32'h00036513 , 32'hFFFE3975 , 32'hFFFE5ECB} , 
{32'h0000BA51 , 32'h0000AC58 , 32'h0003FAE5 , 32'h00011A2D , 32'h0005432D , 32'hFFFE673F , 32'hFFFFD290 , 32'h00004A39 , 32'h00005094 , 32'h00026ADB , 32'h000341B0 , 32'hFFFCCBBC , 32'hFFFFDD8D , 32'hFFFD10AF , 32'h0000C1C9 , 32'h00032CDF , 32'h000283D1 , 32'hFFFFA50C , 32'h000188A2 , 32'hFFFE2162 , 32'hFFFE9C05 , 32'h00055ACF , 32'hFFFB9431 , 32'h0000229E , 32'h0000E84A , 32'h0000BB45 , 32'hFFFBBA00 , 32'h0001255F , 32'h0000DADE , 32'h0003363F , 32'h00005065 , 32'hFFFE75DC , 32'h0001CDA1 , 32'hFFFF6051 , 32'hFFFFCEB1 , 32'hFFFAF153 , 32'hFFFDCC5F , 32'h0004FE81 , 32'h00003848 , 32'hFFFEBBE6 , 32'h0002E74E , 32'h0000E72E , 32'hFFFE3732 , 32'h0001CE9B , 32'hFFFABD81 , 32'hFFFE03CA , 32'h000317F4 , 32'h00015B49 , 32'h00024FC4 , 32'h00036EFD , 32'hFFFE2E64 , 32'h0000CA25 , 32'hFFFAEBE6 , 32'h00026B3D , 32'hFFFF75A0 , 32'hFFFFC155 , 32'h0002398A , 32'h000021AC , 32'h000287E4 , 32'h00020A3E , 32'hFFFCA2CA , 32'hFFFE98D0 , 32'hFFFFD228 , 32'h0001CED1 , 32'hFFFEB5EB , 32'h000078F0 , 32'h0001C7E3 , 32'h00035F4C , 32'h000100D3 , 32'h0004E07F , 32'h0001D3EA , 32'h000200EF , 32'hFFFEEB3D , 32'h0000E09E , 32'hFFFC4812 , 32'hFFFFD9BD , 32'h00021153 , 32'hFFFE235E , 32'h0001524D , 32'h0001A9F0 , 32'h00003A83 , 32'hFFFF93E1 , 32'h0003E1BD , 32'hFFFDF842 , 32'hFFFE58D1 , 32'h000194B3 , 32'hFFFFD5C4 , 32'h00035B0B , 32'hFFFD8275 , 32'hFFFF8114 , 32'hFFFE1C4C , 32'h0000DF9D , 32'h000218E9 , 32'h000051AD , 32'h00030421 , 32'hFFFCF999 , 32'h00028E94 , 32'hFFFCF746 , 32'hFFFEC74A , 32'h000439BE} , 
{32'h04917CA0 , 32'h00C58C55 , 32'h06980740 , 32'hF9381690 , 32'hF06EB840 , 32'hEED44300 , 32'hF0F287B0 , 32'hFE119E54 , 32'hF4631FE0 , 32'hFCA45700 , 32'h07FEC838 , 32'hF4846770 , 32'hE849F5C0 , 32'h07829948 , 32'hFA1CE1A0 , 32'hF6E9DA80 , 32'h0340F308 , 32'hFA715DC8 , 32'h034B5A30 , 32'hFF3CD746 , 32'h04651798 , 32'h07E8AEC8 , 32'h007C8ADA , 32'h02353C9C , 32'h045E4250 , 32'h078ADB58 , 32'hFC398AF4 , 32'h022BD128 , 32'hFD1FDD58 , 32'hFD06D99C , 32'hFB6BD2F8 , 32'h0635BE28 , 32'h04D7A5C0 , 32'hFD9A9314 , 32'hEFC4AE20 , 32'hFA858B58 , 32'hFD681FFC , 32'hFB513668 , 32'hF6044380 , 32'h031A4FD8 , 32'h01C57498 , 32'h06587B50 , 32'h0FF85350 , 32'h04FF3C90 , 32'hF5F95560 , 32'h0382397C , 32'hF62C7520 , 32'hFF923C06 , 32'hFD4E3B8C , 32'hFB93ADD0 , 32'h018D2504 , 32'hFEA29EF0 , 32'hFEDAAF34 , 32'h063AFCD8 , 32'hFC12A7D0 , 32'hF9E20810 , 32'hFFFD5CD0 , 32'h015C5870 , 32'hF6AA55F0 , 32'h06449700 , 32'hF8588FA0 , 32'h0425D7F0 , 32'h09F705F0 , 32'h0B073C50 , 32'h07BD5030 , 32'h038F6D50 , 32'h016381A4 , 32'hFFE377B7 , 32'h01888020 , 32'h04BF8D30 , 32'h022E002C , 32'hF9B1A558 , 32'hFA87E498 , 32'h00A289DD , 32'h02CE2280 , 32'h02F121F4 , 32'hF9EC56A8 , 32'hFCEDF23C , 32'hFF2D3FE6 , 32'hFFF9CC71 , 32'h01AB5D6C , 32'hFE28559C , 32'hFB3A0AC8 , 32'h02C7BF5C , 32'hFB6A94F0 , 32'hFF2F5756 , 32'hFF4BFEF9 , 32'h026FCE88 , 32'h00F8FD96 , 32'hFFFC43AC , 32'h000238FE , 32'h0001AB6B , 32'hFFFF94F1 , 32'hFFFF40BE , 32'h0000AAB3 , 32'hFFFFF4B5 , 32'hFFFF451A , 32'h000415BF , 32'h000148E9 , 32'hFFFF536C} , 
{32'hB4FECD00 , 32'hDCF3A600 , 32'hE42CC080 , 32'hF0FD1C00 , 32'h4076C700 , 32'h0847ABF0 , 32'hCA46DE80 , 32'h01A5DD7C , 32'h04B02878 , 32'hEC753080 , 32'h03FFFBBC , 32'h1A8838C0 , 32'hF4636FF0 , 32'h1929B040 , 32'h0C6A3820 , 32'h08A1E7B0 , 32'h1CE42760 , 32'h0E9A70E0 , 32'hFEDBE3A8 , 32'hFF97C858 , 32'h12A66D40 , 32'hF24A22A0 , 32'hF3FA18E0 , 32'h05EA6BD8 , 32'h03AFF8AC , 32'h0E27D3A0 , 32'h06F95748 , 32'h088CEAC0 , 32'h08CA8390 , 32'hFC680400 , 32'h180FA1E0 , 32'h0166D058 , 32'hF835D3E0 , 32'hF5CD51A0 , 32'h0B64B710 , 32'h06CB12E8 , 32'hFD6B7C68 , 32'hFA2F5048 , 32'hF555D470 , 32'hF594BCA0 , 32'hFF8EE021 , 32'hF58E1FF0 , 32'h085FE920 , 32'h0BB96570 , 32'hF9327460 , 32'hF98B5000 , 32'hFF609A5F , 32'h048D2618 , 32'h0261A9D8 , 32'hF1A998E0 , 32'hFE9E276C , 32'hFE0FB100 , 32'hF3F82F40 , 32'hFFF8ADD3 , 32'h00FDF677 , 32'h03F7F19C , 32'h00FDFB77 , 32'hFCE957BC , 32'hFE2F867C , 32'h042F5548 , 32'hF99C6798 , 32'hFB789CB8 , 32'h01BBC350 , 32'h00C38AD7 , 32'hFDD2BDF8 , 32'h004E7DB1 , 32'hFCEDB1C8 , 32'hFD4D40CC , 32'h033944C8 , 32'h0397C940 , 32'hFB7BC980 , 32'h040BCDB0 , 32'hFF62D76B , 32'hFFED75DA , 32'h0155EED0 , 32'h032BBDD0 , 32'h01A102B0 , 32'hF48DFCC0 , 32'hFE9449F0 , 32'h022FF594 , 32'h016EC2CC , 32'hFD0442E8 , 32'hFAB2FBB0 , 32'hFD434CC0 , 32'h0140083C , 32'hFE9C1134 , 32'h005483BE , 32'hFA7D56C0 , 32'hFF9817CE , 32'hFFAC1BCE , 32'hFFFD3C17 , 32'hFFFF1B21 , 32'hFFFFE745 , 32'h00024EF2 , 32'hFFFE968A , 32'hFFFF325B , 32'hFFFDA538 , 32'hFFFF7F94 , 32'hFFFF1C7B , 32'hFFFFF7E9} , 
{32'hDA426F40 , 32'h8127E980 , 32'h3FEC9F40 , 32'h26D93D40 , 32'hFBF85738 , 32'hF9F8B8C0 , 32'hFDB6520C , 32'hFB8E6FA0 , 32'hFEB41D58 , 32'h01244104 , 32'h076D5390 , 32'h2215DC40 , 32'h0AA7AA10 , 32'hEE28C720 , 32'hFE55C444 , 32'hF6E2CEE0 , 32'hF32D7F80 , 32'hEA8852E0 , 32'hF1BFD380 , 32'hF4CB9B50 , 32'h0DF974A0 , 32'h15B218E0 , 32'hF07088C0 , 32'h1EA32BC0 , 32'hF5E0D6F0 , 32'hF846E7A0 , 32'h06C1C978 , 32'h08E16710 , 32'hF4B09C70 , 32'h0D8F09A0 , 32'h144CC860 , 32'hF6D02A20 , 32'h0EC0E6D0 , 32'hE69B0700 , 32'h02C31EA4 , 32'hF2485640 , 32'h05ED97D8 , 32'hF64B61F0 , 32'h03A132E4 , 32'hF07B30A0 , 32'h0976F230 , 32'h04B52E60 , 32'hFE475ED0 , 32'hF40DF730 , 32'h0112F330 , 32'h00294EA5 , 32'h0147C6F4 , 32'h091D6560 , 32'hFF549F71 , 32'h0FB6AAA0 , 32'hFE9A4314 , 32'hFD911538 , 32'hFDF41074 , 32'h0768ED28 , 32'h032A0B04 , 32'hFC642CC4 , 32'hFE2A1F2C , 32'h04348300 , 32'h07757560 , 32'hFBB32AB8 , 32'hFF585988 , 32'hFE8B0440 , 32'h0280C088 , 32'hFA787D28 , 32'h049B48D0 , 32'hF646B820 , 32'hFE60AEB8 , 32'h00F5EC68 , 32'hF9C31490 , 32'hFE883DD4 , 32'h000ED460 , 32'hFF05B69B , 32'hFD72E380 , 32'hFEB615AC , 32'h059DC708 , 32'hFF49BBC9 , 32'hFF1E14B6 , 32'hFB00B208 , 32'h0043ED57 , 32'hFC80EEF4 , 32'hFF401077 , 32'hFF2B3D4B , 32'hFF5CA557 , 32'h03D5A9A0 , 32'hFECB0630 , 32'hFF19A944 , 32'hFF7C42CF , 32'hFF41138A , 32'h01D8DB80 , 32'h00D2FF5D , 32'h000018A0 , 32'hFFFBFE5F , 32'hFFFF43D7 , 32'h000201BB , 32'h000073BF , 32'h0001367C , 32'h0000C58C , 32'hFFFFB39D , 32'h0000A434 , 32'h0001ACF4} , 
{32'hE67F4E60 , 32'h21904540 , 32'h22969640 , 32'h29587280 , 32'h00160624 , 32'hE9505CC0 , 32'h083F93A0 , 32'hFA348A30 , 32'h050343D8 , 32'h11EB4700 , 32'h1EE5DF60 , 32'hFFEDF57A , 32'hFF6177AA , 32'hF46B2630 , 32'h154C7F40 , 32'h06CB9570 , 32'h029C2AC0 , 32'hF3A78210 , 32'hFB921788 , 32'hFFBBB924 , 32'hFAF02588 , 32'h0E5B2E30 , 32'h04B85F38 , 32'h02048FC0 , 32'h147CA1E0 , 32'h15C3FA40 , 32'hE9B383C0 , 32'h01C7F2D0 , 32'h0CBBEBB0 , 32'h0191B03C , 32'hFC1DE074 , 32'hF9FFA0F8 , 32'hF5A967D0 , 32'h0A80D890 , 32'h0D3315C0 , 32'hFF80B0E5 , 32'h03997270 , 32'hF8A4A980 , 32'h06A9A4A0 , 32'hF198F650 , 32'hFC998CD4 , 32'hF691B800 , 32'hFAB90140 , 32'hF7804EC0 , 32'hEF4835A0 , 32'hFE54E5E8 , 32'h0FA94400 , 32'hF946B8B8 , 32'h041E3EA8 , 32'hF2323780 , 32'hFF1172DD , 32'hFC3A17CC , 32'hF9015300 , 32'hF82C2700 , 32'h012E34C4 , 32'h06669AF0 , 32'h0B7581E0 , 32'hFE2A7BCC , 32'h09B87330 , 32'hFD52C640 , 32'hFBD90E10 , 32'h0C566180 , 32'hF9339768 , 32'h028F82E8 , 32'h0054B19C , 32'h0223C228 , 32'hFE57FFE0 , 32'hFD66E5B0 , 32'h06DD3FA8 , 32'h024DE054 , 32'h0094AB13 , 32'hFE6475D0 , 32'h01712AFC , 32'hF7512250 , 32'h07911028 , 32'hFD89F858 , 32'hFE4682CC , 32'h00C0D146 , 32'hFD830E00 , 32'hF71B3510 , 32'hFE8B9AD0 , 32'h01CDF9F4 , 32'hFDF1D940 , 32'hFEA5B580 , 32'hFF491644 , 32'hFF2A6C95 , 32'hFFE0E87E , 32'hFFB8464A , 32'hFEF3E3F0 , 32'hFF9D497C , 32'h0001E335 , 32'h0000FA0E , 32'hFFFF9212 , 32'h0000C72A , 32'h00004935 , 32'hFFFDB5DE , 32'h00019214 , 32'h000016E8 , 32'h00017C2D , 32'hFFFF409A} , 
{32'hFFFD6E10 , 32'h0001880C , 32'hFFFEF133 , 32'h00022624 , 32'hFFFB4391 , 32'h00005FAA , 32'hFFFAE3D3 , 32'h000037C9 , 32'hFFFEB2A7 , 32'hFFF98DC5 , 32'hFFFB8952 , 32'hFFF94AF2 , 32'h00032A87 , 32'h0005CBB9 , 32'hFFFD37F8 , 32'h0003AF63 , 32'h0001B514 , 32'h00026848 , 32'h000086FD , 32'h0004ACEB , 32'h00043FB8 , 32'hFFFEF891 , 32'hFFFA020A , 32'hFFFD6DC0 , 32'h0004936F , 32'hFFFE29D2 , 32'hFFFF6C80 , 32'hFFFFCE45 , 32'h0002BA38 , 32'h000762E2 , 32'h00001CAD , 32'hFFFE21B3 , 32'hFFFF8F01 , 32'h00059605 , 32'h000092DA , 32'h00010C50 , 32'h0002A8A9 , 32'h0002B056 , 32'h0005523B , 32'hFFF90071 , 32'hFFFC0687 , 32'hFFFF7740 , 32'h0004F743 , 32'hFFFF3B93 , 32'h0006114B , 32'hFFFCA479 , 32'h0000F9D4 , 32'hFFFEA205 , 32'hFFFD1E77 , 32'h0006E6FF , 32'h00021663 , 32'h00048F7B , 32'hFFFD555D , 32'h00037C0F , 32'h000087A5 , 32'h00036559 , 32'hFFFFDE8A , 32'hFFFD5273 , 32'h00006D0C , 32'hFFFD91F0 , 32'h000178AF , 32'h00005B3D , 32'h0000A738 , 32'h000185DC , 32'h000119B1 , 32'h0000B423 , 32'hFFFECF1F , 32'h000604B1 , 32'hFFFEA82F , 32'h000156D7 , 32'hFFF9C670 , 32'h0001C5C7 , 32'hFFFEE974 , 32'hFFFEDB75 , 32'hFFFCF8EF , 32'hFFFB54A5 , 32'hFFFAFB12 , 32'h0000E422 , 32'hFFFDA477 , 32'hFFFD659E , 32'h00000B1B , 32'h0005DE42 , 32'h00024090 , 32'hFFFDF298 , 32'hFFFC8D9C , 32'hFFFFD4FF , 32'hFFFD1AE5 , 32'hFFFEFCD0 , 32'h00046CDA , 32'h0000DCEB , 32'h0004F153 , 32'h000216C5 , 32'hFFFD9F7F , 32'hFFFFDCEC , 32'h0000CAFA , 32'h0000228D , 32'hFFFF2C36 , 32'h0003466B , 32'hFFFE3041 , 32'hFFFFFB7E} , 
{32'h1F3836E0 , 32'hECC95A40 , 32'h04C85D28 , 32'h0C119EB0 , 32'hF2EC1C50 , 32'h233E2940 , 32'hF3E8D0C0 , 32'hEB2B3580 , 32'hFB06B998 , 32'hE9FAB040 , 32'h0B4336C0 , 32'h069BCE00 , 32'h0630AFA8 , 32'h057FCDF8 , 32'h031197AC , 32'h050B2778 , 32'h09F34000 , 32'h04B6FF20 , 32'hFB438E50 , 32'h12B2E8E0 , 32'h084021A0 , 32'hFB7BE090 , 32'hFFBAE1F5 , 32'h05B445A8 , 32'h16FA1480 , 32'hF5E815E0 , 32'hECBDF3A0 , 32'hFA0E03F0 , 32'h0ACBD3F0 , 32'h0A246D50 , 32'hF75DB4B0 , 32'hFDFF1DC4 , 32'h075E3A40 , 32'h03E33DC8 , 32'h08CA1770 , 32'h0D30C1D0 , 32'hF9353D48 , 32'hF57564F0 , 32'hFD04E3A0 , 32'hF93235F8 , 32'h082C8360 , 32'h06EEAB28 , 32'hF5214380 , 32'hF8DDC508 , 32'h12A50560 , 32'hFB634DD0 , 32'hFBA4BEF0 , 32'h055BFB38 , 32'h02BF0F48 , 32'h025D569C , 32'hF7BC45F0 , 32'hFC54C17C , 32'h00B2E49F , 32'hEC1A8D60 , 32'h039D3268 , 32'h064467C0 , 32'hFC4AB840 , 32'hEF5F8D00 , 32'hFADF6CE8 , 32'h0C44A7D0 , 32'hFF1C38CF , 32'h00FC8A78 , 32'h08102540 , 32'h04E08B78 , 32'h049FE6C8 , 32'hFCA64E24 , 32'hF982E288 , 32'h0B005320 , 32'h075FB908 , 32'hFF77FD5F , 32'hFB105F20 , 32'hF94F6BF0 , 32'hFBB10E78 , 32'hFE0D9508 , 32'h0528DB48 , 32'hFBC9E290 , 32'h0142F528 , 32'h019B1CCC , 32'h06BF5850 , 32'hFED0B80C , 32'h039F4F6C , 32'hFFD80168 , 32'hFD71E5D8 , 32'hFF920412 , 32'hFF7BAA95 , 32'hFDC34378 , 32'h0139DC94 , 32'h005B528E , 32'h0079773D , 32'h002D9B80 , 32'hFFFE4D32 , 32'h000041F1 , 32'h00014AC5 , 32'h000189B4 , 32'h00024E0B , 32'h0000CE6D , 32'hFFFE9F0F , 32'h000006EF , 32'hFFFF783D , 32'hFFFF3993} , 
{32'hEA0BE9E0 , 32'h194B4E00 , 32'h3939F5C0 , 32'hF3111C40 , 32'h168F9CC0 , 32'hDDBDA0C0 , 32'hEB3FA600 , 32'h060CB1F8 , 32'h00F5DB58 , 32'hED2D3AE0 , 32'h142798C0 , 32'hF9650B08 , 32'h0611FA28 , 32'hEE74D4C0 , 32'h01572D20 , 32'hDDDEF580 , 32'hFBE06830 , 32'hEEE19320 , 32'h03E4FA30 , 32'hF7FA9800 , 32'h035D5E24 , 32'hEA4330A0 , 32'h030508B8 , 32'hF59FC9F0 , 32'h091E2F90 , 32'hF9983398 , 32'hFBB696F0 , 32'hE6F75900 , 32'h0035BBD2 , 32'hE0DC2AA0 , 32'hF22DE820 , 32'h06764FD8 , 32'h03111FD0 , 32'h01FDF140 , 32'h0F2DC680 , 32'hEB5AF7C0 , 32'h043BA4A8 , 32'h0ED94630 , 32'hFD0CABD8 , 32'h02CB1240 , 32'h00440AE9 , 32'hF5A6EC70 , 32'hFB59C130 , 32'hFFB1B6FC , 32'h03C3CA20 , 32'h0128DAF8 , 32'h0B716230 , 32'h05554E00 , 32'hF62C9C70 , 32'hFAFB6DE0 , 32'hFF50423A , 32'h0C0C9EB0 , 32'hFA37E608 , 32'hF662EA50 , 32'h0B55CC20 , 32'hF8ED5DE8 , 32'hFDED177C , 32'h000E655E , 32'hFDC0A05C , 32'hFA7A5410 , 32'hF346C080 , 32'h00837686 , 32'h06464BB8 , 32'hFB1EC960 , 32'h000A9140 , 32'hFFA08DCE , 32'hF76DB5A0 , 32'hFF4451A5 , 32'h0357A6B4 , 32'h0A2E6A60 , 32'h00E96B09 , 32'hFC119434 , 32'h03B10954 , 32'h03BCE49C , 32'h033BFD4C , 32'h04128E50 , 32'h04028680 , 32'h053A6018 , 32'h0306B36C , 32'h054B7AB0 , 32'h0190EBF0 , 32'hFE05AC1C , 32'hFC4A53E8 , 32'h009BA9EB , 32'hFCA2170C , 32'hFDC6C59C , 32'h035F0AD0 , 32'h016C87B0 , 32'h00561367 , 32'hFF8805C5 , 32'hFFFFC1CE , 32'h0000643B , 32'hFFFF28D7 , 32'h000021E9 , 32'hFFFD2008 , 32'h0001BB35 , 32'h0000903D , 32'hFFFE2E19 , 32'hFFFE8148 , 32'h00017CCD} , 
{32'h0183BAD8 , 32'hFF9B6427 , 32'hFE31DB24 , 32'h00DF8619 , 32'hFFB621CC , 32'hFE660270 , 32'hFD032EDC , 32'hFD48B7B0 , 32'hFE61BAEC , 32'h002BA310 , 32'h01D98C10 , 32'hFD529BF0 , 32'hFF4B2DD6 , 32'hFE1F6460 , 32'h0133E158 , 32'h0067993A , 32'hFE833288 , 32'h049CCCD8 , 32'hFFAE39FC , 32'hFE16DF00 , 32'h00CDC4A9 , 32'h03EB35E4 , 32'h0421C4C0 , 32'h00980BAB , 32'hFF870A1D , 32'hFE62E05C , 32'hFFE39D46 , 32'h00594AA5 , 32'hFCA61FDC , 32'hFCFB9B40 , 32'h04159EF0 , 32'hFFF82F2F , 32'h0110CA08 , 32'hFDB72A18 , 32'hFC4ECD6C , 32'h011E1E94 , 32'hFBD1F0D8 , 32'h0300E42C , 32'hFECB7094 , 32'hFD549074 , 32'h02C150B8 , 32'h040A5DE8 , 32'h05DA5798 , 32'hFEFF42F8 , 32'h0004F52B , 32'h016256F8 , 32'hFD24D1F8 , 32'h01DC8D30 , 32'h04EE8088 , 32'h00ACA44B , 32'h03679D4C , 32'hFF0F3322 , 32'hFFDAFB68 , 32'hFCB76F68 , 32'hF9653458 , 32'hFD59A444 , 32'h00AD17A1 , 32'hFC74FAD0 , 32'hFE468E78 , 32'hFDB9E7C0 , 32'h02229B60 , 32'hFC9363F0 , 32'h017DCCE0 , 32'h0279F0C0 , 32'h0177DC80 , 32'h01F0D930 , 32'hFDD14300 , 32'hFDA0EE90 , 32'hFF801AB2 , 32'h005E07E5 , 32'hFCF1D258 , 32'h00C69CB1 , 32'h02002564 , 32'hFDCEFF54 , 32'hFD4E7C50 , 32'h00881761 , 32'h0049D12D , 32'h0075A3EF , 32'h02042A94 , 32'h0006B3DE , 32'h01AAF6B4 , 32'hFFBE8234 , 32'h0064E010 , 32'h00AF6481 , 32'hFE2A8D44 , 32'hFFA6DE39 , 32'h0102024C , 32'hFE973550 , 32'h00AFE6F1 , 32'hFFF43BA0 , 32'hFFFBF5E9 , 32'h00000783 , 32'hFFFCD969 , 32'hFFFC8A7C , 32'h0000F519 , 32'h00027D74 , 32'hFFFDA922 , 32'hFFFE6B75 , 32'h00014B9C , 32'h000197ED} , 
{32'hFFFF2CCB , 32'hFFFDBFE9 , 32'hFFFD1ADD , 32'h000232D0 , 32'h00027DF1 , 32'hFFFD1586 , 32'hFFFEBBE7 , 32'hFFFCE87F , 32'h000068C6 , 32'h0001A0E2 , 32'hFFFFBAAB , 32'hFFFEE8A3 , 32'hFFFDF472 , 32'hFFFECFD3 , 32'hFFFEC3FF , 32'hFFFF4D67 , 32'h000507DD , 32'h00048634 , 32'h00016B59 , 32'hFFFD3A0B , 32'hFFF65489 , 32'h00008DDD , 32'hFFFE8502 , 32'h00005A9F , 32'hFFFFEF38 , 32'hFFFDC6CA , 32'h00005308 , 32'hFFFD9FEA , 32'hFFFE6464 , 32'h0001D6BF , 32'h0000BF75 , 32'hFFFE9494 , 32'h000594A6 , 32'h0002793A , 32'hFFFEE41A , 32'h0001E036 , 32'h00001FF7 , 32'hFFFF43BC , 32'hFFFD8E4C , 32'h0001DD87 , 32'h0002D032 , 32'h00032FCC , 32'h00045413 , 32'hFFFD8740 , 32'h00032202 , 32'hFFFBD97B , 32'hFFFEE513 , 32'hFFFD2F02 , 32'h00007EF8 , 32'h00029DEF , 32'h0001061B , 32'h00019B37 , 32'h00019D8D , 32'h00023FA6 , 32'hFFFD849E , 32'h0002470F , 32'h0000B93F , 32'hFFFFA07F , 32'hFFFE2961 , 32'hFFFF6EAC , 32'h0004DB84 , 32'h00027540 , 32'h0003DCDE , 32'hFFFFB78B , 32'h000210D7 , 32'h000049BF , 32'hFFFF9D3D , 32'hFFFB8314 , 32'h00034401 , 32'hFFFA57BE , 32'hFFFD2BAD , 32'h0001A9D0 , 32'hFFFE0ED8 , 32'hFFFF6501 , 32'hFFFA25ED , 32'hFFFCC6F7 , 32'hFFFF7FC8 , 32'h00035692 , 32'hFFFFADE0 , 32'hFFFF0A79 , 32'h0002285F , 32'h000194DE , 32'hFFFB2009 , 32'h000055FF , 32'hFFFC0378 , 32'h0003B9A4 , 32'h00002162 , 32'h00022D45 , 32'h0001259E , 32'hFFFC54E7 , 32'hFFFACF42 , 32'hFFFB7C72 , 32'hFFFDE771 , 32'hFFFF838D , 32'hFFFEBF97 , 32'h000064E1 , 32'hFFFE12E0 , 32'hFFFD5BCA , 32'hFFFBFBB1 , 32'h00038A6E} , 
{32'hF28F2420 , 32'hFB0BD4C0 , 32'hF30AE590 , 32'h1172DD60 , 32'hFB3BD738 , 32'h0FAAEAA0 , 32'hF7BCDB00 , 32'h072C7DA0 , 32'h05292FD0 , 32'hFE5030DC , 32'hF11D5530 , 32'hF739D140 , 32'h00646B9E , 32'hFB7E6428 , 32'h0592C148 , 32'hF874FFC0 , 32'h0AEDBD50 , 32'hFB2A6FA0 , 32'hFF2A578D , 32'h02DC8C70 , 32'h0435F278 , 32'h01A1A9C0 , 32'h05789BC8 , 32'hFB553378 , 32'h09049140 , 32'h0A830040 , 32'hF60C37C0 , 32'h0DED3950 , 32'hF8226730 , 32'hF4D36850 , 32'h0947DE00 , 32'h089F5580 , 32'h0311A278 , 32'h0884A820 , 32'h023FB2CC , 32'h0491EAD8 , 32'hFFCDA206 , 32'hFAC74150 , 32'hFC30ACA4 , 32'h0C9915E0 , 32'hF9E2FC00 , 32'h0071362E , 32'hFC393404 , 32'h028E73F8 , 32'hF59757E0 , 32'h04E2B538 , 32'h040B7260 , 32'hFDA88B3C , 32'hF8236AE0 , 32'h07503440 , 32'h0C015620 , 32'hFE5934C8 , 32'hFD1B4AF8 , 32'hFE1E1148 , 32'hFF8A1CA1 , 32'hF6750360 , 32'hF77F2650 , 32'hF7DB12D0 , 32'hF7EB3610 , 32'h067FCE10 , 32'h023A03B4 , 32'hFC48A6C0 , 32'h004A904C , 32'hFA50EA98 , 32'hFE295554 , 32'h0393260C , 32'hFE37E14C , 32'h01C65CDC , 32'hF862DFA0 , 32'h00B41AAF , 32'hFF15F8BC , 32'h02DCEF1C , 32'hFD0E893C , 32'hF9E91B50 , 32'h03D5AAB4 , 32'hFF2318C7 , 32'h02C71DA4 , 32'h018347D8 , 32'hF6B6AFE0 , 32'h0063663D , 32'hFE2413A0 , 32'h02530704 , 32'h037DF350 , 32'h00C344D1 , 32'hFF4D5D83 , 32'hFC8F9E74 , 32'h03E6C12C , 32'h01180A20 , 32'hFE8B86C8 , 32'hFFD09E78 , 32'hFFFEA985 , 32'h00023215 , 32'hFFFED30E , 32'h00023A15 , 32'hFFFF8337 , 32'hFFFFA20E , 32'h00016F10 , 32'h00000161 , 32'h00015254 , 32'hFFFE8A86} , 
{32'h0BBBAA80 , 32'h00607016 , 32'h227D6380 , 32'hFA0F9430 , 32'h140CE180 , 32'h175CC220 , 32'hE2E141A0 , 32'hECC8CEE0 , 32'hF1C1C1D0 , 32'hF92613C0 , 32'hF4E991D0 , 32'hF54F33A0 , 32'hF865E890 , 32'hEA35BBA0 , 32'hFAEE7ED8 , 32'h01799138 , 32'h040DEC08 , 32'h10694DE0 , 32'h05DBB070 , 32'hF6DFB030 , 32'hF7109200 , 32'hF6C484E0 , 32'h03026F2C , 32'h0600DE10 , 32'hF89A7D90 , 32'h01E43BA0 , 32'hF3D48850 , 32'h11B63760 , 32'h1CE94BE0 , 32'hFF6BA718 , 32'hF6BCF390 , 32'h01507F94 , 32'hFF074EC7 , 32'hFA43E448 , 32'hFC94E2FC , 32'hE8D0F340 , 32'h195A6580 , 32'hEA5DA580 , 32'h03620E8C , 32'h0AAC0230 , 32'h091D8530 , 32'h0FBC8520 , 32'h030B7284 , 32'hFE99D62C , 32'h05A12678 , 32'h0A7876B0 , 32'hFD6A053C , 32'h0127BCF4 , 32'h07168028 , 32'h062CEFE8 , 32'h016EB430 , 32'h14BEB680 , 32'h086A01A0 , 32'hF42FC940 , 32'h06637B48 , 32'h0813BF50 , 32'h006157FD , 32'h048DC710 , 32'h06C5A1B0 , 32'hF50A0BF0 , 32'hFB3AB4E0 , 32'h023164BC , 32'h02F7B44C , 32'h01755DD0 , 32'hFD5662E0 , 32'hFEB9ACC4 , 32'hFE7BD3E0 , 32'hF9CD5E20 , 32'h023C176C , 32'hF4148B40 , 32'h014AA914 , 32'h033210E4 , 32'hFF0144A3 , 32'hFC7A0044 , 32'hFA7488A8 , 32'h011F99E8 , 32'hF90B6C50 , 32'hFB60D810 , 32'hFBA7C400 , 32'h04FF1A60 , 32'h01B580FC , 32'h00B12D38 , 32'hFCE0A50C , 32'hFAB9E4A0 , 32'h053C2CB8 , 32'hFFDD9345 , 32'hFF46E687 , 32'hFED528D4 , 32'hFFC2AC14 , 32'hFF836B7B , 32'h00010269 , 32'h0000CF34 , 32'h0001F6E9 , 32'hFFFE84E9 , 32'h00014E66 , 32'h00021610 , 32'h0000A02F , 32'hFFFE6EF9 , 32'hFFFF126D , 32'hFFFE64C6} , 
{32'hFB1F59A0 , 32'hF7CED1B0 , 32'hE4E5D940 , 32'h1C6B3F40 , 32'hEFFD7A20 , 32'h156230C0 , 32'hE706A260 , 32'h078FDAF0 , 32'hE669E660 , 32'h041B62E8 , 32'h00BA273D , 32'hE8A833A0 , 32'h23809400 , 32'h072F0830 , 32'h06530BE0 , 32'h060FD230 , 32'hF5DF5170 , 32'hF32D5FD0 , 32'hFB9A7C88 , 32'hFF7B4359 , 32'hF9E15E40 , 32'h025134C4 , 32'h01FB7FCC , 32'hF61BFDE0 , 32'h02BAEED0 , 32'h12E0EA60 , 32'h02E64364 , 32'h0DD9EC10 , 32'hF10A1280 , 32'hFCB5CC98 , 32'hFE1EFD84 , 32'hF2BC8B20 , 32'h05BE2D38 , 32'hFFD66E42 , 32'hF5009DC0 , 32'h009EFADF , 32'h05FE4F70 , 32'h00BF057A , 32'hFF69D0BB , 32'hFBBBBB40 , 32'hF3AF72C0 , 32'hF7776C40 , 32'hFFCB8307 , 32'h025FE874 , 32'hFFDE2253 , 32'hF9F9B800 , 32'hFCCA75F4 , 32'hEE417640 , 32'hE8C01420 , 32'h04A30D68 , 32'hF88C6E38 , 32'h0CB52D10 , 32'h00156B42 , 32'hFB368478 , 32'h01B6C000 , 32'h00237572 , 32'hFF4DEF1C , 32'hFEB2CFF8 , 32'h00DE959E , 32'h02CBA1C8 , 32'h0120AFA0 , 32'hFE7A6C58 , 32'h05A56820 , 32'h09C09800 , 32'hFB4DB9E0 , 32'h03B09FC0 , 32'h04130F78 , 32'hFFE1815D , 32'hFD38E678 , 32'h03CA12B8 , 32'hFA187AC8 , 32'h095F38E0 , 32'hFDDA402C , 32'h04BE4220 , 32'hFEFCA254 , 32'hFD2D9780 , 32'h03FA3A8C , 32'hFCEE9CB0 , 32'h0411DD58 , 32'hFDD8B19C , 32'h00BFC9E5 , 32'hFF61D889 , 32'hFB46EC98 , 32'hFF7BB426 , 32'h01E13FDC , 32'h03AAE170 , 32'hFC138458 , 32'hFEC1AB8C , 32'hFF7493B8 , 32'hFF5BEEE9 , 32'hFFFF6203 , 32'hFFFEE54E , 32'hFFFDCAB6 , 32'h000150A7 , 32'hFFFDB8AC , 32'hFFFF82F4 , 32'hFFFF5A03 , 32'hFFFC2D51 , 32'hFFFFFB94 , 32'h00010D8E} , 
{32'hFFFBE665 , 32'hFFFE5099 , 32'hFFFB8596 , 32'h00027B18 , 32'hFFFE8764 , 32'hFFFBD8ED , 32'h0000F591 , 32'hFFFFB578 , 32'hFFFA4524 , 32'h00033D15 , 32'h00034345 , 32'h00014C50 , 32'h0001DFDA , 32'hFFFFC9C2 , 32'h000286AB , 32'hFFFDD66B , 32'hFFFA303E , 32'hFFFF6FCB , 32'hFFF9CAD1 , 32'hFFFC06B2 , 32'h000135DB , 32'hFFFF1F92 , 32'hFFFF6753 , 32'h000077DF , 32'h00007FE8 , 32'hFFFEA08C , 32'h0002517E , 32'h0000E687 , 32'hFFFFC63E , 32'hFFFF31F6 , 32'hFFF9AAA7 , 32'hFFFF7765 , 32'hFFFDE9F0 , 32'hFFF9EDDD , 32'h0003E203 , 32'h00035710 , 32'hFFFDABD9 , 32'h000072EA , 32'h0005A05D , 32'h000402EC , 32'h0005F944 , 32'h0001B0EF , 32'h00019926 , 32'hFFFFB473 , 32'hFFFD2BB5 , 32'hFFFF048A , 32'h00006339 , 32'hFFFE199A , 32'h000311F0 , 32'h00013319 , 32'h0001C8DF , 32'h0000F7E4 , 32'hFFFEE842 , 32'hFFFFFCEB , 32'hFFFE78A4 , 32'hFFFBC8D7 , 32'h00026506 , 32'hFFFDBE12 , 32'hFFFB4951 , 32'h000207C3 , 32'h0002F1A5 , 32'hFFFAC708 , 32'h0000B3DD , 32'h000161F1 , 32'h0000665C , 32'hFFFC89A0 , 32'h0004D341 , 32'h0002770D , 32'h0001C115 , 32'hFFFE5682 , 32'h00004986 , 32'h00055318 , 32'hFFFEA93A , 32'h000430CC , 32'h000308AB , 32'hFFFCFC33 , 32'hFFFF7EBE , 32'hFFFCF926 , 32'h000147C8 , 32'h0001FE29 , 32'h00034818 , 32'h000359C0 , 32'h0003B0E5 , 32'hFFFD1D81 , 32'hFFFD116B , 32'hFFFCBFC3 , 32'hFFFCAB0E , 32'hFFFB8C5F , 32'hFFFE02F4 , 32'h0000585E , 32'hFFFD31F8 , 32'h00005856 , 32'hFFFECEBA , 32'h00023ABC , 32'hFFFF5557 , 32'hFFFB6AC6 , 32'hFFFFACDD , 32'hFFFF36EE , 32'h0001C59D , 32'hFFF98D1F} , 
{32'h07434910 , 32'h05DB6068 , 32'h065FF440 , 32'hFA140160 , 32'hECCF2240 , 32'hFE1B7040 , 32'hF0C478C0 , 32'hFCCBED44 , 32'hFBE378B8 , 32'h01FEDFDC , 32'hFE657504 , 32'h07D34498 , 32'hF793F750 , 32'h07133528 , 32'h09724010 , 32'h0ABC1880 , 32'hFB621258 , 32'h089D6C50 , 32'hF92C81F0 , 32'h0442F100 , 32'hFC06BC80 , 32'hF6D508A0 , 32'hF709AF30 , 32'h0ACB8260 , 32'h03BDC194 , 32'hF68646F0 , 32'hF2459220 , 32'h0035E0B8 , 32'hF8F6A1E0 , 32'hFC86108C , 32'h067C6790 , 32'hFEC84534 , 32'hF66E7F40 , 32'h022A1714 , 32'hFEB02694 , 32'hFEE38AFC , 32'hF9211098 , 32'h03D34F04 , 32'h083323E0 , 32'h020A9558 , 32'hFCBD3AEC , 32'h010F8A88 , 32'hFA591750 , 32'h00669B5C , 32'h035CC8B4 , 32'hFE68A59C , 32'h112351C0 , 32'hF5026240 , 32'hFCA9F57C , 32'h0B62D870 , 32'hFF20F4F6 , 32'hFFDEC4C0 , 32'hFC389E28 , 32'h0136EC64 , 32'h0919A7F0 , 32'hF66DB5A0 , 32'hFAF0B950 , 32'h060EF3F0 , 32'h015E8F0C , 32'hF5135660 , 32'h0C9C3D00 , 32'hFFF0849C , 32'hFE40940C , 32'h01A09A48 , 32'h07B91850 , 32'h05DB17A0 , 32'hF8DA2E10 , 32'hF9141B10 , 32'hFD51D628 , 32'hFC0465C4 , 32'hFF98D562 , 32'h00315C9A , 32'hF7DDC220 , 32'h06FF8A78 , 32'h017D131C , 32'h025AD1D8 , 32'h01A20AA4 , 32'h06D39580 , 32'hF9434880 , 32'h018C61C4 , 32'h07A60860 , 32'h00087DD2 , 32'h01D7B058 , 32'hFF045557 , 32'h00BA6579 , 32'hFE82B808 , 32'hFBCC2930 , 32'hFF4FB6BC , 32'h0167AF00 , 32'hFFC7149B , 32'hFFFF4361 , 32'h00003945 , 32'hFFFE5AF4 , 32'h000032DE , 32'h0000E77C , 32'hFFFF1256 , 32'h00002625 , 32'h00006B1E , 32'hFFFF32C9 , 32'hFFFF24EA} , 
{32'hFFFEC829 , 32'hFFFF2A33 , 32'h0001E6D3 , 32'hFFFFCADA , 32'h0003E98F , 32'hFFFE8E85 , 32'hFFFFADE7 , 32'hFFFF1AE2 , 32'hFFFFFF7A , 32'hFFFF884E , 32'h0001F43B , 32'hFFFA50CD , 32'hFFFD9962 , 32'hFFFFA1E4 , 32'hFFFCB4B0 , 32'hFFFB41BA , 32'h00018503 , 32'h00006388 , 32'hFFFA01E3 , 32'hFFFF367F , 32'h0000DAB0 , 32'h00019476 , 32'hFFFD733C , 32'h0003D587 , 32'h00058BB7 , 32'h00045D90 , 32'hFFFE36F0 , 32'h00017BEF , 32'h00040F3B , 32'h000273BF , 32'hFFFDD2F9 , 32'h00043311 , 32'h0002C4B9 , 32'hFFFD0BBE , 32'h0006EA6B , 32'hFFFEC402 , 32'h0000F9EB , 32'h000287C1 , 32'h000246F9 , 32'h0001FA1B , 32'h000145FF , 32'h00045CF6 , 32'h00056F76 , 32'hFFFFDA3A , 32'hFFFECE4F , 32'hFFFB230E , 32'h0002782A , 32'h000065A1 , 32'hFFFF3897 , 32'hFFFDAE72 , 32'h0000BF60 , 32'h000126EA , 32'hFFFC8E12 , 32'h00011C88 , 32'h0001F87E , 32'hFFFFE88F , 32'hFFFEA824 , 32'h00016546 , 32'h000360AF , 32'h0004B928 , 32'h00016E7C , 32'hFFFE8A2E , 32'hFFFDB5AF , 32'h0001B1DA , 32'hFFFC7574 , 32'h0002C68C , 32'hFFFE8D02 , 32'h000183C4 , 32'h0000FB42 , 32'hFFFD9E4D , 32'hFFFFDE1A , 32'hFFFDA336 , 32'h0003A3A9 , 32'hFFFEFBA0 , 32'hFFFF1F7E , 32'h0000C48E , 32'h000339AF , 32'hFFFCF2A0 , 32'hFFFCAD37 , 32'h00041270 , 32'h0002D763 , 32'hFFFE0D79 , 32'hFFFD5943 , 32'hFFFFAACE , 32'h00044153 , 32'h000088D6 , 32'hFFFDACDE , 32'hFFFF70DB , 32'hFFFD4487 , 32'h000204F0 , 32'h0001B75C , 32'hFFFC218F , 32'hFFFF4584 , 32'hFFFF1B9F , 32'hFFF9CA3A , 32'hFFFFEDB9 , 32'hFFFE93DC , 32'h00008FC7 , 32'hFFFEFFF2 , 32'h0003E521} , 
{32'h00006F2C , 32'hFFFDD25E , 32'h0000727F , 32'h00054FFD , 32'hFFFCF09C , 32'h00023357 , 32'hFFFDD9F9 , 32'hFFFDB5B7 , 32'hFFFDEA15 , 32'h00000DC3 , 32'h00011631 , 32'hFFF9CCCF , 32'hFFFE9290 , 32'h00009E99 , 32'h000490B4 , 32'h0000A891 , 32'hFFFF0C80 , 32'hFFFE82AE , 32'hFFFCAEFC , 32'hFFFF974D , 32'h00026847 , 32'hFFFF723C , 32'h0000D977 , 32'h00002BF5 , 32'h0000D2CF , 32'h0000F551 , 32'h000459EE , 32'h0002212A , 32'hFFFCE432 , 32'h0004F5AF , 32'h0001B84D , 32'hFFFE2479 , 32'hFFFD9812 , 32'h0000610E , 32'h0000D9A8 , 32'h0006BD26 , 32'hFFFE2B33 , 32'hFFFE7266 , 32'hFFFDEEF2 , 32'hFFFF4D38 , 32'hFFFCFAEA , 32'hFFFCE41E , 32'h00045402 , 32'h00028C49 , 32'hFFFC9455 , 32'hFFFE6789 , 32'h00000C94 , 32'hFFFD05D4 , 32'hFFFEFBC7 , 32'hFFFE0224 , 32'hFFF98BCE , 32'hFFFE7156 , 32'h00086336 , 32'h0001219A , 32'hFFF9DDC0 , 32'h0006A872 , 32'hFFFE3CF3 , 32'h0003F3D7 , 32'h00015CDB , 32'hFFFFC96A , 32'h000370DD , 32'h0000B8FC , 32'hFFFF483E , 32'h00039FC7 , 32'hFFFDAB3A , 32'hFFFF91F0 , 32'hFFFFAF2E , 32'h0002EB54 , 32'h0000DA4D , 32'hFFFE37F4 , 32'hFFFFBB1B , 32'h0000EEB7 , 32'h0000EDC6 , 32'hFFFD2904 , 32'hFFFFAE30 , 32'hFFFADAC7 , 32'h0001E2B0 , 32'h00007E16 , 32'hFFFE6194 , 32'hFFF86DE4 , 32'h00022A96 , 32'h0003B4DB , 32'h0002DE39 , 32'h00006E3C , 32'h000008E1 , 32'h00003D3F , 32'hFFFFF9FF , 32'hFFFC7116 , 32'hFFFFC918 , 32'h00032F03 , 32'hFFFFE76A , 32'hFFFE16F7 , 32'hFFFFEDBD , 32'h000321F9 , 32'h00007862 , 32'hFFFC1151 , 32'hFFFF9C9F , 32'hFFFEE8C6 , 32'h00021138 , 32'hFFFF1A1A} , 
{32'h069F18C0 , 32'hF4464F00 , 32'hFCA1D4D0 , 32'h16C52BA0 , 32'hF47ABDB0 , 32'hFCEBF18C , 32'hFF59C90D , 32'h0BC94F20 , 32'hEFE66040 , 32'h09FFBA40 , 32'h01BA16E0 , 32'h0292A52C , 32'h07FA8408 , 32'h0CAA96B0 , 32'hFA394BB0 , 32'hFD18EB20 , 32'h02375074 , 32'h0352F3F8 , 32'h0A766530 , 32'h04288930 , 32'hFD7798A0 , 32'h00A96D1C , 32'hECA321A0 , 32'hF742D6E0 , 32'hF90EB6D0 , 32'hF4EB7D30 , 32'h065B07C0 , 32'hF7CE0350 , 32'hEEF000A0 , 32'h0347CFF8 , 32'hF65067E0 , 32'h02EF3A4C , 32'hFD1AEBF8 , 32'h02A74AE4 , 32'hF82AB1D0 , 32'hFEEB0EF4 , 32'hFCE1EDBC , 32'hF6386030 , 32'hFFFA93CC , 32'hFF6FE839 , 32'h023A8A70 , 32'h047C0CA0 , 32'h05ACDAF0 , 32'hF9953A08 , 32'hFE9FA0F4 , 32'h01A98B34 , 32'hFD4ABA14 , 32'h0114F10C , 32'h01EA5A34 , 32'hF2A0CCC0 , 32'hFB0BED20 , 32'hFABBD540 , 32'hFDB0F054 , 32'h03889B30 , 32'hFC5B27E0 , 32'hF26EEFF0 , 32'hF8443210 , 32'h03EFFE58 , 32'hFB3CA6E0 , 32'hFC0FA018 , 32'hF46A0DD0 , 32'hF61CAFF0 , 32'hFD7B70AC , 32'hF657F600 , 32'hFA395330 , 32'hFDBF2FF8 , 32'h053EA618 , 32'hFC05D040 , 32'h054CE210 , 32'hFC5F5868 , 32'h02975F28 , 32'hFD9A3134 , 32'hFD35B6A8 , 32'h00E09425 , 32'h008798BA , 32'h0324AEC8 , 32'h005104FE , 32'h024EFFCC , 32'hFDE34C08 , 32'hFC82F44C , 32'hFFFCFD05 , 32'h0274E9A8 , 32'hFE2AB134 , 32'hF89901B0 , 32'h034D1320 , 32'hFF3EB843 , 32'h01C96C74 , 32'h0149A04C , 32'h038F600C , 32'hFFDE80A7 , 32'h0005CCA1 , 32'h0002BEC3 , 32'h0000C5B5 , 32'hFFFFB4F3 , 32'hFFFDC990 , 32'h00048626 , 32'h00002841 , 32'hFFFF0095 , 32'hFFFE1245 , 32'hFFFF3143} , 
{32'h01CD6868 , 32'hFD3249F0 , 32'hFB3CD588 , 32'hF5329810 , 32'hFF4B1EF4 , 32'h010289EC , 32'h01620598 , 32'hFEA9DC3C , 32'hFA544488 , 32'h0078355B , 32'hFA7221B0 , 32'h054C7258 , 32'h054CAE70 , 32'hFCF4E30C , 32'hFF023057 , 32'hFEA49B10 , 32'hFDFE41DC , 32'h0312E3BC , 32'hFCD77CA4 , 32'h05743C48 , 32'h011CEE34 , 32'h0115A54C , 32'h01CA9270 , 32'h0066EBA0 , 32'hFEF13AFC , 32'hFCC05F44 , 32'hF8150A80 , 32'h02B7859C , 32'hF9C0E3C0 , 32'h053C14A0 , 32'h025D0F24 , 32'hFD5295D8 , 32'hFE16D8AC , 32'hFDE58164 , 32'hFD3E5A28 , 32'h03E16610 , 32'h045CD270 , 32'h0072E837 , 32'h03F24374 , 32'hFB8B6638 , 32'hFFE1B195 , 32'hFDB76564 , 32'h07DB56C0 , 32'h0130FDE0 , 32'h00A8D812 , 32'hFF33E46A , 32'hF9FA5980 , 32'h037E5070 , 32'h0713CE70 , 32'h0054A554 , 32'h09DACA00 , 32'h01925198 , 32'h01B5B698 , 32'h04DE6080 , 32'hFC31CE2C , 32'hFD50DFD8 , 32'hFD5D65B4 , 32'h01755420 , 32'h03E8DFA0 , 32'hFE62C120 , 32'hFE844658 , 32'hFE8C5D70 , 32'hFAE28248 , 32'h0562C0A0 , 32'hFCE20120 , 32'h05B7D0A0 , 32'hFE908DB8 , 32'h01E70B4C , 32'h02741834 , 32'hFBBB72D0 , 32'h04BE5358 , 32'hFA8AAB20 , 32'h037F269C , 32'hFBB92798 , 32'h027D474C , 32'hFFBDB1AF , 32'h013237C4 , 32'hFF4B082D , 32'h013D6A04 , 32'h02DBF2EC , 32'hFC9F0B58 , 32'hFD420598 , 32'hFC6F1074 , 32'h0034AC54 , 32'h02B7C9E8 , 32'h00872031 , 32'h01633634 , 32'hFB766620 , 32'hFCD35C3C , 32'h0000E187 , 32'h0002774E , 32'h000104BD , 32'hFFFC5BA5 , 32'hFFFFFF59 , 32'hFFFF3B75 , 32'hFFFDB528 , 32'h00038254 , 32'h0000B486 , 32'h00019B3A , 32'h00034853} , 
{32'hFE4AE920 , 32'hFF98C92A , 32'hF83FE230 , 32'h0B5D0160 , 32'h012B95F8 , 32'h1FCA2EC0 , 32'hF9ACC488 , 32'hFE33BE78 , 32'hF78841E0 , 32'h010F9A38 , 32'h01FA1A00 , 32'h0EE42250 , 32'h05C9A5B8 , 32'hFB3B8000 , 32'h07CE7898 , 32'hFEFCF678 , 32'hF2A42240 , 32'h048069D0 , 32'hEE5D3620 , 32'hF4E264B0 , 32'hF919B1D0 , 32'h122E5D00 , 32'hED791900 , 32'h00E4BAC4 , 32'hF6C2D520 , 32'hFCE7C008 , 32'h01C9A7CC , 32'hEF6FF140 , 32'hF723BF80 , 32'hEFA007C0 , 32'hF06D2920 , 32'h00772565 , 32'hF5C8F260 , 32'hFE06A478 , 32'hF9D04850 , 32'hF8A96F90 , 32'h0A877530 , 32'hFE4F5B3C , 32'hF53FC0B0 , 32'h01019268 , 32'hF284BE90 , 32'h0AAB6B90 , 32'hFED4AB70 , 32'hF492D540 , 32'hFF4FB182 , 32'hF1D09310 , 32'hF6D30700 , 32'hFA58F3C8 , 32'h05FBC050 , 32'hF8521D00 , 32'hF943C310 , 32'hFEC890B4 , 32'hEFED2980 , 32'hF896E138 , 32'h057CD400 , 32'h015388B8 , 32'hFEFA3C44 , 32'h0A1107F0 , 32'h0468F760 , 32'h09EE6BA0 , 32'h03014708 , 32'hF9853F70 , 32'hFC933234 , 32'hFD9D86B4 , 32'hFA6DCD98 , 32'h0AA1F890 , 32'hFA47D868 , 32'h00038E97 , 32'h019DBC94 , 32'h01A54D64 , 32'h0195E970 , 32'hFE32A1E4 , 32'hFF2D3CCD , 32'h04227550 , 32'h0053503F , 32'hFF1C0C2C , 32'h0121A8B8 , 32'hFF37EEBA , 32'h04F10988 , 32'hFA46A8D8 , 32'hFED75F68 , 32'h02E9FB70 , 32'h0128BD74 , 32'h033699D8 , 32'h009DE30C , 32'h00E3B788 , 32'hFEA8DCA8 , 32'hFC7040C8 , 32'hFEE0023C , 32'hFFD6022B , 32'hFFFF178A , 32'h00005EC0 , 32'h000129F1 , 32'hFFFDDD98 , 32'hFFFFA92E , 32'h00000295 , 32'h00021472 , 32'h0001A99A , 32'h000093BE , 32'hFFFE8205} , 
{32'h235AD140 , 32'hF0DA6BC0 , 32'hE66A8740 , 32'hE4F0D940 , 32'h2BB58CC0 , 32'hE2167040 , 32'h28E42540 , 32'hEA7F4120 , 32'hFD6F0B20 , 32'h0952F480 , 32'h23A7F600 , 32'h146ED620 , 32'h1DF03560 , 32'h214A73C0 , 32'h1588C280 , 32'h04E037E0 , 32'hEA8FC460 , 32'h0C48B530 , 32'h0EA06660 , 32'h003688D0 , 32'h0FDB7770 , 32'hFEEE4904 , 32'hF6CB8990 , 32'hEB902EE0 , 32'hF7054D70 , 32'hFA417038 , 32'h09772870 , 32'hED946EA0 , 32'h01B9E2C0 , 32'h03AB5170 , 32'hF12517E0 , 32'hF392D0F0 , 32'h0148CB54 , 32'hF390FC50 , 32'hFF73DF21 , 32'hFFF8AECF , 32'h09DD75A0 , 32'h01774BFC , 32'hFBC3C630 , 32'h045295A8 , 32'h02D59F24 , 32'hFBADFDF0 , 32'h03BEB518 , 32'h09989750 , 32'h02C21CC0 , 32'h0BBFB320 , 32'hF67607F0 , 32'h09317D00 , 32'hF4EA2B10 , 32'h0B888F90 , 32'hF0A2B610 , 32'h02586568 , 32'h037DE118 , 32'h027ED6EC , 32'hFFC09168 , 32'hF6D545C0 , 32'h014C4590 , 32'h0286C490 , 32'h05CF42A0 , 32'h00F45D59 , 32'hFE5F9E1C , 32'hFD19443C , 32'h008A5D50 , 32'hFFF360F4 , 32'h02C37838 , 32'h008C5ADB , 32'hFC6870CC , 32'h04776B60 , 32'h06510408 , 32'h006C0C88 , 32'hF5433770 , 32'hFCE4CF08 , 32'hFCC25178 , 32'hF96E45D0 , 32'hFCF95888 , 32'hFFCB54C9 , 32'hF99689B8 , 32'h0189F410 , 32'hFCB7823C , 32'hFAE26B68 , 32'h00513931 , 32'h02D83A54 , 32'h04348948 , 32'h00519EAB , 32'h00DDE366 , 32'hFFFB611A , 32'hFFEC507F , 32'hFD844C70 , 32'hFE2368F4 , 32'hFFB744BC , 32'hFFFFF946 , 32'hFFFF75B5 , 32'hFFFE7C3E , 32'h000354BF , 32'h0000ACB9 , 32'hFFFE4685 , 32'hFFFFBC66 , 32'h0001460B , 32'hFFFF627C , 32'hFFFE3ED0} , 
{32'hFFFE3D83 , 32'h0001442B , 32'hFFFB3D91 , 32'h00004177 , 32'hFFFC2849 , 32'hFFFCB29C , 32'h00007899 , 32'hFFFA50D3 , 32'hFFFF191F , 32'h0001E7C3 , 32'hFFFFF038 , 32'hFFFE16F9 , 32'h000044FA , 32'h0001371B , 32'h0004FCB3 , 32'h00021584 , 32'h00005AF8 , 32'hFFFD060D , 32'hFFFFDF1F , 32'hFFFFD541 , 32'h00021BC7 , 32'h00037E53 , 32'h0000C1FA , 32'h000337D7 , 32'hFFFFCD0F , 32'h00018672 , 32'hFFFE7C3A , 32'hFFFE942A , 32'h0002E9B2 , 32'hFFFE1CDD , 32'hFFFF8174 , 32'h0001C772 , 32'h0002839C , 32'hFFFE360D , 32'h00007839 , 32'h00026DBA , 32'h00005CD8 , 32'hFFFC89CB , 32'hFFFC1820 , 32'hFFFC1519 , 32'h000541E4 , 32'hFFFF5DD5 , 32'hFFFE106F , 32'hFFFF370A , 32'hFFFE41B6 , 32'h0005804E , 32'hFFFE6172 , 32'hFFFAFACC , 32'hFFFBBC0B , 32'h00014380 , 32'hFFFD61B3 , 32'h00027BBE , 32'h000096A6 , 32'h00018905 , 32'hFFFEB671 , 32'hFFFE8627 , 32'h0004F849 , 32'h0001AE43 , 32'hFFFB1416 , 32'h00010A9C , 32'h0001974D , 32'hFFFEDD99 , 32'h0004DD2A , 32'hFFFD4E9C , 32'hFFFC2319 , 32'hFFFB9037 , 32'hFFFC97EF , 32'hFFFF7808 , 32'hFFFEF1AC , 32'h000230FB , 32'h00022FE4 , 32'h000366A5 , 32'h00000C3D , 32'hFFFEFDAD , 32'hFFFB26C7 , 32'h0003B08A , 32'h00004D6C , 32'hFFFE3F29 , 32'h0000F39F , 32'hFFFE52C0 , 32'h00002A5B , 32'h0002E572 , 32'h0001AB74 , 32'h0001FCD4 , 32'h00081464 , 32'hFFFF4822 , 32'h000044F9 , 32'hFFFD9605 , 32'h00034DFB , 32'hFFFDBD5E , 32'hFFFBAB96 , 32'h0002E5F6 , 32'hFFFF2606 , 32'h000186A1 , 32'hFFFC43CA , 32'hFFFD9B07 , 32'h0002082A , 32'hFFFB923D , 32'h000139AB , 32'h000422B2} , 
{32'hB987A880 , 32'h1DFEFD20 , 32'hD599BAC0 , 32'h33A63E80 , 32'hE3772D60 , 32'h376D8B80 , 32'hF6017220 , 32'h3ECC7CC0 , 32'hF82F4A88 , 32'h0D226580 , 32'h32F74F00 , 32'h30FAD9C0 , 32'hF0EDB930 , 32'hF0657240 , 32'h055EADB0 , 32'hF6250170 , 32'hE5F62C60 , 32'h0BEA6A80 , 32'h089F7E80 , 32'h19F47DC0 , 32'h15512940 , 32'hF29F1770 , 32'h06D65168 , 32'h0C401E20 , 32'hF96E4B38 , 32'hFDBC11FC , 32'hFA4436E8 , 32'h05BF0A68 , 32'hEEE52500 , 32'hF25FC700 , 32'hFDD0E284 , 32'hF1980390 , 32'hFC2222FC , 32'h01B58E20 , 32'hE7678B80 , 32'h0C0291E0 , 32'hFCA1FE4C , 32'hF8657068 , 32'h01F2C2AC , 32'h010C22E0 , 32'h03BFC838 , 32'h03E06D84 , 32'hFDAE9CF4 , 32'hFDC974E0 , 32'h05408B48 , 32'h017EBD20 , 32'hFED71514 , 32'hFEFFB924 , 32'hF72E97D0 , 32'hF53AB160 , 32'h08DDC800 , 32'hFD1A7410 , 32'h10F998A0 , 32'hFF8BFAD5 , 32'hF66C9B60 , 32'hFC82F2DC , 32'hFBD62A80 , 32'hFDF8927C , 32'hFEC9C06C , 32'hFDFC28D8 , 32'hFA90E480 , 32'h07CA60B0 , 32'h059F21A8 , 32'h016D0984 , 32'hF9B50198 , 32'h03CBBE88 , 32'h0248314C , 32'hFDED7124 , 32'h05D7EE08 , 32'h0030E1ED , 32'h02B6FF5C , 32'hFC00E454 , 32'h04B58D50 , 32'h0440B1C8 , 32'hFD46BAB8 , 32'hFED1B500 , 32'hFA831BE8 , 32'h018E4DEC , 32'hFF4D9FF1 , 32'h04C9C8E0 , 32'hFD6132F8 , 32'h03FECCD4 , 32'h00378D41 , 32'h0240DF5C , 32'hFC9296AC , 32'hFC4EF3BC , 32'hFF60C041 , 32'h007213F7 , 32'h00F6215C , 32'hFFE6CE84 , 32'hFFFFC8CC , 32'hFFFD0465 , 32'hFFFF3DCE , 32'hFFFE594F , 32'h000009A7 , 32'hFFFF522A , 32'hFFFD8B9B , 32'hFFFF760B , 32'hFFFCADD2 , 32'hFFFEE638} , 
{32'hFFFD5BC5 , 32'hFFFBB110 , 32'hFFFFF83A , 32'hFFFDEBB8 , 32'hFFFAED28 , 32'h0001CBDF , 32'hFFF9C19F , 32'hFFFFF7C8 , 32'h00029C17 , 32'hFFFF3CA4 , 32'h00036E37 , 32'hFFFD8BC2 , 32'h00007E23 , 32'hFFFD2C12 , 32'h00002D0E , 32'h0000C569 , 32'h0004FEE7 , 32'h0002ABB8 , 32'h00035A0F , 32'h0001D11B , 32'h0002CCC1 , 32'hFFFE61C9 , 32'hFFFEB770 , 32'h00032F0D , 32'h0006F85A , 32'h00018A47 , 32'h000256EC , 32'h000300AB , 32'hFFFEF727 , 32'h000171D5 , 32'h0001539A , 32'hFFFD1780 , 32'h0002F2C1 , 32'hFFFC563B , 32'h0004C6B3 , 32'h00033ED4 , 32'hFFFDC578 , 32'h0001285A , 32'hFFFEB4AA , 32'hFFFF30D6 , 32'hFFFFF11D , 32'hFFFFABFC , 32'hFFFE2356 , 32'h0002379F , 32'hFFFC6198 , 32'h00047039 , 32'hFFFFE3BE , 32'hFFFDA6C8 , 32'h00010203 , 32'hFFFB6B64 , 32'hFFFFC9C4 , 32'h0000EC84 , 32'h00059BA7 , 32'h00045EAD , 32'h00019480 , 32'hFFFEB68E , 32'hFFFF5448 , 32'h0000EC68 , 32'h0000381E , 32'hFFFF1322 , 32'h00034EAD , 32'hFFFEC021 , 32'hFFFF5EB1 , 32'hFFFEB08C , 32'h00014E5C , 32'hFFFEE17A , 32'h00008AD5 , 32'h000376DF , 32'h00013B70 , 32'h0000B349 , 32'h0002B0DD , 32'h0006B901 , 32'hFFFF45D6 , 32'h0000EF44 , 32'hFFFDAFFA , 32'hFFF84DAE , 32'hFFFC6F11 , 32'hFFF9C860 , 32'h000086A0 , 32'hFFFE8B97 , 32'hFFFA8965 , 32'hFFFF9C1E , 32'hFFFD429B , 32'h0001672E , 32'hFFFFBE8F , 32'hFFFFA99C , 32'hFFFBF721 , 32'hFFFB46BF , 32'hFFFFDE8F , 32'hFFFE7E84 , 32'hFFFB96E0 , 32'hFFF6A3A3 , 32'hFFFC9420 , 32'h0002CB2D , 32'hFFFD29B4 , 32'h000141AC , 32'h0004E4E2 , 32'h00006275 , 32'h000053DD , 32'hFFFFA515} , 
{32'hEE1BA700 , 32'h3444C940 , 32'h2C3C50C0 , 32'h4F034200 , 32'hFA84E898 , 32'hF4E86D80 , 32'h03FA3820 , 32'hD1008C00 , 32'hE42A2280 , 32'h0B743930 , 32'h06E4F148 , 32'hFA94E7F0 , 32'hF731B2A0 , 32'hFD6AC484 , 32'h09E63B80 , 32'h1FC66420 , 32'hE7A05040 , 32'h009EAEDA , 32'hF696C500 , 32'hFC36F8C8 , 32'hF2E6DB50 , 32'hEA84AAE0 , 32'h060CF2C0 , 32'h0D4B5530 , 32'h22C99C00 , 32'hF23E7020 , 32'h0710B350 , 32'hFE03EED0 , 32'h0EDB9400 , 32'hFDB51044 , 32'h05B3DB08 , 32'hEC392CE0 , 32'hF6B76E60 , 32'hF1EE2BA0 , 32'hFDE86DB4 , 32'h0A9E2A90 , 32'h023AEF38 , 32'hF9894B60 , 32'hF74E80D0 , 32'hF6DD8260 , 32'h0193600C , 32'hF88468E8 , 32'hFD7D21C0 , 32'hFE5BE07C , 32'hF9D8FD00 , 32'h06B7FB10 , 32'hFDE587BC , 32'h0F89C250 , 32'hFE2A13E8 , 32'hFC3C7944 , 32'hFF202D3C , 32'hFCA9B69C , 32'hF8A67578 , 32'h0167F2F0 , 32'h0399F970 , 32'hFEE78DF4 , 32'hF8CB4678 , 32'h05766420 , 32'h026A7BE4 , 32'h004E4F65 , 32'hFD744730 , 32'h051ADFA0 , 32'hFE84A574 , 32'h00B049B3 , 32'h02C628B0 , 32'hFEE1BAF8 , 32'h05830880 , 32'hFD114C88 , 32'h02DBF350 , 32'hFA274D40 , 32'hFFE98399 , 32'h05A58390 , 32'hFC1F6034 , 32'h042473E0 , 32'h04864F98 , 32'h03C81508 , 32'h04806258 , 32'hF5D42B50 , 32'h013FDF00 , 32'h038723BC , 32'hFD5DFAAC , 32'h036C579C , 32'h03A60B24 , 32'h03C0EFAC , 32'hFD0B5680 , 32'hFE6A3438 , 32'h05ED7158 , 32'h0151E3A8 , 32'hFF54090F , 32'h0044A4A2 , 32'hFFFDCCAD , 32'h0001E4BA , 32'h00004EBA , 32'hFFFEC863 , 32'h00005D30 , 32'h0000AD13 , 32'h0000ABF8 , 32'hFFFDA538 , 32'h0000BE0E , 32'h0001796E} , 
{32'h02EE95E8 , 32'hF7D85630 , 32'h0038EE1D , 32'h05551F78 , 32'hF353B020 , 32'hFE81161C , 32'hED3E87A0 , 32'hF8023018 , 32'h0ED8C140 , 32'hF13F71E0 , 32'h06D6C608 , 32'hFF802D9A , 32'hF86545D0 , 32'hF8784E50 , 32'hFCF68634 , 32'hFA0462C0 , 32'hFEF802F8 , 32'h00B79C56 , 32'hF600E4F0 , 32'h039CA0E4 , 32'h010F3510 , 32'hFBC87D48 , 32'hFA736518 , 32'h04E6ACE0 , 32'h0128EAF8 , 32'hFB432270 , 32'h012FF048 , 32'h01792C68 , 32'hFF90D74C , 32'hFD7E4844 , 32'hFF488EAE , 32'hF8EB1400 , 32'hF717DB40 , 32'h01CFF810 , 32'h01E64778 , 32'hFE07230C , 32'hF9B3EE40 , 32'h013321D4 , 32'h086F7E20 , 32'hFE56D190 , 32'h078AB298 , 32'hF7EE61B0 , 32'hFE7EA7AC , 32'hFA080930 , 32'h04142F68 , 32'h026EE8F8 , 32'h0CBEEB50 , 32'hFB1E7E88 , 32'h0C123D00 , 32'h0654A980 , 32'hF60BDF50 , 32'hFCEF68EC , 32'h01FAE60C , 32'h0016F70C , 32'hFF0D274F , 32'hF7FCF680 , 32'h025CFDF8 , 32'h046043E0 , 32'hF95B4358 , 32'h03F1CF20 , 32'h02E62010 , 32'h066E95A8 , 32'hFA99F800 , 32'hF7FB2BC0 , 32'h02A18E80 , 32'h0082077B , 32'h0118772C , 32'h0463DDB8 , 32'h054058D8 , 32'h00DEFC1E , 32'hFF426620 , 32'h031E3F84 , 32'hF7904F00 , 32'h037B9934 , 32'hFFC3B109 , 32'h087DDC30 , 32'h056822A8 , 32'hFB7554D8 , 32'h01FDDD74 , 32'h012C0374 , 32'h0180CF08 , 32'h03AFF1EC , 32'h00F1365B , 32'hFE5329D4 , 32'h0025D87D , 32'hFF0A05BC , 32'hFE449FDC , 32'hFF620079 , 32'hFEE368CC , 32'hFFBD8020 , 32'hFFFFFBA6 , 32'h0002CA33 , 32'h00002350 , 32'h00023682 , 32'h0000F6BF , 32'h00010E33 , 32'h00015335 , 32'h00000B38 , 32'h00018291 , 32'hFFFF29A3} , 
{32'hFFFFCCEA , 32'h00020C43 , 32'hFFFD21FD , 32'h000168A0 , 32'h0001AA75 , 32'hFFFEEE71 , 32'hFFFFF451 , 32'hFFFE3ADA , 32'hFFFA8B84 , 32'hFFFED2DD , 32'hFFFF55BF , 32'hFFFFE9F7 , 32'hFFFD958B , 32'h0000204B , 32'hFFFA3F85 , 32'h00008A9D , 32'h00072D81 , 32'h0000715F , 32'hFFFB29BA , 32'h00038170 , 32'hFFFC5A6B , 32'h0003591D , 32'hFFFFCAAD , 32'hFFFF9D3F , 32'h000125BA , 32'h0002C596 , 32'hFFFCE691 , 32'h00014FA4 , 32'h0002FC4E , 32'hFFFF76CB , 32'hFFFA7C77 , 32'h0001F88E , 32'h0001726F , 32'hFFFF19ED , 32'h000004F4 , 32'hFFFFE8BA , 32'hFFFFECED , 32'h0005B8F5 , 32'hFFFF51D2 , 32'h00005092 , 32'hFFFD7393 , 32'h0002C722 , 32'h000099FA , 32'hFFFFD76F , 32'h0004E290 , 32'h0003B2DD , 32'h000511AA , 32'h000253A4 , 32'hFFFE63D5 , 32'hFFFB8594 , 32'hFFFE6617 , 32'h0006F986 , 32'hFFFBB28F , 32'h0001AB3B , 32'hFFFB2935 , 32'h00018734 , 32'h00001561 , 32'hFFFBDA8B , 32'h00001FA0 , 32'h00026ADB , 32'h00040CF8 , 32'hFFFF3241 , 32'hFFFEF66E , 32'h00010001 , 32'h00019125 , 32'h000164B8 , 32'hFFFDDB73 , 32'hFFFF2149 , 32'h00024CFA , 32'hFFFCE616 , 32'h00044A20 , 32'hFFFED5C3 , 32'h0002B514 , 32'hFFF920A0 , 32'h0000B6BE , 32'hFFFEB9BA , 32'hFFFF4E54 , 32'h0001842A , 32'hFFFE5CC1 , 32'h0000D6F1 , 32'hFFFFC52C , 32'h00024074 , 32'h00037815 , 32'hFFFEEDD7 , 32'h0000618C , 32'hFFFCCA7C , 32'hFFFEC705 , 32'hFFFD46D2 , 32'hFFFDD326 , 32'h0000583F , 32'h0001DFD2 , 32'h000475EA , 32'h0000AD31 , 32'h00014532 , 32'h00012871 , 32'h0000CA30 , 32'h00058060 , 32'h000012B0 , 32'hFFFDBB62 , 32'hFFFEB2F5} , 
{32'hA5BC0D80 , 32'hF465A480 , 32'hDE63F400 , 32'hECE35EC0 , 32'h1E520340 , 32'hD2FF37C0 , 32'h026C8DC8 , 32'h159B3E20 , 32'h21D92580 , 32'h1FB5F1C0 , 32'h04E84978 , 32'hF9110BD0 , 32'hF9492C60 , 32'hF6882910 , 32'h08ED8310 , 32'hF66FFB60 , 32'hF5F11F50 , 32'h0550B120 , 32'hDE117580 , 32'hF7A0FB50 , 32'hFA16A588 , 32'h0074546F , 32'hF9D9DB40 , 32'hF08BC050 , 32'h0C8DC240 , 32'hFF404EE3 , 32'h2A3A0A00 , 32'h09FEB2F0 , 32'hFA6BF800 , 32'hE81E1A00 , 32'h06C9A630 , 32'h002CC55E , 32'hFCEC75CC , 32'h04FBA060 , 32'h011659B0 , 32'hF54B35D0 , 32'hFF938145 , 32'hF535EBD0 , 32'hF4F999E0 , 32'hF431F240 , 32'h008AF7C5 , 32'hFED6D094 , 32'h0126D834 , 32'hFC53D068 , 32'h14C79B40 , 32'h0484AF78 , 32'h034628AC , 32'h015AA190 , 32'h01E11BEC , 32'h052E8A48 , 32'h0083BA73 , 32'hFFDCA237 , 32'hFDC444B0 , 32'h007CA297 , 32'hFD11D56C , 32'h061EE7E8 , 32'h00DE6ED6 , 32'h05BC7138 , 32'hFAAB0840 , 32'h04A76E60 , 32'h01643C50 , 32'h012378C0 , 32'hFFCC03CC , 32'hFFAE3DDC , 32'h04A28548 , 32'hFDC8BF1C , 32'h09CED100 , 32'h0064AA53 , 32'h0638B858 , 32'hFBB61CD8 , 32'h04F8F210 , 32'hF8D9B000 , 32'h002590E2 , 32'h02AAB420 , 32'h026847CC , 32'h01F91C24 , 32'hFE82F2B0 , 32'h01899868 , 32'h07B956E8 , 32'h057480D0 , 32'h02FFA998 , 32'hFC03D11C , 32'h015FD500 , 32'h02242FA0 , 32'h02201D70 , 32'h00EDC4C8 , 32'hFF4690C3 , 32'hFFD34CEA , 32'hFE601D90 , 32'hFF7C0E77 , 32'h00006F58 , 32'h00021314 , 32'hFFFFC8D9 , 32'h0001B162 , 32'hFFFF9014 , 32'h0000515D , 32'h000165DB , 32'hFFFF98E7 , 32'h00020865 , 32'hFFFF0BAE} , 
{32'hD4857240 , 32'hDC84DD80 , 32'h1AF0D540 , 32'hD5F47340 , 32'hD08C2200 , 32'hE9DBA560 , 32'hE2DCD660 , 32'hF3FFD3C0 , 32'h2808E3C0 , 32'h2F12D540 , 32'h19378BC0 , 32'hFB46B190 , 32'hFF98FA4D , 32'h1AC5C8E0 , 32'h0F812750 , 32'h14F8F280 , 32'h02F81E74 , 32'hF455ED80 , 32'h1ECFBCE0 , 32'h0714F518 , 32'hFE3493C0 , 32'h0257F560 , 32'h0B6A8870 , 32'h0BBA34F0 , 32'hFE4AFEA4 , 32'hE98B9F80 , 32'h0082C43F , 32'hF53723E0 , 32'h001154E8 , 32'hF48CB830 , 32'hF87EBC50 , 32'h0A56BFF0 , 32'h0387F504 , 32'hFC768940 , 32'h066D6FD0 , 32'h0BB50D60 , 32'hFDB7B88C , 32'hF5F7B750 , 32'h02B93A8C , 32'h06C35260 , 32'hEF8E1E60 , 32'hFE08E4BC , 32'h06624B78 , 32'hFD85D7D0 , 32'h04693270 , 32'hF50E1240 , 32'h00632B13 , 32'h06DAABA0 , 32'h0738CE80 , 32'hFFAB9A98 , 32'h061BF2B0 , 32'h039E5F84 , 32'hFEC78B20 , 32'hFC6290AC , 32'h037C5C08 , 32'hFB239850 , 32'hFCE560A4 , 32'hFE6C7BDC , 32'h0256093C , 32'hF9382468 , 32'hFE109EA0 , 32'hFA9D2540 , 32'hFA3550B8 , 32'hFF48114D , 32'hFD76174C , 32'hFE034EE4 , 32'hF702EDA0 , 32'h057D6980 , 32'h04F14938 , 32'h03420F58 , 32'h056D27A8 , 32'h032D5DBC , 32'hFFB20B85 , 32'h02427F20 , 32'h0237A33C , 32'h033E548C , 32'hFAFC9DC0 , 32'hFF5F8DA3 , 32'hFA715370 , 32'h02045A00 , 32'hFDB9606C , 32'hFD1E3B0C , 32'hFC4E2288 , 32'h006B818E , 32'h0195DEE8 , 32'hFE81D264 , 32'h00B7A7EB , 32'hFF6E8BCA , 32'h014A21FC , 32'h017F89D0 , 32'hFFFFED2C , 32'h00011579 , 32'h000039DE , 32'hFFFB723F , 32'hFFFE31B9 , 32'hFFFCBC25 , 32'hFFFDB522 , 32'hFFFF0668 , 32'hFFFEFE1D , 32'hFFFFAE2B} , 
{32'hEAD14460 , 32'hF8198DA8 , 32'hD3E91700 , 32'hF59A05B0 , 32'h1BE2D800 , 32'h01154C98 , 32'hF22CC5E0 , 32'h07D118F8 , 32'h14021100 , 32'hFBBBCFF8 , 32'hF85E6AF0 , 32'hFC8E65C0 , 32'h048629E8 , 32'hEB3D05A0 , 32'h04D2B018 , 32'h01365788 , 32'hFC2E9F24 , 32'hF66580F0 , 32'hEDC2C380 , 32'h053FF060 , 32'h0064D7D8 , 32'h0C0FD520 , 32'h044480A8 , 32'hF800F630 , 32'h07FA92F8 , 32'hF796C760 , 32'h10747AA0 , 32'hF2717DA0 , 32'h0741D8F8 , 32'hF8279F20 , 32'hFC657F1C , 32'hE7D5C920 , 32'hFE6DDA1C , 32'h00DEFC7B , 32'hFFA4DA22 , 32'hFDE2CE98 , 32'h116A1E40 , 32'hFDE3A268 , 32'h02097120 , 32'hFD1758AC , 32'h0F07F4C0 , 32'h004F1F57 , 32'h03614A18 , 32'h0BA7DAF0 , 32'hFBA29568 , 32'h0390BD04 , 32'hFFDC4B0B , 32'hFFBDB798 , 32'h06BBC180 , 32'hFD541EB4 , 32'hF906C5C0 , 32'hFE2B19FC , 32'hF88486E0 , 32'hF9887A80 , 32'hF9DAAEC8 , 32'h036CA3C0 , 32'h06253268 , 32'hF8F99508 , 32'hF882C0B0 , 32'h05246970 , 32'hFC372398 , 32'hF86CD260 , 32'hFA583F08 , 32'hF8660BC8 , 32'h0385E354 , 32'h01228DDC , 32'h03EECD24 , 32'hFB9F4A80 , 32'hFD836564 , 32'hFF1529EB , 32'h0170F3A4 , 32'hFFE5D0E4 , 32'h007C1792 , 32'hFC91FC4C , 32'h0AA35110 , 32'hFC53F550 , 32'hFEEFAF5C , 32'h03A602D8 , 32'h00CB9CDC , 32'hFE913F8C , 32'hFB3DFEE0 , 32'h067EC350 , 32'h008930CC , 32'hFFAE39C0 , 32'h00D9FC05 , 32'h08EDCDB0 , 32'h01DFFAD8 , 32'hFFF91C0D , 32'h00F1D49C , 32'hFFD56D28 , 32'h0001643D , 32'h00019FAB , 32'hFFFC8739 , 32'hFFFEB0E7 , 32'h000108D9 , 32'hFFFCC2B6 , 32'hFFFE7A38 , 32'h0001E158 , 32'hFFFB1C74 , 32'hFFFE786D} , 
{32'h0001D9B4 , 32'h00008BBB , 32'hFFFE3D06 , 32'hFFFE6505 , 32'hFFFFD5B1 , 32'hFFFCC4CE , 32'h0002198C , 32'h0002F0DB , 32'hFFFF5FA3 , 32'hFFFD4823 , 32'hFFFF900C , 32'h000406E6 , 32'h0000BC1A , 32'h000031BE , 32'hFFFEEC71 , 32'hFFFC8170 , 32'h00004BDA , 32'hFFFC6350 , 32'h00016B2F , 32'hFFFF03D8 , 32'h0002CEDD , 32'h0001E6EE , 32'hFFFF4393 , 32'h00005506 , 32'hFFFF24E8 , 32'hFFFFEBBF , 32'h00043E48 , 32'hFFFC13EF , 32'h0001C378 , 32'h0000DDBB , 32'h0000693A , 32'h00007C6D , 32'h00014DD1 , 32'hFFFF3571 , 32'hFFFC7B6C , 32'h0000FC9B , 32'hFFF966E0 , 32'h00012E28 , 32'hFFFFBF08 , 32'h00036310 , 32'hFFFE60F0 , 32'hFFFB49D3 , 32'h000328FF , 32'h000117DC , 32'h0000EE78 , 32'hFFFE7A26 , 32'hFFFC06DA , 32'h00019E95 , 32'hFFFCEEED , 32'h0000D3C7 , 32'h0000C914 , 32'hFFFDA985 , 32'hFFFF3DB8 , 32'h00012CFA , 32'h0001FEA2 , 32'hFFFFA529 , 32'hFFFF433E , 32'hFFFDCBAD , 32'hFFFF9B6B , 32'hFFF89A30 , 32'h00018CA8 , 32'hFFFF163A , 32'hFFFFD71C , 32'hFFF8BBDE , 32'hFFFEB2C5 , 32'h0002C8DB , 32'hFFFDF5C8 , 32'h0002D6B6 , 32'h00001ED9 , 32'hFFFDD6EF , 32'hFFFFC554 , 32'h00027F60 , 32'hFFFE1F2B , 32'hFFFEDAC2 , 32'h0002E0EB , 32'h00050CDA , 32'hFFFD4AA6 , 32'h00012177 , 32'h000010E1 , 32'h0001656B , 32'h00047554 , 32'h0000FBE1 , 32'h00014B36 , 32'hFFFC79AA , 32'hFFFFC1D8 , 32'h00014495 , 32'h00047D8D , 32'hFFFE6F71 , 32'h00017F69 , 32'hFFFE45EC , 32'h0005D924 , 32'h00003D15 , 32'hFFFCCD38 , 32'hFFFF0705 , 32'hFFFA5D1C , 32'h000138E4 , 32'hFFFDA1C6 , 32'hFFFF6C2A , 32'hFFFC4709 , 32'hFFFD6659} , 
{32'h00001AA1 , 32'hFFFFE5F4 , 32'h000015D5 , 32'h0000C224 , 32'hFFFE4416 , 32'hFFFCFADE , 32'hFFFEDA7C , 32'h00048455 , 32'hFFF699CF , 32'hFFFB6397 , 32'hFFFCD969 , 32'h00024808 , 32'hFFFDEB01 , 32'h000119C6 , 32'hFFFF3CFB , 32'hFFFFEE6C , 32'hFFFEF1D9 , 32'h0002FFB4 , 32'hFFFAF371 , 32'h0002FCC2 , 32'hFFFF84C1 , 32'hFFFDFC05 , 32'hFFFD2B33 , 32'hFFFDDD64 , 32'hFFFFFFB3 , 32'h00017792 , 32'h00037D8F , 32'h0000E93F , 32'hFFF8186E , 32'hFFFE50D9 , 32'h0001145E , 32'hFFFADD0A , 32'hFFFD4A9B , 32'hFFFCB587 , 32'hFFFF146C , 32'h00015032 , 32'hFFFD9A12 , 32'hFFFE2501 , 32'hFFFED4CA , 32'hFFFBFEF2 , 32'hFFFD2494 , 32'h00040838 , 32'h00034D2E , 32'h00002008 , 32'h0001582A , 32'h00022134 , 32'hFFFC608E , 32'h00016640 , 32'hFFFF579D , 32'hFFFF57D5 , 32'h00005039 , 32'h0004D1AF , 32'h000084A9 , 32'hFFFC4CE0 , 32'hFFFE0F1F , 32'hFFFEFC4F , 32'hFFFB98CE , 32'h0001A06A , 32'h0001D7ED , 32'h00001B1A , 32'hFFFD7B68 , 32'hFFFC3011 , 32'hFFFEDB1A , 32'h00001704 , 32'h0001CB27 , 32'h00061FA2 , 32'h0001CFDE , 32'h00026205 , 32'hFFFC441D , 32'h00012818 , 32'h0004DF3C , 32'hFFFAA607 , 32'hFFFF268A , 32'hFFFEA58A , 32'h00042AB7 , 32'hFFFBA1FE , 32'h00024854 , 32'hFFFF0C1D , 32'hFFFD5936 , 32'h00031C95 , 32'h00003360 , 32'hFFFCE53A , 32'h00034CBF , 32'h00073922 , 32'h0001F222 , 32'h00048E2D , 32'hFFFA322B , 32'h00012AD4 , 32'hFFFCFD3B , 32'h0000BFDF , 32'hFFFFBE5C , 32'h000132A8 , 32'hFFFE93EC , 32'hFFFF619A , 32'hFFFF1EB9 , 32'hFFFFF596 , 32'h000031FE , 32'h00032AE2 , 32'h00009A39 , 32'h000108DF} , 
{32'h0004B32D , 32'hFFFE960F , 32'h0000AD64 , 32'hFFFEA575 , 32'h000152DC , 32'h000185BF , 32'hFFFDB988 , 32'hFFFE064A , 32'h0000C91B , 32'hFFFD3914 , 32'h0000E1C1 , 32'hFFFA72E6 , 32'hFFFE9C23 , 32'h0002994B , 32'hFFFD770A , 32'hFFFE1D75 , 32'hFFFF9569 , 32'h0002AE6E , 32'hFFFF21FE , 32'hFFFF55E1 , 32'hFFFFE494 , 32'h00016714 , 32'hFFFFA3BD , 32'hFFFC8C61 , 32'h0001526F , 32'hFFFFCDE2 , 32'hFFFE381C , 32'h000061F0 , 32'h00032EBA , 32'h0004731D , 32'h0002041B , 32'hFFFE494C , 32'hFFFE0C77 , 32'h00015AAB , 32'hFFFEF287 , 32'h00007328 , 32'h0000127E , 32'h000125AA , 32'h00010699 , 32'h0004654B , 32'h00017546 , 32'hFFFE0325 , 32'h000162D7 , 32'hFFFE5079 , 32'h00007E40 , 32'hFFFFC6F6 , 32'hFFFB7ECA , 32'h000219A2 , 32'hFFFEC0DB , 32'h00024D9B , 32'h00021682 , 32'hFFFECF39 , 32'h000158CC , 32'hFFFCE418 , 32'hFFFED43B , 32'h00008BAD , 32'h0001B3B6 , 32'h00007B7F , 32'h00052195 , 32'hFFFCEA51 , 32'hFFFC3C81 , 32'h00000EA8 , 32'h00008FF1 , 32'h00012310 , 32'h00028E36 , 32'hFFFD5B17 , 32'hFFFC8884 , 32'h000350D3 , 32'h000417B0 , 32'hFFFF99E0 , 32'h0001D191 , 32'h0000A17F , 32'h00007F36 , 32'hFFFE2BDF , 32'h00028F9B , 32'h0000B68F , 32'h0001ED85 , 32'hFFF92E75 , 32'h0000DE05 , 32'h0002E21F , 32'h0000025A , 32'h0000E88B , 32'hFFFEF2D6 , 32'hFFFD2AD3 , 32'h0000A8F9 , 32'h0000289F , 32'hFFFA80E9 , 32'h0002A482 , 32'hFFFFED6C , 32'hFFFFF673 , 32'hFFFED1A9 , 32'h00011BD6 , 32'h00017AFB , 32'h0003A5F4 , 32'h000252BF , 32'h000312F8 , 32'h0002D662 , 32'h0001E48D , 32'hFFFD3067 , 32'hFFFC127C} , 
{32'h1EC7C560 , 32'hDB5FB200 , 32'h059B1EA8 , 32'hCC74C680 , 32'hC9C233C0 , 32'hFD158A94 , 32'h0D648AB0 , 32'h0A2B1E50 , 32'hE39E1E00 , 32'h04360250 , 32'h0A706E40 , 32'hDF131580 , 32'hE6E5F340 , 32'hEBB2C700 , 32'hFD980860 , 32'h1B1BA460 , 32'hFDED1D64 , 32'hDDBA0440 , 32'hF2A1E740 , 32'hF8FF01A8 , 32'hE6C784C0 , 32'hFF7BD4A4 , 32'hEC067640 , 32'h09306360 , 32'hF71B4150 , 32'hF0B05550 , 32'hFF263CA9 , 32'h097E21D0 , 32'hFD4026F4 , 32'h0289C514 , 32'h0003F9D4 , 32'h01245774 , 32'hFF42EAD7 , 32'hEFD9B6E0 , 32'hE377B440 , 32'h0E857F00 , 32'h06F41FB0 , 32'hFE5D42F4 , 32'h051FA2D8 , 32'h109FC340 , 32'h11691040 , 32'hF549EDC0 , 32'hFEA17CF8 , 32'hFD9E1E14 , 32'hF858A080 , 32'hFF274F75 , 32'h0B5CC260 , 32'h07C9DBB8 , 32'hF84CA988 , 32'hF08DD0C0 , 32'hFF993884 , 32'h03CF2A4C , 32'hF3D02190 , 32'hF438BA40 , 32'hFD6DF560 , 32'h0707C060 , 32'h00221145 , 32'hFB3BE2F8 , 32'hFCB96414 , 32'h03268774 , 32'hFD2A3448 , 32'h035CD498 , 32'h034AA1D0 , 32'hFF3A856E , 32'h042F7820 , 32'hFCC29520 , 32'h011E6558 , 32'h0101B830 , 32'h000D2D80 , 32'h00B8BA6D , 32'hFC646AC8 , 32'hFA87B848 , 32'h030DBEAC , 32'h06445AB0 , 32'hFBFA0058 , 32'h008A9DD9 , 32'hFE0E04F4 , 32'hFDEBED18 , 32'hFBE8A5D0 , 32'hFCB60F84 , 32'hFC98C544 , 32'h00654672 , 32'hFC397040 , 32'h00592489 , 32'h044FF970 , 32'h0225E59C , 32'h010ABA44 , 32'hFF36DDD7 , 32'hFD7EED18 , 32'hFF8FF831 , 32'hFFFF3F77 , 32'h0000E8F6 , 32'hFFFD5FE7 , 32'h0002129E , 32'h0000CB20 , 32'h00008772 , 32'h0000375F , 32'h00009E33 , 32'hFFFEB176 , 32'hFFFEBD8D} , 
{32'h0066A103 , 32'h0DDF0A80 , 32'hFF0B0EA3 , 32'h00EADE60 , 32'h0AC7ED40 , 32'h0A2021A0 , 32'h0FA58950 , 32'hFB75D720 , 32'h20B6F4C0 , 32'hFF095319 , 32'hFB335E88 , 32'hFAFD4DA8 , 32'h0AF6ACD0 , 32'h1145D460 , 32'h00646EC6 , 32'h0B9F4550 , 32'hE85B9D00 , 32'h07041590 , 32'h0AD524D0 , 32'hF91479B0 , 32'hFDEFFA24 , 32'hFA8838D8 , 32'h02824ADC , 32'hF407F6A0 , 32'h00CA880D , 32'hF961F7C8 , 32'hED5FB8E0 , 32'h03C4BC14 , 32'hFA5C21E8 , 32'hFAEC7DD8 , 32'h0CD2F540 , 32'h02A6C3D4 , 32'h153E0840 , 32'hFCFBF79C , 32'hFD81E9FC , 32'hF25D6FF0 , 32'hF750DD90 , 32'h02731680 , 32'h0B647180 , 32'h00FE4C5A , 32'h03440470 , 32'hFCD43694 , 32'hFDCE1EF0 , 32'h049516C0 , 32'hEF251FC0 , 32'hFACBDF10 , 32'h0121976C , 32'h036CC5C4 , 32'hF87EE0A8 , 32'h0D36CAE0 , 32'h0763AD78 , 32'hF8535378 , 32'hFB22F1C8 , 32'h03BF9200 , 32'hFA337490 , 32'h092D9F90 , 32'h0524AAD0 , 32'hFFB3D1E3 , 32'hFF55940B , 32'h020D655C , 32'h029A6848 , 32'h02083CE4 , 32'hFB4D19C8 , 32'hF8CD94C8 , 32'hFAA37A68 , 32'hFC54AA94 , 32'hFDD02D1C , 32'h015B7E58 , 32'h03486FF8 , 32'hF9C857A8 , 32'hFD851F70 , 32'hF67A3C40 , 32'h05D79450 , 32'h0357E57C , 32'h04E6DE48 , 32'h061E24B0 , 32'hFEDE4904 , 32'h01B54118 , 32'h019098DC , 32'hF9D1AA18 , 32'hFF6299BD , 32'h00CC544E , 32'hFE57AB24 , 32'h023B0D40 , 32'hFE6C0AC0 , 32'hFB8E8980 , 32'h01E2C314 , 32'h021ADA18 , 32'h025C8D50 , 32'hFF260CA6 , 32'hFFFE9801 , 32'hFFFC9373 , 32'h00015249 , 32'h00007503 , 32'h000154D9 , 32'hFFFFA071 , 32'h0002BD4E , 32'h0001FF64 , 32'hFFFF164E , 32'hFFFFAF54} , 
{32'hFFFCCA18 , 32'h0002D5A3 , 32'hFFFC947A , 32'hFFFF879E , 32'h000352FB , 32'h00011D27 , 32'h00035ABD , 32'hFFFDEE65 , 32'h0000159A , 32'h0000144F , 32'hFFFEC0B2 , 32'h00020B70 , 32'h00002CF9 , 32'h00018570 , 32'h000128DE , 32'hFFFE8AE1 , 32'h000463AD , 32'hFFFDB5D5 , 32'hFFFF86A1 , 32'hFFFFB7A4 , 32'h000027C6 , 32'h00006B78 , 32'h00023064 , 32'hFFFFF29B , 32'h00029CD0 , 32'h000344C1 , 32'h0000BF4E , 32'hFFFF76B4 , 32'hFFFF7E28 , 32'h00017B7C , 32'h0004D5AF , 32'h00021AA7 , 32'h00003DFF , 32'h00014220 , 32'hFFFE1EEF , 32'h000373EE , 32'hFFFF9F85 , 32'hFFFB52DA , 32'h00007508 , 32'h0003898A , 32'h00024E1D , 32'hFFFD04B9 , 32'hFFFFF9D3 , 32'h00021330 , 32'h00011C28 , 32'hFFFF0966 , 32'hFFFFA311 , 32'hFFFE4CEE , 32'hFFFCEAF4 , 32'hFFFB0E2C , 32'hFFFEB23E , 32'hFFFE2400 , 32'hFFFE9829 , 32'hFFFF4CC0 , 32'h00002318 , 32'h00027DBB , 32'h0001F0D3 , 32'hFFFF6937 , 32'hFFFCEA37 , 32'h000184A6 , 32'hFFFDC34D , 32'h00038A79 , 32'hFFFC95B6 , 32'hFFFEDC74 , 32'h00020758 , 32'hFFFF6966 , 32'hFFFF4EB2 , 32'hFFFFB317 , 32'h0000325E , 32'hFFFE82A3 , 32'hFFFF12D6 , 32'h000160D9 , 32'h0003F824 , 32'h0000EDEE , 32'h000222BB , 32'h0004FC8C , 32'hFFFED47E , 32'hFFFC2B16 , 32'h0003FFEE , 32'h0000E4DA , 32'hFFFE1D13 , 32'h0001CE9A , 32'hFFFF09FB , 32'h00026248 , 32'h0000D3E9 , 32'hFFFF1D62 , 32'hFFFE62CC , 32'hFFFD6B36 , 32'hFFFA4774 , 32'h00032D23 , 32'h00005729 , 32'hFFFF2735 , 32'h0000FF65 , 32'hFFFE9A87 , 32'hFFF6B5CF , 32'h000046A1 , 32'hFFFF913D , 32'hFFFFB523 , 32'h00026E61 , 32'hFFFBD0A9} , 
{32'h3F570680 , 32'hA9EC3F80 , 32'h445FF800 , 32'h1E0D3040 , 32'h265439C0 , 32'hE07E10A0 , 32'hFB7DFAD0 , 32'h25FFAF00 , 32'hF904D410 , 32'h063E96F8 , 32'hE69D1220 , 32'hEE55E380 , 32'hE478DB20 , 32'h010E6E2C , 32'hDB089A00 , 32'h1F1CB740 , 32'h1168F620 , 32'h0279E254 , 32'h0380014C , 32'h00E7EDFD , 32'h01FE3848 , 32'h108F2F60 , 32'h1041B5E0 , 32'hE9990DA0 , 32'hF8DC39B8 , 32'h17378AE0 , 32'h1781BDC0 , 32'hF91BE798 , 32'hFF1EDE03 , 32'h07008D38 , 32'h0C6BAB40 , 32'h08F599A0 , 32'hEC654A80 , 32'hFF90CFFE , 32'hEFD19EC0 , 32'hF060F780 , 32'h0ED58220 , 32'h06C9CED8 , 32'hF8C6E878 , 32'hFB822CD0 , 32'hF6736220 , 32'hF0C27130 , 32'hFF1BDD59 , 32'h013894BC , 32'hF83291A8 , 32'hF6A992A0 , 32'h078C7AA8 , 32'h0306181C , 32'hFFE79443 , 32'h003F0896 , 32'hFEA27B80 , 32'hF780A1D0 , 32'h08B5C3E0 , 32'hFD6ED474 , 32'h02848AC4 , 32'hFE3DDC78 , 32'h010229D8 , 32'hFBC8ABB8 , 32'hFBF2FA10 , 32'hFF0785F8 , 32'hFAAF4998 , 32'hF8D95F10 , 32'hFAE9BF40 , 32'h00100CB9 , 32'hF8B44A58 , 32'h02B72018 , 32'hFD45F6F0 , 32'h061A9510 , 32'h02562410 , 32'h0139B7BC , 32'hFD4176F4 , 32'hFF5C2D0A , 32'hFE9DC12C , 32'h01AE07EC , 32'h02917008 , 32'hFB9E1D88 , 32'hFF137ABD , 32'h0001E53E , 32'hFBCBC700 , 32'h00653F92 , 32'hFFA56C44 , 32'hFF92B55C , 32'h0299D2A0 , 32'h002186EF , 32'hFA098D78 , 32'hFBB94CE0 , 32'hFE8D6690 , 32'h02B0FAB8 , 32'h00D1F36E , 32'hFF985ADA , 32'hFFFEF6F9 , 32'h00004EFE , 32'h000126A9 , 32'hFFFE39BA , 32'h000166D7 , 32'h000025D2 , 32'hFFFEC447 , 32'hFFFE543D , 32'hFFFED539 , 32'hFFFF757F} , 
{32'hFD216300 , 32'h0375D80C , 32'h00C2AEF4 , 32'h0185C878 , 32'hF6F3C130 , 32'h02E42988 , 32'h00753E2A , 32'hF2177B60 , 32'h010C5A88 , 32'hFB0B4C50 , 32'hF94AF9E0 , 32'hF9FD3AE8 , 32'hF9B2FB88 , 32'hFF72B74E , 32'hFDB37B40 , 32'h00364285 , 32'h0872EBC0 , 32'hFBACCE80 , 32'h0195C0EC , 32'h01F86264 , 32'h0121DF54 , 32'hFB04FD68 , 32'h06F93378 , 32'hFC146954 , 32'hFF510EA1 , 32'hFECECFF0 , 32'h08BC0330 , 32'hF9A2BAC8 , 32'hFDF78B68 , 32'hF8B0C9A0 , 32'hFBC9F328 , 32'h02F2E3FC , 32'hFFCFAD92 , 32'hFF93BF60 , 32'h0A086C50 , 32'h028D6718 , 32'hFA651478 , 32'h0AF1BD50 , 32'h02F82D68 , 32'hF8852128 , 32'h02E00194 , 32'hFDA81148 , 32'hF9761528 , 32'hFEEB867C , 32'hFB1DCAE0 , 32'h034A1248 , 32'h02B14D10 , 32'h06E897D0 , 32'hFCF133B0 , 32'hFC6EC6B0 , 32'h081328E0 , 32'hFAC51060 , 32'hFFDB9C48 , 32'h04342D90 , 32'h04E11068 , 32'h045DB450 , 32'hFF7B4230 , 32'h03ADE228 , 32'h0244D938 , 32'hFF24DB66 , 32'h02417450 , 32'hFD9C9BA4 , 32'h035D8BE8 , 32'h0B00ADB0 , 32'hFCF9D35C , 32'h0510FAA0 , 32'h054E0498 , 32'hF9367158 , 32'h0346C180 , 32'hFAD52850 , 32'hFC673D14 , 32'hFA92A068 , 32'h00A6C406 , 32'h05016FC8 , 32'hFF497202 , 32'hF793AA70 , 32'h000352D1 , 32'hFE9F8B2C , 32'h055E6B70 , 32'h0414FB80 , 32'hFC1BBFDC , 32'hFDD406C4 , 32'hFE6FA3CC , 32'hFEC7C46C , 32'h02AD2090 , 32'h03F6D860 , 32'hFF3921D1 , 32'h018D2A7C , 32'hFEF24D6C , 32'hFF8E3FC7 , 32'hFFFF6A7D , 32'hFFFD0D8C , 32'h0002F1B8 , 32'hFFFBB35D , 32'h00007CDA , 32'h0004AE61 , 32'hFFFF663F , 32'h00016780 , 32'h0000F0F8 , 32'h0000CB66} , 
{32'hFFFE314A , 32'hFFFD9BAB , 32'hFFFECB37 , 32'hFFFF57B1 , 32'hFFFC6A02 , 32'h000143F7 , 32'h0005B848 , 32'hFFFE8414 , 32'hFFFBAFA1 , 32'hFFFD6479 , 32'h00025B72 , 32'hFFFC4A85 , 32'h00027CD6 , 32'h00008E49 , 32'h0001F1C7 , 32'h000377A2 , 32'h00001489 , 32'h0002FB28 , 32'hFFFCD2E1 , 32'h00033670 , 32'h00005F02 , 32'hFFFD829A , 32'hFFFE637E , 32'h00011CD5 , 32'hFFFDA23D , 32'h0001336E , 32'h000274F8 , 32'hFFFD77A8 , 32'hFFFEFD4B , 32'h0000CB42 , 32'h00002181 , 32'hFFFEDA89 , 32'hFFFF40C2 , 32'hFFFEA730 , 32'h00012A28 , 32'hFFFA3254 , 32'hFFFBFEF5 , 32'h0001C8A5 , 32'hFFFF9FB4 , 32'h00022C91 , 32'h00027653 , 32'hFFFFEC81 , 32'hFFFCBA09 , 32'hFFFFE04D , 32'h00016746 , 32'h0002CD53 , 32'h0000FD82 , 32'h0000357A , 32'h0002B811 , 32'hFFFA6074 , 32'hFFFE7B87 , 32'h0000E063 , 32'hFFFC8D8A , 32'hFFFE7C15 , 32'h0000E964 , 32'hFFFF3767 , 32'h00024AA9 , 32'h0004C705 , 32'h00006B1B , 32'h000197C6 , 32'hFFFF3D39 , 32'hFFFC67D9 , 32'h0002EDF7 , 32'h0002C33C , 32'hFFFE7036 , 32'h00014DFB , 32'h0001A801 , 32'hFFFC3176 , 32'h00010AE9 , 32'hFFFD5AB0 , 32'h0000523C , 32'h00019501 , 32'hFFFD2A51 , 32'h00001011 , 32'h0001C8B5 , 32'h00032EA6 , 32'hFFFDD919 , 32'hFFFFD3DB , 32'hFFFE44A6 , 32'hFFFF7555 , 32'h00023B7E , 32'h0001E137 , 32'hFFFE70D7 , 32'h000173B6 , 32'h0002499B , 32'hFFFF8149 , 32'h000472E0 , 32'hFFFF1C2E , 32'hFFFDDD3D , 32'h00038D20 , 32'hFFFDAF49 , 32'h000175ED , 32'h00033E86 , 32'h0000CAF4 , 32'hFFFF451E , 32'h00011DF5 , 32'h00019C77 , 32'hFFFCA7EC , 32'h00003E60 , 32'hFFFEDF17} , 
{32'hEADA4640 , 32'hA51D0680 , 32'h310FA700 , 32'h0DC0E2D0 , 32'h1F322500 , 32'h03C6359C , 32'hE4719A60 , 32'hD701A080 , 32'h0AEED700 , 32'h120C88E0 , 32'hF61F1480 , 32'hEF79D1C0 , 32'h0D6B4CE0 , 32'hE66E4340 , 32'h0F33A730 , 32'h11549680 , 32'hF6A13B70 , 32'hF6D5CD10 , 32'h174E9AC0 , 32'h0592E4D8 , 32'hFF001377 , 32'hE54A4A00 , 32'hFE0DEDF8 , 32'h02D287EC , 32'hF0CC9B80 , 32'h014660F0 , 32'h08D5E3E0 , 32'h145738C0 , 32'h071A2E20 , 32'hEA99C8A0 , 32'hF34F5A10 , 32'h09C9BCF0 , 32'hF226A7E0 , 32'hFC9B40E4 , 32'hFCCA22AC , 32'hFCA2D6DC , 32'h033A0DA4 , 32'hF8002D08 , 32'h09DC4080 , 32'hFE9F9890 , 32'hF2727A60 , 32'h1B559E40 , 32'h02FBE22C , 32'hFC9EAB80 , 32'h0DAEAFA0 , 32'h0BECF1B0 , 32'h09D96EB0 , 32'hFD2EF344 , 32'hF3A08070 , 32'hFD581D90 , 32'h056F1438 , 32'hFCD4C008 , 32'h0C060430 , 32'h007C74F6 , 32'hFFE04175 , 32'h0410CB08 , 32'h051C1798 , 32'hFABBD460 , 32'hFA2212C8 , 32'h06928898 , 32'hFE7A6F3C , 32'hFB935D20 , 32'hF14937F0 , 32'h07B08A98 , 32'h035F5A58 , 32'hFE7FF5B8 , 32'h046619E0 , 32'h03411450 , 32'hFE0B3EC0 , 32'h070BB948 , 32'hFE395D88 , 32'hFD20296C , 32'h01423E4C , 32'h040DCF08 , 32'hFF6F2BC0 , 32'h00CB51E9 , 32'h02A971B0 , 32'hFFC2C2CB , 32'hFD8D918C , 32'hF89EFDF8 , 32'h00284BE2 , 32'hFD728A88 , 32'h02C0A514 , 32'h0181E444 , 32'h00E99CEB , 32'hFEABB724 , 32'h008D570C , 32'hFF46E692 , 32'hFF3F17C0 , 32'hFFA10451 , 32'h000019CF , 32'hFFFE8C96 , 32'h0000F5A7 , 32'h000135F8 , 32'hFFFF99D4 , 32'hFFFF562B , 32'hFFFFF852 , 32'h0000BB9A , 32'h0000F779 , 32'hFFFFA991} , 
{32'hF1422950 , 32'hFFBD62F2 , 32'hD37AEE00 , 32'hFC150F18 , 32'hFEBAC9DC , 32'hF3B79850 , 32'hFE7D6BB8 , 32'hF7AA0FC0 , 32'hECC05780 , 32'hF5B1B630 , 32'h0F2EEEB0 , 32'hFC9016B0 , 32'h09D629B0 , 32'hF3CB3170 , 32'hF9006818 , 32'hFA1E5428 , 32'hF9A21D70 , 32'h02B265C0 , 32'h08E74E20 , 32'h036C16B8 , 32'h112DD080 , 32'hF9444C10 , 32'hF302EB30 , 32'hFB7C7A60 , 32'hF5ADEC50 , 32'h042941C0 , 32'hFFA07B5B , 32'hFDD3FEA8 , 32'h0A61AE40 , 32'h0C4DF1F0 , 32'h056E9D40 , 32'h017A2134 , 32'h05ED7880 , 32'hFEA3B250 , 32'hF5F5A6A0 , 32'hFD65DEC0 , 32'h011FD4B8 , 32'hFF39FBCA , 32'hFDD8A520 , 32'h07FC3CD0 , 32'hF9544C68 , 32'hF20A8080 , 32'hF0575FB0 , 32'hF1AC5AF0 , 32'h00059B80 , 32'hF5CE7890 , 32'hF141AF80 , 32'h03FEAC0C , 32'hFFBD219E , 32'hFE6639B8 , 32'hFA08DF50 , 32'h033A7E3C , 32'hFD278518 , 32'h072ADBA8 , 32'hFB05F6D0 , 32'hF7837D00 , 32'h06C7DED8 , 32'h00C56FB2 , 32'hFB4ACBD8 , 32'hFA96FF78 , 32'hFF4093A5 , 32'hF7486130 , 32'h015FFBA0 , 32'hFC720C90 , 32'hFE3E0800 , 32'hF8E18E08 , 32'hFB68BB80 , 32'hFCEB8954 , 32'hFE41A968 , 32'hF9D03BA0 , 32'hFCABEF0C , 32'hFCCA2470 , 32'h02C6A4E8 , 32'h02D00120 , 32'h005DD5FD , 32'h000104A0 , 32'h06276A38 , 32'h00964CB6 , 32'hFAE97E70 , 32'h02A07FE0 , 32'hFC9826D0 , 32'hF8C97D18 , 32'h0352F5B8 , 32'h007320BA , 32'hFE4102F0 , 32'h00C96C95 , 32'h013B7710 , 32'h01DBE914 , 32'hFF04C018 , 32'h0054FD1C , 32'hFFFFC86A , 32'h00020D41 , 32'hFFFC6774 , 32'hFFFD6164 , 32'h0001EF32 , 32'hFFFF5588 , 32'hFFFE1F7E , 32'hFFFF6E08 , 32'h00019207 , 32'hFFFCE0D4} , 
{32'h00023080 , 32'hFFFE9E70 , 32'hFFFB34D0 , 32'h000454D0 , 32'hFFFF8E13 , 32'hFFFA56A8 , 32'h00031569 , 32'hFFFBFEBD , 32'hFFFAC85F , 32'hFFFE9198 , 32'hFFFCE514 , 32'hFFFF942B , 32'hFFFE3D5D , 32'h00040AB3 , 32'hFFFEFD2C , 32'h000252B9 , 32'hFFFEBD31 , 32'hFFFF9ED7 , 32'hFFFFE453 , 32'h0000F4EA , 32'h00052B44 , 32'hFFFD2070 , 32'hFFFFB547 , 32'hFFFF82AB , 32'h00020A6A , 32'hFFFF8492 , 32'h00023312 , 32'hFFFC0A30 , 32'h0004EAE8 , 32'h00049FE6 , 32'hFFFF2304 , 32'h0000E82B , 32'hFFFF5D70 , 32'hFFFF1AEF , 32'hFFFEB15C , 32'hFFFEDFF3 , 32'hFFFFC3AE , 32'hFFFE4867 , 32'h00026B49 , 32'hFFFEE4EA , 32'h00041CDA , 32'hFFFDF26B , 32'hFFFECAC9 , 32'hFFFB56EE , 32'h00012508 , 32'h00001AEC , 32'h000255CB , 32'h00015845 , 32'hFFFA90CC , 32'hFFFDFD50 , 32'hFFFDD81C , 32'hFFFE6BCC , 32'h0001DA45 , 32'hFFFC346C , 32'hFFFEFA54 , 32'h00018CA2 , 32'hFFFD8B98 , 32'hFFFDCED9 , 32'h0000BD8F , 32'h0004C843 , 32'hFFFE499A , 32'h00026FE9 , 32'h000057F9 , 32'hFFFEF2B0 , 32'hFFFFE07A , 32'h0000F7AA , 32'h00007BC0 , 32'hFFFC9CF3 , 32'hFFFE35EC , 32'h00006EB4 , 32'hFFFB1B19 , 32'h00034435 , 32'hFFFE7A87 , 32'hFFFD1A15 , 32'h0000EDA7 , 32'h00011340 , 32'hFFFD5FEC , 32'h0003BED5 , 32'h00010D06 , 32'h00022AA0 , 32'hFFFAB5E0 , 32'hFFFECEAD , 32'hFFFE6FD1 , 32'h0003CE71 , 32'hFFFD96DF , 32'h00021141 , 32'hFFFE14D5 , 32'hFFFD28C6 , 32'h000106F8 , 32'hFFFCC222 , 32'h00013114 , 32'h000175C3 , 32'h00046874 , 32'hFFFF895F , 32'h00042FAB , 32'hFFFE7987 , 32'hFFFEB613 , 32'h0001A3A2 , 32'hFFFE18DB , 32'h0001194A} , 
{32'hEC63FDE0 , 32'h0AED0830 , 32'h1879AD80 , 32'hE08AE660 , 32'hF7C4DAE0 , 32'hFF9FB67E , 32'h0415E6C0 , 32'hF318EBA0 , 32'h20B31540 , 32'hF692C410 , 32'hFEC5B384 , 32'h0A28F0F0 , 32'hFA858598 , 32'hFE94F3D8 , 32'h03F63F74 , 32'hFD9BDAFC , 32'hF52D5E40 , 32'hFEA565B0 , 32'hFD5BCFE4 , 32'h02241700 , 32'hF9C538B8 , 32'h0CC4DBF0 , 32'hFA9EC400 , 32'h071C84F0 , 32'h040583C0 , 32'h0F705FE0 , 32'h0150D988 , 32'h006E9331 , 32'h0284B8B0 , 32'hF4FC1840 , 32'h06203E28 , 32'h043CFCD8 , 32'h0229311C , 32'hF1D38520 , 32'hF81E6A20 , 32'h07936450 , 32'hFCED19C0 , 32'hF879CB78 , 32'hFFB4C78D , 32'hFC3CF85C , 32'h039D0F84 , 32'hF8929850 , 32'hF791F2A0 , 32'hF3DA5AC0 , 32'hFBEC62D0 , 32'hFA94DA98 , 32'hFE28CB74 , 32'hFF70D78A , 32'h019DA270 , 32'h00B3C208 , 32'h001FF9D4 , 32'h0180FB08 , 32'hFFE8071E , 32'hF7DE0D90 , 32'hFDA67D54 , 32'h00D9C90F , 32'hF954E140 , 32'hFD953CF4 , 32'h0497A068 , 32'h00BE17BF , 32'h032BE214 , 32'hF9F69578 , 32'h037F7BC0 , 32'h035F6104 , 32'h0842B7B0 , 32'h0809E2E0 , 32'hFC907094 , 32'h03E6B1A8 , 32'h01457F9C , 32'hFCDAD7C0 , 32'hFD8D66CC , 32'hFC14BAC8 , 32'h03FBB1D0 , 32'h0A60E530 , 32'h03164188 , 32'h0094B565 , 32'hF6A11B80 , 32'h04DF1F70 , 32'hFEA57734 , 32'h001F746B , 32'h00D05D24 , 32'h0495A1B8 , 32'h048D8A00 , 32'hFD921670 , 32'hF9E2D098 , 32'h01EC3828 , 32'hFD767A54 , 32'hFE321FFC , 32'hFFEEEDA7 , 32'hFFE1BFF8 , 32'h00023762 , 32'h00029B7D , 32'h00034C73 , 32'hFFFEC270 , 32'hFFFCE4C3 , 32'hFFFD2578 , 32'h0000C7D7 , 32'h00005FE4 , 32'h00010358 , 32'h0002B4D1} , 
{32'hE264E040 , 32'h1E687E20 , 32'hF595C110 , 32'h0DBC9A30 , 32'h1DFFCDA0 , 32'hE8965D40 , 32'hEBCB7040 , 32'h04DC3590 , 32'hF29F0390 , 32'hDD4AF580 , 32'h05659B38 , 32'h0A7E4480 , 32'h0F162D40 , 32'h1AFA23A0 , 32'h0A683160 , 32'h0D80A810 , 32'h0F8C57F0 , 32'hFA15A738 , 32'h065531E0 , 32'hF4F22DB0 , 32'hF75F5890 , 32'h00660902 , 32'h10FECA40 , 32'hF83D2708 , 32'hF53DD4E0 , 32'hF1AC9D80 , 32'h107691A0 , 32'h1E1DFE20 , 32'hF8558C50 , 32'h12010520 , 32'h00DC701C , 32'h033CF43C , 32'hFF5822A1 , 32'h141BC800 , 32'hF99A6C68 , 32'h094D7DE0 , 32'h0C6939D0 , 32'h096BD170 , 32'hF4A4D820 , 32'h07B3C6B0 , 32'h03FA1570 , 32'h04022D18 , 32'h06922B48 , 32'hF9CEBAD8 , 32'h06BD9910 , 32'h08FC4180 , 32'h015B20B4 , 32'hF962F3A8 , 32'h04202160 , 32'h040208E8 , 32'h0D5D7AF0 , 32'h013150C4 , 32'hF859CF30 , 32'h06A04FA8 , 32'h070A5D80 , 32'h05656690 , 32'hF9522188 , 32'h02F66CBC , 32'h09171BF0 , 32'hFA794C48 , 32'hFB0B5188 , 32'hFD02AC60 , 32'h0C760570 , 32'h034EEEE0 , 32'hFC8C9DD0 , 32'h01AB3578 , 32'hFEDE14D4 , 32'h08BE9E90 , 32'h006F8A18 , 32'hFC536CF8 , 32'h023A4D20 , 32'hFED128B0 , 32'h045B9F08 , 32'h048C3CD0 , 32'h0722D0C0 , 32'hFC444524 , 32'hF9E79CD0 , 32'h04628268 , 32'h06207228 , 32'hFB9954C8 , 32'h01543ADC , 32'h0350D540 , 32'hFCA6F7DC , 32'hFDFA61C4 , 32'hFEE63284 , 32'h008D00E2 , 32'h010DEC00 , 32'hFE8E8358 , 32'hFFAAB1B3 , 32'hFFED5FD5 , 32'hFFFA75C3 , 32'h00012E88 , 32'h00012872 , 32'hFFFD5111 , 32'hFFFFF363 , 32'h0000453A , 32'h000043B2 , 32'hFFFF9079 , 32'h0001AB28 , 32'hFFFEC89F} , 
{32'h0A02F860 , 32'hFE332B8C , 32'h0F59F050 , 32'hF0295A70 , 32'h0006D94B , 32'hE6FF9B60 , 32'hF28F8650 , 32'h0868EFC0 , 32'hFC8D54D4 , 32'hF4AF8690 , 32'hFE678E64 , 32'hE8D78260 , 32'h0174EB6C , 32'hFF88EC4F , 32'hF8A3F828 , 32'h04BD40F8 , 32'h0C7AF550 , 32'h03BE1B00 , 32'hFDDD71DC , 32'h0852F240 , 32'h037F8818 , 32'hE9923340 , 32'h0BFE2230 , 32'hFE73E950 , 32'h041C8C98 , 32'hFF098E3B , 32'h05871C58 , 32'h00D46F4F , 32'h08A9F850 , 32'hF7A5ABC0 , 32'h06154538 , 32'hF594E6A0 , 32'h12A2B020 , 32'hFF75ACC7 , 32'h000E4DD8 , 32'h064583B0 , 32'h095473A0 , 32'h0006C3C7 , 32'hFFE2DE74 , 32'hFE024A0C , 32'h0B590B40 , 32'hFA700980 , 32'hF9B54400 , 32'h01A5C3C4 , 32'h045C2340 , 32'h02505784 , 32'h07C19F78 , 32'hFE9C8A28 , 32'hED38A000 , 32'h071A53B8 , 32'hF5C06550 , 32'hFA9A9EE8 , 32'hF5815B90 , 32'h00E74708 , 32'hF90B1E40 , 32'hF51AB9F0 , 32'hFCC57088 , 32'h0017DADE , 32'h09B71E70 , 32'hFAB3D5B0 , 32'hFE4F63B4 , 32'hF8A5CAC0 , 32'hFB740700 , 32'h00863C44 , 32'hFF87A20F , 32'hFD5DAE10 , 32'hFFE5B35D , 32'hFBDDCBE0 , 32'h0493DED8 , 32'h05C7C8A8 , 32'h0A331140 , 32'hFD940430 , 32'h0A0EC510 , 32'h02E87104 , 32'hF97A9120 , 32'h02A0E27C , 32'hFBCEF828 , 32'hFD4D0ECC , 32'h03647314 , 32'h006EF783 , 32'h002B4FC3 , 32'hFC3EC8E0 , 32'h0375AC58 , 32'h0360F438 , 32'hFE157770 , 32'h03DBAA2C , 32'h0158E084 , 32'h003CEB60 , 32'h017519D8 , 32'hFFA37393 , 32'hFFFDAEC9 , 32'hFFFEC69B , 32'h00005D99 , 32'h00010CFB , 32'h0003B440 , 32'hFFFD76A1 , 32'h00019756 , 32'hFFFFC15B , 32'hFFFEDE2C , 32'hFFFF3BF8} , 
{32'hFFFE7E8F , 32'hFFFF2843 , 32'h00014415 , 32'h00033D2D , 32'h00009D42 , 32'h0000EB49 , 32'hFFFF7514 , 32'hFFFEF5C6 , 32'h00034147 , 32'h00047F34 , 32'h0000FD63 , 32'h0001ECF5 , 32'h0003BD8A , 32'h0000A98D , 32'h000552BA , 32'hFFFD40D6 , 32'h00041EB3 , 32'hFFFFADE0 , 32'hFFFDEDC0 , 32'h00029601 , 32'hFFFCAD3F , 32'h000226BD , 32'hFFFEAF4F , 32'h0001DDBD , 32'hFFFE6552 , 32'hFFFF64E4 , 32'h00033599 , 32'h000799C3 , 32'hFFFCAE71 , 32'hFFFD7363 , 32'hFFFE24E2 , 32'hFFFDDDF4 , 32'hFFFE0D17 , 32'h0000CC2A , 32'hFFFF2DD0 , 32'h00023CB7 , 32'hFFFFBD3D , 32'h0005851B , 32'h000010F4 , 32'h0001FBE6 , 32'h00018A09 , 32'hFFFEFB7D , 32'h00039A7E , 32'h0002F93B , 32'h0001B093 , 32'hFFFECE6A , 32'h0001A235 , 32'hFFFDE244 , 32'hFFFBFD18 , 32'h0004A191 , 32'h00022164 , 32'hFFFCCCBD , 32'hFFFB3468 , 32'h0001B759 , 32'h00000503 , 32'hFFFBE990 , 32'hFFFDE8FC , 32'h000192ED , 32'h0000123C , 32'hFFFD4410 , 32'hFFFF3C46 , 32'hFFFCF4D9 , 32'h000094B8 , 32'hFFFD8407 , 32'hFFFDD709 , 32'h000254A4 , 32'h00002F81 , 32'hFFFE5ED0 , 32'h00022578 , 32'hFFFE6A54 , 32'hFFFB7E68 , 32'hFFFE675D , 32'h00025B5C , 32'h0000A2E2 , 32'h00006395 , 32'h00011A30 , 32'h0001C64B , 32'hFFFA3CC9 , 32'hFFFBEF2E , 32'hFFFE3951 , 32'h00016A15 , 32'hFFFE4466 , 32'hFFFF6F90 , 32'h00042919 , 32'h0001713F , 32'h0000BB81 , 32'hFFFC8BF8 , 32'hFFFFA254 , 32'hFFFE93D3 , 32'hFFFEFA35 , 32'hFFFFD6F6 , 32'h00024BDA , 32'h00003C3D , 32'hFFFCBB31 , 32'h000037A0 , 32'hFFFC68BF , 32'h000174BA , 32'h0004E375 , 32'hFFFF48F4 , 32'h0000C7D4} , 
{32'h0004BCFE , 32'hFFFF4630 , 32'h000157C8 , 32'hFFFF92D6 , 32'hFFFFDFBF , 32'h00038266 , 32'hFFFCD621 , 32'hFFFE3F42 , 32'h00007B62 , 32'h000431B9 , 32'hFFFF8AC9 , 32'hFFFF7EA4 , 32'h0000660D , 32'h0000A5D3 , 32'hFFFC8667 , 32'hFFFF8A8A , 32'hFFFDAE65 , 32'h0002B5FA , 32'h0001095C , 32'hFFFB17EA , 32'h00024C82 , 32'h0002966A , 32'hFFFEB7F0 , 32'h0003EBA3 , 32'h00051405 , 32'h0001F2E9 , 32'hFFFDF7D2 , 32'hFFFE36C8 , 32'h000442F4 , 32'h00044169 , 32'hFFFD69D1 , 32'hFFFFC715 , 32'hFFFEF0AA , 32'h0004AE06 , 32'h00044136 , 32'hFFFEF227 , 32'h0000065F , 32'hFFFEE47D , 32'h00016C20 , 32'hFFFE73C4 , 32'hFFFFDC19 , 32'h000110F7 , 32'hFFFE1A0E , 32'h00003E98 , 32'hFFFE5566 , 32'h00006984 , 32'hFFFE64E5 , 32'hFFFE5660 , 32'h000120C8 , 32'hFFFE4FE7 , 32'hFFFD1243 , 32'h0001D0EE , 32'h00010374 , 32'hFFFDA64D , 32'h00004D9B , 32'hFFFEFB0B , 32'h00001A2C , 32'hFFFAC889 , 32'h00015652 , 32'hFFFFE86B , 32'h00027477 , 32'h000052F7 , 32'hFFFEF1DF , 32'h00047298 , 32'h000285BE , 32'h000132BE , 32'hFFFFBF5A , 32'h000467C4 , 32'hFFFCAAF2 , 32'hFFFBDF42 , 32'hFFFB053D , 32'hFFFF44EA , 32'h00038963 , 32'h0001408D , 32'h0001BEF3 , 32'h00059868 , 32'h00039B1C , 32'hFFFB8484 , 32'h0002E28A , 32'hFFFCF96F , 32'hFFFD94E9 , 32'h00062046 , 32'h0001AA22 , 32'hFFFEF350 , 32'hFFFF4BFA , 32'hFFFE7652 , 32'hFFFF55EF , 32'h000348AE , 32'hFFFD20AB , 32'hFFFF896E , 32'h0003D1FD , 32'hFFFF751E , 32'hFFFD41F5 , 32'hFFFBBCFD , 32'hFFFDBA53 , 32'hFFFB3821 , 32'h0001D85F , 32'h0000D4AE , 32'h000552F2 , 32'hFFFFC75D} , 
{32'hF6A625F0 , 32'hE9AD5F60 , 32'hE87665A0 , 32'h3FEF6B40 , 32'hC5E03B00 , 32'h0C42E4C0 , 32'hCCB39700 , 32'hEB3D1460 , 32'hDD08AFC0 , 32'h16AF48A0 , 32'hEF30C9A0 , 32'hE4C91AE0 , 32'h164FD620 , 32'h06311628 , 32'hFCD949C0 , 32'hEBD8A080 , 32'h03FDE934 , 32'h101DAC40 , 32'h0BB119D0 , 32'hF9CEA390 , 32'hEE976040 , 32'h13FDEF80 , 32'h084BA620 , 32'h0D7C4EA0 , 32'h03475520 , 32'h17C0AC20 , 32'hF6636F10 , 32'h0D03F550 , 32'h04DA2FF0 , 32'hFA87F428 , 32'hF6C3F3A0 , 32'h0A1AC570 , 32'h13F46580 , 32'hF5C2EC50 , 32'h0211ED74 , 32'hF9D05508 , 32'h111A1C80 , 32'h09F362E0 , 32'hE9C725E0 , 32'h01288840 , 32'h05471B60 , 32'h02BDFD54 , 32'h0A925620 , 32'h0863D730 , 32'hFFD022CE , 32'h09E57E20 , 32'h09A21600 , 32'h0A0CBE40 , 32'h004233CA , 32'h01D981DC , 32'hFA421B30 , 32'hEE28EBE0 , 32'hF1ADB320 , 32'h04CAC998 , 32'hFCEF1C10 , 32'hF09148A0 , 32'h04366EF8 , 32'h056F9900 , 32'hFEA8852C , 32'hF92CFBF8 , 32'h054F6340 , 32'h004B6E62 , 32'h0863E600 , 32'h052C8088 , 32'h02C1A230 , 32'h05365E08 , 32'hFB05E208 , 32'h00847D05 , 32'h06173B88 , 32'h01338F54 , 32'hFFE6EDF9 , 32'h01E419C8 , 32'h04E7DCB0 , 32'hFFF2B7C9 , 32'hFDE5E228 , 32'h02183B50 , 32'hFDD6F380 , 32'h030103D0 , 32'h00CD42E9 , 32'hFFD3FDFB , 32'hFD28B55C , 32'h0481AA50 , 32'h01E7BDE0 , 32'h00200816 , 32'h0186D630 , 32'hFF463F3C , 32'h00C28F6D , 32'h003A2B35 , 32'hFFEC36BC , 32'h005766A6 , 32'h0001083A , 32'hFFFDB050 , 32'h0001A0BF , 32'h00027D99 , 32'hFFFFE484 , 32'hFFFE0FB2 , 32'hFFFFD2AE , 32'h00014C05 , 32'hFFFFAF40 , 32'h00003561} , 
{32'hFFFB6C4B , 32'hFFFE369F , 32'h00033305 , 32'hFFFDD454 , 32'hFFFEACF9 , 32'h0003471B , 32'hFFFCB303 , 32'h000014FF , 32'hFFFE8D10 , 32'h000426BB , 32'h00011136 , 32'h0002566F , 32'h0001E3F3 , 32'h000223E9 , 32'hFFFF53B5 , 32'h000252B9 , 32'h0002711A , 32'h0004A3B5 , 32'hFFFDFF0E , 32'h0002A477 , 32'h0000A290 , 32'hFFFE7BF0 , 32'hFFFF005A , 32'h00031054 , 32'h0000BCF3 , 32'hFFFD24C3 , 32'h0000138E , 32'h0000A4AE , 32'hFFFE5832 , 32'h0003448A , 32'hFFFF7156 , 32'h00012747 , 32'hFFFF31AA , 32'hFFFAEF30 , 32'h00009273 , 32'hFFFCD49C , 32'h00045DAC , 32'hFFFC8EA3 , 32'hFFFC8FE3 , 32'h0001CA22 , 32'hFFFA18A3 , 32'h00038ACD , 32'h000598CC , 32'h000374B1 , 32'h000142D0 , 32'hFFFC79C7 , 32'h0005262B , 32'hFFFF73DC , 32'h0001C2B7 , 32'h000132BE , 32'h00027CAF , 32'h0001FFBC , 32'h0001D256 , 32'hFFFBB373 , 32'hFFFF134E , 32'hFFFFB2F0 , 32'hFFFF709D , 32'h0001A812 , 32'h0001E5D1 , 32'hFFFD498F , 32'h00011C52 , 32'hFFFF1D5A , 32'hFFFDE86B , 32'h000180F8 , 32'h0001E8DB , 32'hFFFECF77 , 32'h0001C1F7 , 32'hFFFD3E39 , 32'hFFFFAB9B , 32'hFFFFD0CE , 32'hFFFFFA34 , 32'hFFFFF9DA , 32'h00004B59 , 32'h000196EA , 32'h0000EDFE , 32'h0001DB21 , 32'hFFFCA4D1 , 32'h0000AEDA , 32'h0004661F , 32'hFFFE5DA7 , 32'hFFFEA0BE , 32'hFFFF2248 , 32'h00065FC1 , 32'hFFFE1EAD , 32'h00024DB7 , 32'hFFFB0F2A , 32'hFFFDDEA3 , 32'h0001C52A , 32'hFFFDA220 , 32'h00025342 , 32'h00036A72 , 32'h0008620D , 32'hFFFEDB3A , 32'hFFFB6E24 , 32'h00006CD5 , 32'h0002DB48 , 32'h0003CC14 , 32'hFFFCA60F , 32'hFFFEB774 , 32'hFFFF7BD7} , 
{32'hE9927140 , 32'h05262C40 , 32'h09347960 , 32'hEFDE75A0 , 32'h12B76340 , 32'h1D5DF000 , 32'hFC48061C , 32'hEE4ED4C0 , 32'h12F63BA0 , 32'hFA1D1AA8 , 32'h0D3ABA10 , 32'h080AB150 , 32'hF4FA8140 , 32'h09B65B40 , 32'hF0ECF5A0 , 32'hFD14915C , 32'h00912E8F , 32'hF504CDB0 , 32'hF6C26F20 , 32'hF6D67270 , 32'h00BD871B , 32'hFA948A30 , 32'h15105180 , 32'h07378688 , 32'hF8DA96F8 , 32'hFDD1FCCC , 32'hEFAA6F20 , 32'hF66342D0 , 32'hF9FA9D58 , 32'hF5743890 , 32'h0D1545C0 , 32'h06EFE708 , 32'h08BD4B40 , 32'hF8AA1868 , 32'hF5BE8730 , 32'hFE813CDC , 32'h0A5975E0 , 32'hF8764E88 , 32'hF8DD0968 , 32'hFB3DDF30 , 32'h094A1230 , 32'hFCDB6118 , 32'h03F844E8 , 32'h00AA3E79 , 32'h06ABCAA8 , 32'hFCBE57C8 , 32'h07A6E9D0 , 32'hEA96BE60 , 32'hFA5E8748 , 32'hFC1A83DC , 32'hFF36A9B2 , 32'h08F63F30 , 32'hFB650EB8 , 32'hFD752310 , 32'h07A3AC18 , 32'hFC6BCBD0 , 32'h05039FE0 , 32'hF8A42160 , 32'hFDEAB97C , 32'h01695F70 , 32'h02A9DC44 , 32'hF6881870 , 32'hF80393B0 , 32'hFF231E0C , 32'h000D45A7 , 32'h03F3B044 , 32'h016853D4 , 32'hFD32FA08 , 32'h02804004 , 32'hFB148958 , 32'h01E20D28 , 32'hFEA802B8 , 32'hFFC03892 , 32'hFCF7155C , 32'h024BE234 , 32'hF3EFA100 , 32'hFE5F6E70 , 32'hFA90CD30 , 32'hFE54EE54 , 32'hFE1B4CE4 , 32'hFFFDB357 , 32'h00BC3797 , 32'h02CC321C , 32'h034C051C , 32'hFE9BD058 , 32'hFFFF1464 , 32'hFC3DB82C , 32'h005EAD2B , 32'h00B53A14 , 32'hFFC9A9CA , 32'h00017F24 , 32'hFFFFD20A , 32'hFFFDF584 , 32'h00000DF6 , 32'hFFFF3D40 , 32'h00046E7E , 32'hFFFFFF11 , 32'hFFFF3357 , 32'hFFFEB077 , 32'h0002FC0C} , 
{32'h0000668A , 32'hFFFFF589 , 32'hFFFE1476 , 32'h000324D3 , 32'hFFFEB3AF , 32'hFFFEABE3 , 32'h0001C739 , 32'h00033CD2 , 32'h00026FA2 , 32'h0001820B , 32'h000014C6 , 32'hFFFDE073 , 32'hFFFF3F4C , 32'hFFFD4A3D , 32'h00013C9D , 32'h00003B40 , 32'h0000728B , 32'h0002BCD8 , 32'hFFFC3CA8 , 32'h00004E9F , 32'h00029EED , 32'h0000326D , 32'h000448A8 , 32'h0000922D , 32'h00008C9F , 32'h0003263A , 32'h000157DB , 32'h0002104A , 32'hFFFAD2D6 , 32'hFFFFF1D2 , 32'h0001A9DB , 32'hFFFEFCFE , 32'hFFFD8434 , 32'hFFFCA2AF , 32'hFFF9D6A1 , 32'h000578F0 , 32'h00029F38 , 32'h00057FA8 , 32'h00035940 , 32'hFFFEF058 , 32'hFFFDF59D , 32'h000404C6 , 32'hFFFF512C , 32'hFFFD199E , 32'h00024476 , 32'hFFFCEAC8 , 32'h0000707A , 32'h00042E7A , 32'h00036A77 , 32'h0001C18E , 32'h0002B109 , 32'hFFFCC2F6 , 32'h00021B0C , 32'hFFFF7166 , 32'hFFFC5671 , 32'h00034940 , 32'h0003EAF1 , 32'h0000D5A3 , 32'hFFFB6857 , 32'h0000F64F , 32'hFFFC44CE , 32'hFFFEC4B1 , 32'hFFFE181D , 32'h0003C296 , 32'hFFFF48E6 , 32'hFFFCF8D8 , 32'h0002A83B , 32'hFFFFFCE2 , 32'h000082DC , 32'h000207BB , 32'h0002F3F7 , 32'hFFFCCB46 , 32'hFFFE5AFB , 32'h000103D4 , 32'h00013C95 , 32'hFFFE9775 , 32'h0003B42A , 32'hFFFCB896 , 32'h00027A53 , 32'h00003C86 , 32'hFFFF3B6E , 32'hFFFCAA74 , 32'hFFFF59C7 , 32'hFFFD1052 , 32'hFFFF6509 , 32'hFFFF228D , 32'hFFFD0A95 , 32'h00047E73 , 32'hFFFD9FFB , 32'h0000B138 , 32'hFFFD78BC , 32'hFFFDFC4E , 32'hFFFC3BBB , 32'h0000652C , 32'hFFFFA115 , 32'hFFFFE719 , 32'h00024CC9 , 32'hFFFECE0F , 32'hFFFF2462 , 32'hFFFE6E6A} , 
{32'hF037C2E0 , 32'hF9297918 , 32'hE5D891E0 , 32'h14F2C4A0 , 32'h1E8DA880 , 32'h09E7DEC0 , 32'hF8154988 , 32'h046DB948 , 32'hEA28FA00 , 32'hFFD12344 , 32'hF8E205C0 , 32'h0E742B60 , 32'hFA5EBF08 , 32'h094EBAF0 , 32'hF38EB2D0 , 32'hFAF75A70 , 32'hEE4A0580 , 32'hFC115C4C , 32'h10F91480 , 32'h066A4E08 , 32'hF1406350 , 32'hF98C8770 , 32'h03A37D18 , 32'h0B70D2B0 , 32'h0E7CB2C0 , 32'hF83A9F80 , 32'hFA9A14A8 , 32'hFEA5FE78 , 32'h020183A4 , 32'hF9D95A40 , 32'h1D327E00 , 32'h0148635C , 32'hF995ED40 , 32'hFFEFAF41 , 32'hF9B5F7E0 , 32'hF98BD6A8 , 32'h0D812060 , 32'h07511BB0 , 32'h086D6620 , 32'h02CC2A8C , 32'h04F988E0 , 32'h08F40A70 , 32'h01000E60 , 32'h08BB1200 , 32'hFDA7E3B8 , 32'h04EF5F80 , 32'h07B3DF90 , 32'h01361EF8 , 32'h0053E66D , 32'hF575D770 , 32'hFF79AE14 , 32'h02797F54 , 32'h0542B910 , 32'hFFD085A7 , 32'h0A341030 , 32'h06E4C198 , 32'h06D16EE0 , 32'hFECE16F4 , 32'hF9232860 , 32'h02FC4A98 , 32'h065237E0 , 32'hFD4043FC , 32'hFDE5162C , 32'hFCC22B68 , 32'hFB2AD198 , 32'hFD07875C , 32'hFC7296C8 , 32'h09161F20 , 32'h01599028 , 32'h019AA8C0 , 32'hF28ACB30 , 32'hFD40B1E8 , 32'hFFAFBC60 , 32'h001A0702 , 32'hFAFABCE0 , 32'h07792330 , 32'hFA8EB3D8 , 32'h0190ADC8 , 32'h07100D00 , 32'h05B59678 , 32'hF86F7938 , 32'h004C126F , 32'h03D64598 , 32'h01E2FFF0 , 32'h02A27E18 , 32'h019102A8 , 32'hF9DB3350 , 32'hFED2DB60 , 32'h04060570 , 32'h00617585 , 32'h00013C75 , 32'h0003F1F1 , 32'h00023CC8 , 32'hFFFCB6EF , 32'hFFFEE52B , 32'hFFFEA091 , 32'h00040434 , 32'hFFFF37A6 , 32'h0001B95A , 32'hFFFE38F9} , 
{32'h01CD4214 , 32'h01C09FE8 , 32'h019F83F8 , 32'h019E0334 , 32'h034C8124 , 32'h0453C810 , 32'h0197871C , 32'h0070C677 , 32'hFF48A0C3 , 32'hFFE289EE , 32'hFF8CEE7B , 32'h012BE61C , 32'hFFC946C7 , 32'h00BD35BB , 32'h01FE89C0 , 32'h01DE9E48 , 32'h020BAB58 , 32'hFF1EF8EF , 32'hFBA28B20 , 32'h02E671E8 , 32'hFF11ACEF , 32'hFD86F748 , 32'hFE317F9C , 32'hFE9EDCC0 , 32'h0220F40C , 32'hFFD3E404 , 32'h014397FC , 32'h0172514C , 32'h00A26829 , 32'hFDB48688 , 32'hFD686F9C , 32'hFF25A2E8 , 32'h02594880 , 32'hFEC3DD38 , 32'hFDC5EBB0 , 32'hFF3D1DD0 , 32'hFFCE31B5 , 32'h00ABB351 , 32'h0082AAD2 , 32'h009A5446 , 32'h015D57F8 , 32'h0082EC5A , 32'h022736F4 , 32'hFDE74114 , 32'hFE7C8B18 , 32'h02468E30 , 32'hFF930C6C , 32'h01D535D0 , 32'h0078E66F , 32'hFEA06B64 , 32'hFF5BF6CF , 32'hFFFD701E , 32'h008356B3 , 32'hFFA70E46 , 32'hFF423AFD , 32'hFF3643C9 , 32'hFEA86864 , 32'h00B0AB64 , 32'hFFB092E6 , 32'hFF9E05AD , 32'h0086D734 , 32'h0302AC08 , 32'hFFC3659F , 32'h0037983F , 32'h01607A9C , 32'h02E01F1C , 32'hFD265978 , 32'h01C9FCB4 , 32'h00F6A19F , 32'h014F2374 , 32'h006D2341 , 32'hFF40D25D , 32'hFED1F984 , 32'hFF9543EC , 32'hFDB934AC , 32'hFEFC3E44 , 32'hFE6AF4E4 , 32'hFE77A8A4 , 32'hFFA1D7DB , 32'hFFACB86A , 32'h01F974FC , 32'hFE7CA4CC , 32'h00A5E7FD , 32'hFE806288 , 32'hFFDF927F , 32'h00FBD5AE , 32'hFE21DF10 , 32'hFF5CC79E , 32'hFF322810 , 32'hFFDF4DB7 , 32'hFFFFFD9B , 32'h00018203 , 32'hFFFB8493 , 32'h00012CD0 , 32'h0002F17B , 32'hFFFC9817 , 32'hFFFD7ECF , 32'hFFFFC076 , 32'hFFFF4C6E , 32'h0000B1A2} , 
{32'hFFFF736B , 32'hFFFF7D38 , 32'h00000E90 , 32'h0003C0D5 , 32'h00033790 , 32'hFFFE8774 , 32'h00017647 , 32'hFFFDA82A , 32'h00020B34 , 32'hFFFD11FD , 32'h0001FDC5 , 32'h0001E9A8 , 32'h0001F0C7 , 32'hFFFD92F9 , 32'h000322B0 , 32'h00002172 , 32'h00011391 , 32'h00001451 , 32'h0002E0C1 , 32'hFFFE3C62 , 32'hFFFF28FC , 32'h00006B93 , 32'h00018C58 , 32'hFFFF1BF3 , 32'h0000EF43 , 32'hFFFE9328 , 32'hFFFEF6DE , 32'h000027C6 , 32'h00011345 , 32'hFFFF8707 , 32'hFFFC52A3 , 32'h0000ECEB , 32'h00028EF4 , 32'h00015790 , 32'hFFFB201A , 32'h0003FBCE , 32'h0000285F , 32'hFFFF2602 , 32'hFFF861F8 , 32'h0003F99B , 32'h0004D726 , 32'h0001E816 , 32'h00011ED4 , 32'hFFFD4D17 , 32'hFFFD99E8 , 32'hFFFE7C6B , 32'h0000018D , 32'h0002EC35 , 32'h0001F639 , 32'h0002FDF9 , 32'hFFFF957F , 32'h000269E5 , 32'hFFFCC7A6 , 32'h0000CC59 , 32'h0003CD04 , 32'hFFFBD39A , 32'h000288B4 , 32'h00002446 , 32'h00004026 , 32'h00011D9A , 32'hFFFF89AF , 32'hFFFFC2A9 , 32'h00040DF7 , 32'hFFFFFDA4 , 32'hFFFB849A , 32'h0003F63D , 32'h0000AA00 , 32'hFFFE19CA , 32'h000427A3 , 32'hFFFCDA8B , 32'hFFFD7BE0 , 32'h0000B4B5 , 32'h0005AD9B , 32'hFFFCDA25 , 32'h0003BC0B , 32'hFFFDC567 , 32'hFFFC356F , 32'hFFFF06C6 , 32'h0000B011 , 32'hFFFC6DA2 , 32'h00054825 , 32'hFFFF69D4 , 32'h00018CF5 , 32'h0006F1A9 , 32'hFFFECBAE , 32'hFFFD7B32 , 32'h0000B837 , 32'h0000424B , 32'h0000B6C1 , 32'hFFFFE6D4 , 32'hFFFC3EEA , 32'h000100E7 , 32'h0000E35D , 32'hFFFDFB77 , 32'hFFFF1BAF , 32'hFFFCD914 , 32'hFFFFCCAF , 32'h0000235C , 32'h0002391B , 32'hFFFCB89D} , 
{32'h00042EC6 , 32'hFFFF7781 , 32'hFFFBD9B7 , 32'hFFFE86E3 , 32'hFFFA7069 , 32'h00051348 , 32'hFFFE5917 , 32'h00007090 , 32'hFFFCCA60 , 32'hFFFE0556 , 32'hFFFEB05C , 32'h0000C98C , 32'hFFFFF418 , 32'hFFFE9EB3 , 32'h00012BB0 , 32'hFFFED834 , 32'h00033C9C , 32'h0003190B , 32'hFFFC4351 , 32'hFFFE1D7A , 32'h0003B8C8 , 32'h000609C7 , 32'hFFFF9354 , 32'hFFFDC194 , 32'hFFFE57EB , 32'hFFFA0CFC , 32'hFFFE67A1 , 32'hFFFD2A4B , 32'hFFFDC334 , 32'h0000041C , 32'h0000C0E5 , 32'hFFFF60FC , 32'h00027D1E , 32'hFFFF2237 , 32'hFFFCB610 , 32'hFFFDB340 , 32'hFFFF43DD , 32'h00042B3E , 32'h00012C30 , 32'h0003430A , 32'hFFFEF2C8 , 32'h0001B082 , 32'hFFFE2969 , 32'hFFFB8E54 , 32'h0000E3F6 , 32'hFFFE44DE , 32'hFFFEE25B , 32'hFFFD5F66 , 32'hFFFF7288 , 32'h0005C28C , 32'h0000BDF1 , 32'h000347C8 , 32'h0000FED7 , 32'h0001034B , 32'hFFFC82D6 , 32'h000225F2 , 32'hFFFEF794 , 32'h0000C265 , 32'hFFFF8F33 , 32'hFFFF0B34 , 32'h000077B3 , 32'h00029EBA , 32'hFFFE55ED , 32'h00036E06 , 32'h00004B82 , 32'h0002361E , 32'h000169BD , 32'h00007B5C , 32'hFFFE547D , 32'hFFFF8005 , 32'h0002EAE8 , 32'h0002AC8E , 32'hFFFF42FC , 32'hFFFA464E , 32'h00028CEE , 32'h00040F62 , 32'h00024966 , 32'hFFFE5526 , 32'h00049D04 , 32'hFFFB709A , 32'hFFFFFD2E , 32'hFFFDBD61 , 32'hFFFFB973 , 32'hFFF7E96D , 32'hFFFF5BB8 , 32'h0000DA26 , 32'hFFFD8D18 , 32'h00028F8C , 32'hFFF90B8F , 32'hFFFD2000 , 32'h0003BD9C , 32'hFFFFD3F9 , 32'hFFFF2B1D , 32'hFFFEA812 , 32'h00025B7C , 32'hFFFE6E45 , 32'hFFFBED69 , 32'hFFFDFC68 , 32'hFFFD5E91 , 32'hFFFDF6F1} , 
{32'hFFFCD678 , 32'h0004B4CC , 32'hFFFCBBE0 , 32'h00002795 , 32'h00019272 , 32'h00013C7A , 32'h0003A446 , 32'hFFFAC8DD , 32'hFFFFC990 , 32'h0000B94F , 32'hFFFC4F20 , 32'hFFFE088F , 32'hFFFF2CD5 , 32'h00011466 , 32'h000163FB , 32'hFFFCFEF3 , 32'hFFFF14A6 , 32'hFFFEB22D , 32'h00018EF3 , 32'h00028A9A , 32'h00015818 , 32'hFFFB6D22 , 32'h0001DFD9 , 32'hFFFDAF8D , 32'h0001A574 , 32'h0000F044 , 32'hFFFFD585 , 32'h0002CB92 , 32'hFFFDB8E3 , 32'hFFFE9EF6 , 32'hFFFEE756 , 32'h00011863 , 32'hFFFDE245 , 32'h000217B8 , 32'hFFFFDC28 , 32'h000168B4 , 32'hFFFFC2AB , 32'h0003ADF9 , 32'h0001A6DB , 32'hFFFF1D68 , 32'h000078C2 , 32'h00012899 , 32'hFFFFEEEA , 32'h00020C8F , 32'h0001BED3 , 32'hFFFCB7BC , 32'hFFFE7511 , 32'h00001670 , 32'hFFFF0D1C , 32'hFFFE6384 , 32'h00032257 , 32'hFFFFD047 , 32'hFFFE7DE5 , 32'hFFFE30EC , 32'hFFFE0039 , 32'h000549B5 , 32'h00002F25 , 32'h0001AA9D , 32'hFFFEB890 , 32'hFFFE4ADC , 32'hFFFD3573 , 32'hFFFEA85C , 32'h0001DAB2 , 32'h00007CBF , 32'hFFFF6B60 , 32'hFFFFF1D7 , 32'hFFFE088C , 32'hFFFFA0E6 , 32'h00015E15 , 32'h000272A5 , 32'hFFFC01BD , 32'h0000315E , 32'hFFFEA6A6 , 32'hFFFC92C7 , 32'h00017774 , 32'h0001436A , 32'hFFFD5C21 , 32'hFFFF791F , 32'h00044355 , 32'h0004CCCB , 32'hFFFB0426 , 32'hFFFDF4EF , 32'hFFFED0E8 , 32'h0002C8EF , 32'hFFFF8DD7 , 32'h00020564 , 32'hFFFD74AF , 32'hFFF7095A , 32'h00010963 , 32'hFFFC65FE , 32'hFFFEF5EA , 32'hFFFCF995 , 32'h0001267E , 32'hFFFF196C , 32'hFFFD0EB3 , 32'h0004DC06 , 32'h00033C3D , 32'hFFFC8579 , 32'hFFFB8C9F , 32'hFFFFC535} , 
{32'h0002BE65 , 32'h0005E665 , 32'h00062C34 , 32'h00013863 , 32'h0001A3F3 , 32'h00015601 , 32'h0002B5B4 , 32'hFFFE45DA , 32'hFFFC9311 , 32'hFFFB5D9D , 32'hFFFE1DCC , 32'hFFFFC4C4 , 32'h00052891 , 32'h0001E2E4 , 32'h0001DB2F , 32'hFFFFE4ED , 32'hFFFBC896 , 32'hFFFE7220 , 32'hFFFE5FFA , 32'h0003880D , 32'h00023795 , 32'h0002E567 , 32'h00011860 , 32'h00014F52 , 32'h00003731 , 32'hFFFFCD17 , 32'hFFFAFE50 , 32'h00014A12 , 32'hFFFF3D80 , 32'hFFFFA7F4 , 32'h000422FB , 32'h00022F54 , 32'hFFFED9F3 , 32'h0000BFCA , 32'hFFFE9EF3 , 32'hFFFF319F , 32'hFFFEA620 , 32'h00034A76 , 32'hFFFDFA11 , 32'hFFFBEDEB , 32'h0001DF3D , 32'h00015951 , 32'h0001AD03 , 32'h00026CCC , 32'h00008594 , 32'hFFFA49FE , 32'h00026B87 , 32'h00046807 , 32'h0000D2DA , 32'hFFFBCE54 , 32'h0002502E , 32'h0001F229 , 32'h0000BF89 , 32'hFFFF565F , 32'hFFFC98ED , 32'hFFFF471A , 32'h0001AE19 , 32'h0005E25B , 32'h0000A213 , 32'h0002BF35 , 32'hFFFDC928 , 32'h0002AEC2 , 32'h0002B0F9 , 32'h0004B6EB , 32'h0002FF9B , 32'h0000943F , 32'h000077AA , 32'h00030F1C , 32'hFFFF36EF , 32'hFFFA4F25 , 32'hFFFE6795 , 32'hFFFE67BD , 32'h00043ED1 , 32'h0001B994 , 32'hFFFFCD16 , 32'h0002F0F1 , 32'hFFFD54EC , 32'hFFFC8AD7 , 32'hFFFE5897 , 32'hFFFF25A0 , 32'h0000421D , 32'hFFFF2B6F , 32'hFFFF53D0 , 32'hFFFF2CB1 , 32'hFFFEC2FA , 32'h0001032B , 32'h000189A3 , 32'h0001E0E9 , 32'hFFFE654A , 32'hFFFF9997 , 32'h0001CD54 , 32'hFFFB620E , 32'h00015F8E , 32'hFFFE8D7B , 32'h0001F943 , 32'h0001452C , 32'h0003570A , 32'h000263CC , 32'h0000CA15 , 32'hFFFE3404} , 
{32'hFB6CB248 , 32'h0DE52F50 , 32'h13939D20 , 32'hE9217C00 , 32'h0E7C4B00 , 32'h1101A0E0 , 32'h0DB9E0A0 , 32'hEE916600 , 32'h14F1F540 , 32'hF7DE6560 , 32'h23B0D4C0 , 32'hECD424C0 , 32'hF580D6F0 , 32'h100DA6C0 , 32'hFE1E2598 , 32'h0DA4BB00 , 32'hE5B06F40 , 32'hFF908FD4 , 32'hF6989800 , 32'h022F9EB8 , 32'hFB961A20 , 32'hF82C93B8 , 32'h0421B910 , 32'h080269C0 , 32'hFC481310 , 32'h17BE1BE0 , 32'hFDDC7D54 , 32'hF3A99790 , 32'hF3305200 , 32'h0BAF7AC0 , 32'h0E345AE0 , 32'h05482480 , 32'h07B470B8 , 32'h0A0A97A0 , 32'hF7A0EA00 , 32'h0831CB60 , 32'h07A1E490 , 32'h007D097C , 32'h061D1128 , 32'hFE53506C , 32'h018DE1B4 , 32'hFFADA78E , 32'hFFF27734 , 32'hF2A87FF0 , 32'hFAEB6B20 , 32'hF448D6D0 , 32'h03832EB4 , 32'h05EA1AB8 , 32'h08E206C0 , 32'hFB4FEB50 , 32'hF5501170 , 32'h07F3F1A0 , 32'h0B21CDE0 , 32'h08CE3E30 , 32'h055495E0 , 32'hFE11F86C , 32'hFE8A981C , 32'h003B5244 , 32'h0B883ED0 , 32'h08D6DD30 , 32'hF91AF108 , 32'hF0FC6440 , 32'hF917A460 , 32'h08643620 , 32'h00FC6F6D , 32'h02E1D1B0 , 32'h009F573F , 32'hFF075F3C , 32'hFDB8EFF4 , 32'hFEEB5814 , 32'hF8012A58 , 32'hFEED0B24 , 32'h0237E3F4 , 32'hFF6238AB , 32'h003119DA , 32'h068E2398 , 32'h00DF900A , 32'h003FED72 , 32'hFF6B4F88 , 32'h00C22013 , 32'h008D2B67 , 32'h070E0650 , 32'hFE95F000 , 32'hFD9E6494 , 32'h011582C8 , 32'hFF799624 , 32'h0344236C , 32'h0066B9E0 , 32'hFE775CCC , 32'hFFDC107D , 32'h0001EE38 , 32'hFFFD727A , 32'hFFFF268C , 32'hFFFF8231 , 32'hFFFE35DE , 32'h00006C93 , 32'h0000926D , 32'hFFFF62D8 , 32'h0001F295 , 32'h00007381} , 
{32'h0E824DA0 , 32'h0309BA1C , 32'h07722970 , 32'hE39B5280 , 32'h06EB3EB8 , 32'hF43571A0 , 32'hFD7057B8 , 32'hFF125C3C , 32'h08341670 , 32'hF9238D08 , 32'hFEB5F950 , 32'hFBF01E90 , 32'h07B09D10 , 32'hFA3C8EE8 , 32'hFF893691 , 32'h061E69D0 , 32'h07740B40 , 32'h1511D160 , 32'hF03D6E70 , 32'h08CB7330 , 32'hF14FB150 , 32'hF5219360 , 32'h0E7FA660 , 32'h0B056D80 , 32'h01F64D1C , 32'hFEBB9A10 , 32'h00FC1E90 , 32'h00D4503B , 32'h02593570 , 32'h1720B920 , 32'hFD7AD924 , 32'h03701B0C , 32'h0BD650B0 , 32'hF49CD110 , 32'hF6D1C430 , 32'h0C4F1930 , 32'hFFE18ED4 , 32'hF43D07C0 , 32'h01AAC9BC , 32'h05EBA348 , 32'hF8F6F940 , 32'hF5CAF610 , 32'h01A3470C , 32'h0291EB3C , 32'h0894E640 , 32'h055A8BD8 , 32'h0200DE10 , 32'hF85915C0 , 32'hFDC6D950 , 32'h004BB004 , 32'hFD0EBA80 , 32'hFEC58CF4 , 32'h004CD07E , 32'hFA9A7680 , 32'hE8803820 , 32'hFD81F700 , 32'h0137974C , 32'hF5B05A10 , 32'h099D18B0 , 32'h03B7F20C , 32'h000BD0EF , 32'hFFBDD78C , 32'hFD25CF20 , 32'hFD5D2F2C , 32'h00340A7A , 32'h010BD8C0 , 32'h07F71510 , 32'h0334BDC0 , 32'h000F2C71 , 32'h03BCB24C , 32'hFF42D41C , 32'h07A2B728 , 32'h03F355C0 , 32'h00502B0F , 32'h0410C050 , 32'hFFBDF1B8 , 32'hFB4B75B0 , 32'h01C3FD60 , 32'hFD4285E4 , 32'h00F69B99 , 32'hFDFC76F4 , 32'hFFD18F09 , 32'h0148F9B0 , 32'h034FB9C0 , 32'hFEC32E74 , 32'hFE63148C , 32'h01816138 , 32'hFAE1FF78 , 32'h03E10F6C , 32'h00A067C2 , 32'h00029675 , 32'h0001E4E3 , 32'h00027AF8 , 32'hFFFF3E17 , 32'hFFFF9A70 , 32'h00017A38 , 32'h00009010 , 32'hFFFD6C28 , 32'h000043FD , 32'hFFFFFD1B} , 
{32'h0001A408 , 32'hFFFC4D73 , 32'hFFFC4056 , 32'h00024675 , 32'hFFFEC902 , 32'hFFFDF490 , 32'h000313E0 , 32'h000110A6 , 32'h0002AEE7 , 32'h00008111 , 32'hFFFFC36C , 32'hFFFF35ED , 32'hFFFED43F , 32'h00047BD0 , 32'hFFFF7F92 , 32'h00022C93 , 32'hFFFCEF1E , 32'h00000A5B , 32'hFFFEB279 , 32'hFFFF9337 , 32'h0000C4CB , 32'h0001F41E , 32'hFFFC5D5A , 32'h0000B240 , 32'hFFFC97AB , 32'h00066665 , 32'hFFFB0B69 , 32'hFFFDC30C , 32'h0008BAAC , 32'h000292C3 , 32'hFFF9DDB5 , 32'hFFFD1B1C , 32'h000256B3 , 32'h000334F4 , 32'hFFFF7CAE , 32'h0003F6DB , 32'h0000FAA5 , 32'hFFFDBD8B , 32'hFFFED512 , 32'hFFFB792B , 32'h000240BB , 32'h0001A5ED , 32'hFFFC872B , 32'hFFFC04A3 , 32'h00005586 , 32'hFFFFD948 , 32'hFFFDE278 , 32'hFFFFC777 , 32'hFFFBD562 , 32'h000101AF , 32'h0000108B , 32'hFFFDF300 , 32'h00069687 , 32'h00013DB2 , 32'hFFFDF53E , 32'hFFFDABB0 , 32'hFFFE8E82 , 32'hFFFD2526 , 32'h0001DFB4 , 32'h00001C34 , 32'h00041554 , 32'h0002FA85 , 32'h00025BE5 , 32'h0004EBE9 , 32'hFFFD9F1C , 32'h00005C0B , 32'h0000F09A , 32'h0001AC0A , 32'h00031AEB , 32'h00005042 , 32'h00065A01 , 32'hFFFF1AC6 , 32'h0002EBC3 , 32'h0000398C , 32'h00011294 , 32'h000063A2 , 32'hFFFD7F32 , 32'hFFFE47F7 , 32'h0000FD86 , 32'hFFFC9649 , 32'h00030A16 , 32'hFFFD83C9 , 32'h000286CE , 32'h00013831 , 32'h00012B79 , 32'h0005B9CC , 32'h000413B2 , 32'h0001CA0F , 32'h0002CE08 , 32'hFFFE0BFA , 32'h00008258 , 32'hFFFD7326 , 32'hFFFF4005 , 32'hFFFEAB2D , 32'h0000C025 , 32'h00029FA6 , 32'hFFFAD9EF , 32'h00039AF7 , 32'h00030A2D , 32'h000186FF} , 
{32'h0B3C2230 , 32'hF5DD7FB0 , 32'h01492908 , 32'hE84CFF60 , 32'h2C0225C0 , 32'h28E70FC0 , 32'h0D885760 , 32'hFBC19228 , 32'hFB77E510 , 32'hFAD78780 , 32'h26E2FC00 , 32'hEB4D1100 , 32'h08BDF660 , 32'h187C8A80 , 32'hFD19F300 , 32'h044539D8 , 32'h08E78560 , 32'h0B90B310 , 32'hFBE39D48 , 32'hF34F28C0 , 32'h03C60720 , 32'hE87369C0 , 32'hFCDD7D04 , 32'hF9341938 , 32'hF2BEEA80 , 32'hF75E7230 , 32'hFD5EA9BC , 32'hF8AB2F60 , 32'hFC18E1D4 , 32'h05012690 , 32'hFBD28738 , 32'h032CF3E0 , 32'hF55854B0 , 32'hF6830750 , 32'h08B514E0 , 32'hF84A2690 , 32'hF4D42A50 , 32'hF2B28C60 , 32'h05BDC080 , 32'hF1D4D8A0 , 32'hF86FB030 , 32'h0F2E4450 , 32'h0F329D70 , 32'hFF3C0005 , 32'hF8F457F8 , 32'hF7E74920 , 32'h04A14858 , 32'hF40263C0 , 32'hFB3C0418 , 32'hFD26F950 , 32'hFE140910 , 32'hEF7A5B40 , 32'hF3AFF450 , 32'hFB334E40 , 32'h04AB3E90 , 32'hFC939E58 , 32'h07BFCBE0 , 32'h0851FC10 , 32'h00716B3A , 32'hFC8DE090 , 32'h016A17B4 , 32'h04852478 , 32'h091218F0 , 32'h0470FC78 , 32'hF6290D00 , 32'hF95AA620 , 32'hF93E43F8 , 32'hFC837880 , 32'h00B13BE2 , 32'h03A91400 , 32'hFCF6483C , 32'hFD13716C , 32'h00BEBFB6 , 32'h005EA86B , 32'h049AD2B0 , 32'hFF4BB201 , 32'hFA4DAEB0 , 32'h01B4DAA8 , 32'hFE33D538 , 32'h07D69E40 , 32'hF92DF1A0 , 32'h061078D0 , 32'h01BDC0CC , 32'hFE3DF908 , 32'h037C5894 , 32'h0063EAFD , 32'h0177D5F4 , 32'h00DE3359 , 32'hFD270690 , 32'hFF83EA95 , 32'hFFFFD793 , 32'h0000E085 , 32'hFFFF3A3C , 32'h0002319D , 32'h0001CADA , 32'h00003541 , 32'h000048FB , 32'hFFFEDACB , 32'hFFFFF6AD , 32'h000126B7} , 
{32'hD4A5D580 , 32'hCF0ADE00 , 32'hD47ED500 , 32'hF46C2430 , 32'h2094D180 , 32'hF4096580 , 32'hF56B6BD0 , 32'h04D24EC8 , 32'hF90E20D8 , 32'hEC70A2C0 , 32'h0481DD98 , 32'hEAAF2BC0 , 32'hE9B10800 , 32'h125E8D20 , 32'hC2192240 , 32'h03523CD0 , 32'hFA7CD8D8 , 32'hFD1BF548 , 32'hE9384480 , 32'hFD26F084 , 32'hFC967328 , 32'hF27F3770 , 32'hF3B20930 , 32'hF6003FA0 , 32'h0ABF7310 , 32'hF0D65630 , 32'h0A2917B0 , 32'hF9943B88 , 32'h19101420 , 32'hF736E080 , 32'hF0608F10 , 32'h09961180 , 32'hFF6AB940 , 32'h0794F3F8 , 32'hF1815F80 , 32'h15C2E7A0 , 32'h03EA7834 , 32'hF8D792D0 , 32'h02BB4258 , 32'hF72B47D0 , 32'h001E99C7 , 32'hFCFC35C8 , 32'h01A42AF4 , 32'h009DB21D , 32'hF4466720 , 32'hFFFBA0F8 , 32'h044C1158 , 32'h093FDF60 , 32'hFDDEE504 , 32'h0D2AF860 , 32'h076230D0 , 32'hFBEE23C8 , 32'h0EBA6AA0 , 32'hF0AE67E0 , 32'hFA0505A0 , 32'hFF75DE8D , 32'h04BEE290 , 32'h05D228D8 , 32'h013EF2B8 , 32'hF12E37E0 , 32'hFE9236F0 , 32'h03A54024 , 32'h071B3080 , 32'hFECEB21C , 32'h00DBED7E , 32'h040F9430 , 32'hFAF8F310 , 32'h04AAFF98 , 32'hFCAFBA9C , 32'hFF313FB3 , 32'hFD937390 , 32'hFCFF4258 , 32'hFB92BBA0 , 32'h0044D1EA , 32'hFDFD76E8 , 32'hFC59EFE0 , 32'h01E2A1E4 , 32'hFE7BB814 , 32'h054C15D8 , 32'hF9201580 , 32'h032F89F4 , 32'h0330EA44 , 32'hFD644DF4 , 32'hFEAAC744 , 32'h02F8453C , 32'h012C883C , 32'h009957F2 , 32'h014A74A4 , 32'hFF91BB75 , 32'h01431A6C , 32'h0002A315 , 32'hFFFD01EA , 32'hFFFEF545 , 32'hFFFF1240 , 32'hFFFDE7D3 , 32'hFFFC4B94 , 32'hFFFF0DB5 , 32'hFFFEFA4C , 32'h0000E44C , 32'h00012986} , 
{32'h0F5D3A00 , 32'h04EFA280 , 32'h1E22A700 , 32'hF475CE90 , 32'h08B05DA0 , 32'hEECF3F20 , 32'hF547C640 , 32'hFC9BBA64 , 32'hF29393A0 , 32'hF3269000 , 32'h151F9100 , 32'h01DFDB94 , 32'h08661850 , 32'h0C84F510 , 32'hFA728A10 , 32'hF8F14038 , 32'hFCE26B5C , 32'h04583400 , 32'hF8BE1050 , 32'hFD44E988 , 32'hFC05121C , 32'hFC94352C , 32'hED9AD860 , 32'h0640CB20 , 32'h00F7B4E1 , 32'hF7AD5BD0 , 32'h0E8A58C0 , 32'hF067C950 , 32'h000200DF , 32'hFE66DDE0 , 32'hF9C46628 , 32'h022E5280 , 32'h15B89060 , 32'h00B63E9C , 32'h07178240 , 32'h049FFD88 , 32'h01791984 , 32'hFBCFE250 , 32'h009B7F59 , 32'hF64E8400 , 32'hF77B2350 , 32'hFAE984D8 , 32'hF91B9398 , 32'h0821C280 , 32'h0C213D60 , 32'h00302843 , 32'h068426C0 , 32'hFC20B8AC , 32'h025451F0 , 32'hFB51B9A0 , 32'h0273421C , 32'hF8C94980 , 32'h05566770 , 32'hFB8542A0 , 32'hFC12501C , 32'h0821DDC0 , 32'hFCE4CAE0 , 32'h04E97C10 , 32'hFE9BFBB8 , 32'h038A6694 , 32'h03F85120 , 32'hF5FF1930 , 32'hFCA19FB0 , 32'h01932D08 , 32'h00BBE23E , 32'h03E924E4 , 32'hFEE37990 , 32'hFD067FB0 , 32'h0143E290 , 32'h020D9368 , 32'hFB0D3908 , 32'h047DB5F8 , 32'h039E1608 , 32'hFFD33E3D , 32'h00776ADE , 32'hFD327480 , 32'hFFEFE336 , 32'hFEF7B5B4 , 32'hFD50CA4C , 32'h060C7690 , 32'hFF7D1677 , 32'h036F0228 , 32'h017DBB30 , 32'hFD362848 , 32'hFB2B23F0 , 32'h016639D8 , 32'h006F4483 , 32'hFECF098C , 32'hFE8810E8 , 32'h01413290 , 32'hFFFFAA97 , 32'hFFFDF781 , 32'h00007AF4 , 32'h0002EC11 , 32'hFFFF6BC2 , 32'h0001B7D3 , 32'hFFFE958A , 32'h0002C848 , 32'hFFFFEDC6 , 32'hFFFEC16F} , 
{32'h0005B3B2 , 32'h0002629C , 32'hFFFFE327 , 32'hFFFECBD4 , 32'hFFFD4D13 , 32'hFFFE1702 , 32'hFFFDA7E7 , 32'h0000C4B5 , 32'h00000E8B , 32'hFFFDB9E5 , 32'hFFFDC127 , 32'h0001FDF9 , 32'h0000D2B1 , 32'h00011B4F , 32'hFFFDF965 , 32'h0001A69D , 32'h000232E7 , 32'h0000B22D , 32'h00034A53 , 32'h0004ADDC , 32'hFFFF2008 , 32'h00028C50 , 32'h0003B94A , 32'h00006F38 , 32'hFFFDE178 , 32'hFFFAC30A , 32'hFFFF1D0B , 32'h00001F74 , 32'hFFFA0EE9 , 32'hFFFD2D3F , 32'h00010A1E , 32'h00017112 , 32'hFFFE808B , 32'hFFFF4208 , 32'h0000942A , 32'hFFFF1033 , 32'h0003DD89 , 32'hFFFBE8BB , 32'hFFFDE6BA , 32'hFFFD5996 , 32'h00027DEB , 32'hFFFFB7E0 , 32'h000089A2 , 32'h0003BE97 , 32'h00025C76 , 32'h0003026F , 32'hFFFF829C , 32'h00002FC9 , 32'h0002AE6A , 32'hFFFDB71C , 32'h0001BD56 , 32'h00002CED , 32'h00034E8E , 32'hFFFDC101 , 32'hFFFC1ADF , 32'h0002B6C5 , 32'h00004AA9 , 32'h000596EF , 32'h00027642 , 32'h00020144 , 32'hFFFCE256 , 32'hFFFB404B , 32'hFFFEEA7F , 32'hFFFF575C , 32'h0004A647 , 32'h00017B1A , 32'h00006F37 , 32'hFFFD9528 , 32'h0001F016 , 32'h0000E107 , 32'hFFFECCE2 , 32'h00027FC8 , 32'hFFFBCA1F , 32'hFFFEBD3F , 32'h00002AEF , 32'hFFFCF491 , 32'h00013487 , 32'hFFFF5C69 , 32'h0000450B , 32'h0001B1A5 , 32'hFFFE6789 , 32'hFFFBFAF6 , 32'hFFFE5C84 , 32'h00016770 , 32'hFFFBFD86 , 32'h00009F24 , 32'h0001DD57 , 32'h0001EE72 , 32'h0007DE3A , 32'h0003090E , 32'hFFFE3EA3 , 32'h0000245F , 32'hFFFE54B9 , 32'h0001C41A , 32'hFFFF76AD , 32'h000405D2 , 32'h000029D9 , 32'hFFFD3F96 , 32'hFFFC6A5F , 32'hFFF9D132} , 
{32'hFFFF9DA3 , 32'hFFFF1A04 , 32'h0000EF02 , 32'hFFFED041 , 32'hFFFEE931 , 32'hFFFE523F , 32'hFFFF099F , 32'hFFFFB7B9 , 32'h0001A609 , 32'h0000E906 , 32'hFFFEDF05 , 32'hFFFD8052 , 32'hFFFFD628 , 32'h0000705A , 32'hFFFFCD54 , 32'hFFFFE616 , 32'h000082DD , 32'h000026DB , 32'hFFFF75F9 , 32'hFFFDF057 , 32'h00005940 , 32'h00020FDB , 32'hFFFF9759 , 32'hFFFE62B2 , 32'hFFFF2FA1 , 32'h00000892 , 32'hFFFD38EC , 32'hFFFEB6FC , 32'h0000E42A , 32'hFFFEA987 , 32'hFFFE6DE1 , 32'h00027BBD , 32'h0002508B , 32'hFFFEE576 , 32'hFFFD1CD8 , 32'h0000391F , 32'hFFFD6422 , 32'h00003259 , 32'hFFFF6170 , 32'hFFFFFEA1 , 32'h00006F37 , 32'h00009A8E , 32'hFFFD1B8F , 32'h000026AE , 32'h00013833 , 32'hFFFFB4BC , 32'h00009312 , 32'h0000EDE6 , 32'h000116CE , 32'hFFFFC322 , 32'h000201B8 , 32'hFFFFACD1 , 32'hFFFE857F , 32'h00002AB8 , 32'hFFFD9663 , 32'h0002A19E , 32'hFFFDBC80 , 32'h000050AA , 32'h00008A9C , 32'hFFFEC6C5 , 32'h00016E60 , 32'h00002C40 , 32'hFFFE71C3 , 32'h00013B97 , 32'h0000CB7C , 32'hFFFF44E3 , 32'hFFFF6039 , 32'h0000BBD6 , 32'h0000AB8D , 32'h00017264 , 32'hFFFD810E , 32'hFFFE8DB2 , 32'hFFFF29FC , 32'h00012846 , 32'hFFFFF71C , 32'hFFFCE33F , 32'h0000098E , 32'h00007976 , 32'h0000BFE5 , 32'h00007F97 , 32'h000109EE , 32'h0000E0C3 , 32'hFFFD185A , 32'h0000FA6E , 32'hFFFFCDA3 , 32'h0001282C , 32'hFFFE0BA8 , 32'h000063F9 , 32'hFFFED357 , 32'h00016E0C , 32'h0000ABC8 , 32'hFFFCA5D0 , 32'h00072E62 , 32'h000227B8 , 32'hFFFD7B38 , 32'hFFFDCDDC , 32'hFFFF6908 , 32'hFFFD0034 , 32'hFFFFF573 , 32'hFFFD9FAF} , 
{32'hFFFC7412 , 32'hFFFC3A70 , 32'h00008CF8 , 32'h00009B9F , 32'hFFFF3C23 , 32'hFFFF6F1D , 32'hFFFF4C25 , 32'hFFFF116C , 32'hFFFF3613 , 32'hFFFED158 , 32'hFFFBE08B , 32'hFFFB9542 , 32'h00003205 , 32'hFFFA12C7 , 32'hFFFD5AA1 , 32'hFFFE6645 , 32'h0001FD16 , 32'h00014FF6 , 32'hFFFEB109 , 32'hFFFB89EA , 32'h00026360 , 32'hFFFD63C7 , 32'hFFFF2261 , 32'hFFFE5B1A , 32'hFFFFF5F4 , 32'hFFFBBAB8 , 32'h0001FDA2 , 32'h0001D143 , 32'h0001CE7E , 32'hFFFF6FF2 , 32'hFFFD40FB , 32'h00035EFE , 32'h0001D841 , 32'hFFFEED37 , 32'h00029D54 , 32'hFFFEE593 , 32'hFFFFC1E3 , 32'h00054E20 , 32'hFFFE1A5E , 32'hFFFE9A88 , 32'hFFFEB465 , 32'h00044857 , 32'h0001D329 , 32'hFFFE4A59 , 32'h0005AE1E , 32'h00007306 , 32'hFFFFA9D3 , 32'h00023C62 , 32'h0002B3C2 , 32'hFFFE4D1B , 32'h0000E784 , 32'h00014E09 , 32'hFFFBDF5A , 32'h000245BC , 32'h0002CDDD , 32'h0005848D , 32'hFFFDE494 , 32'hFFFAFE0F , 32'hFFFCB852 , 32'hFFFB419C , 32'hFFFD4B07 , 32'h00030EAA , 32'h0002002B , 32'h0003632D , 32'hFFFD1EF4 , 32'hFFFB882B , 32'hFFFEF952 , 32'hFFFEC4C3 , 32'h0001AE0F , 32'h0003D9C4 , 32'hFFFEB035 , 32'h00001DE5 , 32'h0004DF30 , 32'h00003B39 , 32'hFFFB8001 , 32'h00013B65 , 32'hFFFE88AD , 32'hFFF5EE3F , 32'hFFFF21D0 , 32'h0003E7CC , 32'h0000BC14 , 32'hFFFF1C44 , 32'h00036088 , 32'hFFFE5BCC , 32'h0002D182 , 32'h00033D78 , 32'h00054171 , 32'hFFFD3E4B , 32'hFFFBB105 , 32'h0001A72A , 32'hFFFEE600 , 32'h0000E8E0 , 32'hFFFC9F24 , 32'hFFFF72BE , 32'hFFFD7549 , 32'hFFFE8C63 , 32'hFFFEAC86 , 32'hFFFE8EB1 , 32'h0000DA1D , 32'h00004A9A} , 
{32'hEDAA8780 , 32'h0400D9C0 , 32'hFD25BA70 , 32'hF5177360 , 32'hE3196D20 , 32'hFD580E64 , 32'h1969B1A0 , 32'hF40085D0 , 32'h10DDA7E0 , 32'h04A01878 , 32'hF5273F50 , 32'h13460940 , 32'hEDF50100 , 32'h0D89F6B0 , 32'h08E9F450 , 32'hF1B278A0 , 32'h065A8B98 , 32'hF4A8DD20 , 32'hF2807980 , 32'hFD87E624 , 32'h091C4550 , 32'hEE87CC60 , 32'h095EAEB0 , 32'hE82012E0 , 32'hF7BCD7E0 , 32'h06A9A8B8 , 32'h00057022 , 32'h02FF2510 , 32'h02072A10 , 32'h08318260 , 32'hF36AF410 , 32'h1073CD20 , 32'hF014A620 , 32'hDD846740 , 32'h004C764A , 32'hF9708428 , 32'hFB544F40 , 32'h0CC8ADA0 , 32'h03673C40 , 32'hFC4A30F4 , 32'h08D3E5C0 , 32'hF133CE00 , 32'h02F2A10C , 32'h007E885A , 32'h04BBA9B0 , 32'hFC3A1C9C , 32'h01C88FB8 , 32'hFEB29D3C , 32'h06AB3DC8 , 32'hFFB4F2A8 , 32'h0FC21F70 , 32'hFCB5F1F4 , 32'hFC6A0040 , 32'hF5B0B030 , 32'hF7EB74B0 , 32'hFED328A4 , 32'hFD4B061C , 32'hF9BFF968 , 32'h056CEC78 , 32'h09A3B700 , 32'hFFFF018B , 32'hFB523C80 , 32'h02B62A74 , 32'h08C70ED0 , 32'h00DE9D22 , 32'h02DE7574 , 32'hFB715328 , 32'hFB590B78 , 32'hF8171850 , 32'hFC338DB4 , 32'hFABBB688 , 32'h02EA04BC , 32'h017BF860 , 32'hFA2FFDF8 , 32'hFF300708 , 32'h04675D50 , 32'h000BD91B , 32'hFE3FD4D8 , 32'h025525CC , 32'h00764183 , 32'hFFCB2159 , 32'h0385FD20 , 32'h01AC50AC , 32'hFF9EEB36 , 32'h02DCB150 , 32'hFEF1F6D8 , 32'h002D6B97 , 32'hFFF5EEC0 , 32'h02B8CFF4 , 32'h005CE7B0 , 32'hFFFE1595 , 32'hFFFF2441 , 32'h00009984 , 32'hFFFF85D6 , 32'h000212CF , 32'hFFFF383D , 32'h00039551 , 32'h00020C1F , 32'hFFFE0FB5 , 32'hFFFE04CD} , 
{32'hFBBF9900 , 32'h201CBC00 , 32'hE92A0E00 , 32'hFA72AF40 , 32'hE2602F20 , 32'h195111C0 , 32'h07E0D6B0 , 32'hC638D480 , 32'h2BA8E800 , 32'h0597D6B8 , 32'hEE5519E0 , 32'hFD4CE7AC , 32'h1BD26780 , 32'hF9033C58 , 32'h096402C0 , 32'hFFF801E9 , 32'h06D69EC0 , 32'h21D53D80 , 32'hEA8BB5A0 , 32'hF6A38AB0 , 32'h0E11D1A0 , 32'hF1402070 , 32'hEA532BA0 , 32'h0C6DF430 , 32'hE4A3AF80 , 32'hF1471F20 , 32'h02B31594 , 32'h05099B80 , 32'hE85D5620 , 32'h0148A1C4 , 32'h01F6BF4C , 32'h228BFE00 , 32'hF66C5460 , 32'h0C2BB3D0 , 32'h000C0C5D , 32'hFAD41EC0 , 32'h16A88A80 , 32'h024BDA74 , 32'h0312E164 , 32'hE835B060 , 32'hFC21F7E4 , 32'hFAD4C5C0 , 32'h04564E78 , 32'hFF0E404F , 32'hFBC02FA0 , 32'hF7C6D090 , 32'hF5BFC790 , 32'h11353340 , 32'hF4E19AB0 , 32'h015C0630 , 32'hF5F8BC10 , 32'h01260B00 , 32'h02887204 , 32'hFB362650 , 32'h01713DB0 , 32'h08774580 , 32'hF0F199F0 , 32'hF0F07DB0 , 32'hF95D3B20 , 32'hF2F23E10 , 32'h028EFB14 , 32'h088DB000 , 32'hFB43A7A0 , 32'hFF0A13E3 , 32'hFF87043A , 32'h034F4C84 , 32'h05223FD0 , 32'hFBBF8460 , 32'hFDE0BF68 , 32'h02357D74 , 32'h026294B0 , 32'h0007C924 , 32'h00A84E7B , 32'h01A5D088 , 32'hFF8B1A86 , 32'hFB5EAC70 , 32'hFD098AAC , 32'hFC58AFE4 , 32'hFE0317D8 , 32'hFF9FF87E , 32'h017DEDF8 , 32'h03FFBAE8 , 32'hFDAE2388 , 32'h019C553C , 32'hFE0C0200 , 32'h024367A8 , 32'hFFE35932 , 32'h02FC72D4 , 32'hFF697167 , 32'h009E75C2 , 32'hFFFF927A , 32'h00021DBA , 32'h0000FBA9 , 32'hFFFFDC15 , 32'hFFFFF6D3 , 32'hFFFE757D , 32'h00007EF7 , 32'h00004DCB , 32'h00008885 , 32'hFFFEEF7D} , 
{32'hFFFF833E , 32'h000187BA , 32'hFFFE2E78 , 32'hFFFC8DEB , 32'h00035C59 , 32'h000097FE , 32'h0003AE56 , 32'hFFFC59F7 , 32'hFFFE036F , 32'h0001D7BB , 32'h0003496E , 32'h0000FEC2 , 32'hFFFBF633 , 32'h0000C233 , 32'hFFFDAAEB , 32'h00003624 , 32'h000134C4 , 32'h0001B3C2 , 32'hFFFF65EA , 32'hFFFDAD0A , 32'h0002636F , 32'h000137EB , 32'hFFFEBAF2 , 32'h0003C38E , 32'hFFFCAF1D , 32'h000045D4 , 32'h0001A245 , 32'hFFFFFBAB , 32'hFFFD258C , 32'h00030F96 , 32'hFFFEE203 , 32'hFFFCBDC9 , 32'h00016E4A , 32'h00022A71 , 32'h0001AB5B , 32'hFFFC00E3 , 32'h00029D7B , 32'h0001AAB6 , 32'hFFFE4E7D , 32'h0001676F , 32'h000263FE , 32'h0000A68B , 32'hFFFF7456 , 32'hFFFEFD7E , 32'h0001B3D1 , 32'h0001C003 , 32'hFFFEBCBA , 32'h00051620 , 32'h0001CEED , 32'hFFFF9CCE , 32'h00004C3F , 32'hFFFF34E0 , 32'h00034AE4 , 32'h0002708C , 32'h00033E60 , 32'h0001813F , 32'h0000682F , 32'hFFFC4E6A , 32'h000072A8 , 32'hFFFD255A , 32'h0001FE93 , 32'hFFFF03DC , 32'hFFFFEF09 , 32'hFFFE2B21 , 32'hFFFA6EFE , 32'hFFFAA278 , 32'hFFFD8DE4 , 32'h0000EF51 , 32'hFFFBF787 , 32'hFFFED574 , 32'h000078CF , 32'hFFFF22EC , 32'h00042EFA , 32'hFFFA0016 , 32'hFFFD1AC9 , 32'h0002B4CB , 32'h00019DD2 , 32'hFFFACC4F , 32'hFFFDDD8D , 32'h0003470E , 32'h00045C2E , 32'hFFFDA7E5 , 32'hFFFE6078 , 32'hFFFC001B , 32'h00023B65 , 32'h00014CB0 , 32'hFFFB0030 , 32'hFFFF534E , 32'hFFFEB1B3 , 32'hFFFE7F43 , 32'h000107E7 , 32'hFFFEFB51 , 32'hFFFEAFDF , 32'hFFFA59BD , 32'h0004FE8A , 32'hFFFF3705 , 32'h00023C75 , 32'h00007B11 , 32'hFFFF38D5 , 32'hFFFE7EC5} , 
{32'hC0AF1180 , 32'h09E21AE0 , 32'h2D068440 , 32'h2F9E4E40 , 32'h3C835880 , 32'hD89E4000 , 32'h05C75690 , 32'hFD71CF3C , 32'h06B63BC0 , 32'h03B8272C , 32'h34088BC0 , 32'h245D0940 , 32'hF9976258 , 32'h0F8CC490 , 32'h024B0A68 , 32'h0872F5E0 , 32'h1910D940 , 32'hF1F94BB0 , 32'h0875B2D0 , 32'h20AC9F00 , 32'hE2301D40 , 32'hF9EBA248 , 32'hFA4A9F00 , 32'hFA163290 , 32'hEFCE2860 , 32'h0A4C20B0 , 32'hF7F86EE0 , 32'h00F3F0C5 , 32'hFFABC351 , 32'h04990B90 , 32'hE9E336A0 , 32'h14F48C00 , 32'h04564FD8 , 32'hF9C93658 , 32'hFAC0C958 , 32'h0BB99E30 , 32'h0554A258 , 32'h0C034520 , 32'hF2BFAC10 , 32'h07F3A1E0 , 32'h035EC33C , 32'hFB8BAC10 , 32'hF7964390 , 32'hF8DD44F0 , 32'hF726EFA0 , 32'h077F2738 , 32'hF55F7DB0 , 32'hFBBE54B0 , 32'h01FA14C8 , 32'h038FAA98 , 32'h076FE170 , 32'h03E05F44 , 32'hFA8AB680 , 32'h0383A880 , 32'h01BC81E4 , 32'hFD2DD564 , 32'h0103DFB8 , 32'hF5C34600 , 32'hFEAB724C , 32'hF7F66860 , 32'h030321E4 , 32'h0372DFB4 , 32'hEFC90660 , 32'hFE5D7CE8 , 32'h06E4B408 , 32'hFB13A370 , 32'hFBF299D0 , 32'h03BD90C8 , 32'hFCE7358C , 32'hFBA458B8 , 32'h0138555C , 32'hFE3C288C , 32'hFBB65750 , 32'hFFBE62ED , 32'hFDE56884 , 32'h01CCBDA8 , 32'h03BC50B4 , 32'h00B074E7 , 32'h02ADCB1C , 32'h03244DB8 , 32'h02A2A43C , 32'h0267F2FC , 32'h02EFE758 , 32'hFD813904 , 32'h0092AB71 , 32'h03653BF4 , 32'hFE4E2CDC , 32'h0106E78C , 32'hFD67A5F8 , 32'h00ADED61 , 32'hFFFE1188 , 32'hFFFFC4B8 , 32'h0000797D , 32'h00011AC2 , 32'h000043DA , 32'h0002685E , 32'h00006372 , 32'hFFFFA300 , 32'hFFFF42EE , 32'hFFFF336C} , 
{32'h0003DE90 , 32'h00027B8B , 32'hFFFE03AA , 32'hFFFEB947 , 32'h00004A2C , 32'h000242DB , 32'hFFFE8034 , 32'hFFFDF746 , 32'h00001CE0 , 32'hFFFDEAB3 , 32'h0003E193 , 32'hFFFE0043 , 32'h000001BB , 32'hFFFEDF6B , 32'hFFFED6B7 , 32'h0002D08D , 32'h000004A5 , 32'h0002AC64 , 32'h00021AD7 , 32'hFFFB1BDD , 32'h00002745 , 32'h000172FA , 32'h00008EDD , 32'hFFFD299A , 32'hFFFDE63A , 32'hFFFCE56A , 32'h00034185 , 32'h0003333D , 32'h0001961B , 32'h00023C5E , 32'h0001823C , 32'hFFFF4450 , 32'hFFFBDACB , 32'hFFFEBA97 , 32'h000008FF , 32'h0001A60B , 32'hFFFC258B , 32'h0001BEC7 , 32'h00019449 , 32'hFFFC4505 , 32'h0004338F , 32'h0000C164 , 32'hFFFAF8F3 , 32'h0000B2EE , 32'hFFFE4A43 , 32'h00002174 , 32'hFFFDC012 , 32'h00000F89 , 32'hFFFE4B1C , 32'h00025538 , 32'h00030F33 , 32'hFFFF770D , 32'hFFFAAB2E , 32'h0003CB54 , 32'h00035CDB , 32'h0000629E , 32'h00004AEF , 32'hFFFD3E86 , 32'hFFFB22C6 , 32'h0001AF67 , 32'hFFFF2ECF , 32'hFFFD0135 , 32'h0005D2C0 , 32'hFFFF0E25 , 32'hFFFCF2CD , 32'h000459AB , 32'h000189B8 , 32'h00028262 , 32'hFFFE5615 , 32'h0006095E , 32'hFFFE6A62 , 32'h00003846 , 32'hFFFE8B5F , 32'h0001F397 , 32'hFFFFCC14 , 32'hFFFEFFFE , 32'h00004710 , 32'hFFFF7609 , 32'hFFFA4CB3 , 32'h00005D7D , 32'hFFFE24E4 , 32'h000376E9 , 32'hFFFBDE14 , 32'h00004D5A , 32'hFFFEF6D5 , 32'hFFFF0649 , 32'hFFFA9428 , 32'h0000AF9B , 32'hFFFBE4C8 , 32'h0002663B , 32'h0005F053 , 32'h000134BF , 32'h0002FF10 , 32'h00060CC6 , 32'hFFFE7604 , 32'h00018A0F , 32'hFFFF44C2 , 32'h0001F32E , 32'h0003D722 , 32'h0001416F} , 
{32'hFFFDB31A , 32'h00005AAE , 32'hFFFB0F4B , 32'hFFFFB3BF , 32'h00005FD1 , 32'hFFFC58F0 , 32'hFFFE34BC , 32'hFFFCC0E1 , 32'hFFFD3D25 , 32'h0000D8BA , 32'hFFFBDB2B , 32'hFFFD9BD1 , 32'hFFFEF167 , 32'h0000A002 , 32'hFFFF5A3A , 32'hFFFFAF45 , 32'h0001C1A3 , 32'hFFFBD3E7 , 32'hFFFE4891 , 32'hFFFC2276 , 32'h0004A412 , 32'h00033152 , 32'h0001231E , 32'hFFFCB062 , 32'hFFFFFE82 , 32'hFFFFD0AF , 32'h0000E7AF , 32'h00010087 , 32'h0001D7A3 , 32'hFFFF8CA2 , 32'hFFFD7F7D , 32'h000285AB , 32'hFFFEC73C , 32'hFFFC80F7 , 32'h0002C45D , 32'hFFFF1C8A , 32'h0000F6B9 , 32'h00013E75 , 32'hFFFE3D88 , 32'hFFFE964F , 32'h000116EF , 32'hFFFE958F , 32'h00002C88 , 32'h0000CEC6 , 32'h00060F3D , 32'hFFFD3A26 , 32'hFFFD6FA2 , 32'h0000D80B , 32'hFFFE50A3 , 32'hFFFF483A , 32'hFFFE7D3A , 32'hFFFF3EB6 , 32'h000320B4 , 32'h000019F1 , 32'hFFFEC0CE , 32'hFFFD937E , 32'h00006708 , 32'h000172A3 , 32'hFFFF0C07 , 32'h00008DFA , 32'hFFFE90FC , 32'h0001A276 , 32'hFFFE7E1C , 32'h0002EB5B , 32'hFFFD982B , 32'h0001CB46 , 32'hFFFED893 , 32'hFFFFE405 , 32'hFFFF4F4C , 32'hFFFF3CEE , 32'hFFFD7FC4 , 32'h0000F640 , 32'hFFFF34C6 , 32'h00041E21 , 32'h0005582A , 32'hFFFC8C7D , 32'hFFFEAC4A , 32'h000223E8 , 32'hFFFE3FA3 , 32'h000111C3 , 32'h0002E8D4 , 32'hFFFECB24 , 32'hFFFC21C1 , 32'h00036934 , 32'hFFFCF265 , 32'h0000A83E , 32'h0000913F , 32'h000123CA , 32'h000097FC , 32'h000076C8 , 32'h00073E13 , 32'h00013E5C , 32'h0002782A , 32'h0004FE2B , 32'h00025B93 , 32'h00028DCC , 32'h0000DC97 , 32'h0002C966 , 32'h0000BE46 , 32'h000100C6} , 
{32'hEC789540 , 32'h29A1CD00 , 32'hEF803F40 , 32'h07D83328 , 32'h07811080 , 32'h22FD8040 , 32'h1B5F7720 , 32'h1556DA20 , 32'h0ED58C80 , 32'h05AFC4F8 , 32'hF2BB5970 , 32'hF275D890 , 32'hE9FFD9C0 , 32'h1014AD80 , 32'hF32B9280 , 32'h316ACF80 , 32'hF28CBCB0 , 32'h0A8C3C20 , 32'hFF9D7169 , 32'hE874F380 , 32'h0E5720B0 , 32'hED725220 , 32'hF4704CC0 , 32'h01697190 , 32'hF4C3CCF0 , 32'hEFB6F480 , 32'hF4B42500 , 32'h1393DAA0 , 32'hF73797D0 , 32'hFF066D7B , 32'h0D99AB40 , 32'h0B7EF5C0 , 32'h14D19F40 , 32'hF5F14690 , 32'h196EE720 , 32'hF4FF5FF0 , 32'hF9630498 , 32'hFD322400 , 32'hFFDB6385 , 32'hFFD78ABC , 32'h03038CD8 , 32'h043ECF90 , 32'hF38C3340 , 32'hF7149C00 , 32'hF8627CD8 , 32'h0A4FD460 , 32'hF42B6BF0 , 32'hFC096130 , 32'h07B93D40 , 32'hFF8B1AEC , 32'h113FA3C0 , 32'hFF3FEF26 , 32'h02A4AC54 , 32'hF3F321D0 , 32'hF9562968 , 32'hFDAC7638 , 32'h043C5438 , 32'h01B1E504 , 32'h02A9AB58 , 32'hFFBE103E , 32'h043DCD50 , 32'h063338C8 , 32'hFFD2BF95 , 32'hFE06D26C , 32'h03627758 , 32'h0357654C , 32'hFC30D9E0 , 32'h0227C4A8 , 32'h07D9FDD8 , 32'h01666624 , 32'hFEF91BFC , 32'h0357A38C , 32'h06433EF0 , 32'h04922B30 , 32'hFED49358 , 32'h00676C8C , 32'h059C5488 , 32'hFF0B5D55 , 32'h011E502C , 32'hFBCA5C48 , 32'hFBFB6080 , 32'hFA4EDCD8 , 32'h0344372C , 32'hFE59CA30 , 32'hFD33FA10 , 32'h025DE188 , 32'h00D1F92B , 32'h004CF203 , 32'h00A145CF , 32'hFFDD7FC9 , 32'h0000E9D2 , 32'hFFFF9CF5 , 32'hFFFEC7E7 , 32'h000178BB , 32'hFFFE5057 , 32'hFFFF1DDD , 32'hFFFEF688 , 32'hFFFF56DD , 32'hFFFEF2F6 , 32'h000018D1} , 
{32'h1098D020 , 32'hF3309440 , 32'h05622088 , 32'hF3C56AF0 , 32'h09CCEC40 , 32'hFCD12254 , 32'hF5F27CD0 , 32'h0C3D99C0 , 32'hFC982278 , 32'hFE03790C , 32'hFBD8CC98 , 32'hEF496DE0 , 32'hF16BAAC0 , 32'hFF542E19 , 32'hF6820FB0 , 32'h0037E0FF , 32'h00C89FA1 , 32'h072D3250 , 32'hFB6A44B0 , 32'h037AF4D4 , 32'h0396ED0C , 32'hFECC1814 , 32'hFFEB58A5 , 32'hFE818410 , 32'hFF1FA8CF , 32'hF6568450 , 32'h0171345C , 32'h0F9D23D0 , 32'hFBAAA970 , 32'hF8C17D40 , 32'h00C6FA5D , 32'h0345AF6C , 32'hFBC2AAA0 , 32'hFF0A71C1 , 32'hF8BD2258 , 32'hFBA7DD88 , 32'h0C01B490 , 32'hFF7666E4 , 32'h050E1058 , 32'hFCE75558 , 32'h03146F3C , 32'h00803D80 , 32'hF9D24C28 , 32'hFF0DD6FD , 32'h03CD61F0 , 32'hFD6C1C6C , 32'hF6F38760 , 32'hF711AE00 , 32'h01D7FE60 , 32'h081E33B0 , 32'hFCFF0CB8 , 32'hF7E4C850 , 32'hF8B2D3C0 , 32'h00F87714 , 32'hFB6D8720 , 32'hFD7FC8AC , 32'hFAC26388 , 32'hFE53A99C , 32'h0CF9C910 , 32'h07A7EC70 , 32'h02E78B70 , 32'hF96D0330 , 32'h002BCDAF , 32'h018146DC , 32'hFFD4C22E , 32'h0946F850 , 32'hFE45DA8C , 32'hFDF0BE54 , 32'h04B8BE70 , 32'hFF1AE7F7 , 32'h063C6B80 , 32'hF3F3D340 , 32'h01B7C5D4 , 32'hFB05CD40 , 32'h07E68328 , 32'h04F6E090 , 32'h03F7A410 , 32'hFF138638 , 32'hFC61681C , 32'h0173B5B8 , 32'h016C9FF4 , 32'hFF15BEA3 , 32'h02679904 , 32'h031F6B24 , 32'h0460F038 , 32'hFDCEC944 , 32'hFFB0F46B , 32'h023CA474 , 32'hFEC7E780 , 32'h002B4019 , 32'h0002D2BB , 32'h000276BD , 32'hFFFD8762 , 32'hFFFFCCBB , 32'hFFFE94F7 , 32'h000169A4 , 32'h00003F0F , 32'hFFFE0FF9 , 32'hFFFFEA20 , 32'h000051AC} , 
{32'hFE2D95F8 , 32'h00319C4A , 32'hF781ECE0 , 32'hFF029AD7 , 32'hFA43DF20 , 32'hFEAB6F1C , 32'h0B4D14A0 , 32'h002019EB , 32'h01DC46C0 , 32'hFDA70A84 , 32'h038C5228 , 32'h03A1BCBC , 32'hFD5CB86C , 32'h081C3F70 , 32'hF74BC0B0 , 32'h05C460C8 , 32'h00C58DD1 , 32'h0AC39050 , 32'h0237D240 , 32'hFE6895BC , 32'hFDADE678 , 32'hF526A2A0 , 32'hFCF800F8 , 32'h03FA8ACC , 32'h072F6FE0 , 32'hFF70D5BA , 32'h05B1B748 , 32'h05848630 , 32'hFB116C70 , 32'hFCD12EB8 , 32'h00562036 , 32'h03C0BAC4 , 32'hFBDA9EA0 , 32'hFAF7B1F8 , 32'hFB458160 , 32'hF6B349B0 , 32'h040E8680 , 32'h072789B0 , 32'hFAD48A98 , 32'hF6698700 , 32'hFAADA8E8 , 32'hF9D780A0 , 32'h007D7EA3 , 32'h06008CB0 , 32'h07696528 , 32'hFA8B47D0 , 32'hF6B47250 , 32'h0039F78C , 32'h06075D88 , 32'h04796170 , 32'h030DE5B8 , 32'h028FF7A0 , 32'hFAF6EE60 , 32'hFF96F8AC , 32'h069C8DA8 , 32'hFA445128 , 32'hFF2C5039 , 32'hFBB9AC50 , 32'hFB1D56C8 , 32'h02C56CE8 , 32'hFA8DE208 , 32'h03F5093C , 32'h0753E1A0 , 32'h0265C440 , 32'h002F0C4A , 32'h06284A10 , 32'h025E2FDC , 32'h07B35F90 , 32'hFB39E628 , 32'h06213B00 , 32'hFD745454 , 32'hFAB38E18 , 32'hF824B1F0 , 32'h0106E768 , 32'hFD10E2A0 , 32'h04D79908 , 32'hFB9F92E0 , 32'hFB69C450 , 32'hFB53CF40 , 32'h01191314 , 32'hF7CF7200 , 32'hFFCEAC0C , 32'hFE3C2518 , 32'hFFD66DA3 , 32'hFA86C860 , 32'hFEB76830 , 32'h0030B985 , 32'hFDD098A0 , 32'h00382059 , 32'h0112F0D0 , 32'h00005EF9 , 32'h000036BB , 32'hFFFCFF3D , 32'h0003B78A , 32'h000054E3 , 32'h0000D3C6 , 32'hFFFFC938 , 32'hFFFED1D0 , 32'h0000BC32 , 32'hFFFF1BC5} , 
{32'hFFF8BFB1 , 32'h0000ABA4 , 32'hFFFE8192 , 32'hFFFEED0F , 32'hFFF895A9 , 32'h0003AED1 , 32'h0004F0E6 , 32'h00003EEE , 32'h00043836 , 32'hFFF9CB0A , 32'hFFFF359D , 32'h0001DDB4 , 32'hFFFDD995 , 32'h0002AF47 , 32'hFFFFCFD2 , 32'hFFFF74F8 , 32'hFFFF3C9C , 32'hFFFB5A1A , 32'hFFFD4284 , 32'hFFFEB8F5 , 32'hFFFF492F , 32'hFFFF1D7B , 32'h00005B2A , 32'h000301CA , 32'hFFFE99D1 , 32'h00014180 , 32'h0004C69F , 32'hFFFF3168 , 32'h00003444 , 32'hFFFE6777 , 32'hFFFEBD93 , 32'hFFFF2437 , 32'hFFFBC678 , 32'hFFFE4E3D , 32'h0000D0BE , 32'h000093FA , 32'h000064AA , 32'hFFFA5A93 , 32'h0002E10A , 32'hFFFCFE55 , 32'hFFFD025A , 32'h00021693 , 32'h00003C8C , 32'h0001D18F , 32'hFFFA356E , 32'hFFFC9EE9 , 32'hFFFF6C45 , 32'hFFFD1890 , 32'hFFFC6529 , 32'h0001135F , 32'h00023BB6 , 32'hFFFC8C9C , 32'hFFFE72CA , 32'h0002C032 , 32'hFFFE2438 , 32'hFFFD0870 , 32'hFFFFE1AB , 32'hFFFDB413 , 32'h00005D68 , 32'hFFFF906E , 32'hFFFE9290 , 32'hFFFC97DC , 32'hFFFD4845 , 32'hFFF886B9 , 32'hFFFE9DA8 , 32'h000606B1 , 32'hFFFFFFF2 , 32'hFFFA488E , 32'hFFFDE4D9 , 32'hFFFE8759 , 32'hFFFE27D1 , 32'hFFFFB073 , 32'h00035F33 , 32'h0003AEAB , 32'hFFFF3A3F , 32'h0001E29E , 32'h00075D60 , 32'h0000B251 , 32'h00027AC2 , 32'h00053464 , 32'h00063FA7 , 32'hFFFF08C0 , 32'h0001B3B4 , 32'h00000970 , 32'h0001FA07 , 32'h0007482C , 32'h0001E6D4 , 32'hFFFB406B , 32'h0003B5FB , 32'h000357BE , 32'h0001A6AC , 32'h00017D63 , 32'h0000186E , 32'hFFFA3908 , 32'h00081AAD , 32'hFFFF072B , 32'h00013767 , 32'h00002274 , 32'h00004DE1 , 32'h0000EC19} , 
{32'h09D049D0 , 32'h08606840 , 32'h137E2FA0 , 32'hF712FB60 , 32'h30843940 , 32'h12CBF7C0 , 32'hE71D9240 , 32'h11F89360 , 32'hEF6DC8A0 , 32'hFA6F9828 , 32'hF938A2F8 , 32'hF8181FE8 , 32'hFAFEB0F8 , 32'h07F0DFB8 , 32'h183D1E60 , 32'hFAD9A358 , 32'hFD2514A8 , 32'h02517CC8 , 32'hFD99C6E4 , 32'h0A96F380 , 32'h0E8FD360 , 32'hED092A60 , 32'hFB964EA0 , 32'hED4674E0 , 32'h01D69F2C , 32'h10234520 , 32'hF33A5B10 , 32'h14D27100 , 32'hFC87280C , 32'hFA158BC0 , 32'hFA38CA28 , 32'h00EEA53E , 32'h05488200 , 32'hF9291188 , 32'hF529B1A0 , 32'hF6F674F0 , 32'hF74CC4E0 , 32'hF71D8720 , 32'h005FEAFD , 32'hF89BD8D8 , 32'h0BC664B0 , 32'hED842140 , 32'hFD990038 , 32'hFB2F2050 , 32'h0B3EC2A0 , 32'h073BDAA8 , 32'hF9A73798 , 32'h03E6E9B0 , 32'h105B2920 , 32'h03A667A8 , 32'hF7912C10 , 32'h0A05B2D0 , 32'hF20D51D0 , 32'hFFC1B12E , 32'hFF8CE1BE , 32'hFA7F4B28 , 32'hFFA49C54 , 32'hFEE10214 , 32'h01E9231C , 32'hF832E4C8 , 32'h0B45A9A0 , 32'h011D6B00 , 32'hFA693C38 , 32'hFA21E810 , 32'hFC49587C , 32'h01C76558 , 32'h0DF8B280 , 32'h04020B28 , 32'h0302DC08 , 32'h00F0D988 , 32'hFD28B6B0 , 32'hFFA7B985 , 32'hF8067E18 , 32'h01C0EC8C , 32'hF9718B00 , 32'h01B2DFBC , 32'hFC5D67E0 , 32'h034D4D3C , 32'hFD0EB7C8 , 32'hF98C41B0 , 32'hFB13CB88 , 32'h05EC0BD8 , 32'hFD6567A4 , 32'hFCC56014 , 32'hFDFACCF0 , 32'hFFA27945 , 32'h01A42A44 , 32'h016BD690 , 32'h00B40928 , 32'hFF0C7A46 , 32'h00025D56 , 32'hFFFB8F50 , 32'hFFFF4CB4 , 32'hFFFC3145 , 32'h0001B192 , 32'hFFFEEB88 , 32'hFFFFAD9D , 32'hFFFFE2C5 , 32'h0000BBED , 32'h00007C6D} , 
{32'hFFFECE16 , 32'h00001CFD , 32'hFFFBEE2D , 32'h00044505 , 32'h00004155 , 32'hFFFEFDAC , 32'h00014A18 , 32'hFFFF88A5 , 32'hFFFFBAC0 , 32'h0004A7C5 , 32'hFFFEBE3F , 32'h00004CD7 , 32'h0006BD42 , 32'hFFFCD3ED , 32'h000091FA , 32'hFFFD5796 , 32'h00011FA9 , 32'h00004878 , 32'h0000D016 , 32'hFFFE044C , 32'hFFFFA009 , 32'hFFFC1792 , 32'hFFFEC679 , 32'h00018D4D , 32'h0001936E , 32'h000660E5 , 32'h00014844 , 32'h000409D6 , 32'hFFFAB7E1 , 32'hFFFDE212 , 32'hFFFC4656 , 32'hFFFFB653 , 32'h0000A717 , 32'h00051C30 , 32'hFFFFDD37 , 32'h0006F9B4 , 32'h0000DDC3 , 32'h0000EDD0 , 32'h00029E66 , 32'h0001B35D , 32'hFFFF5CE2 , 32'h0000D175 , 32'hFFFD188C , 32'hFFFD9DC2 , 32'h0002A6C8 , 32'h0001CDFB , 32'hFFFF3E70 , 32'h00012289 , 32'h0003908D , 32'hFFFC0E41 , 32'hFFFE329F , 32'h00017721 , 32'h0004DA16 , 32'hFFFDFDAA , 32'hFFFD6B01 , 32'hFFFFF2E6 , 32'hFFFF9D4A , 32'h0003649D , 32'h0002A7E7 , 32'hFFFEB197 , 32'h0000836A , 32'hFFFDCE17 , 32'h000045A9 , 32'hFFFF0D26 , 32'hFFFD2A33 , 32'hFFFF8F32 , 32'h00013141 , 32'h0000FCB1 , 32'h00009D61 , 32'hFFFC48F2 , 32'h000065A5 , 32'hFFFC790D , 32'hFFFDE605 , 32'h000246EF , 32'hFFFF9981 , 32'hFFFFD55D , 32'hFFFECB97 , 32'h00020906 , 32'hFFFF060D , 32'hFFFD2B06 , 32'h0004FD37 , 32'hFFFE78A6 , 32'hFFFD6566 , 32'hFFFD4552 , 32'h00009BA4 , 32'h0000C1FE , 32'h000181A9 , 32'hFFFC6CAD , 32'h0001855F , 32'h0000046A , 32'h00026802 , 32'h0000898E , 32'hFFFF1339 , 32'h000106D7 , 32'hFFFB8B3F , 32'h00023A80 , 32'h000090A0 , 32'h0000E5ED , 32'h0001EA47 , 32'hFFFFFDFC} , 
{32'h00045B90 , 32'hFFFE0F2F , 32'h00004490 , 32'h00008F2A , 32'hFFFDB75A , 32'h00019ED6 , 32'h00016FC2 , 32'h0004740E , 32'hFFFC5747 , 32'hFFFEF6A2 , 32'hFFFEFFD7 , 32'hFFFE51CC , 32'h0000967A , 32'hFFFD55B8 , 32'hFFFC5C05 , 32'hFFFEA996 , 32'h00014C59 , 32'h00038830 , 32'hFFFE9F86 , 32'h00019B3A , 32'hFFFBAA8D , 32'h00019D5F , 32'hFFFE6FF8 , 32'hFFFBA49C , 32'h0000281D , 32'h0000E473 , 32'h00049F70 , 32'h00017993 , 32'hFFFEEE21 , 32'hFFFD8A14 , 32'hFFFDADDC , 32'hFFFC2BF6 , 32'h000283FB , 32'hFFFFFEC4 , 32'h0000EF02 , 32'h00031AB9 , 32'h0002B042 , 32'h00049893 , 32'h0002E7AA , 32'h00013940 , 32'h00018D20 , 32'h00014E85 , 32'hFFFD366A , 32'hFFFECD91 , 32'h0000FAE7 , 32'h0000ADD8 , 32'hFFFF34C8 , 32'h00041DB2 , 32'h0000DD63 , 32'hFFFD29A0 , 32'h0002697D , 32'hFFFEF2A8 , 32'hFFFFEFDF , 32'h000016EE , 32'h0000AFFA , 32'hFFFC1920 , 32'hFFFF16E7 , 32'h00039B1A , 32'hFFFFE955 , 32'h0000A1B7 , 32'h0001E83F , 32'h00007F41 , 32'h00005B06 , 32'hFFFF6E56 , 32'hFFFBDDCF , 32'hFFFC56BE , 32'hFFFB82ED , 32'h00060A22 , 32'hFFFE5241 , 32'h00024982 , 32'h00005D73 , 32'h0002633A , 32'hFFFFF253 , 32'hFFFEA360 , 32'hFFFF3A6F , 32'hFFFE2EC4 , 32'hFFFFC494 , 32'h00001B6E , 32'h0004BD47 , 32'h0003C782 , 32'hFFFE0237 , 32'h0002486E , 32'hFFFF56CD , 32'h000066CF , 32'h000347E5 , 32'h0000B65E , 32'h00029BAC , 32'h000019A1 , 32'hFFFBAB79 , 32'h00034362 , 32'hFFFD83B1 , 32'h0000A62C , 32'hFFFE6797 , 32'h00021C2B , 32'h0006535A , 32'hFFFF7107 , 32'hFFFE0137 , 32'h00017E52 , 32'h000276EB , 32'hFFFE9129} , 
{32'hFC7F4778 , 32'h04994708 , 32'h045B8A98 , 32'h0E108720 , 32'h092B61F0 , 32'h007C02A8 , 32'h118CB4A0 , 32'hED8E0B60 , 32'h10317840 , 32'h10D28BC0 , 32'h0994F1F0 , 32'h051CC5E0 , 32'h12D18040 , 32'h0099D645 , 32'h00213070 , 32'hF6EDFC10 , 32'h01D17620 , 32'h09D32ED0 , 32'hFCA9A38C , 32'h01CAE6F8 , 32'h0DFE0FE0 , 32'hFA102998 , 32'h0B717810 , 32'h0A25EF70 , 32'hF6DBA130 , 32'hF8965F50 , 32'hF49AB110 , 32'hF7ADD630 , 32'hFBE91078 , 32'hFD562104 , 32'hFC1604A4 , 32'h067D76A8 , 32'h07C608B8 , 32'h09DAE990 , 32'hFE18B478 , 32'hFCB277AC , 32'h064B6278 , 32'hF6C61560 , 32'h06F8F2A0 , 32'h0B39D9A0 , 32'h020CF400 , 32'hFB008D18 , 32'h027F0D54 , 32'h037DCBE0 , 32'hFEE0E04C , 32'h10B45DA0 , 32'h050E3E80 , 32'h01920C1C , 32'h02B8EAD8 , 32'h02BD1664 , 32'h04E017E8 , 32'hFF840C3E , 32'hF9BDA250 , 32'h05CC1B90 , 32'h00F1E1EF , 32'h06279728 , 32'h12923800 , 32'h08131230 , 32'hEB540DC0 , 32'h03B884D0 , 32'h00FFE3B2 , 32'hF7CE4F30 , 32'hFD5B8D88 , 32'h04F1A428 , 32'h0168BF68 , 32'h001A0955 , 32'h01F04720 , 32'h059DA200 , 32'h04F834B0 , 32'hFA4F18E0 , 32'hFC52F924 , 32'hFE50036C , 32'h0355DC20 , 32'h042AAC60 , 32'h0161E71C , 32'h06EBF728 , 32'h00B90CF2 , 32'hFF1B185B , 32'hFF7DF2B0 , 32'hFF23217F , 32'h07CD9AF0 , 32'h00C57799 , 32'hFD077924 , 32'hFF6FA6CB , 32'hFFB02A96 , 32'h02353140 , 32'h014B8488 , 32'hFF20B82E , 32'h02511CF0 , 32'hFF932F43 , 32'hFFFC76B1 , 32'hFFFFAA9E , 32'hFFFD5C66 , 32'h0001F8A7 , 32'hFFFFD267 , 32'hFFFF746A , 32'hFFFD73EA , 32'hFFFE196A , 32'h00020985 , 32'h0001C5B5} , 
{32'h00018564 , 32'h0000386B , 32'hFFFDC717 , 32'hFFFF0DDD , 32'h000308F8 , 32'h00008CC1 , 32'h0000F3D1 , 32'h00042E44 , 32'h000358FB , 32'hFFFF43D2 , 32'hFFFF3D20 , 32'h00046DD3 , 32'h000199DC , 32'hFFFD9DAB , 32'hFFFFE361 , 32'hFFFDDFF1 , 32'h0001B94C , 32'h0001B134 , 32'h000068A0 , 32'h00017EE1 , 32'hFFFE9F68 , 32'h00016550 , 32'h00007D4E , 32'hFFFDACBF , 32'hFFFE4831 , 32'h0003C169 , 32'h0002B519 , 32'hFFFE46EB , 32'h000069BA , 32'hFFFDD26E , 32'hFFFD9A2F , 32'h0001B7AF , 32'h000039E4 , 32'h00013496 , 32'h00013422 , 32'hFFFB00AB , 32'h0003B67A , 32'h00013315 , 32'hFFFF32D9 , 32'hFFFF26D9 , 32'hFFFD441D , 32'hFFFBE431 , 32'h0001ED63 , 32'hFFFFA55F , 32'hFFFF936A , 32'h0002A5F0 , 32'hFFFD62F8 , 32'hFFFEEEFD , 32'h00007A54 , 32'hFFFF09C7 , 32'hFFFD0FC2 , 32'h0002AA8C , 32'h0000AD88 , 32'hFFFF60CE , 32'hFFFF5165 , 32'hFFFA871A , 32'hFFFDF350 , 32'h00049A6E , 32'h00055B4F , 32'hFFFE1C2E , 32'hFFFD48E3 , 32'h0002C567 , 32'h0001A627 , 32'h0001FA48 , 32'h00017F49 , 32'h000464AA , 32'h000039C1 , 32'hFFFEC029 , 32'h000074DE , 32'h0002F38C , 32'hFFFE91B7 , 32'h0003086D , 32'h00024E35 , 32'hFFFF71E6 , 32'h0005947B , 32'h00026777 , 32'hFFFC2ACE , 32'h00025147 , 32'h00035E6C , 32'h00006B5D , 32'h0001D1A9 , 32'h0000CE4A , 32'hFFFC34D1 , 32'hFFFE5F5B , 32'hFFFDE989 , 32'hFFFEDE3E , 32'hFFFF4123 , 32'hFFFEA327 , 32'h0004179B , 32'h0004470D , 32'h0004A9D9 , 32'hFFFBCCF5 , 32'h0003DCD4 , 32'hFFFE14C7 , 32'hFFFFB290 , 32'h00000790 , 32'h00009ACD , 32'hFFFF9534 , 32'h000241F5 , 32'h0003194B} , 
{32'h0002D81D , 32'h0001D0BE , 32'hFFFDC8C1 , 32'hFFFE1657 , 32'h00031FB4 , 32'h00005D8A , 32'h00018989 , 32'hFFFD8449 , 32'h000140E4 , 32'h000100A9 , 32'h00032786 , 32'h0000DE87 , 32'h000029BC , 32'h0000F4B2 , 32'hFFFD2684 , 32'hFFFD9460 , 32'hFFFFF882 , 32'h00019A1E , 32'h00026B9A , 32'hFFFD67E9 , 32'hFFFF2142 , 32'h00004D0A , 32'hFFFE2B4E , 32'h00001FA8 , 32'hFFFEB9B2 , 32'hFFFD6D90 , 32'hFFFA8619 , 32'h00021F83 , 32'h0000A30D , 32'hFFFCBDFC , 32'hFFFC2420 , 32'h0002E6BE , 32'h0001B40A , 32'h0003691A , 32'h0003255D , 32'h00001730 , 32'h000365D6 , 32'hFFFF7FAB , 32'h00010C27 , 32'h00030D9D , 32'h00004D01 , 32'h00020D36 , 32'hFFFFFBB5 , 32'h00032289 , 32'h00038D7E , 32'hFFFD6B3B , 32'h00017377 , 32'h0002C31A , 32'h0002AEE8 , 32'hFFFF0F6B , 32'hFFFD1045 , 32'h0001A26C , 32'hFFFD4B74 , 32'h0001090F , 32'hFFFE0A62 , 32'hFFFEB7A8 , 32'hFFFAF011 , 32'hFFFF87F2 , 32'h0000988F , 32'h00031021 , 32'h0001396E , 32'hFFFF5784 , 32'hFFFCCAF8 , 32'hFFFD815E , 32'hFFFB059A , 32'hFFFE7088 , 32'h0003FDF5 , 32'hFFFFA8F6 , 32'h00009514 , 32'h00002191 , 32'hFFFEC97E , 32'hFFFF25EC , 32'hFFFE392C , 32'h0001D32F , 32'hFFFE6CB7 , 32'h00040964 , 32'h00022B38 , 32'hFFFC9DC9 , 32'h00002F2D , 32'h000010F8 , 32'hFFFCAE78 , 32'hFFFF9F54 , 32'h0002FAEE , 32'h000615D2 , 32'hFFFFABA2 , 32'hFFFCEF49 , 32'hFFFF3161 , 32'h0002896C , 32'h0003240C , 32'hFFFBFAEE , 32'hFFFFE15A , 32'h0003BBE7 , 32'hFFFE8755 , 32'hFFFFF2DD , 32'hFFFDD5F0 , 32'hFFFD7F5B , 32'hFFFBDC7A , 32'hFFFD8AC3 , 32'hFFFF3F47 , 32'hFFFE9F33} , 
{32'hE30FEE80 , 32'h29A0E8C0 , 32'h09EE57C0 , 32'h0B736780 , 32'h1738DD40 , 32'h0328BCBC , 32'h23FE79C0 , 32'h3FD77C00 , 32'hF0FF1050 , 32'h021B3E74 , 32'h038343DC , 32'hF9FF17D0 , 32'h0E10D9F0 , 32'hFA8C5498 , 32'h0DEC8C10 , 32'h0888A5A0 , 32'h00FAFE09 , 32'h0A87D520 , 32'h12C0F5E0 , 32'h00D10A9E , 32'hFCF6D04C , 32'h0899E520 , 32'hFD609D28 , 32'h0CD0DA40 , 32'h10E17900 , 32'hF3E61250 , 32'h10599BA0 , 32'h0587FD50 , 32'hF43E4EA0 , 32'hFFA72D65 , 32'h0536A9C8 , 32'h06302BE0 , 32'hFAAFED58 , 32'hF20973F0 , 32'hFAE6E9F0 , 32'hFC5FDED0 , 32'h02E7E128 , 32'h032C0DB8 , 32'hF9C7C478 , 32'h07E30F88 , 32'h10863A00 , 32'h0ECB57C0 , 32'hFC9C3CA0 , 32'h0CE086B0 , 32'h008CD736 , 32'hF34EA150 , 32'hFB089880 , 32'hF4D488B0 , 32'hFBB41E98 , 32'h07E0A5B0 , 32'hFDB5E440 , 32'h0168DA3C , 32'h0936E8B0 , 32'hF3C41720 , 32'h02447604 , 32'hFC83AE74 , 32'h00866259 , 32'hFC873FD4 , 32'h02166C50 , 32'h04A8F320 , 32'hFD91E0B4 , 32'h05D0CC00 , 32'hFA5559C8 , 32'h094D6DE0 , 32'hFE683E84 , 32'hF3E74080 , 32'hFF4C5D40 , 32'h021FB6B8 , 32'hFC094AD0 , 32'h0325D184 , 32'h060EA248 , 32'hFC637518 , 32'h000281CB , 32'hFE74C5C8 , 32'hFE181468 , 32'hFF0CD20A , 32'hFFE43786 , 32'hF95C92D8 , 32'hFFC74471 , 32'hFDBC3F44 , 32'h020168E8 , 32'h03333724 , 32'h01DC85E0 , 32'h003CD473 , 32'h01E39E3C , 32'hFD616418 , 32'h0122E5F0 , 32'hFF4EEDEF , 32'hFE9D32B0 , 32'hFF5102A1 , 32'h0000BEBE , 32'hFFFFE9D5 , 32'h00011A9C , 32'h00008A77 , 32'hFFFE65C4 , 32'hFFFFB791 , 32'hFFFE537D , 32'h0000D8BD , 32'h000202CF , 32'hFFFFAAD4} , 
{32'h0425D558 , 32'h0CA451D0 , 32'h00B3BB1D , 32'hE9F7E420 , 32'h02F649D4 , 32'hEA7EEC80 , 32'h2F7907C0 , 32'hD9AB5E40 , 32'h16389D00 , 32'h14E3EB40 , 32'hF4C85CC0 , 32'hFE1865A8 , 32'h03B8413C , 32'hFC176CB8 , 32'hEB2CD340 , 32'hFA125538 , 32'h0C5A62D0 , 32'h1456CF40 , 32'hED058500 , 32'h0790A9B0 , 32'hFF531EFA , 32'hFCB1F980 , 32'hF64579D0 , 32'h10E41C20 , 32'h03426A04 , 32'h0EBEFC30 , 32'h09136070 , 32'hF1A9B340 , 32'hF1CA0730 , 32'h0B862D30 , 32'h0828E6B0 , 32'h081F8B30 , 32'h04211E38 , 32'h167DF8C0 , 32'hF3830F70 , 32'h02312B88 , 32'hF74576A0 , 32'hFB2A5C00 , 32'hFBB457D8 , 32'h007DBA66 , 32'h0F9D5910 , 32'h09943250 , 32'h0DF98EB0 , 32'h07614B58 , 32'hF5CC7450 , 32'h06B01268 , 32'h040CA4E0 , 32'hF4175250 , 32'hFABC9C20 , 32'hF3762430 , 32'h0D6BD940 , 32'hFC838270 , 32'hFAC319E8 , 32'hF32E3D30 , 32'h0FFED920 , 32'hF8CA9E90 , 32'h053CACE8 , 32'h076AA170 , 32'h0B92B5E0 , 32'h031965AC , 32'h0112F394 , 32'hFD7B42E8 , 32'hFD5A1748 , 32'hFF46ACF5 , 32'h0082C9B8 , 32'h04D0C220 , 32'h04B75BF0 , 32'h026D0FBC , 32'hFC1CACF0 , 32'h02371974 , 32'h08A8B4B0 , 32'hFE367A1C , 32'hF59E96E0 , 32'h03615F28 , 32'hFE7E13B8 , 32'h0322986C , 32'h005B42B1 , 32'h0111886C , 32'hFF0F24EF , 32'hFFBB1E4C , 32'hFC4B1CAC , 32'hFB7C8888 , 32'h00EA0EED , 32'hFF74B100 , 32'hFF750879 , 32'h009FDBCE , 32'h03D949B8 , 32'hFD4307DC , 32'h02882EDC , 32'hFF33FEC3 , 32'hFFFBDDC7 , 32'hFFFC5225 , 32'h00013A35 , 32'hFFFDE12F , 32'h00012907 , 32'h0000686C , 32'hFFFD9945 , 32'hFFFEC573 , 32'hFFFED927 , 32'hFFFD31A2} , 
{32'hFFFFE0A1 , 32'h00035A3C , 32'hFFFF338D , 32'h000132DB , 32'h00032FB7 , 32'hFFFCFEED , 32'hFFFC7D82 , 32'hFFFF493A , 32'hFFFED025 , 32'hFFFE5E40 , 32'hFFFE0C77 , 32'hFFFDEAE9 , 32'h0000B217 , 32'hFFFDF9C1 , 32'hFFFFEE69 , 32'h0000306B , 32'hFFFF5D50 , 32'h0003129A , 32'hFFFED08F , 32'hFFFD8642 , 32'h0002E83C , 32'hFFFFCB1A , 32'h0000C875 , 32'hFFFADCA2 , 32'h0000325E , 32'h00032854 , 32'hFFFFF130 , 32'hFFFF964B , 32'h000037EB , 32'h000182D4 , 32'h0000033C , 32'hFFFBDC5A , 32'h00038938 , 32'hFFFFFBFD , 32'h00010FCF , 32'hFFFE11F6 , 32'hFFFEAF86 , 32'hFFFEE0D1 , 32'h000221C7 , 32'h00011BD2 , 32'hFFFEE42C , 32'h00020F6F , 32'h0006D2B1 , 32'h00023D58 , 32'h00044407 , 32'hFFFF9566 , 32'hFFFFE3FD , 32'h0000872F , 32'hFFFF1B6C , 32'hFFFF7E8F , 32'hFFFE78C3 , 32'hFFF72829 , 32'h00009CE0 , 32'hFFFF86B1 , 32'hFFFDF5CD , 32'h00017A70 , 32'hFFFE4D93 , 32'hFFFE0428 , 32'hFFF8F160 , 32'hFFFFF674 , 32'hFFFC348D , 32'h00028340 , 32'h000260F6 , 32'h000443C4 , 32'h00012A98 , 32'h000577A4 , 32'hFFFB1E2F , 32'h0000D8E3 , 32'hFFFEE296 , 32'hFFFA5702 , 32'hFFFFDAB7 , 32'h0002B319 , 32'h0000C482 , 32'h0000C629 , 32'hFFFE17B1 , 32'h0002F6D3 , 32'hFFFF0F13 , 32'hFFFB05B4 , 32'h0004FA1B , 32'hFFFC3679 , 32'hFFFECCA9 , 32'hFFFF57D0 , 32'hFFFEF817 , 32'hFFFF0466 , 32'hFFFD4040 , 32'h00011314 , 32'hFFFDDB2C , 32'h0001065A , 32'h00044CBE , 32'hFFFA5539 , 32'hFFFFB679 , 32'hFFFFCEB7 , 32'hFFFE4171 , 32'hFFFC9623 , 32'h00013E05 , 32'h0000DF5C , 32'h0001F6D9 , 32'hFFFD5C71 , 32'hFFFA3411 , 32'h00000715} , 
{32'hFFFE6C78 , 32'hFFFED531 , 32'h0005213B , 32'h0002B5DF , 32'hFFFEE8C0 , 32'hFFFE91F6 , 32'hFFFF4AAA , 32'h0005FD51 , 32'h00054ACD , 32'h000187BD , 32'hFFFD023B , 32'hFFFEF344 , 32'hFFFE984D , 32'h00046C93 , 32'hFFFC86BF , 32'h00020735 , 32'hFFFAC0F3 , 32'h00009007 , 32'h00000F24 , 32'h000244EF , 32'hFFF9F7D7 , 32'hFFFE5120 , 32'hFFFCBA0D , 32'hFFFDF638 , 32'h0000271E , 32'h0002898C , 32'hFFFCEA0C , 32'hFFFDEF68 , 32'h0001FCD0 , 32'hFFFFA33A , 32'h0000CC34 , 32'h000410D3 , 32'hFFFE4DA3 , 32'h000108F9 , 32'h000288B9 , 32'hFFFD241E , 32'h00017C9B , 32'h0002C731 , 32'hFFFA326E , 32'h000193EC , 32'hFFFBA522 , 32'h00009AF1 , 32'hFFF8B4C4 , 32'hFFF961EE , 32'h0000ADB0 , 32'h0005A7D5 , 32'hFFFEF868 , 32'hFFFE2773 , 32'hFFFE71B9 , 32'h0000545F , 32'h0003324D , 32'h00007BDC , 32'hFFFA337C , 32'hFFFCF2EC , 32'h0003BC25 , 32'hFFFAF7F8 , 32'h0000DBC9 , 32'h0006E996 , 32'h0002D021 , 32'hFFFF824E , 32'hFFFEE493 , 32'h0002F929 , 32'h000295DD , 32'hFFFF0AB4 , 32'hFFFBDBFE , 32'hFFFEFAF0 , 32'hFFFA8801 , 32'hFFFDA44E , 32'hFFFF1C47 , 32'hFFFCD76A , 32'hFFFF2496 , 32'h000170DA , 32'hFFFF211E , 32'hFFFF60CF , 32'hFFFDE0A2 , 32'hFFFC4DAB , 32'hFFFD7E22 , 32'h00052F70 , 32'hFFFE1E8A , 32'h0000D624 , 32'h00020265 , 32'h00060866 , 32'h0004017E , 32'hFFFE4E25 , 32'h000125FA , 32'h00040C59 , 32'h0001D548 , 32'h000302C6 , 32'h0000035A , 32'hFFFC4DBE , 32'hFFFD7BC8 , 32'h00004F7F , 32'h0007ED02 , 32'h0003E16A , 32'hFFFFCECF , 32'hFFFDDF32 , 32'h0001ECF8 , 32'hFFFF2428 , 32'h00012D5C , 32'hFFFFABAA} , 
{32'hFFFD8124 , 32'h0003DAFB , 32'hFFFF706B , 32'hFFFEF1C9 , 32'hFFFE5659 , 32'hFFFE9C7D , 32'h000266F0 , 32'h0000679E , 32'hFFFEA6BE , 32'hFFFD950F , 32'h0002D8AD , 32'hFFFFAD9C , 32'h0001E1FC , 32'h0003C2B9 , 32'hFFFFD674 , 32'h00016A4E , 32'h0000B47E , 32'hFFFDCE65 , 32'hFFFEF291 , 32'hFFFEDD6C , 32'h00037D06 , 32'h0000968A , 32'h00018208 , 32'h0000B795 , 32'hFFFDDFE0 , 32'hFFFD7BB8 , 32'hFFFD1311 , 32'hFFFEFBFD , 32'h00021A3D , 32'hFFFF2CA5 , 32'h0002B063 , 32'hFFFC9015 , 32'hFFFC39CB , 32'h00000E3D , 32'h0001F49F , 32'h000298D4 , 32'hFFFFD10F , 32'h0001B46A , 32'hFFFF4617 , 32'h000156AE , 32'hFFFE27FC , 32'hFFFF3AF7 , 32'h0002174F , 32'h000121CF , 32'hFFFEB5F7 , 32'hFFFC63DD , 32'h00014677 , 32'hFFFC8A52 , 32'h00055DB6 , 32'hFFFF3682 , 32'hFFFE2324 , 32'hFFFDFE52 , 32'hFFFDD13A , 32'h000147F7 , 32'h0000BC50 , 32'hFFFF0312 , 32'hFFFD0D13 , 32'hFFFCDA26 , 32'h0004B343 , 32'hFFFFC3EE , 32'h00007D11 , 32'hFFFD5B3F , 32'hFFFE8458 , 32'h0000911D , 32'h0002FE9F , 32'h00021FC3 , 32'hFFFEBDBA , 32'hFFFDBDB4 , 32'h00013B85 , 32'h00004E20 , 32'h0004353D , 32'hFFFEE937 , 32'h000270AD , 32'h0003C5FF , 32'h000299FC , 32'hFFFBD90D , 32'h00017F78 , 32'h0002C1F4 , 32'hFFFBF122 , 32'h00050C43 , 32'h00023C90 , 32'hFFFD9080 , 32'h00013689 , 32'h000B5B8D , 32'hFFFC9D96 , 32'h00002E64 , 32'hFFFEBD2B , 32'hFFFFF204 , 32'h00003972 , 32'h00017625 , 32'h0000D12D , 32'hFFFF9160 , 32'hFFFB15AD , 32'hFFFF13EC , 32'h000200BE , 32'h00025A42 , 32'hFFFCD430 , 32'h0005202C , 32'h000287D9 , 32'h0001CFB5} , 
{32'h00048E24 , 32'h0001B06E , 32'h00028559 , 32'hFFFC92E6 , 32'hFFFED567 , 32'h0002998E , 32'hFFFC4278 , 32'hFFFD36BC , 32'hFFFD75BB , 32'hFFFDC23C , 32'h000303C1 , 32'hFFFE5A97 , 32'hFFFB864F , 32'h000148EA , 32'hFFFE9702 , 32'h0000467B , 32'h000279DC , 32'hFFFE5A3E , 32'h0000C4F9 , 32'h00031B10 , 32'hFFFF146D , 32'h0002A9E7 , 32'h00001F0A , 32'h00000576 , 32'h0001B2AD , 32'hFFFD4055 , 32'h00009DF5 , 32'hFFFF849F , 32'h0001E19D , 32'hFFFF90C0 , 32'hFFFCD53C , 32'h0000DA8E , 32'hFFFEDE41 , 32'h0000315C , 32'h0002A2EE , 32'h0001501D , 32'h00022CB9 , 32'h0001FF9B , 32'hFFFA5272 , 32'h00060761 , 32'h000127F4 , 32'h0001D891 , 32'hFFFE5B8D , 32'h0001BB04 , 32'h00022934 , 32'hFFFFD3A4 , 32'h00002BF4 , 32'hFFFBE3AD , 32'h0001E053 , 32'hFFFE04A6 , 32'h0003F4E3 , 32'h000379E7 , 32'hFFFE7E10 , 32'hFFFEC8E9 , 32'h00001B68 , 32'h0003CEEF , 32'h0000CDCD , 32'hFFFC6639 , 32'hFFFCD5F8 , 32'h0000B481 , 32'h000374B5 , 32'h000014B2 , 32'h000357C6 , 32'h000040A1 , 32'h0002396B , 32'h0001F232 , 32'hFFFD740C , 32'h0000C06B , 32'hFFFF248A , 32'h000039EB , 32'hFFFCB3B5 , 32'h0001B1BF , 32'h00021A0E , 32'h00017354 , 32'h00035361 , 32'h0002967E , 32'h00036B1C , 32'hFFFF30B8 , 32'h000388E3 , 32'h000142E7 , 32'h00013EBD , 32'hFFFB2B66 , 32'h0000D2FE , 32'h0001167F , 32'h0004036E , 32'h00035CBB , 32'hFFFF31DB , 32'h0001E120 , 32'hFFFD66A4 , 32'hFFFF55AB , 32'h0000ADFE , 32'hFFFDD6D1 , 32'h00049AF6 , 32'hFFFFEDE2 , 32'h0005729B , 32'h00012D56 , 32'h0000C081 , 32'hFFFDC29B , 32'hFFFE1874 , 32'hFFFFD379} , 
{32'hFFFD5DF2 , 32'hFFFAF290 , 32'h0003C056 , 32'hFFFD73BC , 32'hFFFE9D30 , 32'h00032D3C , 32'hFFFDB510 , 32'h0001AFF0 , 32'hFFFF5C12 , 32'h00043600 , 32'hFFFFF6E2 , 32'hFFFEF4E6 , 32'h00033D20 , 32'h0000CDC3 , 32'hFFFFEEE3 , 32'hFFFBEB2D , 32'hFFFFC7D7 , 32'h0002A3F3 , 32'hFFFFB853 , 32'hFFFEE41D , 32'h0002E1D3 , 32'h000129B8 , 32'hFFFF34E3 , 32'h00001788 , 32'hFFFD49EF , 32'hFFFE081D , 32'hFFFB558F , 32'h0003ED1F , 32'h00005851 , 32'h00016388 , 32'hFFFCFB96 , 32'h00027AB8 , 32'h000133A8 , 32'hFFFE42DC , 32'hFFFF792A , 32'h000030F7 , 32'hFFFF1EF5 , 32'hFFFE8B46 , 32'h0005086A , 32'h0000C8DC , 32'h0000A1EB , 32'h0002BD25 , 32'h00028FAB , 32'hFFFE92A1 , 32'hFFFF55E0 , 32'h0001E0AF , 32'h0001E91B , 32'hFFFFC1EB , 32'hFFFF7BED , 32'hFFFB60E5 , 32'hFFFFECED , 32'h00005653 , 32'hFFFF4E27 , 32'hFFF70FCD , 32'hFFFE6985 , 32'hFFFBA403 , 32'hFFF97405 , 32'h000088D6 , 32'hFFFD65D5 , 32'hFFFFAA58 , 32'hFFFC8EFC , 32'hFFFE59C1 , 32'hFFFD085A , 32'hFFFF63B2 , 32'h0001EBC1 , 32'h00007858 , 32'hFFFE851C , 32'h0001FD1D , 32'h0000626F , 32'h0005121A , 32'hFFFF7477 , 32'h0001F465 , 32'h000135B9 , 32'hFFFB102E , 32'hFFFC38E8 , 32'h0002FE1B , 32'h0001D20E , 32'hFFFBBCBE , 32'hFFFF768E , 32'h000055C8 , 32'hFFF9D546 , 32'h00028F31 , 32'hFFFE6B7E , 32'h0002470E , 32'hFFFF37F6 , 32'h0001077C , 32'h0001EE74 , 32'h00021312 , 32'hFFFF3BB1 , 32'hFFFFB256 , 32'h0001BFDB , 32'hFFFB6EDF , 32'hFFFEFAC8 , 32'h0000E9D0 , 32'h00034625 , 32'hFFFEC03A , 32'h00011ED1 , 32'hFFFE7800 , 32'h0002DCA8 , 32'hFFFC788F} , 
{32'hEAB853E0 , 32'h00172B16 , 32'h0B1ED0B0 , 32'hFB9FF570 , 32'hF709D600 , 32'h148E7AC0 , 32'hF1B485A0 , 32'h0CCC37A0 , 32'hEB0B2FE0 , 32'h026D5EDC , 32'hF47A9CC0 , 32'h188FF8C0 , 32'hEEAECB00 , 32'hEC40AF00 , 32'hFDCC5C24 , 32'hFF62013B , 32'hF0E334B0 , 32'hFE48BA28 , 32'h10182AE0 , 32'hFA151010 , 32'hFFE6F9A1 , 32'h05B20D78 , 32'hFBE14980 , 32'h0685F658 , 32'h080DA850 , 32'h0191B04C , 32'h0C42BFC0 , 32'h075ADBD0 , 32'h007324DA , 32'hF7B6F5A0 , 32'hEEFD3F80 , 32'h0721C5C8 , 32'hFD84FF48 , 32'h08298980 , 32'h059F1388 , 32'h04779058 , 32'hF346A080 , 32'h03F1CD20 , 32'h06F6F480 , 32'hFDF69E68 , 32'hF886C258 , 32'hFFDAB6DC , 32'h06FDD260 , 32'hFD47B398 , 32'h075B5758 , 32'hFB81B688 , 32'hF7A2D750 , 32'hFD1CB02C , 32'h04A83F88 , 32'h013F0B24 , 32'hFAFA9930 , 32'hFE0F7B54 , 32'hFE6415DC , 32'hF57CE3C0 , 32'hFF708667 , 32'h023BE858 , 32'h004C2ECE , 32'h0259B084 , 32'h0A01B880 , 32'hFB2C58A0 , 32'h060896D8 , 32'hFA4359E8 , 32'hF9B17B60 , 32'h02A7A3AC , 32'h092AD990 , 32'h01A1884C , 32'h094EE920 , 32'h09ADF6E0 , 32'h0060E6F6 , 32'h061D3140 , 32'hFAA75398 , 32'hFCA858D8 , 32'h017DA808 , 32'h0520C730 , 32'hFE2104D0 , 32'hFD32FA7C , 32'hFD6BD2AC , 32'hFE21B094 , 32'hFF1315F9 , 32'h02EA9A60 , 32'hFF83475D , 32'hFEA5AFB0 , 32'hFA5C2F00 , 32'hFE729100 , 32'hFEF23378 , 32'hFFE463B8 , 32'hFEDAE8CC , 32'h013FF9C8 , 32'h002750ED , 32'hFFF71C65 , 32'hFFFEBA26 , 32'h00017619 , 32'hFFFBC991 , 32'h0003869E , 32'h0002E76E , 32'h00032ED5 , 32'h0000BCD1 , 32'h0001DE7A , 32'hFFFEC4E7 , 32'hFFFEE27A} , 
{32'hEBF18860 , 32'h0DB3E6F0 , 32'h00C33D2A , 32'hF07029B0 , 32'hE49817A0 , 32'hF3AACED0 , 32'h0DC82D60 , 32'hF24173D0 , 32'h004B4FBC , 32'h0D7A5240 , 32'hFD8D40A0 , 32'h130E46E0 , 32'hDFF1C5C0 , 32'h04F83738 , 32'h0FCF3150 , 32'hED7D6400 , 32'hEF900360 , 32'h13013F00 , 32'hF147DE00 , 32'h0A371B10 , 32'h0687D470 , 32'h031EFBC0 , 32'hF3DAFAD0 , 32'hF8415AD8 , 32'hEBDC3D00 , 32'hF2C5D100 , 32'h13B636E0 , 32'h04AF5AA0 , 32'h04BA39A8 , 32'h10BCD000 , 32'h08B69990 , 32'hE4DCDF20 , 32'h0B18E780 , 32'h08D2AC60 , 32'hFB1D76F0 , 32'hF3B22B60 , 32'h0BFECB50 , 32'h10C23D20 , 32'h0397B558 , 32'hFDAFDDA0 , 32'h03D705B4 , 32'h030D9178 , 32'h0B3022C0 , 32'h037C86C0 , 32'h040CE9B8 , 32'hF792F1B0 , 32'h0CDABC90 , 32'hF9FE6790 , 32'hFAEBD628 , 32'hF8CABC90 , 32'h0A52F4A0 , 32'h08C7C2A0 , 32'hEAAFF780 , 32'hFDB1BC0C , 32'hFB093360 , 32'hFF08F877 , 32'hFAAEF8D0 , 32'hFBB44680 , 32'hFE205660 , 32'hFDA2046C , 32'h009E4880 , 32'hFDA02E50 , 32'h02E72254 , 32'h08C39EA0 , 32'h095F8C70 , 32'hFAF62060 , 32'hF840FF88 , 32'h08827A30 , 32'hFEA72734 , 32'h03A43378 , 32'hFD1A96F4 , 32'h02155F24 , 32'hFE37D8A4 , 32'hFEC8D71C , 32'hFEDA4F58 , 32'hFDAF75A4 , 32'h001CE892 , 32'h02CC3020 , 32'h00377C65 , 32'hFE32FAD8 , 32'h03F1BA54 , 32'hFBD3DD28 , 32'h04C880C0 , 32'hF9621F00 , 32'h01E11480 , 32'hFD19F468 , 32'h002D36AE , 32'h03689FE8 , 32'h01A29F90 , 32'h00AD179A , 32'h0004B357 , 32'h0000D7E3 , 32'hFFFE6B31 , 32'h00012C00 , 32'h00009BBA , 32'hFFFE5084 , 32'hFFFF8389 , 32'hFFFDEF13 , 32'h000103E8 , 32'h0001D7F7} , 
{32'hFFFDFC21 , 32'h00008A54 , 32'hFFFF4155 , 32'hFFFF27EC , 32'h00000087 , 32'h0000877F , 32'h000401FD , 32'h00004456 , 32'h00022535 , 32'hFFF9D35E , 32'h00004E0F , 32'hFFFECE2D , 32'h0001A7FA , 32'h00006607 , 32'hFFFF352F , 32'hFFFB6252 , 32'h00056F5D , 32'h0008B7FE , 32'hFFFFEFDE , 32'h0003A7CC , 32'h000073F0 , 32'hFFFBC51B , 32'h00021B1E , 32'h00011B12 , 32'h0000D786 , 32'hFFFFA236 , 32'h00008CB0 , 32'h0000B274 , 32'h00035171 , 32'hFFFF5888 , 32'hFFFBA2A5 , 32'hFFFEE92E , 32'h000592A0 , 32'h00032B8A , 32'h0000A9DC , 32'hFFFB1DA9 , 32'h0000D60A , 32'hFFFA47CD , 32'hFFFF2460 , 32'h0004BB7F , 32'h0003F67C , 32'h0000DA52 , 32'hFFFFC9C5 , 32'h00027B28 , 32'h0001B692 , 32'h00012565 , 32'hFFFCEFEA , 32'hFFFFD3D2 , 32'hFFFD58FC , 32'h00015A33 , 32'hFFFF5EB5 , 32'hFFFE07B2 , 32'h00026CD5 , 32'h00028853 , 32'hFFF74DED , 32'hFFFEF152 , 32'h0004C2E3 , 32'h00039B5C , 32'hFFFF3DBF , 32'h000200B1 , 32'h00060710 , 32'hFFFDEC89 , 32'h00021A4E , 32'hFFFDCF33 , 32'h00019BDB , 32'hFFFEF70E , 32'h0000C88A , 32'h0000652E , 32'hFFFEB210 , 32'hFFFF9BF5 , 32'hFFFC06DB , 32'hFFFDE025 , 32'h0001683B , 32'h000054DE , 32'h0000B963 , 32'h00016BF2 , 32'hFFFF03CB , 32'hFFFB8E8C , 32'h00045F39 , 32'h00042D5B , 32'h000019EC , 32'hFFFE4335 , 32'hFFF93550 , 32'h000170AD , 32'hFFFE6933 , 32'hFFFFF87F , 32'h00002EE0 , 32'h00005B53 , 32'hFFFE2BF9 , 32'hFFFD9A8A , 32'hFFFFA778 , 32'h0000070B , 32'h000412C7 , 32'h0000195F , 32'hFFFF8BCA , 32'h00023242 , 32'h000385AF , 32'h00055074 , 32'hFFFF8C70 , 32'hFFFAFC20} , 
{32'h0001999F , 32'hFFFEC9AD , 32'h0000AC41 , 32'h0000D764 , 32'h000154B0 , 32'hFFFE600F , 32'h00051127 , 32'hFFFFB7D2 , 32'h000562AF , 32'h00001C45 , 32'h0001817B , 32'h0003FDCA , 32'hFFFFAC60 , 32'h0000D526 , 32'hFFFEBC88 , 32'hFFFDDA82 , 32'hFFFB83A7 , 32'hFFFD81E2 , 32'hFFFFE799 , 32'h00002466 , 32'h000337AD , 32'hFFFDD51F , 32'hFFFFE74F , 32'hFFFFB876 , 32'h00038C4E , 32'hFFFE71B6 , 32'hFFFEF90A , 32'h00010535 , 32'hFFFD2649 , 32'hFFFFECE1 , 32'h00036356 , 32'hFFFEBB4F , 32'hFFFE3FBE , 32'hFFFE701A , 32'hFFFDFA40 , 32'h00040617 , 32'h000044EF , 32'hFFFE6EB7 , 32'h000421C1 , 32'hFFFDFA03 , 32'h0001DF86 , 32'h00002F9C , 32'h0000A4F5 , 32'h000021E0 , 32'h0001FC56 , 32'hFFFF3A12 , 32'h0001655A , 32'h00057356 , 32'h0001AB98 , 32'h0001827C , 32'h00028713 , 32'hFFFD39D9 , 32'h0000F80F , 32'h000422E6 , 32'h0002B39D , 32'h0002737D , 32'h00005977 , 32'h00013230 , 32'h00010CA8 , 32'h00018861 , 32'h0000D688 , 32'hFFFBC7CB , 32'hFFFE2F14 , 32'h00005627 , 32'hFFFF70E5 , 32'h00009433 , 32'hFFFE0097 , 32'hFFFEDEF2 , 32'h00024F49 , 32'hFFFFB7A9 , 32'hFFFF4046 , 32'h0005A637 , 32'hFFFEE8DE , 32'hFFFECF5A , 32'hFFFBD976 , 32'hFFFF4CF5 , 32'hFFFE8213 , 32'h0001529D , 32'h00024A82 , 32'h0001C918 , 32'hFFFFF751 , 32'hFFFF0BA6 , 32'h0001CAC9 , 32'h00039AA6 , 32'hFFFBD7A9 , 32'hFFFD8A6F , 32'hFFFDD905 , 32'hFFFF7876 , 32'hFFFEDD16 , 32'h0002C852 , 32'h00025EFF , 32'hFFFCAE71 , 32'h0002766B , 32'h0000B7EE , 32'hFFFEBBF3 , 32'hFFFF712A , 32'h00000D7B , 32'hFFFD7D0E , 32'h000051A0 , 32'hFFFF55D8} , 
{32'h4ABB7600 , 32'h15626900 , 32'h42F0FE00 , 32'h1C8F4C60 , 32'hC4048100 , 32'hFCA6C768 , 32'h0D366B60 , 32'h21178600 , 32'h0BD0F0F0 , 32'hFF22F41E , 32'h0118344C , 32'h0638DDB8 , 32'h1554C340 , 32'h15E57F60 , 32'hFE7881D0 , 32'h0446FBF0 , 32'hE76AFD60 , 32'h0873A4F0 , 32'hF0D93250 , 32'hF217F6E0 , 32'h01D8508C , 32'h08C9C1D0 , 32'h044D5CD0 , 32'hF00600C0 , 32'h046F9C08 , 32'h081703A0 , 32'hFA6433D0 , 32'h08FFBF20 , 32'h10C58800 , 32'hF3E77F00 , 32'hF14E2050 , 32'h114DABC0 , 32'h0F002040 , 32'h010D9E64 , 32'hEF711000 , 32'h081B05E0 , 32'h035DD600 , 32'h0F296150 , 32'h07D75718 , 32'hEDFC4400 , 32'h0A4EE5A0 , 32'h0A467E20 , 32'h00DCF18F , 32'h10A31EA0 , 32'h01D59E84 , 32'hFC40D83C , 32'hFD909B80 , 32'h03324750 , 32'h08378EB0 , 32'h02096764 , 32'h02170220 , 32'h077B5A48 , 32'h04BC0F48 , 32'hFDAFD290 , 32'h099F58C0 , 32'h03C85DE4 , 32'h06FC2CC8 , 32'h022E3BD4 , 32'h02C60DE0 , 32'h054D2108 , 32'hFCE2F370 , 32'h077A6270 , 32'hFAAF3AF0 , 32'hF8A09F80 , 32'h05241880 , 32'h030BF3CC , 32'hFF79D36A , 32'hFDAD36AC , 32'h0287BB7C , 32'h050DB508 , 32'h013E593C , 32'hFE39E670 , 32'hF82F7240 , 32'h0207E798 , 32'h02CFA780 , 32'hFD6D9964 , 32'h009066E6 , 32'h03268334 , 32'h00B8C09F , 32'h05726E58 , 32'h01354AFC , 32'hFCE856F8 , 32'h0220E154 , 32'hFFD622FE , 32'h014FE7A0 , 32'hFF7855C8 , 32'h010A7660 , 32'hFD547290 , 32'h01097344 , 32'h00AED403 , 32'hFFFDACCF , 32'h0000AAC9 , 32'hFFFD9F5A , 32'hFFFE60D0 , 32'hFFFEB998 , 32'hFFFD159C , 32'hFFFF6948 , 32'hFFFF5511 , 32'hFFFFDBBB , 32'h00012015} , 
{32'h1591CB60 , 32'h0F21EF80 , 32'h24196740 , 32'h0DF57010 , 32'hE9EC3B00 , 32'h0B136280 , 32'hF2FEAF10 , 32'h08078A00 , 32'h0DF2AEB0 , 32'hFE0ED4E4 , 32'h0663ED98 , 32'h0DCF64D0 , 32'hF9F3F3F0 , 32'h0A199D70 , 32'h19A21B00 , 32'h02B5F6E4 , 32'h057F1BC8 , 32'hFBF845E0 , 32'h05DE4CB0 , 32'h0DDE8880 , 32'hF33331E0 , 32'hFB240030 , 32'h019ECD40 , 32'h0DC5BFB0 , 32'h04592C10 , 32'hF279DFB0 , 32'h00CD1C64 , 32'hFD604490 , 32'hF98F7058 , 32'h0C617700 , 32'h13433580 , 32'h03F0F6CC , 32'hEF863C40 , 32'hFC02E988 , 32'hFC6207D4 , 32'hF83F7C08 , 32'h02D8EDE8 , 32'h06F2B9C0 , 32'h0498D100 , 32'h02ADA02C , 32'hFB983060 , 32'hF89536F8 , 32'hF88312E0 , 32'h024120D8 , 32'h05101628 , 32'hFB32C940 , 32'h02151ADC , 32'hF91BAC70 , 32'h0074EA22 , 32'h13CF2540 , 32'h0B24C980 , 32'hFB91EB58 , 32'hFE380F8C , 32'hFDA3FBEC , 32'hFB452128 , 32'hFDEFAAEC , 32'h04C08BC0 , 32'h00DB4DD8 , 32'hF5485480 , 32'hF96B0958 , 32'h0ACE8EC0 , 32'hF60E59F0 , 32'h019C92F4 , 32'hF6505110 , 32'hFC4CCE18 , 32'hFE2A33B0 , 32'hFC3D9500 , 32'hFC7F79F0 , 32'hFB516908 , 32'h049CA0F8 , 32'h01045B10 , 32'hFD258EDC , 32'hF9EBE0B0 , 32'hFE20A250 , 32'h02692668 , 32'hFB7B23A8 , 32'hF89D84D8 , 32'hFE01C830 , 32'h09DBC7D0 , 32'hFFE5A24A , 32'hFCB62E2C , 32'hFF882EE1 , 32'hFCF97550 , 32'h019EBC4C , 32'h0448DAA0 , 32'h03D271A0 , 32'h045B7110 , 32'hFDD73DB0 , 32'hFE51DFB0 , 32'hFF05D14B , 32'h000105A8 , 32'h0000C40C , 32'h00015521 , 32'hFFFFA2EE , 32'hFFFF2235 , 32'h0000783F , 32'hFFFCDD19 , 32'hFFFF6860 , 32'hFFFF41B3 , 32'h000030BA} , 
{32'h0001B5E9 , 32'h000047E1 , 32'h0000AD61 , 32'h000179D4 , 32'hFFFF1214 , 32'h0001A253 , 32'h00048A63 , 32'hFFFFA308 , 32'hFFFE30C6 , 32'hFFFEA8AB , 32'h000221C2 , 32'hFFFFE6B7 , 32'hFFFA14DB , 32'h0005B63F , 32'hFFFDFE51 , 32'hFFFC64E3 , 32'h00002EF1 , 32'hFFFB8361 , 32'h00026AC9 , 32'hFFFC00A4 , 32'h000122EE , 32'h00015BEA , 32'hFFFD2EB0 , 32'h00001EF9 , 32'h00020412 , 32'h0003206B , 32'h00006B6D , 32'h000246AA , 32'hFFFE6012 , 32'hFFFE8152 , 32'h00034CA1 , 32'h00045775 , 32'h0001B87F , 32'h000056B6 , 32'h0002A797 , 32'h000004C5 , 32'hFFFF73AC , 32'hFFFCEB0B , 32'h0002FF71 , 32'hFFFFE716 , 32'h00011379 , 32'hFFFFD833 , 32'hFFFD969E , 32'hFFFC2703 , 32'hFFFCAFCE , 32'h0001AC0F , 32'h0002B450 , 32'hFFFC43F3 , 32'hFFFDEDF4 , 32'hFFFE4CBC , 32'hFFFF058C , 32'hFFFE1C3B , 32'h00000612 , 32'hFFFD5615 , 32'hFFFFC4CC , 32'h00014C5E , 32'hFFFDCA72 , 32'hFFF9252B , 32'h000237CB , 32'hFFFC405C , 32'hFFFC8A64 , 32'h00039B50 , 32'h000413BF , 32'hFFFE2457 , 32'hFFFD2087 , 32'h00038B86 , 32'hFFFF0B34 , 32'hFFFDE561 , 32'hFFFBEE47 , 32'h0000295F , 32'hFFFFE59B , 32'hFFFF2643 , 32'hFFFFC0CA , 32'h0002A64A , 32'h0000AAFE , 32'h0001CB48 , 32'h00039078 , 32'hFFFE6F28 , 32'hFFFF9FA1 , 32'hFFFACD0F , 32'h0001EA6B , 32'hFFFF3FDD , 32'h0002B85D , 32'h0002CE3E , 32'h0004835B , 32'h00019318 , 32'h00004024 , 32'h0000DCEC , 32'h00014BB4 , 32'h0001ECB8 , 32'h0000BB1A , 32'h000073AF , 32'h0000F773 , 32'hFFFEEC51 , 32'hFFFEEC64 , 32'h000352A0 , 32'h000151E2 , 32'hFFFF3289 , 32'h00005FD7 , 32'h00001E42} , 
{32'hFFFFDFC7 , 32'hFFFF9141 , 32'hFFFCF334 , 32'hFFFFBEBA , 32'h00001A2E , 32'hFFFC73C8 , 32'h00036706 , 32'h0001AF03 , 32'hFFFD90C5 , 32'h00013A5A , 32'h0001F93B , 32'h0003A251 , 32'hFFFDF478 , 32'hFFFE36A3 , 32'h0003ECE9 , 32'hFFFE38A1 , 32'hFFFE1B64 , 32'hFFFC016B , 32'h0002CDA0 , 32'hFFFE050D , 32'hFFFFC03A , 32'hFFFD10AA , 32'hFFFDB9E7 , 32'h00009FC3 , 32'h00009C5D , 32'hFFFD3C66 , 32'hFFFFE05E , 32'hFFFD8A72 , 32'hFFFD80E0 , 32'hFFFC81E3 , 32'h0003ED38 , 32'h0000240A , 32'hFFFDBC2C , 32'hFFFFB6C1 , 32'hFFFFD3DE , 32'hFFFCBB23 , 32'hFFFF02B2 , 32'h0003E713 , 32'hFFFF9BA1 , 32'hFFFBAFA0 , 32'hFFFFB89C , 32'h0002DE58 , 32'h0003C0B8 , 32'h00003412 , 32'hFFFFF0ED , 32'hFFFCEAF8 , 32'hFFFA5F76 , 32'h00021146 , 32'h000166B4 , 32'h00055A54 , 32'h0001B19F , 32'h0004507A , 32'hFFFE933F , 32'h0003AE78 , 32'hFFFE01E5 , 32'h00047EA7 , 32'h00008A1C , 32'h0001884E , 32'hFFFB6D6E , 32'hFFFA2F50 , 32'h00025C68 , 32'hFFFD302B , 32'hFFFD6BA0 , 32'hFFFE4F75 , 32'hFFFE1FCD , 32'hFFFD0729 , 32'h00019EB1 , 32'h00021023 , 32'hFFFCDBD8 , 32'h0004C39E , 32'h0002D949 , 32'hFFFDC8E9 , 32'h00030DEE , 32'h00014122 , 32'h000223B4 , 32'hFFFBE986 , 32'hFFFFFD27 , 32'hFFFEF3B7 , 32'h00006F35 , 32'h000230A0 , 32'hFFF92FFA , 32'hFFFDE015 , 32'h0002BFDE , 32'h000023D5 , 32'hFFFFC705 , 32'h00002D3B , 32'hFFFD8C1A , 32'h00024FA0 , 32'h0000D2DA , 32'hFFFEADDF , 32'hFFFEC643 , 32'hFFFE7C1F , 32'hFFFE341E , 32'hFFFBCA0C , 32'hFFFEC7FD , 32'h00000F65 , 32'h00032439 , 32'h000107E1 , 32'hFFFDCBD4 , 32'hFFFC5B73} , 
{32'hE5FE0AE0 , 32'h113B3BE0 , 32'h01B8BB94 , 32'h28851D00 , 32'hF392E730 , 32'h06B3CC90 , 32'hFAE365A8 , 32'hF95FDAA0 , 32'h09855860 , 32'hF99F1BE0 , 32'hF85D0BD8 , 32'h0D456940 , 32'h10B24620 , 32'hF3F64D30 , 32'h15C14300 , 32'hF7C937A0 , 32'hFB56CE10 , 32'h11450060 , 32'hF7BCC8B0 , 32'h034D2274 , 32'hF0835E00 , 32'hF763AD70 , 32'h07A108A0 , 32'h0BB98AA0 , 32'hFA231DC8 , 32'h129603A0 , 32'hFB30A908 , 32'hECC81F80 , 32'h00BE46E7 , 32'h09108D70 , 32'hFE1982F8 , 32'hF4460500 , 32'h0DB5B2B0 , 32'h00F8E719 , 32'h0531CE98 , 32'hFF734782 , 32'h11ADBFA0 , 32'h051C0888 , 32'hFC8D90AC , 32'hF22FCCE0 , 32'hF4517C00 , 32'hFFD78182 , 32'hFFACBC74 , 32'h0E53B4F0 , 32'hFB7FD768 , 32'hFF97BE96 , 32'h0033314F , 32'h01322140 , 32'hFDCA41D0 , 32'h00363C5B , 32'h073845B0 , 32'hF7737FE0 , 32'h06526BE8 , 32'hF686A8E0 , 32'hFCF0A630 , 32'h05581F88 , 32'h0B514CD0 , 32'h0254179C , 32'hF9F5AF38 , 32'hFA2D4018 , 32'h00B98BE3 , 32'hFA3F3678 , 32'hF9C57EE0 , 32'h05F9DAE8 , 32'h06DD26F0 , 32'h05D72FE0 , 32'hFF9DDD7B , 32'h0543EEE8 , 32'hFC8D8C6C , 32'hFB342260 , 32'h03E647D8 , 32'hF6D2B770 , 32'h038A8780 , 32'h02E88D44 , 32'hFA1874D8 , 32'h01123B54 , 32'h003587C4 , 32'hFF5054A2 , 32'hFDF80F30 , 32'hFE3E495C , 32'hFE2DDA34 , 32'hFFB0FB63 , 32'hFDE00DB4 , 32'hFE79584C , 32'h01287948 , 32'hFDC2C118 , 32'h00D773A0 , 32'hFF885007 , 32'h003A39B2 , 32'h0042E0E4 , 32'h0003A1FD , 32'h00014990 , 32'hFFFD324C , 32'hFFFE3B53 , 32'h00027D3C , 32'h000415AE , 32'hFFFE1CBD , 32'hFFFF6FC1 , 32'hFFFE141D , 32'hFFFF514F} , 
{32'h0000A203 , 32'hFFFD82B9 , 32'h0003CE1D , 32'h0003900F , 32'hFFFCDB4B , 32'h00007A62 , 32'hFFFED6C8 , 32'h000156EB , 32'hFFFD768F , 32'hFFFD5318 , 32'h0001C1C2 , 32'h0003E257 , 32'h0002EAC4 , 32'hFFFD74E3 , 32'h0000603E , 32'hFFFECF43 , 32'h0002C359 , 32'hFFFE7E71 , 32'h0002BA69 , 32'h000099EC , 32'hFFFD99CC , 32'hFFFCAD99 , 32'h0001C22E , 32'hFFFF0800 , 32'h000641A8 , 32'h00045C39 , 32'hFFFE7F8F , 32'hFFFDBC90 , 32'hFFFEDBCF , 32'h0001FC7B , 32'hFFFE221F , 32'hFFFCDD15 , 32'hFFF95AF0 , 32'h000127A8 , 32'h0003CBE9 , 32'h0000DE20 , 32'h0000C363 , 32'h0000B77D , 32'hFFFF158F , 32'hFFFF2BAA , 32'hFFFCB5B3 , 32'hFFFB87DC , 32'h00049870 , 32'h0001A241 , 32'h000149EF , 32'h00039562 , 32'hFFFD83DA , 32'hFFFF4A34 , 32'h00024749 , 32'h0000766A , 32'h0001E78D , 32'h0003E253 , 32'h0000171C , 32'hFFFE5917 , 32'hFFFEDA31 , 32'h000053EE , 32'hFFFFB99F , 32'hFFFF54B5 , 32'hFFFD7A79 , 32'hFFFED297 , 32'hFFFFE070 , 32'hFFFC1418 , 32'h00016D56 , 32'h00006033 , 32'hFFFD3118 , 32'hFFFF4828 , 32'h00001E87 , 32'h000008B5 , 32'h0000F3A8 , 32'hFFFF94C3 , 32'hFFFD45C1 , 32'hFFFFEA99 , 32'h00023272 , 32'hFFFD2D6A , 32'hFFFD503C , 32'h0002F2B0 , 32'h0002F0CB , 32'h0002BE47 , 32'h00007888 , 32'hFFFD41D7 , 32'hFFFBFBE3 , 32'hFFFED511 , 32'h000019A2 , 32'h0003F508 , 32'h00033738 , 32'h0000B0FF , 32'hFFFFE073 , 32'hFFFF8CFC , 32'h0006B4A1 , 32'h00000C46 , 32'hFFFDB7EA , 32'h0003DA10 , 32'h00000FFF , 32'h00013B9B , 32'hFFFE91CB , 32'hFFFF4BA3 , 32'h00008285 , 32'h00028755 , 32'hFFFC3515 , 32'h00015D50} , 
{32'hFFFEE053 , 32'hFFFE1028 , 32'hFFFEA739 , 32'h0001BA68 , 32'hFFFF54EF , 32'h0001E406 , 32'hFFFB7F05 , 32'h0001904F , 32'h0000DEA0 , 32'h00001808 , 32'h0002C6C7 , 32'h0001117F , 32'hFFFE49AD , 32'h00025752 , 32'hFFFE0F24 , 32'hFFF97842 , 32'h0002D84A , 32'hFFFEBB8E , 32'hFFFDE032 , 32'h000107CF , 32'h000265D8 , 32'h00023B8F , 32'hFFFD8372 , 32'h00008A06 , 32'h00012F68 , 32'h0000FB2C , 32'hFFFFE30D , 32'hFFFEB017 , 32'hFFFCB07D , 32'hFFFF14E6 , 32'h00033075 , 32'hFFFD3592 , 32'h0000FFC4 , 32'hFFFE7F59 , 32'hFFFF6512 , 32'hFFFE4736 , 32'hFFFE92CE , 32'h0005E833 , 32'hFFFE258B , 32'h00019929 , 32'hFFFCE81D , 32'hFFFADCD1 , 32'hFFFB5005 , 32'h00015240 , 32'h0004891E , 32'h00009587 , 32'h00039186 , 32'hFFFE8900 , 32'h0001D120 , 32'hFFFB8301 , 32'hFFFF427E , 32'hFFFCD66B , 32'h0002211A , 32'h00027A29 , 32'h0007B2EF , 32'hFFF778D9 , 32'hFFF8ED6C , 32'hFFFE159C , 32'hFFFA7F8F , 32'h000402FE , 32'hFFFA58C1 , 32'h0004ED4D , 32'h0001BDAD , 32'h00012FB0 , 32'hFFFF002F , 32'h0000417D , 32'h00014183 , 32'hFFFD357F , 32'h0002B376 , 32'h00002E31 , 32'h00029CC2 , 32'hFFFBB597 , 32'h00056708 , 32'hFFFB626D , 32'hFFFD38AE , 32'hFFFD3924 , 32'hFFFE7217 , 32'h00020C5A , 32'hFFFFBECA , 32'h0001904D , 32'h00050FAE , 32'h0001DD0A , 32'hFFFD2242 , 32'hFFFF4385 , 32'h00020BE2 , 32'hFFFCE7ED , 32'hFFFEEB23 , 32'h0000F5A0 , 32'h00009A5D , 32'hFFFB9687 , 32'hFFF850FF , 32'hFFFF6B2F , 32'hFFFE4A17 , 32'h000520E6 , 32'hFFFF604B , 32'hFFFDDC68 , 32'hFFFD4380 , 32'hFFFCD4C5 , 32'h0000353D , 32'hFFFE5701} , 
{32'h029AF8A4 , 32'hF22F42D0 , 32'h05DEC378 , 32'h00CB2F0F , 32'hF96B3408 , 32'h08036A40 , 32'h10590380 , 32'hF579CD10 , 32'hF696B860 , 32'hF51060F0 , 32'h0A0D0900 , 32'hFECE87F8 , 32'h005A31F5 , 32'h089E2250 , 32'hFA9D5268 , 32'hFC80B588 , 32'h038C34A8 , 32'h185100C0 , 32'h0CA85EB0 , 32'hFA150560 , 32'h029D9A38 , 32'hF6FC8BD0 , 32'h0281FF1C , 32'hFF28C8D3 , 32'h0971D130 , 32'h0F733E00 , 32'hFDD53D10 , 32'hFBC6B810 , 32'h015E34A8 , 32'hFFB2DF69 , 32'hFB67FC40 , 32'h057BEB28 , 32'hF82F9560 , 32'h047CA148 , 32'h037A050C , 32'h00E22E56 , 32'h0C01C620 , 32'hFF43093A , 32'h0380C8B8 , 32'h0CB64C70 , 32'h034764BC , 32'h06D8E2A0 , 32'hFBE39338 , 32'hF95EDDC8 , 32'hFE3B83E0 , 32'h024BA92C , 32'h07F88060 , 32'hFF157FF3 , 32'h0A3B4DD0 , 32'h02D65DD8 , 32'h063D8CE8 , 32'h03BAD928 , 32'hF7A65F80 , 32'hFB125F58 , 32'h018B7B08 , 32'hFD974F50 , 32'hFFBF4EC6 , 32'hFCB6838C , 32'h03FCF360 , 32'hFB7B20A0 , 32'hFB7B1E50 , 32'h0587BED0 , 32'h001F4AA5 , 32'h0A6B2810 , 32'h046BCBC8 , 32'h02CFF378 , 32'hFEEF8884 , 32'h06567FF8 , 32'hFC2A8588 , 32'h03C06B20 , 32'hFFFE4DF8 , 32'hFE6CEEE8 , 32'h04EAB2A8 , 32'h01FFCB78 , 32'h0293C850 , 32'h00C1ED90 , 32'h0252EDD0 , 32'hF8934C88 , 32'h0026EF49 , 32'h04887E38 , 32'h0297A3E0 , 32'h013CD1D4 , 32'h05214CA8 , 32'hFF8F291C , 32'hFF428B11 , 32'h03671878 , 32'hFF4D767D , 32'hFD984588 , 32'h025DD78C , 32'hFF61C3EC , 32'h000551E9 , 32'hFFFF3CB6 , 32'hFFFCDF30 , 32'h00024479 , 32'h0000C809 , 32'h00012248 , 32'h000084DA , 32'h000168E6 , 32'hFFFF096E , 32'h0000D35A} , 
{32'hF47AEB30 , 32'hCC259A40 , 32'h0C0E3D00 , 32'h070AFEE0 , 32'h027C5324 , 32'h11290360 , 32'h11C15DC0 , 32'h00CEBF28 , 32'hEF69F140 , 32'hF505B0F0 , 32'hF6ADF260 , 32'h18D81C00 , 32'h0C6B86E0 , 32'h05FEC740 , 32'h05B39650 , 32'hFF9CC494 , 32'hF5868240 , 32'h09745390 , 32'hF08CD4E0 , 32'hF6AF12D0 , 32'hFA34E930 , 32'hF282A570 , 32'h0BEF70B0 , 32'hFED04B18 , 32'hF63AC3B0 , 32'hFAA94380 , 32'h05ADA308 , 32'h0B9F0800 , 32'h038EB268 , 32'h06A41EA0 , 32'h083325F0 , 32'hF9908C80 , 32'h0F005F30 , 32'h0B3685B0 , 32'hF2836A10 , 32'h0054A02C , 32'hFD551048 , 32'h00836E06 , 32'hFE757AD4 , 32'hFE8E3C64 , 32'h0D6B5BF0 , 32'hFC413D48 , 32'hF9034E10 , 32'hF3BC5270 , 32'hF4A77610 , 32'h053E01B0 , 32'h064C1EE8 , 32'hFB874B50 , 32'h081CAD20 , 32'hFA5D73E8 , 32'hFBD59240 , 32'hFBBA7FA0 , 32'h00CB260C , 32'hFB8D5C68 , 32'h07A4A130 , 32'hFD7FE8D8 , 32'h077DBB08 , 32'hF74001A0 , 32'h08A8D880 , 32'hFE2C25D4 , 32'hFE421E88 , 32'hFFD156C3 , 32'h00CB704F , 32'h070F2940 , 32'hFA628B20 , 32'hF6DA63D0 , 32'hF7BE3C50 , 32'hF8EF00F8 , 32'hFE5CEFD0 , 32'h05931870 , 32'h04AC9528 , 32'hFF30A13C , 32'hFF3B430B , 32'h02E299B8 , 32'hF9718A70 , 32'h02E9E430 , 32'hFE42E7C8 , 32'hFFBF0E62 , 32'hFC71E50C , 32'h02CDD0A4 , 32'h021C1A78 , 32'h00E0F30C , 32'hFD668414 , 32'h0337FBB4 , 32'hFE5CD290 , 32'h015FE0E0 , 32'h00FE1B42 , 32'h04A89390 , 32'h0277972C , 32'h0068FBA4 , 32'hFFFEC8A5 , 32'h0005D002 , 32'hFFFF8CA4 , 32'hFFFF6D38 , 32'hFFFBCBC0 , 32'h0000CF97 , 32'hFFFFDDCF , 32'h0001C120 , 32'h00013036 , 32'hFFFEFE74} , 
{32'h090DDA30 , 32'hF9988DD0 , 32'h08AE7F70 , 32'hFD8E4E90 , 32'h00744F75 , 32'h052304B8 , 32'hFB464F30 , 32'h0172FD40 , 32'h026A3018 , 32'h04800A28 , 32'h050A1880 , 32'hFE3577B0 , 32'hFC1190F8 , 32'hFF99E4AD , 32'h058554F8 , 32'hFF4AF098 , 32'h069EBB90 , 32'h0844DFC0 , 32'h05FC9CB0 , 32'hFEDFA498 , 32'hFC32D1B0 , 32'hFF71EAB1 , 32'h06D65508 , 32'hFBAF6CD0 , 32'hFC934774 , 32'hF9EAA608 , 32'hFF9819CC , 32'h03D6B9C0 , 32'h02941FC0 , 32'hFFDE7C50 , 32'hFCBD2C90 , 32'h00F0FB17 , 32'hF927D990 , 32'h04A78D70 , 32'h01D39D98 , 32'hFE710330 , 32'h027A586C , 32'hFF947C15 , 32'hFBF023E8 , 32'hFE90D430 , 32'h008E6A38 , 32'hFEF22AD8 , 32'hFCC6BA4C , 32'h01CA9C80 , 32'hF8FCC5C8 , 32'h061EF5A8 , 32'hFF708480 , 32'hFDE25D84 , 32'h0796C600 , 32'hFFE45105 , 32'hFFF1E33B , 32'h06401D18 , 32'hFF0FFE40 , 32'h04BEC420 , 32'h00D55739 , 32'h0673A2F0 , 32'hFB905708 , 32'hFC30640C , 32'h04C004E8 , 32'h013C2410 , 32'hFEA22CE4 , 32'hFCB6C4A4 , 32'h028ABA54 , 32'hFD02DB2C , 32'h02390548 , 32'h05578AE8 , 32'h020EDB0C , 32'h0254E6C4 , 32'hFECD5898 , 32'hFFCF226C , 32'h01E34798 , 32'hFE60BD14 , 32'h03198714 , 32'hFD4236F8 , 32'h03F91C04 , 32'hFCE7275C , 32'h001915D4 , 32'hFDFC69F4 , 32'hFCA7B8BC , 32'h0157097C , 32'h0142314C , 32'h020F789C , 32'hFF62312F , 32'hFDDD6080 , 32'h027893AC , 32'hFF6E9F58 , 32'hFE2BCF2C , 32'h03ADBF08 , 32'h02A4A54C , 32'h002F1492 , 32'hFFFC1472 , 32'hFFFEDF1E , 32'hFFFFB2C5 , 32'h00023625 , 32'h0003A549 , 32'hFFFF2D70 , 32'hFFFE8210 , 32'hFFFDBCDD , 32'h0001FF32 , 32'h0000235F} , 
{32'h04F31928 , 32'h0828E020 , 32'hF7F0AC30 , 32'h03DBC114 , 32'h01548924 , 32'h0793F540 , 32'hFB659A30 , 32'hFD9AAAC4 , 32'h02329008 , 32'h02D8E3A4 , 32'hFB3D5860 , 32'hFCEF7678 , 32'hFBF82BB0 , 32'hF5DEFC20 , 32'hFFBF3106 , 32'h02C694F0 , 32'h07513D90 , 32'h015D2EF4 , 32'h02CD6F44 , 32'h07EC1160 , 32'h0988AF20 , 32'hFAC809D0 , 32'hFBC382C8 , 32'hF98B9268 , 32'h07B19768 , 32'h02ADB598 , 32'h0012ACB3 , 32'hFE0AB86C , 32'hFA861A58 , 32'hFA17A0B0 , 32'hFEEAF84C , 32'hFFD439A3 , 32'hFD62CE94 , 32'hFA98DA10 , 32'h0068EB2E , 32'hFFE62498 , 32'hFED982C4 , 32'hFE60A194 , 32'hFEBE6160 , 32'h01028AC0 , 32'hFB668FD8 , 32'hFCCDB240 , 32'h0282877C , 32'hFF7CF0FE , 32'hFEAA1054 , 32'h03E97A70 , 32'h0599A700 , 32'h012388FC , 32'h00C2A412 , 32'h007ACF39 , 32'h067AA210 , 32'hFE62653C , 32'hFF327621 , 32'h009116D2 , 32'h0091A784 , 32'h010CB360 , 32'hF9FFED18 , 32'h044169D0 , 32'h004A8850 , 32'h03AE44C0 , 32'hFFD46F63 , 32'hFD4504FC , 32'h0463DAB0 , 32'h03AD3AE0 , 32'hFA76D288 , 32'hFCC5C968 , 32'hFE640934 , 32'h080106C0 , 32'hFB33E950 , 32'h060AB460 , 32'h030E774C , 32'hFEEA5988 , 32'h00AB5C3A , 32'hFE990868 , 32'hFB83EFA8 , 32'hFF2B77AF , 32'hFD15A21C , 32'hFFADE39B , 32'hFF1ADD9D , 32'hF72148B0 , 32'h021FC5A0 , 32'h0295FDBC , 32'h05825020 , 32'h01A45784 , 32'hFF01AC54 , 32'h03492BE0 , 32'hFF92CCFB , 32'h01C73FFC , 32'hFE738A0C , 32'hFFDFE74E , 32'hFFFFB655 , 32'h000416D0 , 32'hFFFF8912 , 32'hFFFE03A8 , 32'hFFFC4979 , 32'h0003119D , 32'hFFFC71C1 , 32'hFFFE25D8 , 32'hFFFD630A , 32'h0003AEDA} , 
{32'hFFFF7454 , 32'hFFFD6A48 , 32'hFFFE6EFF , 32'h00007176 , 32'h00024ABD , 32'h00036BDF , 32'h00037C4A , 32'hFFFE4F01 , 32'hFFFF3309 , 32'hFFFD5CC3 , 32'hFFFF817C , 32'hFFFFC050 , 32'h0001089D , 32'h000142AA , 32'h0003653D , 32'h0000C779 , 32'hFFFED3FB , 32'h00017D15 , 32'hFFFF86E4 , 32'hFFFE8CB3 , 32'h0000388E , 32'hFFFBC6CF , 32'h0003FE1B , 32'hFFFCD237 , 32'hFFFBF1C7 , 32'hFFFE3F5B , 32'h00006C41 , 32'h0002D0AB , 32'h000108AB , 32'h000241B5 , 32'hFFF8606B , 32'h00035432 , 32'h0003936C , 32'h00016B87 , 32'hFFFF747A , 32'h0002E7E3 , 32'hFFFFDA8E , 32'hFFFF81D9 , 32'hFFFF6266 , 32'hFFFF9EDB , 32'h000166ED , 32'h00003A0D , 32'hFFFE245E , 32'h00048FDC , 32'hFFFDDD83 , 32'h0000E1C1 , 32'hFFFF137A , 32'hFFFB888E , 32'h00015037 , 32'hFFFD1D32 , 32'hFFFDC625 , 32'h0002CE40 , 32'h0000A499 , 32'hFFFFCBC7 , 32'h0002AE8C , 32'hFFFEFBB3 , 32'hFFFEFE58 , 32'hFFFBB8F8 , 32'hFFFE2A37 , 32'h0001A85B , 32'h000082D3 , 32'hFFFD4E93 , 32'h00034AE7 , 32'hFFFEF9E9 , 32'hFFFE02FE , 32'hFFFF15DB , 32'hFFFDF1DF , 32'hFFFF4EFD , 32'h00031D2B , 32'h00004401 , 32'h000093A7 , 32'hFFFB1F7B , 32'hFFFF2C64 , 32'hFFFFF803 , 32'h0003E106 , 32'hFFFD336F , 32'hFFFE6C36 , 32'hFFFE4D76 , 32'hFFFEFEB8 , 32'hFFFD2EB5 , 32'hFFFC7313 , 32'hFFFF01C3 , 32'hFFFF8DE1 , 32'h00018970 , 32'h0002982B , 32'h0000426E , 32'hFFFC03D3 , 32'hFFFA3F0A , 32'h0002EB8D , 32'h00038A11 , 32'h00015B27 , 32'hFFFC26BA , 32'h0001E283 , 32'h0000BC61 , 32'hFFFD02B1 , 32'hFFFC668A , 32'hFFFB35E9 , 32'hFFFE4CDE , 32'h00019A07 , 32'hFFFEC40A} , 
{32'h0000EF7F , 32'h00034058 , 32'hFFFD7AE9 , 32'h00047808 , 32'h00023080 , 32'h0000F744 , 32'h000134E8 , 32'h00049BA7 , 32'hFFFD099B , 32'h00005142 , 32'hFFFC70DA , 32'hFFFE2AFF , 32'hFFFD348F , 32'h0002090B , 32'hFFFA95C1 , 32'hFFFEC723 , 32'h000216C4 , 32'h00042B9E , 32'hFFFC5FA0 , 32'h00009B33 , 32'hFFFF58B8 , 32'h00026E97 , 32'h0000EDAF , 32'hFFFEFAF8 , 32'h0000676A , 32'h0001599A , 32'h000160BF , 32'h000096DF , 32'hFFFC731A , 32'hFFF7D180 , 32'h0000B9F2 , 32'hFFF99C49 , 32'h00016A55 , 32'h00026272 , 32'h000017BA , 32'h000220CC , 32'h0000AE79 , 32'hFFFFC95C , 32'h000198F0 , 32'h0001A74C , 32'hFFFE0E03 , 32'hFFFFC5F0 , 32'hFFFEE4E3 , 32'hFFFD9B90 , 32'hFFFCC825 , 32'hFFF9BECE , 32'hFFFCA44C , 32'h00014C6E , 32'h0004E9F3 , 32'h0004248F , 32'h00011EC8 , 32'hFFFC80D5 , 32'hFFFF64FC , 32'hFFFD817A , 32'h0006532A , 32'hFFFD0902 , 32'hFFFE4474 , 32'hFFF824D6 , 32'h00025EEB , 32'h000092C3 , 32'h000285AF , 32'h0001CF39 , 32'hFFFF5134 , 32'hFFFFBD62 , 32'h00049210 , 32'h0000C977 , 32'hFFFE6709 , 32'hFFFF4F2B , 32'h0002F6B6 , 32'hFFFF8ED0 , 32'h000177D5 , 32'h00023B92 , 32'hFFFC4015 , 32'hFFF9F473 , 32'hFFFB679A , 32'hFFFCACF9 , 32'h00013E8C , 32'h00017216 , 32'h00026A63 , 32'hFFFFE9E4 , 32'hFFFBC23D , 32'h00029F2C , 32'hFFFDEE5F , 32'h000425FA , 32'hFFFE8F8B , 32'h00011B57 , 32'hFFFEF616 , 32'hFFFD2FC7 , 32'h00024E74 , 32'h000216F3 , 32'hFFFF655B , 32'h00024E9D , 32'hFFFF7B95 , 32'h00034D14 , 32'hFFFEAB64 , 32'hFFFC4EAE , 32'hFFFF4D06 , 32'h00029A55 , 32'h00048FE6 , 32'hFFFEF291} , 
{32'hF5DF52A0 , 32'hF882A140 , 32'hF5E69FC0 , 32'h0943C840 , 32'h01F3E5B8 , 32'hFD0AF6B8 , 32'hF5E56D00 , 32'h05E2DB20 , 32'hF0437520 , 32'h05084AA8 , 32'hFB6DF538 , 32'hFD342EF8 , 32'h03F41E9C , 32'hF89E2AC0 , 32'h0141A8B4 , 32'h06C67050 , 32'h08DAB1E0 , 32'h05994090 , 32'hF2035250 , 32'h05098640 , 32'h047F6758 , 32'hFBC24ED8 , 32'h03EBD8B0 , 32'hF93D2728 , 32'hFED52704 , 32'h019FE118 , 32'hF60C3C60 , 32'h06B038F0 , 32'hFE287924 , 32'hF9464000 , 32'h031715C8 , 32'hFB644168 , 32'hF7474050 , 32'h03EA0F44 , 32'h0D6D85E0 , 32'hFEB4F52C , 32'hFD0D538C , 32'h07BE2300 , 32'hFF7E4EA4 , 32'h0A7E3F20 , 32'hFD664094 , 32'hFAA71A68 , 32'h003E8441 , 32'hFF4EEA9B , 32'h096E1F70 , 32'h02D87860 , 32'hF6C26600 , 32'h05850698 , 32'h0206A5A4 , 32'h09562E70 , 32'h01F368E0 , 32'h0EC26930 , 32'hFC38F090 , 32'hFDB46F50 , 32'h06597FD0 , 32'h0D361610 , 32'h00825D47 , 32'h072516A8 , 32'hFFDB64C2 , 32'hFEC95CF8 , 32'h0124764C , 32'h01195154 , 32'hFE647EFC , 32'h0847FE70 , 32'hF6987BF0 , 32'h02DE6D3C , 32'hF4DC6860 , 32'hFFED7AAF , 32'hFC6AA308 , 32'hFB04B920 , 32'h0734CE68 , 32'h01E23FEC , 32'hFEFBC708 , 32'hFE9F5F28 , 32'h004CF17D , 32'h03060610 , 32'hFF8E1DD4 , 32'h03213460 , 32'hFAC05E50 , 32'h02884E70 , 32'hFE463BA0 , 32'h04FF4D88 , 32'h025530D4 , 32'h0491C820 , 32'hFB7136F8 , 32'h03AF1A20 , 32'h02E40640 , 32'hFE646E34 , 32'hFEF0E9AC , 32'h00B84E31 , 32'h0002FAB4 , 32'h00022C4C , 32'hFFFE5273 , 32'hFFFFA16C , 32'hFFFDE8D7 , 32'hFFFFB947 , 32'h00002FB9 , 32'hFFFF2500 , 32'hFFFD2DA9 , 32'h00009B0E} , 
{32'h0001010E , 32'h00020756 , 32'hFFFF2BD3 , 32'h000353F4 , 32'hFFFD8194 , 32'hFFFC1F41 , 32'hFFFF1936 , 32'h0001C3E0 , 32'hFFFF5BB5 , 32'h0002AD49 , 32'hFFFF05DA , 32'hFFFDEF64 , 32'h0001604C , 32'h0002B789 , 32'hFFFD7543 , 32'hFFFEE876 , 32'h000339FE , 32'hFFFD87B7 , 32'h00006D1B , 32'h0000EB41 , 32'hFFFF28C8 , 32'h0001D4C8 , 32'h0000ACE1 , 32'h000071ED , 32'h000158FC , 32'h0002D002 , 32'h0003252C , 32'hFFFE8084 , 32'h0000265C , 32'hFFFF6AA2 , 32'h0000B25F , 32'h0003CBAA , 32'h0001B43F , 32'hFFFD5F64 , 32'hFFFF4471 , 32'h00001AB5 , 32'hFFFFBE1B , 32'hFFFA8C2D , 32'h0001527A , 32'h0002D3B0 , 32'h00002099 , 32'h0002B94C , 32'h000236FE , 32'h00081866 , 32'hFFFE133B , 32'hFFFDDA83 , 32'hFFFF36AD , 32'h0002E6FD , 32'h00008264 , 32'h00045FEF , 32'h00005363 , 32'h00049F0C , 32'hFFFAE59E , 32'hFFFC59C1 , 32'h00000D54 , 32'hFFFD8E21 , 32'h0002BEEA , 32'hFFFE31A8 , 32'h0002BBFA , 32'h0001AA70 , 32'h0001BB6D , 32'h00030C9C , 32'h0001C23C , 32'hFFFE5E86 , 32'hFFFF812B , 32'h0002459D , 32'h00009158 , 32'hFFFE25D0 , 32'h00019AF6 , 32'hFFFD5D23 , 32'h00001AAC , 32'hFFFD0FC2 , 32'h0000381A , 32'hFFFBB60F , 32'h00027859 , 32'hFFFECB92 , 32'h000116C2 , 32'h000144E8 , 32'hFFFE1ACC , 32'hFFFBDEE5 , 32'hFFFB4DFF , 32'hFFFC8349 , 32'hFFFF48C7 , 32'hFFFF1A92 , 32'h0001629E , 32'h0000DB08 , 32'hFFFAFB98 , 32'hFFFAC168 , 32'h00018FAA , 32'hFFFF4311 , 32'h0001054B , 32'h0002119E , 32'h0000A2B4 , 32'hFFFE8631 , 32'h0003C50D , 32'h00014AA0 , 32'hFFFB69B2 , 32'h0000E525 , 32'h00017E06 , 32'hFFFF0CFD} , 
{32'hFFFCF58F , 32'hFFFC9551 , 32'hFFFE1AD3 , 32'h00022D4F , 32'h0001D312 , 32'hFFFC285E , 32'hFFFFDDDB , 32'h000286B4 , 32'h000103A7 , 32'h000008B0 , 32'h000213CB , 32'h0002B231 , 32'h000017B2 , 32'hFFFED6B3 , 32'h0002E045 , 32'h000098CD , 32'hFFFBB772 , 32'hFFFF5449 , 32'hFFFF1394 , 32'h0003B065 , 32'h00013C41 , 32'hFFF9F006 , 32'h00015574 , 32'hFFFFC34D , 32'h00024683 , 32'h00005A9D , 32'hFFFFE171 , 32'hFFFDEFB9 , 32'hFFFB6F46 , 32'h0002945A , 32'hFFFCC6F2 , 32'h00061902 , 32'hFFFFF7E1 , 32'h000024D8 , 32'hFFFBC2EE , 32'h000118F2 , 32'hFFFF21C6 , 32'h00020E30 , 32'h0001D13A , 32'h000383DC , 32'hFFFF169D , 32'h00028CAF , 32'h0003F68B , 32'h000294A3 , 32'hFFFE69BF , 32'hFFFFAC17 , 32'hFFFF0753 , 32'h000158C5 , 32'h0001BFBC , 32'h00016FB7 , 32'hFFFD80EF , 32'h00038BEC , 32'hFFFC1BB5 , 32'hFFFC5540 , 32'h0000AF6F , 32'h00015CC4 , 32'hFFFD6C0F , 32'h0003B471 , 32'hFFFDA654 , 32'hFFFC47ED , 32'h000022CC , 32'hFFFB8F98 , 32'h0000FE9D , 32'hFFFE3608 , 32'h00027FE2 , 32'h00010415 , 32'hFFFFC4E7 , 32'h00038A9C , 32'h00055ABC , 32'h00026049 , 32'hFFFFE587 , 32'h0001726D , 32'hFFFF837F , 32'hFFFD3A21 , 32'h00036F4F , 32'h000561A3 , 32'hFFFDED96 , 32'h00026A44 , 32'h000269AC , 32'hFFFDB7C6 , 32'h0000C083 , 32'h00019AA8 , 32'hFFFE9243 , 32'hFFFE8DFD , 32'h000376DD , 32'h00016ABF , 32'hFFFE8FB4 , 32'hFFFF2B3C , 32'h0000D6A6 , 32'h000056FF , 32'hFFFB935A , 32'h00042405 , 32'hFFFF09F7 , 32'h0005B5A3 , 32'hFFFE27D9 , 32'h000112F4 , 32'hFFFD81E3 , 32'hFFFC9B4E , 32'hFFFE9696 , 32'h000195C0} , 
{32'h048BE350 , 32'hF237A820 , 32'h06964388 , 32'hEB32DE80 , 32'h0DAEFC30 , 32'hF23A5560 , 32'hFE8DDE48 , 32'hFFBD7EFC , 32'h0B893AA0 , 32'hFC4D5B50 , 32'h0216FC74 , 32'hFF1B8824 , 32'hF3E0B1E0 , 32'h05245670 , 32'hFF355766 , 32'hFC3A2AC8 , 32'hF4022AF0 , 32'hFB9C4638 , 32'h00E405F8 , 32'hF7386890 , 32'hFB31E060 , 32'h04936850 , 32'hF73B16C0 , 32'h069F9028 , 32'h0BA01320 , 32'hFBCAC2B8 , 32'hFAD06988 , 32'hFBAE1980 , 32'h07180BF8 , 32'h066B36C0 , 32'hF7940C00 , 32'h040F0EF0 , 32'h00D5020A , 32'hFB8F8938 , 32'hF53CE3A0 , 32'hFF0AEBDD , 32'h076F0048 , 32'h08C8B7F0 , 32'h020B01D8 , 32'hFCB4B034 , 32'h06D665E8 , 32'h08A57D90 , 32'hFD8BB9D0 , 32'hF779AE20 , 32'h067E5728 , 32'hFDFC40F0 , 32'h005AB9FD , 32'hFAE3C108 , 32'hFB1F0C50 , 32'h034B1744 , 32'hFB2E5A20 , 32'hFBD69768 , 32'hFA647630 , 32'h010362D8 , 32'h0647EDF8 , 32'hFB4F71C0 , 32'hF9BD7608 , 32'hFFF2B479 , 32'hFCE19B08 , 32'h0364ACAC , 32'h0653A198 , 32'h0109E3F4 , 32'hFCC6811C , 32'hFB97D458 , 32'hFF50D00B , 32'h06C37A60 , 32'hFDE921D8 , 32'hFDFC567C , 32'h045D8260 , 32'hF952FDD8 , 32'h022A73F0 , 32'hFF6133CA , 32'h07CC2138 , 32'hF94DBA80 , 32'hF3C08560 , 32'hF82CB8C0 , 32'hFD45B114 , 32'hFAB09898 , 32'h012B7A1C , 32'h02CD2310 , 32'hFC9AF1F8 , 32'hFF390641 , 32'hFDC15FFC , 32'hFDA95C88 , 32'hFC67F274 , 32'hFDDE7474 , 32'h0091BAEC , 32'hFCC70B54 , 32'h04AD64E8 , 32'h003786BE , 32'hFFFC3B69 , 32'hFFFE6B2E , 32'h00026254 , 32'hFFFF80CC , 32'hFFFF767E , 32'hFFFE90BC , 32'hFFFEBE67 , 32'hFFFF847D , 32'h00002C68 , 32'h00013022} , 
{32'hFFFC6056 , 32'h0002EBE0 , 32'h00017684 , 32'h00042AFE , 32'h00009A8A , 32'hFFFF083E , 32'hFFFFB3BD , 32'hFFFCDFCE , 32'h0000E4C7 , 32'hFFFA70EE , 32'h00023B53 , 32'h00014DE4 , 32'h00039E6F , 32'hFFFB69FE , 32'h0000F415 , 32'h000119DF , 32'h0000BDE2 , 32'h0003832C , 32'hFFFEF176 , 32'hFFFFF400 , 32'h0003FC7E , 32'h0005BCEF , 32'h00016E79 , 32'hFFFFA0D2 , 32'h00051179 , 32'h0001C551 , 32'h00001F6B , 32'hFFFE8453 , 32'h00004750 , 32'hFFFF1DC1 , 32'h000530D4 , 32'hFFFFB87C , 32'hFFFFABDE , 32'h00003E34 , 32'hFFFF7515 , 32'hFFFE2E9E , 32'hFFFD81FA , 32'hFFFBABE1 , 32'h00044E82 , 32'h00030A82 , 32'h000249A5 , 32'h0000D730 , 32'h00006FBB , 32'hFFFECDD7 , 32'hFFFE1C9E , 32'hFFFE482E , 32'h0001B79A , 32'h000247A5 , 32'hFFFC3692 , 32'hFFFE2771 , 32'h000009DD , 32'hFFFC754B , 32'hFFFEA522 , 32'h00003416 , 32'h000238EA , 32'hFFFF5B25 , 32'hFFFE7F0A , 32'hFFFD0997 , 32'hFFFDDD3B , 32'hFFFD3FFD , 32'hFFFF5AA4 , 32'h00019C0C , 32'hFFFE0783 , 32'hFFFEF766 , 32'hFFFF3FEF , 32'h000163AE , 32'h000176CD , 32'hFFF9CF96 , 32'hFFFEA946 , 32'h00013EC9 , 32'h00022AA8 , 32'h00002D9E , 32'h0002060A , 32'h00006CA8 , 32'h00019F2B , 32'hFFFD84E4 , 32'h0003EBF2 , 32'hFFFB5879 , 32'h0007E4B5 , 32'h00014A5B , 32'h0001849D , 32'h00022797 , 32'h0002F53A , 32'h0004585D , 32'h000083A8 , 32'h0000D7E4 , 32'h00001EEB , 32'hFFFE997C , 32'h00016A05 , 32'hFFFCAF23 , 32'h0004EA88 , 32'h0002F5FD , 32'h00009050 , 32'hFFFFAAEB , 32'h000206F5 , 32'h000126CE , 32'h0002C5A9 , 32'h0002F110 , 32'hFFFF9438 , 32'hFFFB8B4C} , 
{32'hFFFBEB47 , 32'h00030A57 , 32'h000082A3 , 32'h00037EBC , 32'hFFFFB286 , 32'h0000D60E , 32'hFFFEAAB2 , 32'hFFFF6FA0 , 32'h0000B22E , 32'hFFFE5CB4 , 32'h0000DA8E , 32'hFFFC013B , 32'hFFFEDBD6 , 32'h0004BD80 , 32'h0003D005 , 32'h00005FCB , 32'h0002873F , 32'h0000F279 , 32'hFFFF1050 , 32'h00036838 , 32'h0001992C , 32'h0001BD32 , 32'h000391DB , 32'hFFFB8886 , 32'hFFF9A483 , 32'h0001838A , 32'h0000B5C3 , 32'h000051B7 , 32'hFFF97A6C , 32'h000217D2 , 32'h0001691B , 32'hFFFF7CC2 , 32'hFFFFD691 , 32'hFFFE5D90 , 32'hFFFEBA39 , 32'h00000657 , 32'h0000A79C , 32'hFFFE815A , 32'hFFFEECA8 , 32'h00004D4E , 32'hFFFBDD74 , 32'h0002927D , 32'h0001802D , 32'hFFFDB23D , 32'h00066588 , 32'hFFFE4326 , 32'hFFFEC2A1 , 32'hFFFF2378 , 32'hFFFEB651 , 32'h00001182 , 32'hFFFF3AC7 , 32'h0003B6FD , 32'h0004A83A , 32'hFFFABA63 , 32'h00004FF6 , 32'h0000230A , 32'h00008FD2 , 32'hFFFF75F4 , 32'hFFFD87FD , 32'h0001E6E9 , 32'hFFFDD906 , 32'hFFFCF6D2 , 32'h0000EC15 , 32'h000249B5 , 32'hFFFB60B9 , 32'h00018410 , 32'h0003FFB2 , 32'hFFFD396B , 32'hFFFF2152 , 32'hFFFF0269 , 32'hFFFEAB17 , 32'hFFFBD60A , 32'hFFFF65B5 , 32'hFFFE7C0C , 32'h0003B978 , 32'h00050B5A , 32'hFFFDC67F , 32'hFFFBDCC3 , 32'hFFFC336A , 32'hFFFE972A , 32'hFFFAC2F9 , 32'hFFFF239D , 32'h000420F6 , 32'h000081D0 , 32'hFFFF2AFC , 32'h0004FB40 , 32'hFFFD485E , 32'hFFFDAC3E , 32'hFFFF0B9F , 32'hFFFFF4F4 , 32'hFFFEF4E9 , 32'hFFFACC59 , 32'h00044632 , 32'hFFFF8363 , 32'hFFFA41D7 , 32'hFFFF9EEF , 32'hFFFFFD4C , 32'h000119B8 , 32'h00003828 , 32'hFFFE7481} , 
{32'h0F478820 , 32'hFC959DA8 , 32'hF48E04B0 , 32'hCB5DED40 , 32'h1E15A480 , 32'hFE1A7804 , 32'hFBF7F010 , 32'h0EF62ED0 , 32'h0157D690 , 32'hFBB8C8D0 , 32'hFF240733 , 32'h0DB49FB0 , 32'hF8456950 , 32'h08C80530 , 32'hF7EE9770 , 32'h1C1529A0 , 32'hF2291DF0 , 32'h019C6C98 , 32'h144686C0 , 32'hF97E7788 , 32'hF98F34D0 , 32'hF54A44A0 , 32'hFF4B8320 , 32'hFC1CA398 , 32'hF1501670 , 32'hF4278BC0 , 32'hFC3B818C , 32'hFF194E80 , 32'h072FA308 , 32'hFB827700 , 32'h0EEF13F0 , 32'hFAC46E28 , 32'hF87A4A28 , 32'h01F02284 , 32'h01BE3800 , 32'h0A6B7AC0 , 32'h0B3518D0 , 32'h10E42E60 , 32'h099C1B50 , 32'hED51B5C0 , 32'h0807EC70 , 32'h10EC19C0 , 32'h0095DBEC , 32'hF5FC9C90 , 32'hF7D060E0 , 32'h0F080BC0 , 32'hFBBF1138 , 32'h037954B4 , 32'hF6007FF0 , 32'hFF9420BE , 32'hF9B29430 , 32'h00CC2F1E , 32'hFB62A490 , 32'hFA27E310 , 32'hFF2C2FE5 , 32'hF52CC060 , 32'h0296F92C , 32'h06EBCB58 , 32'hF80E95C8 , 32'h037C0F94 , 32'h07BAE808 , 32'h001EAA4C , 32'h02E86398 , 32'hFF8BBC30 , 32'hF9D0CD60 , 32'h021D8B00 , 32'h0395A118 , 32'h06D84F40 , 32'h06AD8180 , 32'h03DF00B4 , 32'h0AFB1710 , 32'h04193228 , 32'hFF41C078 , 32'hFCC96124 , 32'h04A78970 , 32'h055E8DC8 , 32'h014D9E44 , 32'h022AEEF4 , 32'hFD4CDFA0 , 32'h0243E2F0 , 32'h00853DB8 , 32'hFECBBFA8 , 32'hFE92C274 , 32'hFE6EDA64 , 32'h02045538 , 32'hFDF0FD98 , 32'hFFDC7882 , 32'hFF1F0E88 , 32'hFCB90E94 , 32'h00C8F99D , 32'h0001E8D7 , 32'hFFFE5F21 , 32'hFFFECB62 , 32'hFFFF75B3 , 32'h0002191E , 32'h0002251B , 32'h0000FE1A , 32'h00015BD6 , 32'h00010C75 , 32'h0001941F} , 
{32'h0000C6C6 , 32'hFFFC67FB , 32'hFFFDA3C6 , 32'hFFFFFA70 , 32'hFFFA763C , 32'h0000FC7D , 32'h00043C6A , 32'h0003471E , 32'hFFFF7637 , 32'h0002940C , 32'hFFFFFD8C , 32'hFFFD6F58 , 32'h00045AFC , 32'h000044FA , 32'hFFFE9D9D , 32'h00018991 , 32'hFFFFF5D8 , 32'h00029137 , 32'hFFF8A983 , 32'h00005406 , 32'h0000F9AD , 32'h0000CCFA , 32'hFFF90A67 , 32'hFFFFF47C , 32'h0002A189 , 32'hFFFAABEA , 32'h0001F918 , 32'hFFFBF175 , 32'hFFFF7399 , 32'h0002CC1D , 32'hFFFEAF93 , 32'hFFFEB21D , 32'hFFFD19B2 , 32'hFFFDF653 , 32'h0007DBBA , 32'h0003D765 , 32'h0000AED2 , 32'h000032F0 , 32'hFFFEC700 , 32'hFFFC19C1 , 32'hFFFB243C , 32'hFFFFCAD0 , 32'hFFFFD265 , 32'hFFFA1A3E , 32'hFFFEDE84 , 32'hFFFEA4BF , 32'hFFF9990B , 32'h0002BD73 , 32'hFFFFFF9C , 32'h000452F9 , 32'hFFFDF4DF , 32'h0002D752 , 32'h0001EDC0 , 32'hFFFC1C63 , 32'h0004E566 , 32'h00012FFA , 32'h00026410 , 32'h0000A596 , 32'h000473C1 , 32'hFFFBC48F , 32'hFFFCC89E , 32'h00011919 , 32'h00048A48 , 32'hFFFBF1E8 , 32'hFFFC7FC3 , 32'hFFFD6B99 , 32'hFFFC4327 , 32'hFFFD7AA2 , 32'hFFF9C6B4 , 32'h000238B8 , 32'h00039176 , 32'hFFFD84DA , 32'h00029E07 , 32'h0000488C , 32'hFFFC61A5 , 32'hFFFC2B22 , 32'hFFFEA748 , 32'h0001F3B2 , 32'h00009749 , 32'hFFFFCC9E , 32'h00063518 , 32'h000000D0 , 32'hFFFF8ACB , 32'hFFFC9D28 , 32'hFFFF0883 , 32'h0001C346 , 32'h0000A53E , 32'h00050B6B , 32'h000443E2 , 32'h0003BE72 , 32'h00011493 , 32'hFFFE0CD1 , 32'h00007751 , 32'hFFFF51B5 , 32'h00038DEA , 32'hFFFD8FB9 , 32'h00001B96 , 32'hFFFEF3F3 , 32'hFFFF4E3E , 32'h0003EC49} , 
{32'h2255E080 , 32'h0AF7B020 , 32'hFE490558 , 32'hF5ACDA80 , 32'h0002496C , 32'hDF8DAE80 , 32'hF61312A0 , 32'h0830C550 , 32'h18D06800 , 32'hF733DC60 , 32'hF989D618 , 32'h061E11F0 , 32'h01F96048 , 32'hE8FB5680 , 32'hF01B09A0 , 32'h04AFBE78 , 32'hF391AF50 , 32'h1F6A6200 , 32'h044B2C50 , 32'h16C56460 , 32'h11287D40 , 32'hF0F2E230 , 32'h0D34B730 , 32'hFFCD69F5 , 32'h0A4D0AF0 , 32'h0650D868 , 32'h0332B5C4 , 32'h09E8A1C0 , 32'hF17B8A10 , 32'hFBC93EA0 , 32'hFFA76716 , 32'hFC76F96C , 32'h0ED48E10 , 32'h03F0A664 , 32'h00595B8E , 32'h030FEB3C , 32'h04ED94A8 , 32'hFE7440EC , 32'h0466DE90 , 32'hFF7B75BC , 32'h0AEF75E0 , 32'h0074B9D8 , 32'hFE5CFEC8 , 32'h01F17C24 , 32'h01B0A42C , 32'h029FA08C , 32'h022BA494 , 32'h1986DA60 , 32'h00BE067D , 32'hFE8A3300 , 32'h04CFDA38 , 32'h012F5380 , 32'hFA032430 , 32'h0AB3DEE0 , 32'h034E3D3C , 32'hFE10E028 , 32'h04CC1650 , 32'h04A3F230 , 32'h0E3A5530 , 32'h00342A9F , 32'hFB0200A8 , 32'h0366B200 , 32'hF3234510 , 32'h028A6088 , 32'hFC27B6B4 , 32'h00A82532 , 32'hFCC397C8 , 32'hFF947C0F , 32'h04EF7DA8 , 32'h06DE1E68 , 32'hFE3D2FF4 , 32'h09371D50 , 32'hFE7641EC , 32'hFD229224 , 32'h006BB9BC , 32'hFB52E100 , 32'hFF0EF11B , 32'h05164D50 , 32'h0308A6B0 , 32'hFB4B6388 , 32'hFEB8D6A8 , 32'hFE75E238 , 32'hFDBD1504 , 32'hFD884FB4 , 32'hFF3A7A88 , 32'h0277FAD4 , 32'hFCF1D1F0 , 32'hFED39728 , 32'hFE677558 , 32'hFF79DD75 , 32'h00010986 , 32'h00031ECE , 32'h000097E5 , 32'h00023013 , 32'hFFFD8701 , 32'h00024066 , 32'hFFFEBCF1 , 32'h0000D552 , 32'hFFFFE9F6 , 32'hFFFFD2A3} , 
{32'h03376058 , 32'h02A1C838 , 32'hFF3DA661 , 32'h0086D5C7 , 32'h0547F158 , 32'h063B9640 , 32'h026899D8 , 32'hF90D2E20 , 32'h043D46E8 , 32'h02187A24 , 32'h02A006AC , 32'hFD9FAE8C , 32'h029F944C , 32'h0393EB2C , 32'h0081A4BD , 32'h00F95568 , 32'h008C41CD , 32'h0053A6B0 , 32'hF77204B0 , 32'h00165FAB , 32'h03D47F24 , 32'hF68DF870 , 32'hFF13867F , 32'hFE8CCF54 , 32'hFF30FA56 , 32'h00724F2B , 32'hFD039B38 , 32'h004B8668 , 32'hFA9F3E60 , 32'h0073EC1A , 32'h021CE944 , 32'h01B5E358 , 32'h053A4188 , 32'h006E9CC7 , 32'hF9110A08 , 32'hFA0DE318 , 32'h00A71BD2 , 32'hFA7ACB28 , 32'hFE7E9E9C , 32'h0079F52F , 32'h0276F608 , 32'hFFDC2D86 , 32'h0181018C , 32'hFD95AD68 , 32'hFDB24F00 , 32'h06A2DE08 , 32'hFFC8B78C , 32'h03C13990 , 32'hFF59C6EF , 32'hFF1A8699 , 32'hFF69F777 , 32'h019FBFF8 , 32'hFAD0F968 , 32'h00349B4C , 32'h030FBB64 , 32'h014CBB80 , 32'h01C0D574 , 32'h04E82440 , 32'hFB8E5AF8 , 32'h02263C04 , 32'h02B9E6B8 , 32'hFF20C2EF , 32'h01922A20 , 32'hFD70D1B0 , 32'hFEEF7AB8 , 32'h01507ECC , 32'hFB332FD8 , 32'h00AFD535 , 32'h01F07DD4 , 32'hFF89BD8F , 32'h00A773DF , 32'hFB0E3678 , 32'h00D48B01 , 32'hFF466066 , 32'hFFB8CABC , 32'hFDA490EC , 32'hFEE2B16C , 32'h00A13C19 , 32'h0415C9A8 , 32'hFE4E9DC4 , 32'h02A4999C , 32'h0294F754 , 32'hFF70759C , 32'hFE6628E8 , 32'h0017A060 , 32'h0047A545 , 32'hFD7D48B0 , 32'h01D6A7FC , 32'h003990BC , 32'hFF8FF7CA , 32'hFFFE18A6 , 32'h000127DC , 32'hFFFF3A84 , 32'hFFFF1908 , 32'hFFFD20BA , 32'hFFFEC085 , 32'h0002FA90 , 32'hFFFE834E , 32'h0000276E , 32'hFFFE5849} , 
{32'hFFFBE8C8 , 32'hFFFD245A , 32'hFFFDA808 , 32'h0003FC15 , 32'hFFFE034A , 32'h0001CADE , 32'h00004504 , 32'hFFFE95B1 , 32'h00063669 , 32'h0000D041 , 32'hFFFDBED3 , 32'h0000170D , 32'h00018A7E , 32'hFFFE4CBF , 32'hFFFC6E62 , 32'h00001B99 , 32'h000327A8 , 32'h0001C6F7 , 32'h00035824 , 32'h00008C4C , 32'hFFFEFCD2 , 32'h0000AA1E , 32'h0001311F , 32'h0001BD93 , 32'hFFFC1982 , 32'hFFFDF8DB , 32'hFFFEE8B1 , 32'h00007B6F , 32'h00008A44 , 32'hFFFE7DDA , 32'hFFFF0146 , 32'h00056BA7 , 32'h00037FB2 , 32'h000061DA , 32'h0004CDEF , 32'h00002A3B , 32'hFFFE6E33 , 32'h0001C3DF , 32'hFFFD3AC6 , 32'hFFFC4521 , 32'h000158E8 , 32'h0002E8CB , 32'hFFFE939C , 32'hFFFF22F6 , 32'h0000132A , 32'h0001FD9D , 32'h0003938D , 32'h0001473B , 32'hFFFFE669 , 32'hFFFC8E2E , 32'h00013E74 , 32'h00035BE3 , 32'h0003413F , 32'h0001B0E4 , 32'h00011960 , 32'hFFFE88D8 , 32'h000271F6 , 32'hFFFF8FE6 , 32'h00017D0F , 32'h000098F8 , 32'hFFFE36C4 , 32'hFFFE2DAF , 32'h000157E9 , 32'h0001F0F2 , 32'h000224A9 , 32'h0001931F , 32'hFFFE4EBB , 32'h00006D7C , 32'h0001D9A7 , 32'h0002500C , 32'hFFFE3388 , 32'h00012EA8 , 32'hFFFAC4DE , 32'h00006102 , 32'h0000FE2D , 32'hFFFA3E3B , 32'hFFFCFC89 , 32'h000253F9 , 32'hFFFED1E1 , 32'h00005BCD , 32'h0002ACCA , 32'hFFFE7583 , 32'hFFFE7582 , 32'hFFFE84DF , 32'hFFFDDB0F , 32'h00023EC6 , 32'h00024994 , 32'hFFFDD630 , 32'hFFFE2075 , 32'h000222B4 , 32'h000418B7 , 32'hFFFE2C91 , 32'h000074ED , 32'h000037C1 , 32'hFFFEA32A , 32'h0003C4F8 , 32'hFFFBAB30 , 32'hFFFBD71E , 32'h0001E405 , 32'hFFFF362D} , 
{32'h0001C1CD , 32'hFFFDCBC8 , 32'hFFFD3649 , 32'h000035DC , 32'h000302F9 , 32'hFFFE6CA0 , 32'hFFFE6226 , 32'hFFFE4970 , 32'hFFFE1A3D , 32'hFFFB2E54 , 32'h00000FC1 , 32'h000263D8 , 32'hFFFE0764 , 32'h000087A7 , 32'h0002B872 , 32'hFFFF7E4B , 32'h0002B463 , 32'hFFFDDB47 , 32'hFFFC1FA0 , 32'hFFFFDAFF , 32'h00031E33 , 32'hFFFFD1A0 , 32'h0002964C , 32'h00017833 , 32'h00038F8B , 32'h0001D168 , 32'h000333A0 , 32'h00017E0A , 32'h0000B987 , 32'hFFFDA1DC , 32'h00002C0A , 32'hFFFF03C6 , 32'hFFFB6EB7 , 32'h0003F3BC , 32'hFFFCC4A0 , 32'h0001E215 , 32'hFFFCA1D8 , 32'hFFFFBDDF , 32'hFFFE4273 , 32'h00002146 , 32'hFFFBBB09 , 32'hFFFE2399 , 32'h0002340B , 32'hFFFF336E , 32'h0000C360 , 32'hFFFE3E38 , 32'hFFFEF3F6 , 32'hFFFD140E , 32'h00009144 , 32'h0002BC83 , 32'h00000094 , 32'hFFFF6EE2 , 32'hFFFF2FBD , 32'h0000B1C6 , 32'h0000D818 , 32'h0004193A , 32'h000286D8 , 32'hFFFBA139 , 32'h000083B8 , 32'h0001A08B , 32'hFFFF8093 , 32'h00052F68 , 32'hFFFDCD77 , 32'hFFFE310E , 32'h0000B7BD , 32'h00056523 , 32'hFFFE033B , 32'hFFFF8EF2 , 32'h00012446 , 32'hFFFE15CC , 32'hFFFAAE32 , 32'h0000788A , 32'hFFFF3691 , 32'hFFFE64D7 , 32'hFFF83216 , 32'hFFFE013B , 32'h000145EA , 32'h00000159 , 32'hFFFC5D50 , 32'h00007AE4 , 32'h0001BD24 , 32'hFFFDEC4A , 32'h0003FBCB , 32'h00018221 , 32'h00002687 , 32'hFFFBC324 , 32'hFFFFADB7 , 32'hFFFF7109 , 32'h0003355A , 32'h0000AF69 , 32'h0003D063 , 32'h000138F4 , 32'h0001F2E4 , 32'h00024EE2 , 32'h0000DEE0 , 32'h0000C2F7 , 32'h00040F1B , 32'hFFFE4086 , 32'h0002BF75 , 32'hFFFEFFB0} , 
{32'hFFFDB542 , 32'hFFFBFD0B , 32'hFFFEE485 , 32'h00020E77 , 32'h000553CE , 32'hFFFF9251 , 32'hFFFF9854 , 32'hFFFD5BEF , 32'hFFFEBB2E , 32'hFFFF7CC5 , 32'h00051D28 , 32'hFFFEBC8E , 32'hFFFD6117 , 32'hFFFE0435 , 32'h00018617 , 32'h00006B84 , 32'h0002CFD1 , 32'h0001A77A , 32'hFFFE6839 , 32'h0002F6E0 , 32'h00014822 , 32'hFFFF0982 , 32'hFFFF995C , 32'hFFFDB95D , 32'h0003817E , 32'h0000B5A3 , 32'hFFFD9D9D , 32'hFFFFF738 , 32'hFFFA5079 , 32'h0002B357 , 32'hFFFDDCEB , 32'h00009EE6 , 32'hFFFFAEEC , 32'hFFFFDAE9 , 32'h0000F72D , 32'h0000FEF7 , 32'hFFFEEA5A , 32'hFFFF548B , 32'hFFFA6E29 , 32'hFFFF8219 , 32'h000253DF , 32'h0000A7A4 , 32'hFFFF7A2E , 32'hFFFF4A59 , 32'h0000651E , 32'h00024E37 , 32'h0001023C , 32'hFFFE0C85 , 32'h00015C7E , 32'hFFFECB6E , 32'hFFFFA7F4 , 32'h0001481D , 32'h0002FB3C , 32'h0000EBB0 , 32'hFFFEAA71 , 32'hFFFF83ED , 32'h000241FD , 32'hFFFF099C , 32'hFFFE3412 , 32'hFFFE724A , 32'hFFFED09B , 32'hFFFE8F3F , 32'hFFFC6BBD , 32'h0002D7DC , 32'h0007FFCC , 32'h000414E9 , 32'hFFFE056D , 32'h00021FBD , 32'h000463C4 , 32'h0003B17C , 32'h0002B01E , 32'h00035453 , 32'hFFFAAD47 , 32'h00041CF5 , 32'h0000E750 , 32'h00005651 , 32'h00010A93 , 32'hFFFFB910 , 32'h00003A0A , 32'h0000D740 , 32'h000099B5 , 32'h0000B326 , 32'hFFFFC605 , 32'hFFFDDC09 , 32'hFFFFC387 , 32'hFFFF96B9 , 32'hFFFE9585 , 32'hFFFFA522 , 32'h00010CBA , 32'hFFFA446C , 32'h000713E6 , 32'h00007524 , 32'h0004653B , 32'hFFFDAEF9 , 32'h00011ABF , 32'h0004B4A2 , 32'hFFFFDFD3 , 32'hFFFD4502 , 32'hFFFDAE8F , 32'h00018DA6} , 
{32'h30E92840 , 32'h0CFD6D70 , 32'h18CBB0A0 , 32'hDAAA68C0 , 32'h1C7D1580 , 32'hF1829020 , 32'hEE5EA920 , 32'hE6495200 , 32'h03D24704 , 32'hF9362538 , 32'h0BC85BA0 , 32'h215EE2C0 , 32'hFB813AC8 , 32'h01F61E74 , 32'h04CC4A58 , 32'h0A50C2D0 , 32'hECDC7B20 , 32'h0A7DE440 , 32'h05621610 , 32'hFCCE5E0C , 32'hFEEBBB48 , 32'hFE5BD77C , 32'h17F55100 , 32'hFEEB7C9C , 32'h0AEFD560 , 32'h040641A0 , 32'hFC384C40 , 32'hFF3A7084 , 32'h00243752 , 32'hECF4DE20 , 32'hFCCBF07C , 32'h00DC84DA , 32'hFE61018C , 32'h063CA590 , 32'h0A8EABA0 , 32'h0397D06C , 32'h199B9280 , 32'h07841D98 , 32'h070E9540 , 32'h062D5A58 , 32'hF36910F0 , 32'hF4D96210 , 32'h014258B8 , 32'hF2C9C3B0 , 32'hF41AAB40 , 32'hF949F2F8 , 32'h05A08E10 , 32'hF9FB9898 , 32'hFEC14F64 , 32'hFEAA15AC , 32'hFE96A120 , 32'hFC2D65D8 , 32'hFFB8970D , 32'hFC24FA58 , 32'h00507BD8 , 32'h0572BAF0 , 32'hF860D7D0 , 32'h031819DC , 32'h09281B70 , 32'h07910A18 , 32'h0930D170 , 32'h03C3FA90 , 32'h0B949100 , 32'h0018FA87 , 32'hFD930C00 , 32'hFDE49D24 , 32'h0EF163F0 , 32'hFE34021C , 32'hF774A620 , 32'hFFE286EC , 32'h015B4238 , 32'hFE6FBA0C , 32'h011CE0DC , 32'hFDB27E78 , 32'hFFE6E2F1 , 32'h051AB4E8 , 32'h03251318 , 32'hFEC64B48 , 32'h00DF972C , 32'hFED925B4 , 32'hFE1579A8 , 32'hFDDF66B0 , 32'h02C4ACAC , 32'h016603F8 , 32'h04249CD0 , 32'hFF804B0C , 32'h00B2E30B , 32'h00AEB396 , 32'h0216C854 , 32'h00E0FD76 , 32'h0002D8FB , 32'hFFFEAC4D , 32'hFFFF4264 , 32'hFFFF95CD , 32'hFFFDEBAD , 32'hFFFECB88 , 32'hFFFC4D3A , 32'h00013155 , 32'hFFFE1B9D , 32'hFFFF8344} , 
{32'hE8D0A6E0 , 32'h09A95350 , 32'hEFA82500 , 32'h07915E68 , 32'hEB446620 , 32'h188DC860 , 32'hFF95F35D , 32'hFCAC9B18 , 32'h10CA1BC0 , 32'hEF757D80 , 32'hE74C9FA0 , 32'h08126070 , 32'hE7F76940 , 32'hF10074B0 , 32'hF809B520 , 32'hEA4DAA20 , 32'hFB559E10 , 32'h0311EF34 , 32'hF163CB90 , 32'hFEC86744 , 32'h008C31E5 , 32'hF8627F88 , 32'h061010A0 , 32'hF8A9BD68 , 32'hF493B800 , 32'hFA4EC8C0 , 32'hF51F5B50 , 32'hF9F4CEB0 , 32'h005B4DA9 , 32'h1200CC40 , 32'hF45FEBE0 , 32'hFFC0C102 , 32'hF87D02C0 , 32'hF957D478 , 32'h002AC691 , 32'h029A476C , 32'h10BCC2C0 , 32'h02879E70 , 32'h0BEBF0E0 , 32'hFE48DAC0 , 32'hFD979834 , 32'hFF3F5E29 , 32'hF693ED40 , 32'hF55AFE00 , 32'h06529FC0 , 32'hFE432AEC , 32'h074CB6F0 , 32'h093195E0 , 32'hF1A50B00 , 32'h005B6A30 , 32'h03C7FE18 , 32'h0695C4F8 , 32'hFBD91A30 , 32'h03EF8D5C , 32'hF9A419D0 , 32'hF7322B50 , 32'h039E701C , 32'h01FA8CB4 , 32'h03B717D0 , 32'h0305C710 , 32'h01D32ED0 , 32'h012572C0 , 32'hFD02BF40 , 32'h03F67B78 , 32'hFA0EDD98 , 32'hFD0AB8C0 , 32'hFBB2D8C8 , 32'h06C26490 , 32'h076FE560 , 32'hFE24AA54 , 32'h01D20DEC , 32'hFFDEA2C6 , 32'hFF32C98B , 32'hF8E36970 , 32'h074B6060 , 32'h03C72E74 , 32'hFD0A0300 , 32'hFF08D272 , 32'h02EBDD60 , 32'hFEC23734 , 32'hFE23672C , 32'hFC64CBF8 , 32'h006408F0 , 32'h0155A720 , 32'hFFCA7034 , 32'h008C2153 , 32'hFF3FDC4E , 32'h0123F1C8 , 32'hFD43047C , 32'hFFFE2E0B , 32'hFFFBDF68 , 32'h0000E354 , 32'h00017352 , 32'hFFFF7C42 , 32'hFFFF4E60 , 32'h0001E8A6 , 32'hFFFE6FC1 , 32'hFFFFDDC0 , 32'hFFFFC407 , 32'hFFFC3D4F} , 
{32'hF289C060 , 32'h01708D24 , 32'h0A1C9E60 , 32'hEE95AB60 , 32'hF1E1FA50 , 32'hFE604BE0 , 32'hFECF38F0 , 32'hFA0E6000 , 32'h0C525C80 , 32'hF3478920 , 32'hF9BD44E0 , 32'h12B98080 , 32'hF5D45E00 , 32'hF2D26E70 , 32'hEFFD4AA0 , 32'h16D49700 , 32'h0A65C010 , 32'h00A07B6C , 32'hED82D200 , 32'hF65833E0 , 32'h09F1D1E0 , 32'h084C1790 , 32'h068B92F8 , 32'hF7880EB0 , 32'h0C67CFE0 , 32'h012768AC , 32'hE6776000 , 32'h056EA658 , 32'hF9CB2048 , 32'hF3D7ADB0 , 32'hFACC2538 , 32'hF7321170 , 32'h07B5DF08 , 32'hFD57D39C , 32'hF61E4500 , 32'h084A0080 , 32'h069E9908 , 32'h05BF74E8 , 32'hFC75709C , 32'h019C4CB8 , 32'h03C9C930 , 32'h03EC6304 , 32'h0581C300 , 32'h016DC82C , 32'hFC7D6D24 , 32'hF4050F10 , 32'h023165B8 , 32'h05854680 , 32'hFE44E378 , 32'h0D3DDCD0 , 32'h0BC8E6D0 , 32'h080615B0 , 32'h01B19E78 , 32'h0AB7AA20 , 32'h094656D0 , 32'hF90A92A0 , 32'h02710ACC , 32'h07BBD618 , 32'hFAA1F938 , 32'h01979868 , 32'h02002DE4 , 32'hFBF1CEF8 , 32'h035BF400 , 32'hFF6C82AB , 32'h028478C8 , 32'hF87A1020 , 32'h0328C3D8 , 32'h083BB4B0 , 32'hFDC4E408 , 32'h0394986C , 32'h007F58E6 , 32'h03D669FC , 32'h03F8CBC8 , 32'h06A15A78 , 32'h050CFE18 , 32'hFC535F34 , 32'hFD918734 , 32'hFF4B478B , 32'hFAF5DDF8 , 32'h0487F620 , 32'h002C83B2 , 32'h03BF3FA0 , 32'hFE4C3B2C , 32'hFFCC6142 , 32'h011C9E7C , 32'hFE683088 , 32'h001C890E , 32'hFDEB847C , 32'hFD4D9D8C , 32'hFF96B632 , 32'hFFFFF15C , 32'hFFFE819E , 32'hFFFEC3E2 , 32'h00022B3F , 32'h0001CE27 , 32'h00023E7E , 32'h00010C89 , 32'h000256DD , 32'hFFFE9579 , 32'hFFFDCD27} , 
{32'h0AD28B30 , 32'h005F74EC , 32'h161780E0 , 32'hDA166640 , 32'h0E67DE00 , 32'hFAD41010 , 32'h1F6096C0 , 32'hFC313840 , 32'hEB3161E0 , 32'h016AF8D8 , 32'h080E66B0 , 32'h0A832070 , 32'hFADC8D00 , 32'h0C31AE80 , 32'hFA95D600 , 32'h07281D08 , 32'h021EB0F0 , 32'hF81E78F8 , 32'h0AB3A8B0 , 32'h03E4F22C , 32'h19121DA0 , 32'h0613D898 , 32'hFEFE5B48 , 32'hF2CAC420 , 32'h136F7B60 , 32'hFA906F68 , 32'hFD24C290 , 32'hFA598E98 , 32'hF98C1DF8 , 32'h02121594 , 32'hF8AB7108 , 32'h0CAA82A0 , 32'h044A26C0 , 32'hF20EF270 , 32'hFDCF0954 , 32'hEF632720 , 32'hF9E8A7E0 , 32'hFAA1FB18 , 32'h02F5973C , 32'hF4E44900 , 32'h020F60DC , 32'h10C0ADC0 , 32'h064EDA60 , 32'hFA3DD018 , 32'hFC2AFC7C , 32'h01F113C4 , 32'h085E7B40 , 32'h0377A074 , 32'h039419E8 , 32'hEF9AD160 , 32'h002E3D40 , 32'hFBBBB378 , 32'hF92EFE60 , 32'h0889AFF0 , 32'hFEA67200 , 32'h07421068 , 32'h02ABC680 , 32'hF7E27650 , 32'hFE3A0404 , 32'hFF1A5D90 , 32'hFDA5B3F4 , 32'h0532F7F8 , 32'hFA6C4400 , 32'h04B53AE0 , 32'hFEF96214 , 32'hFFFBDD75 , 32'h03B4BAE8 , 32'h03C41E7C , 32'hFC8E4638 , 32'hF62EF040 , 32'hFEE6A56C , 32'h08C1AE40 , 32'hFE211114 , 32'h05FCDBC8 , 32'hFA8293E0 , 32'hF9E06CD0 , 32'hF990D510 , 32'h079A0C18 , 32'h0587C8C8 , 32'h01C7DFF0 , 32'h0540B8A8 , 32'h01491758 , 32'h0087089F , 32'h07F9F5E0 , 32'h0109E9EC , 32'h0040484F , 32'h058AD868 , 32'h0206D618 , 32'h00356681 , 32'hFFA0152B , 32'h000199DD , 32'h00008EAF , 32'hFFFE5110 , 32'h0002058C , 32'h0000F244 , 32'h00003E70 , 32'hFFFEB0E6 , 32'hFFFEC4A4 , 32'hFFFF15E0 , 32'hFFFF5EFD} , 
{32'hFFFE13EF , 32'hFFFE58C8 , 32'hFFFF26EA , 32'h0003AE67 , 32'hFFFB5F09 , 32'h0002EC3B , 32'h000338C4 , 32'h0001077B , 32'hFFFD713F , 32'hFFF7542F , 32'h0004BD28 , 32'h00000B7B , 32'h0000FBD4 , 32'h00035BC0 , 32'hFFFBFEDA , 32'hFFFB6BD1 , 32'h0003EC4C , 32'h00004502 , 32'hFFFF54C0 , 32'h00028C14 , 32'hFFFE4417 , 32'h000163AF , 32'h00006888 , 32'h0004EE1F , 32'h0003835B , 32'hFFFD1319 , 32'hFFFF8840 , 32'h00033530 , 32'h0000E45B , 32'h00003D62 , 32'h0003391C , 32'hFFFD378B , 32'h00035881 , 32'hFFFF2108 , 32'hFFFE6B11 , 32'hFFFEFCFD , 32'h0001C63A , 32'hFFFD694C , 32'hFFF7387E , 32'hFFFBC93E , 32'hFFFF3523 , 32'hFFFD7467 , 32'hFFFFAA7F , 32'hFFFA9B4F , 32'h0001091D , 32'hFFFAFCD7 , 32'hFFFD72E2 , 32'hFFFEC828 , 32'hFFFCCC3D , 32'hFFFF2BEC , 32'h00034A11 , 32'hFFFDC132 , 32'h000505A4 , 32'hFFFF71D5 , 32'hFFFE20E1 , 32'hFFFC7668 , 32'h000337C9 , 32'h00000A25 , 32'hFFFAD5F8 , 32'hFFFD5C18 , 32'hFFFE9CB1 , 32'hFFFF09DD , 32'h0001AACA , 32'h000259BB , 32'h0001407B , 32'h00011FC8 , 32'hFFFF3F95 , 32'h0001F216 , 32'h00011F85 , 32'hFFFEF661 , 32'h00015E96 , 32'hFFFD5706 , 32'hFFFEAD93 , 32'hFFFCEBFE , 32'hFFFFBB04 , 32'h0002E9E7 , 32'hFFFC723C , 32'hFFFAF0DE , 32'hFFFFD19B , 32'h0002E576 , 32'h00016D99 , 32'h00056A65 , 32'hFFFE5238 , 32'h000465E4 , 32'hFFFE0FC6 , 32'h0003C66C , 32'hFFFBD213 , 32'h000298D6 , 32'h0000CEAC , 32'hFFFF59FF , 32'hFFFF8A6F , 32'hFFFF7662 , 32'h00014547 , 32'h00007447 , 32'hFFFCB254 , 32'h0002F29D , 32'h0001099C , 32'h0001A00A , 32'hFFFEF278 , 32'hFFFE15A1} , 
{32'hE6E99800 , 32'h3DD22480 , 32'h3FA6E100 , 32'h53CB2080 , 32'hF5BA4B80 , 32'hCB87C580 , 32'hB0FC3E80 , 32'h05C17B58 , 32'hF148F530 , 32'hFF6E11DF , 32'h0CAF8610 , 32'hEDB643C0 , 32'hD9020E40 , 32'h1739EFA0 , 32'h0F37BD00 , 32'hF2895870 , 32'hF68B4220 , 32'h05B66760 , 32'hF074AC10 , 32'hF1C53870 , 32'h0E729550 , 32'h011D025C , 32'h1337F320 , 32'hF7B1C620 , 32'hE3260620 , 32'h02A401E8 , 32'hF5E9B420 , 32'hE6D29680 , 32'hF43C8360 , 32'h07336410 , 32'h09BC4E10 , 32'hF8805E88 , 32'hF9A20CA8 , 32'hF3A8F4A0 , 32'h02FC0A58 , 32'h05823CB0 , 32'hF2948CE0 , 32'hFDA00B64 , 32'h05E26090 , 32'h068CA700 , 32'h0CC14560 , 32'h1A4BEBE0 , 32'h027ABF54 , 32'hF9C77CB0 , 32'hFE36A1D8 , 32'h04818D40 , 32'hFA177838 , 32'h010ED9D0 , 32'hFF901E06 , 32'hFF6C448A , 32'hF9946DB0 , 32'hF9CD4DC0 , 32'h046E15B8 , 32'hF8B585B0 , 32'h01180FC0 , 32'h0AA11B30 , 32'h0034739B , 32'h01BAF56C , 32'h00812777 , 32'h00F5B3D4 , 32'hFE8D4264 , 32'hF950EF50 , 32'h03A697A0 , 32'h010C5118 , 32'hFDD94BE8 , 32'h00110B34 , 32'h098A3710 , 32'h06007830 , 32'hFE2B7D54 , 32'hFD7EDB40 , 32'h02B36E84 , 32'hFC60388C , 32'hFFACE669 , 32'hFDCE3AD4 , 32'hFF1E9B42 , 32'hF9E80EB0 , 32'hFFB0C808 , 32'h027D76C4 , 32'hF7B65870 , 32'hFDAE5CF8 , 32'hFDCA0334 , 32'hFB174560 , 32'h007A0BE3 , 32'hFD95E2C4 , 32'hFE3184BC , 32'h058C3E70 , 32'h007C8094 , 32'hFFDB178E , 32'hFE48CDBC , 32'h00785FAD , 32'hFFFEAF6F , 32'h00022D42 , 32'h0000B947 , 32'h0001D243 , 32'hFFFFA97D , 32'hFFFCFE85 , 32'h0000D820 , 32'h00002473 , 32'h00012600 , 32'hFFFEB87F} , 
{32'h000516E9 , 32'h0003DE6E , 32'hFFFDC2B7 , 32'hFFFD5E6E , 32'h0000E80E , 32'h00015E19 , 32'hFFFD3556 , 32'h00034880 , 32'hFFFB0C77 , 32'hFFFDF246 , 32'hFFFAF693 , 32'h0004EF89 , 32'hFFFCC2E9 , 32'h0001AA62 , 32'h00039B1C , 32'hFFFC9048 , 32'hFFFF6E4E , 32'h00005897 , 32'h0004BCCD , 32'h0001462D , 32'hFFFCFBFF , 32'h0002BA6D , 32'h00013D0E , 32'h00022A33 , 32'hFFFCFA12 , 32'h000194BF , 32'h000333C7 , 32'hFFFDAE55 , 32'hFFFAE9C1 , 32'h00043265 , 32'hFFFF5E73 , 32'h00035654 , 32'h0001F6B0 , 32'h00010662 , 32'h00029279 , 32'hFFFD066F , 32'hFFFEBF65 , 32'hFFFAA4D6 , 32'hFFF932FC , 32'hFFFE6325 , 32'hFFFE9B9F , 32'h000066E9 , 32'h0002F23A , 32'hFFFA4C4D , 32'h0001A105 , 32'hFFFFAEC5 , 32'hFFFFDC7B , 32'h0000BF70 , 32'hFFFEC621 , 32'hFFFEC880 , 32'hFFFE40A9 , 32'hFFFEF197 , 32'hFFFE821D , 32'h0001B787 , 32'hFFFF216C , 32'h00029344 , 32'h0002E5D8 , 32'hFFFF9EE7 , 32'h0001A94C , 32'h0001FBD7 , 32'hFFFFF783 , 32'h00034E1D , 32'hFFFEA2DF , 32'hFFFE65FB , 32'hFFFD8ED2 , 32'hFFFFFA46 , 32'h0003B7C9 , 32'h0002773D , 32'hFFFFFF16 , 32'h0003C812 , 32'h00017C77 , 32'hFFFEB0B5 , 32'hFFFCC392 , 32'hFFFE1B8B , 32'h0002AD24 , 32'h00006A8C , 32'hFFFE4006 , 32'hFFFD7E55 , 32'h0000CD48 , 32'h000469C0 , 32'h0001DD93 , 32'hFFFE4D4B , 32'h000003EB , 32'h00022021 , 32'h0001C896 , 32'h00026CBD , 32'h0000A46E , 32'hFFFE662C , 32'h0001C37E , 32'hFFFB3C00 , 32'hFFFE6A6A , 32'h00067B79 , 32'h00005E90 , 32'hFFFB6D21 , 32'hFFFFB0C1 , 32'h0000ED7A , 32'hFFFF5E34 , 32'h00032F55 , 32'h0000A304 , 32'h00033418} , 
{32'hFFFF313E , 32'h00010478 , 32'h00063827 , 32'hFFFD1D02 , 32'h00004A5C , 32'hFFFC9AC7 , 32'hFFFDBBDA , 32'h00029333 , 32'h0004EF04 , 32'hFFF9B2A5 , 32'h000070A3 , 32'h000033B4 , 32'hFFFFBED6 , 32'h000018CD , 32'hFFFFD4B4 , 32'hFFFFF0E6 , 32'hFFFF7018 , 32'hFFFEB885 , 32'h0001ECE2 , 32'h00017A23 , 32'hFFFE31F8 , 32'h0002D1D6 , 32'h00006E01 , 32'hFFFF883B , 32'hFFFD5F1C , 32'hFFFD798D , 32'h000396F5 , 32'h00020148 , 32'hFFFE9B2E , 32'hFFFD1C25 , 32'hFFFCD247 , 32'hFFFA0CBC , 32'hFFFFFD9C , 32'hFFFD3088 , 32'h0003D6E9 , 32'hFFFB5684 , 32'hFFFB1B09 , 32'h00030AA5 , 32'h000034FF , 32'h00001B39 , 32'hFFF91E8B , 32'hFFFED585 , 32'hFFFB5047 , 32'h00027D4F , 32'hFFFC19BC , 32'hFFFDFD8A , 32'hFFFF7A05 , 32'h00021CD5 , 32'h00014EEB , 32'hFFFFDF9F , 32'h00031C02 , 32'hFFFE6499 , 32'hFFFF1ED7 , 32'h0000C1D5 , 32'hFFFACD21 , 32'hFFFFE632 , 32'h00035121 , 32'hFFFF5021 , 32'hFFFEE8F1 , 32'hFFFF03D6 , 32'h00002879 , 32'h0004BE84 , 32'hFFFED0E3 , 32'h0000392C , 32'h0002D32B , 32'hFFFC5D8B , 32'hFFFDAFA8 , 32'hFFFE5B1F , 32'hFFFE5DEF , 32'hFFFE4DAE , 32'hFFFFE798 , 32'h0003BE33 , 32'hFFFE87CC , 32'h0001BF94 , 32'hFFFFBA44 , 32'hFFFDFE0D , 32'h00035810 , 32'hFFFD40C3 , 32'hFFFD935D , 32'hFFFCF2EC , 32'h0002C940 , 32'h00021D3E , 32'h00002A85 , 32'hFFFD8162 , 32'hFFFE1E21 , 32'h000171C0 , 32'hFFFA0267 , 32'hFFFC4EE4 , 32'hFFFF56C0 , 32'h00016039 , 32'hFFFD878E , 32'h00005495 , 32'h000283FB , 32'hFFFA2941 , 32'hFFFF038E , 32'hFFFF75D2 , 32'h000440DA , 32'h000303F6 , 32'hFFFCDBE8 , 32'h000154E6} , 
{32'h3110E700 , 32'hF2E5C360 , 32'h0083CE9B , 32'hE7F435C0 , 32'h38EE5980 , 32'h15540F00 , 32'hEB585840 , 32'hFD2D3AB8 , 32'hEF60F060 , 32'h162E2E00 , 32'h0E5FA710 , 32'hF8B1F300 , 32'hFF452171 , 32'hDBF4F5C0 , 32'h128C2220 , 32'hFF8DCF83 , 32'h09D1DCF0 , 32'h0C0F69C0 , 32'hFF6551F0 , 32'hEA45C700 , 32'h0B354760 , 32'h083F9FE0 , 32'h0C93A7D0 , 32'h05BCF0A8 , 32'hF66BEEE0 , 32'h13B8FCA0 , 32'h0529B5C8 , 32'hFEB432C4 , 32'hF5D9AE90 , 32'hFC9F9070 , 32'h04044A60 , 32'hF1E0A730 , 32'hFBFD55A8 , 32'h08D6D6E0 , 32'hF8BA5F98 , 32'hF45F0E70 , 32'hE75B8760 , 32'hFADF7478 , 32'hFAF728E8 , 32'h0A58F6D0 , 32'h067F3EA8 , 32'hFBA16E30 , 32'hF6734D30 , 32'h050BA678 , 32'hFE353748 , 32'hF5935500 , 32'h03824794 , 32'h06B39128 , 32'hFDB5186C , 32'h06EC23B0 , 32'h0BF5EDA0 , 32'hF6701020 , 32'hFC9FF690 , 32'hFFA8D475 , 32'h11556400 , 32'hFAF7FCD8 , 32'h00995C93 , 32'hF1758760 , 32'h06112300 , 32'hFEB1C41C , 32'h023278A8 , 32'h04DD72B8 , 32'hFB2B05C0 , 32'hF94DE830 , 32'hFC8F1B64 , 32'h04E1A450 , 32'hFDF47038 , 32'h05D9E828 , 32'h08B580E0 , 32'hFE422B60 , 32'hFBC92030 , 32'hFD673A64 , 32'h02E17984 , 32'h05373B00 , 32'hFE6B56D4 , 32'hFEF87C04 , 32'hFE934080 , 32'hFE749044 , 32'h05C3A210 , 32'hFDFCD4F4 , 32'h019511F4 , 32'hFE1EF1C0 , 32'h0056482B , 32'h017F9B90 , 32'h05AF5938 , 32'h02D8A898 , 32'h01F1DF84 , 32'hFFDCF53C , 32'hFEC01BE8 , 32'h04344800 , 32'h00014AF5 , 32'hFFFF60D1 , 32'hFFFEFF75 , 32'hFFFFEEF3 , 32'h00015E23 , 32'h0000414E , 32'h000023B6 , 32'h0000DE42 , 32'hFFFF6847 , 32'hFFFF5304} , 
{32'h08B7F7C0 , 32'hFC28A238 , 32'hF6B91C30 , 32'hEC3508A0 , 32'hF77D9900 , 32'hF9A706D8 , 32'h01E1E8BC , 32'hF5CFB2A0 , 32'hF3526E70 , 32'h06700B28 , 32'h0B6ABEC0 , 32'h0744ED10 , 32'h041DEF00 , 32'hEE65B040 , 32'hFF67CE14 , 32'h08D418B0 , 32'h01F27044 , 32'hFDA463D4 , 32'hF2CD4DB0 , 32'h046F1B10 , 32'hF061BEB0 , 32'h03CC7790 , 32'hF7C71500 , 32'h00B9A322 , 32'h04A442F0 , 32'h0D747740 , 32'hFCD873DC , 32'h0259B410 , 32'hF8B87E70 , 32'h0415A1B8 , 32'hFDDF17D8 , 32'hFE419D84 , 32'hFE9735DC , 32'hFE34A090 , 32'h0740AF98 , 32'hFE206D1C , 32'h04A6AC78 , 32'hFC051050 , 32'hFF46735F , 32'h00C3F6FD , 32'h01360748 , 32'h02758A24 , 32'hF9C201E0 , 32'h085AFD00 , 32'hFD4DF070 , 32'h008ACCD9 , 32'hFD769B40 , 32'hFE529158 , 32'hFA879B68 , 32'h0285F65C , 32'h00FDC5A3 , 32'h0057164A , 32'h04E283E0 , 32'hFE8F0B78 , 32'hF99ACC18 , 32'h04DD9CC8 , 32'h02ECA9B8 , 32'h02546DC4 , 32'hFECB2290 , 32'hFA9AB8D8 , 32'h0343247C , 32'hFA8F72B8 , 32'hFF8B3C47 , 32'hFAB893F0 , 32'h0075DBD3 , 32'h046E5390 , 32'hFA6B85C8 , 32'h0DE0F380 , 32'h070AD7D8 , 32'hFFB2A0AB , 32'h011BF714 , 32'hFECD7A4C , 32'h06BFDEA0 , 32'hF9A84BA8 , 32'hFC56BA50 , 32'hFBD34360 , 32'h0361A140 , 32'h0155520C , 32'hFBB40F38 , 32'h05BBA938 , 32'hFDC5AF34 , 32'hFEEF7970 , 32'hFA4C8D10 , 32'hFFF53482 , 32'hFD98635C , 32'h00E1FCCE , 32'h03EA0564 , 32'h0002489B , 32'h0042A799 , 32'hFFCFBFA2 , 32'h0002A57F , 32'hFFFE43D4 , 32'h0000200A , 32'hFFFFF380 , 32'hFFFD0105 , 32'h00008363 , 32'h00029303 , 32'hFFFE5022 , 32'h000111A9 , 32'h00010FA2} , 
{32'h0962CCB0 , 32'hF902BD70 , 32'hFDBBCE30 , 32'hEF6C76C0 , 32'h09283E10 , 32'hEDF07720 , 32'hFCC91E8C , 32'hF11F5690 , 32'h0759DE10 , 32'h045AEAB8 , 32'hFDFF90A8 , 32'h0997F840 , 32'h0C1F4E80 , 32'hF16C0130 , 32'hF8ADAE90 , 32'hF203AEE0 , 32'h06356D88 , 32'hFA1CB680 , 32'hF2440640 , 32'h03A75F50 , 32'hF7FAEC00 , 32'hF63F6CA0 , 32'h0CC16550 , 32'hFFE38513 , 32'h03FFB12C , 32'hFD1B93DC , 32'hFFE68E96 , 32'hFEFC01D4 , 32'h081ABB30 , 32'h0B467360 , 32'hF42D40F0 , 32'h0149C164 , 32'hF65FE950 , 32'hEE988460 , 32'hF9AA9080 , 32'h0BA15690 , 32'hECE4EF00 , 32'hFFAF1ACE , 32'h01BFB158 , 32'hFE555B1C , 32'h02B4D5D0 , 32'hFE053C6C , 32'h013CA810 , 32'h0919DFB0 , 32'hF7C916A0 , 32'h03BB4AD4 , 32'hFFFA8707 , 32'hFA2F8C08 , 32'hFB7D2650 , 32'hFFB94ECA , 32'hFC9A52B4 , 32'hF8941230 , 32'h09FDC580 , 32'hFBB89A20 , 32'h020E3D70 , 32'hFFEC6409 , 32'hF92B6940 , 32'h052DE8E8 , 32'h058D1B58 , 32'hFA28C410 , 32'hFF95AB75 , 32'h00AF956D , 32'h02303210 , 32'hFC20E204 , 32'hFCCF7C78 , 32'hFDEE3794 , 32'hFEC9356C , 32'hF9238A10 , 32'h0251736C , 32'hFDA6A870 , 32'h01321300 , 32'hFB2BE4C0 , 32'hFE4AF2E8 , 32'hFEC2F6C8 , 32'h03EA5678 , 32'h062773A0 , 32'hFDA33C54 , 32'h01B1C304 , 32'hFF57FAF2 , 32'hFEC62090 , 32'h00C5BA69 , 32'hFCEC71EC , 32'hFF8396E4 , 32'hFDD19188 , 32'hFEE02944 , 32'h02500B84 , 32'hFF1EA09A , 32'h00621C6E , 32'h00CC4815 , 32'hFFE9CDF0 , 32'hFFFFCB88 , 32'hFFFFCE3F , 32'hFFFF53B8 , 32'h00042071 , 32'hFFFE2886 , 32'h0002697E , 32'hFFFFE774 , 32'hFFFF74E8 , 32'hFFFFA34A , 32'h0000AE65} , 
{32'hFFFBB7CA , 32'hFFFF6F9A , 32'hFFFF0872 , 32'hFFFF87FF , 32'hFFFFCBF0 , 32'h0003AAE5 , 32'h0000FF8F , 32'h0000178B , 32'h0000BB91 , 32'hFFFF1C93 , 32'hFFFD0E3D , 32'h00011442 , 32'hFFFCC302 , 32'hFFFE467E , 32'hFFFEAD29 , 32'hFFFD4E62 , 32'hFFFD45E9 , 32'hFFFF1141 , 32'h0000D59D , 32'h00035C33 , 32'hFFFC22EE , 32'hFFFF7A25 , 32'hFFFCB761 , 32'hFFFDCD6B , 32'h0003F88A , 32'hFFFD41AF , 32'h000183B0 , 32'hFFFD1E1F , 32'h00013DC4 , 32'hFFFF5ABF , 32'hFFFC3FBD , 32'hFFFDDE3E , 32'h00024EB9 , 32'hFFFEE83F , 32'hFFFDBBDC , 32'hFFFFE73D , 32'h0003F0B3 , 32'h0002AC5F , 32'h00021D8B , 32'hFFFEA733 , 32'h00007552 , 32'h00002A0D , 32'h0002577E , 32'h0001ADE2 , 32'h0002E7E2 , 32'h0000B16A , 32'h00012F9C , 32'hFFFF0D24 , 32'h0000E16C , 32'hFFFE8358 , 32'h0008EC41 , 32'h000284E0 , 32'hFFFE7986 , 32'h00002C0A , 32'hFFF9BBEC , 32'hFFFF7200 , 32'hFFFE26BF , 32'h0001842A , 32'h0000D59A , 32'hFFFEF190 , 32'hFFFCAA9A , 32'h00007781 , 32'hFFFD75F1 , 32'hFFFDFB13 , 32'hFFFE44FE , 32'h0001063C , 32'h0005DA04 , 32'h00015528 , 32'hFFFE070B , 32'hFFFBBEAC , 32'hFFFD2C0D , 32'hFFFB000B , 32'hFFFACA15 , 32'h00036B58 , 32'hFFFDDC4D , 32'h0000A9EE , 32'hFFFECBB7 , 32'hFFFFAED9 , 32'h0000C73C , 32'hFFFFBE6B , 32'h0002A8C7 , 32'h00016661 , 32'hFFFEF837 , 32'h0000E2B9 , 32'hFFFC8773 , 32'h00006CE0 , 32'h00024155 , 32'hFFFEFFBF , 32'hFFFD2659 , 32'h00001437 , 32'hFFFE79F4 , 32'h00013080 , 32'hFFFAC9BA , 32'h0002ACCA , 32'hFFFB0C89 , 32'h0000E379 , 32'h000059C5 , 32'h0001B6BE , 32'hFFFFB99F , 32'h000240F1} , 
{32'h3B2B6FC0 , 32'h1B1B9920 , 32'h4AF0D580 , 32'h0ED58830 , 32'hE2866BC0 , 32'h00E25FE7 , 32'hFD938AEC , 32'h212681C0 , 32'hFD82B730 , 32'hC1775000 , 32'h15A55840 , 32'hE3C44D80 , 32'hFD595670 , 32'h0CB58990 , 32'h04BB8B70 , 32'hFEA620C0 , 32'h125AE580 , 32'hEE98A580 , 32'hF01CB410 , 32'h0A443070 , 32'h167ED120 , 32'h12CC56A0 , 32'hF0936C50 , 32'h0A4EEEB0 , 32'hE8762520 , 32'hF2756660 , 32'h02582AB4 , 32'h0413E4D8 , 32'hEF236060 , 32'hF4A60BE0 , 32'h118A9160 , 32'hFD92F928 , 32'hFB914B00 , 32'h0858B930 , 32'h1488C660 , 32'h023B8448 , 32'h01D677D4 , 32'hEF0DCFC0 , 32'hF766EC10 , 32'h082B5EE0 , 32'h05E86890 , 32'hF668BB20 , 32'h06A2E3E8 , 32'hFE8DCB98 , 32'hFF3D7EBA , 32'h00BB420E , 32'h09C91940 , 32'h0CA020B0 , 32'hF9216CB8 , 32'hFCF3CDF8 , 32'hFBA46C68 , 32'hF5AE4990 , 32'h04E8DFA0 , 32'h026F52D0 , 32'hFC6161C4 , 32'h0072A540 , 32'h05CA8530 , 32'h0232C9BC , 32'h01AD13F8 , 32'hF85EB060 , 32'h06228E68 , 32'h02E6C870 , 32'hF8A0B6F0 , 32'h0688C140 , 32'h03540194 , 32'hFE6AD2D8 , 32'h035F9C94 , 32'h0114A340 , 32'hFACE3070 , 32'h0397D140 , 32'h004E7E01 , 32'hFDBEC6D8 , 32'hFEE366E4 , 32'hFADE15A8 , 32'hFBEDF180 , 32'h08C5D8C0 , 32'hFDAFEA48 , 32'hFCE9D554 , 32'h04D0FB98 , 32'h03B95750 , 32'h017DBABC , 32'h01612D54 , 32'h00EF37DA , 32'hFE29B56C , 32'hFFEBC8DF , 32'h00C7440D , 32'hFE5B2C20 , 32'hFC920CA0 , 32'h01972EB0 , 32'h00368DC8 , 32'h0000DEAD , 32'hFFFEA401 , 32'hFFFDF6F5 , 32'hFFFD7F05 , 32'hFFFEF745 , 32'h00003E3A , 32'h000013A1 , 32'h00020657 , 32'hFFFFFB5B , 32'hFFFF99DA} , 
{32'h120DCBA0 , 32'h0014C44A , 32'hF8B33560 , 32'hEE77C140 , 32'h09D49400 , 32'hF5AC2D90 , 32'h04513BB8 , 32'hFDB8DA88 , 32'h09F74870 , 32'h04F3D1A8 , 32'h124160A0 , 32'h09F16E10 , 32'h013D0AA8 , 32'hF05F7AD0 , 32'hFD4849B0 , 32'h0DB49D80 , 32'h01338DFC , 32'hFE039D6C , 32'h01D73748 , 32'hFDB85A18 , 32'hF9DFFAC0 , 32'hFC36B984 , 32'h072B83A8 , 32'h05771960 , 32'hFF9B0FA3 , 32'h0CEDEB00 , 32'h04C114D0 , 32'hFBA5A698 , 32'hFF6D2407 , 32'h0B63EB90 , 32'hFD66B960 , 32'hFA1368D0 , 32'h09AEB7D0 , 32'hFBA295C0 , 32'h03FB4020 , 32'h018DEBE0 , 32'h010D7860 , 32'hFD97A938 , 32'hFFE217A6 , 32'h02287A78 , 32'hFF18B253 , 32'h029439B8 , 32'hFD496320 , 32'h04051620 , 32'hFE66C61C , 32'h086B8160 , 32'h0144978C , 32'hF7DBD2C0 , 32'hFA34B680 , 32'h098E43B0 , 32'hFDD98F84 , 32'hFAAA0288 , 32'h09E34640 , 32'hF6DFF910 , 32'hFF90DFB3 , 32'hF7025B30 , 32'hFB9FAF70 , 32'hFE9E6F0C , 32'h03D9E5F0 , 32'hFF57FFC2 , 32'h023A1680 , 32'h0263BB50 , 32'hFDD6176C , 32'h02575C98 , 32'h02262EC4 , 32'h02564DD4 , 32'h03F96864 , 32'h007CE645 , 32'hFFCA5DFD , 32'h02AE2570 , 32'hFFBBD839 , 32'h00EE3F7B , 32'h008AAFFA , 32'hFFEEE611 , 32'hFF5E555E , 32'h00CCF1A5 , 32'hFC745508 , 32'h011C9144 , 32'h01864E88 , 32'h04728E50 , 32'h018F9EA4 , 32'h04ADFF38 , 32'h02FCA0A4 , 32'h01676FDC , 32'h014E0048 , 32'h0062B2BA , 32'hFD8C44E4 , 32'hFF51B184 , 32'hFDF51DC8 , 32'hFF762BDD , 32'hFFFB13FF , 32'h0003BC3E , 32'hFFFD9A4A , 32'h000286FA , 32'hFFFFE648 , 32'hFFFD0E6E , 32'h00056ADE , 32'hFFFDF948 , 32'h00028009 , 32'h000047FE} , 
{32'h1F47ABE0 , 32'h06CA8808 , 32'h1ED68D60 , 32'h0CDB7160 , 32'h26005F40 , 32'hFE844B10 , 32'h16A5EE00 , 32'hF6BC5050 , 32'h06EDE7E8 , 32'h031B9100 , 32'hF17EF520 , 32'h02BCC9D8 , 32'hFB5BF2B8 , 32'hF3DEE700 , 32'h039EBA84 , 32'hF9A6B538 , 32'h1D20C7E0 , 32'hED92C020 , 32'h032610E4 , 32'h070AD788 , 32'hDF40E200 , 32'hFF567460 , 32'hF04E4E00 , 32'h017C6BF8 , 32'hF22F6330 , 32'hFA2DCAF0 , 32'hECBCBA40 , 32'hED7D9820 , 32'hF3A40F70 , 32'hFC99EACC , 32'h1878FBA0 , 32'h0AB1D500 , 32'hFA762AC0 , 32'h054F96A0 , 32'hFCF171D8 , 32'h0C5C8C30 , 32'h06A010E8 , 32'h04EF04B8 , 32'hE4EDE220 , 32'hF8261E58 , 32'hFE1721FC , 32'h0A573420 , 32'hFAAD8B70 , 32'hFAE59F30 , 32'h177C80A0 , 32'h09A8F9C0 , 32'hFF0017D3 , 32'h09AE2E00 , 32'h098C6300 , 32'h05F937A8 , 32'hFFC0FB9C , 32'hFF360F0F , 32'hFBBCA2F8 , 32'hFE397B00 , 32'hF5AF12B0 , 32'hF9F4DDB0 , 32'hFF6604FC , 32'h08F3CA80 , 32'h074D8560 , 32'h11E54220 , 32'h018DB354 , 32'h07CC6640 , 32'h0013FE40 , 32'h046319D0 , 32'h02ADE974 , 32'hFF1D1819 , 32'hFFC2C24D , 32'hFE392DB0 , 32'h02394A78 , 32'h01A7F19C , 32'h02387920 , 32'hFEBAA374 , 32'h005E037E , 32'h01B58DFC , 32'hFAC6C2F0 , 32'hFC6773A0 , 32'h0367F790 , 32'h03E88FC4 , 32'h02E80B9C , 32'hFECC9CEC , 32'hFB9DCF60 , 32'h020C377C , 32'hFAEA83D0 , 32'hFF39F5E6 , 32'h00B9F68F , 32'hFA90DD40 , 32'h0081DCD0 , 32'h03865284 , 32'h00BC3FAF , 32'h00673544 , 32'h0000C3D5 , 32'h000127F0 , 32'hFFFD506D , 32'h0000CE92 , 32'hFFFF46D4 , 32'hFFFD3358 , 32'h000092BD , 32'hFFFE3BF2 , 32'hFFFE6228 , 32'h000020CF} , 
{32'hFAAF4BD0 , 32'h1E2F1A80 , 32'h456AE480 , 32'hD55B0F00 , 32'h09D02CD0 , 32'hE4C374E0 , 32'hF89B0CD8 , 32'h067C0088 , 32'hF0A495F0 , 32'hE93CD580 , 32'h05D71B78 , 32'h14C6DD40 , 32'h028BFD0C , 32'hFD288494 , 32'hEE804320 , 32'h03C92CCC , 32'hE5801CC0 , 32'h28380E00 , 32'hF9424EB0 , 32'h0EDC8100 , 32'hEA2AA4A0 , 32'h03499714 , 32'hFC6A9C38 , 32'h16C87800 , 32'h028D09A4 , 32'hF7EDB450 , 32'hEFFDE960 , 32'h06B659D8 , 32'h012E0FE4 , 32'h08E068D0 , 32'hF5185180 , 32'hFE9F18FC , 32'h0B27A810 , 32'hFA9C39F8 , 32'hF295D6D0 , 32'hED394B80 , 32'hF252E6C0 , 32'hF71F2D50 , 32'hF2287FA0 , 32'h04B86A80 , 32'hF56D2860 , 32'hEDFAEA60 , 32'h10BF6FA0 , 32'h041BBE98 , 32'h0E47C3D0 , 32'hFCCC6A80 , 32'hFFE4A121 , 32'h090B7B00 , 32'hFAEBCAA8 , 32'hF67FB1C0 , 32'h06BC4BC0 , 32'hFB636C20 , 32'h00D3124B , 32'h003D33FB , 32'hFC868F10 , 32'h0A3C1090 , 32'h07957450 , 32'h01E806AC , 32'hF7E7EA60 , 32'h0290B068 , 32'hF58A6930 , 32'h01AC1328 , 32'h03927BE4 , 32'hF9CB6BF0 , 32'hF5268280 , 32'h009247FA , 32'h04303268 , 32'hFD90B06C , 32'hFDBC42DC , 32'hFFE3492E , 32'h065C26D8 , 32'hFBE30840 , 32'hFE247CC8 , 32'hFD5DE6C0 , 32'h03EE2088 , 32'hFF42F29D , 32'h040A65E8 , 32'hFF0166FA , 32'hFFDB6C7A , 32'hFFC5F4BF , 32'h00C49E6A , 32'h00A4473C , 32'h03F88064 , 32'hFE3F193C , 32'h03569A24 , 32'hFE9B8CE0 , 32'hFC08AD9C , 32'h0118A3C4 , 32'hFE843B9C , 32'h009A510A , 32'hFFFFA080 , 32'hFFFF69C9 , 32'hFFFF46B8 , 32'h0000C122 , 32'hFFFFA916 , 32'hFFFE0796 , 32'h00032F05 , 32'hFFFEACDA , 32'hFFFF9D6E , 32'h0000C780} , 
{32'hFB27EC00 , 32'hD863F740 , 32'hF473A510 , 32'h0D4BA290 , 32'h11CF0180 , 32'h102B2600 , 32'hDD220440 , 32'h3049C4C0 , 32'h0CF2F4E0 , 32'h11BA6F80 , 32'h0E0B6FC0 , 32'hF937E690 , 32'h09337BC0 , 32'h04C1DCE0 , 32'hFA747690 , 32'hF427C7B0 , 32'h0BB69240 , 32'h05FBEBF0 , 32'hEAD73360 , 32'hEC598BE0 , 32'hDA2FE980 , 32'hF691E2B0 , 32'hF6C6FF20 , 32'hDF86E680 , 32'h141F9780 , 32'h08314F70 , 32'h09EC7250 , 32'hE9D244C0 , 32'h04B750C8 , 32'h0889C490 , 32'hFE08D4C8 , 32'hF3C3D8D0 , 32'h0EC6FA00 , 32'hF6633750 , 32'h0D62A3D0 , 32'hFEBCE398 , 32'h003C8146 , 32'hEBEB9A40 , 32'h0B288320 , 32'h0C68C0D0 , 32'h0DC04350 , 32'h0A0D3490 , 32'h05A53CE8 , 32'hF5CC0800 , 32'hFD84CD1C , 32'hF5CFCC90 , 32'hF22E11E0 , 32'h034F2BF8 , 32'h01F2F134 , 32'h04688F80 , 32'h0EE2F6C0 , 32'h02F08C48 , 32'hF72A9A50 , 32'h030543FC , 32'hFE1EBD08 , 32'h031152B8 , 32'h033B87C4 , 32'hFAA1E678 , 32'hFB64FB90 , 32'hF8143288 , 32'h0F4E4670 , 32'h03334284 , 32'hFA8B45C8 , 32'h08AD3470 , 32'hFA9D7BF0 , 32'h041E9748 , 32'h0706FC80 , 32'hFA8351E8 , 32'hFBAE9160 , 32'h056E0708 , 32'h02E21ADC , 32'h00DEF5D6 , 32'h0042AAA6 , 32'h01961B08 , 32'hFF33A33B , 32'h0423E618 , 32'h026A19C8 , 32'h011CE100 , 32'hFFA967D4 , 32'h00C7B564 , 32'h01F1C6FC , 32'h02EA5A70 , 32'hFE0BDBA0 , 32'h02A6E678 , 32'hFD5C5884 , 32'hFAFCB088 , 32'hFD845394 , 32'h000D354C , 32'h022D3D48 , 32'h00A5C9EE , 32'hFFFF6DFD , 32'h000200A4 , 32'hFFFFCDDC , 32'h0001095F , 32'hFFFF4D10 , 32'h00000290 , 32'hFFFE6EC9 , 32'hFFFFB5D6 , 32'h00001196 , 32'hFFFF0034} , 
{32'h93F75900 , 32'hF99DEE28 , 32'h35B30140 , 32'hC5D5A980 , 32'hD357A680 , 32'h0E29A4B0 , 32'hE9446440 , 32'h0FD23290 , 32'h1E8E4EC0 , 32'h12C795E0 , 32'hFDBB2FEC , 32'hF35B73A0 , 32'h1BD7C180 , 32'h0E94C270 , 32'hF2DE7000 , 32'h127CEB40 , 32'hFCAD0DDC , 32'h1394DA40 , 32'h1BBA4400 , 32'h01F77AC4 , 32'h0BD680B0 , 32'h2B7EF580 , 32'h01BA74F8 , 32'hE89F9020 , 32'h01AACCBC , 32'h01C13A58 , 32'hF5047600 , 32'hFA507E20 , 32'hF4B6E360 , 32'h0BCBF020 , 32'hFB3B5448 , 32'hEF29A160 , 32'hE74D6520 , 32'h0777FCD0 , 32'hF14ABAD0 , 32'hFA84FBB0 , 32'hF7161AC0 , 32'h080D2020 , 32'hF62A10B0 , 32'hF8EC1A60 , 32'h02F34280 , 32'hFB25D7B0 , 32'hF9D5EE48 , 32'hFAEAF700 , 32'hF0E0E670 , 32'h0FF92EC0 , 32'h06D80320 , 32'h06816100 , 32'h084B40C0 , 32'h071CC688 , 32'hF8D00BE0 , 32'hFF3A7BCE , 32'h06559720 , 32'h013C1944 , 32'hF8740F78 , 32'h0280D430 , 32'h0652F9B8 , 32'hF8AC5328 , 32'hFFB3D553 , 32'h04FDF288 , 32'h06889C90 , 32'h040CAFF0 , 32'h02C11D8C , 32'hFF4CD15C , 32'h014F63A0 , 32'h06FFE688 , 32'hFD61FB38 , 32'hFF5BAF29 , 32'hFDAA0730 , 32'hFC598EA4 , 32'h05B74F00 , 32'h00CDA52E , 32'h02B68F20 , 32'h01BC8F4C , 32'hFE66A4CC , 32'h029C6B08 , 32'h008CE5CB , 32'hFAE22F48 , 32'h040454D0 , 32'h02E177D4 , 32'hFEC560DC , 32'hFEE54470 , 32'hFEBC6F00 , 32'hFF4C2627 , 32'h006C5ABA , 32'h021F58A4 , 32'h015572B8 , 32'hFEEC4884 , 32'h00D07400 , 32'hFFE1F19F , 32'hFFFFF70D , 32'h0001B917 , 32'hFFFE3BAC , 32'h00035E6C , 32'h00001477 , 32'h0001EF93 , 32'h0000A711 , 32'hFFFD9A42 , 32'hFFFFB781 , 32'hFFFF631B} , 
{32'h00F31C9B , 32'h08476630 , 32'hFD18C06C , 32'h03A1D23C , 32'hFD18FF0C , 32'h01C0FB18 , 32'hFCB90D30 , 32'h04B19A58 , 32'h02E6F3C8 , 32'h0424F220 , 32'h02AC18A4 , 32'hFD138A80 , 32'hFD851608 , 32'hFD0F40B8 , 32'hFBEE59B0 , 32'h05A14D80 , 32'hFCAF0C6C , 32'h01350C18 , 32'h035C0270 , 32'h06CD9AB8 , 32'h08F2EFA0 , 32'hFE88A824 , 32'hF93C76E8 , 32'h012B9858 , 32'h0382A80C , 32'h011B9E28 , 32'h039758F0 , 32'hFD237BA8 , 32'h0206BAB8 , 32'h02102B4C , 32'h01619818 , 32'hFF176975 , 32'h01CB51D4 , 32'hFA990D58 , 32'h0601AA60 , 32'hFE1CFEB8 , 32'h0573F5F0 , 32'h0020211F , 32'hFB866A20 , 32'hFD280348 , 32'h04441F90 , 32'hFF00CA12 , 32'hFDE03D84 , 32'h008A2E60 , 32'hFF98F472 , 32'hFD55CAA0 , 32'h00525B36 , 32'hFBE8A280 , 32'h04721518 , 32'hFE464DA0 , 32'h08F42B70 , 32'h05BAC9F8 , 32'hFE8338B4 , 32'hFF3A6562 , 32'hFECE85FC , 32'h0043F7E3 , 32'h059B2D18 , 32'hFE7AA768 , 32'hFE0AD7F4 , 32'hFE588964 , 32'hFEB664B4 , 32'hFC012ED8 , 32'h01CF3E24 , 32'hFD3D06D8 , 32'h034CA014 , 32'h03771284 , 32'hFEEA30E0 , 32'h04152318 , 32'hFE28E99C , 32'h01B256FC , 32'h04897300 , 32'hFE9B8F78 , 32'hFE7C13AC , 32'h004D0D85 , 32'hFF7C80CA , 32'hFEB1640C , 32'h008DC28E , 32'h00057CE5 , 32'h0046CAEF , 32'h01C4D87C , 32'h01557D68 , 32'hFF65409F , 32'h006DFF93 , 32'h010FBF70 , 32'h014C2570 , 32'h01A6B764 , 32'h02CAD094 , 32'h00066E2D , 32'hFF7DC233 , 32'hFFEEDAFE , 32'h00048793 , 32'hFFFFCFBA , 32'h000787D5 , 32'hFFFF6377 , 32'h00010990 , 32'hFFFFD0C2 , 32'h00021E83 , 32'hFFFF1C96 , 32'h0002C4E7 , 32'hFFFEE35A} , 
{32'hD6504540 , 32'h1BC544E0 , 32'hF66DEF80 , 32'h0EB35700 , 32'h0666AC20 , 32'hEE7061E0 , 32'hF5DD5680 , 32'hF4E8D030 , 32'hFEA489B4 , 32'hFDCD7250 , 32'hF0CD67F0 , 32'hFDE7153C , 32'hEA0BAE40 , 32'hF9215DC0 , 32'hFD2F5410 , 32'hFE4E5C04 , 32'h07F141B8 , 32'h08047470 , 32'hF20907D0 , 32'h14E6ED20 , 32'h0653F928 , 32'hF74A6880 , 32'hF2BB40F0 , 32'h08A91740 , 32'h005351E3 , 32'h08628580 , 32'hFDCBB154 , 32'hF7D27430 , 32'hF24937C0 , 32'h08B3CF10 , 32'hF89623B8 , 32'h06BFB298 , 32'hF21A3310 , 32'hF0224EF0 , 32'hFB1876C0 , 32'hFD497A10 , 32'h0449B118 , 32'h0BB00F00 , 32'h07362A78 , 32'h0A82BF00 , 32'hF37B2070 , 32'h0E9E8360 , 32'h07653618 , 32'h07320C50 , 32'hFB3EB088 , 32'h03799AFC , 32'hFBFE7430 , 32'h0C94D6A0 , 32'h00743DEE , 32'h0786D678 , 32'h018C8460 , 32'hF71E8760 , 32'h0675EF80 , 32'h06340630 , 32'h03B5E160 , 32'hFD960C04 , 32'h094A5990 , 32'h0636B438 , 32'h0C6F9C30 , 32'hF8CE4C28 , 32'h00C2E1CE , 32'h0148D9A4 , 32'h015ACCB4 , 32'h037B2768 , 32'hFDF96D04 , 32'hFC731C94 , 32'h02082100 , 32'hF96A5298 , 32'hFE567810 , 32'h025E4E08 , 32'hFB0C5268 , 32'h01F439D4 , 32'h04654C70 , 32'h026F0EC0 , 32'h045AC0C0 , 32'hFB406778 , 32'h02E1BCE8 , 32'hFEE83434 , 32'h04E58948 , 32'h0036B827 , 32'h02D12F8C , 32'h041A7FF8 , 32'hFFCF69F6 , 32'h04171EF0 , 32'h019C7E98 , 32'hFAC13B20 , 32'h01BC97B0 , 32'hFF40A28D , 32'h021871BC , 32'hFFCBB475 , 32'h0003A18B , 32'h00019A6B , 32'hFFFCCD03 , 32'hFFFFC5C7 , 32'h000103B2 , 32'hFFFD2366 , 32'h00005B3B , 32'hFFFFEF48 , 32'hFFFFE6F9 , 32'hFFFF6ACD} , 
{32'h00019068 , 32'h0002D5AD , 32'h0000A139 , 32'h0001EE9C , 32'hFFFF3E49 , 32'hFFFCF2B7 , 32'h00002EE2 , 32'h00035E9A , 32'h00035726 , 32'h00001142 , 32'hFFFFB827 , 32'h0000B56D , 32'h00008D0F , 32'h00023690 , 32'h000136DD , 32'hFFFBB5D0 , 32'h00013DE1 , 32'hFFFD53A4 , 32'hFFFD76E8 , 32'h0001F671 , 32'hFFFF141B , 32'h000009B2 , 32'hFFF9EAB0 , 32'h0003C1C2 , 32'hFFFE91DC , 32'hFFFFC8E2 , 32'h0001D8D4 , 32'hFFFC877D , 32'hFFFAE9FE , 32'hFFFEB28B , 32'hFFFCEC2C , 32'hFFFEF226 , 32'hFFFD7083 , 32'h0001F43C , 32'hFFFFCD90 , 32'h00032A9E , 32'hFFFFC387 , 32'hFFFC5AE1 , 32'hFFFAF668 , 32'hFFFFB911 , 32'h000567BD , 32'h00007CF4 , 32'h0001A2CA , 32'h0002AAF0 , 32'h000176B8 , 32'h000262DC , 32'hFFFFC7DA , 32'hFFFFD727 , 32'h0003CD73 , 32'h0003B926 , 32'hFFFCBD38 , 32'hFFFECCDA , 32'h000045DE , 32'hFFFFEB71 , 32'hFFFC8F33 , 32'h00012D81 , 32'h000028F1 , 32'hFFFC2040 , 32'hFFFCA2C3 , 32'h00039ADF , 32'h000177D2 , 32'hFFFF54D7 , 32'hFFFB4CBF , 32'h00016F55 , 32'h00034295 , 32'hFFFF3699 , 32'h0004A330 , 32'h0002D7E0 , 32'hFFFC5D46 , 32'hFFFD2318 , 32'hFFFCD1BE , 32'h0000C1AB , 32'hFFFE9F70 , 32'h0001B47D , 32'h0003B440 , 32'hFFFCBD7F , 32'hFFFDC01B , 32'h000360F5 , 32'hFFFFAF44 , 32'hFFFE4420 , 32'hFFFE445B , 32'h0001DA02 , 32'h0000861C , 32'hFFFFCB2F , 32'hFFFFE52A , 32'hFFFC46DF , 32'h00002EFB , 32'hFFFEB6E0 , 32'hFFFFD23A , 32'hFFFE3D9F , 32'h00005E72 , 32'hFFFF9B4E , 32'h00023C63 , 32'h000165A1 , 32'h000157EA , 32'hFFFF6739 , 32'hFFFC3C8C , 32'h00009142 , 32'hFFFF90F7 , 32'h000052DD} , 
{32'h0000D3F8 , 32'hFFFE5DB4 , 32'hFFFFC1F6 , 32'h0000D999 , 32'hFFFF1414 , 32'h00014E14 , 32'h000269C6 , 32'hFFFEAF8C , 32'hFFFEBE11 , 32'h0001B42C , 32'h00015D8E , 32'hFFFDB7E2 , 32'hFFFBF654 , 32'h00010C18 , 32'h000389B2 , 32'hFFFE759E , 32'hFFFDEBF6 , 32'hFFFEE14F , 32'h0001A8A4 , 32'hFFFE6A35 , 32'hFFFE5AF2 , 32'h0005F36A , 32'h000026BA , 32'hFFFD609B , 32'h00052019 , 32'hFFFBC124 , 32'hFFFCCA6A , 32'h00049621 , 32'hFFFD0955 , 32'h0000567C , 32'hFFFF5AF7 , 32'hFFFF0E3F , 32'h00013F8D , 32'h00021A95 , 32'hFFFF9DC6 , 32'h00009430 , 32'hFFFEEAB4 , 32'h0000B0BD , 32'h0005DEF2 , 32'hFFFB5AAF , 32'h000330C0 , 32'h0000A81A , 32'hFFFD8036 , 32'hFFFF59A1 , 32'hFFFDB241 , 32'h00003C29 , 32'hFFFB9177 , 32'h000568E6 , 32'hFFFCEAF4 , 32'hFFFE7C31 , 32'h000134CD , 32'hFFFDA3F9 , 32'hFFFD2CA5 , 32'h00016035 , 32'hFFFB7188 , 32'hFFFB25DB , 32'h00014DC8 , 32'h0000C8C9 , 32'h000106A3 , 32'hFFFBD9D0 , 32'h0003FFBB , 32'hFFFFD141 , 32'hFFFF9E74 , 32'h000054E6 , 32'hFFFD7288 , 32'h00019FF3 , 32'h0004DFDD , 32'h00016A5E , 32'h00044CDD , 32'h00045FC0 , 32'h00023403 , 32'h0002E050 , 32'hFFFF10C6 , 32'hFFFCFB40 , 32'h000290A9 , 32'h00034035 , 32'hFFFE8A65 , 32'hFFFDD1E7 , 32'hFFFF2FDD , 32'h000229A4 , 32'h0000BB18 , 32'hFFFFBD3B , 32'h0003C090 , 32'hFFFFDF4F , 32'h00000E69 , 32'h000406A1 , 32'h0003308F , 32'hFFFE1467 , 32'hFFFCAB42 , 32'hFFFEA165 , 32'hFFFF8190 , 32'hFFFEFC8D , 32'hFFFF8103 , 32'h0000470D , 32'h00028473 , 32'h0002DC9D , 32'h00015288 , 32'h0000D617 , 32'hFFFFE0C0 , 32'hFFFDF6CD} , 
{32'hFFFFD94C , 32'hFFFB1A4C , 32'hFFFFA5A6 , 32'h00023E33 , 32'h000172B5 , 32'h0000B32D , 32'h00003676 , 32'hFFFC1647 , 32'hFFFBCE0C , 32'h00061DB0 , 32'h0006AB38 , 32'h0000EA7B , 32'h00002ED9 , 32'h000280A3 , 32'h0001203F , 32'hFFFFB110 , 32'h0000DA18 , 32'h0002BED8 , 32'h0000D2F9 , 32'h000473D0 , 32'hFFFDB9B2 , 32'hFFFE09B3 , 32'hFFFE77B0 , 32'h0000471F , 32'hFFFF70E1 , 32'hFFFCBF9B , 32'h000013E1 , 32'h00023A31 , 32'hFFFD0078 , 32'hFFFE9D83 , 32'hFFFECE3F , 32'h0004934F , 32'hFFFC4F89 , 32'hFFFE5E47 , 32'hFFFFE644 , 32'hFFFFC372 , 32'h00010BE2 , 32'hFFFDB73C , 32'hFFFD0EAB , 32'h00010286 , 32'h0001605C , 32'hFFFF0196 , 32'hFFFFBA65 , 32'hFFFCD2E4 , 32'h00066540 , 32'h00000C30 , 32'hFFFE94FF , 32'h000095EF , 32'h00000C40 , 32'hFFFEA049 , 32'hFFFE4E68 , 32'hFFFE4EB9 , 32'h00020B57 , 32'h00017452 , 32'hFFFC5E04 , 32'h00010146 , 32'hFFFFA3BA , 32'h00024329 , 32'hFFFC230E , 32'h0000C1E6 , 32'hFFFF1F0B , 32'h000261F6 , 32'h00005E54 , 32'hFFFDCEEE , 32'hFFFB4E75 , 32'h0002A03C , 32'hFFFB6BCF , 32'hFFFCFE3D , 32'h00033540 , 32'h0002ACDD , 32'h0004627A , 32'h000036FB , 32'h0002658D , 32'hFFFCEB5F , 32'hFFFA2360 , 32'hFFFBC7D3 , 32'hFFFB38CF , 32'h0000B281 , 32'h0001E9A2 , 32'hFFFA9A6E , 32'hFFFDD4B7 , 32'h0002935F , 32'h00005FBD , 32'h00048911 , 32'hFFFEDADE , 32'hFFFCD0BE , 32'h0004348B , 32'h00041914 , 32'hFFFF2F01 , 32'h00006120 , 32'h000393A8 , 32'h00012FCB , 32'h00066C53 , 32'h00014804 , 32'h0000D38E , 32'h0002140C , 32'h0002A93C , 32'hFFFEF88D , 32'hFFFD5273 , 32'h00039003} , 
{32'hEEF984A0 , 32'h01AC5E28 , 32'hE93BC5C0 , 32'hFBA227F8 , 32'h0D6DD570 , 32'h018CE630 , 32'hF671EF30 , 32'hFE115AC8 , 32'hF3851FD0 , 32'h10235240 , 32'hF94983D8 , 32'h00E40A02 , 32'hF814E8E8 , 32'hFB46B290 , 32'hF661E2E0 , 32'h07E3A980 , 32'hF20B6610 , 32'hFA4CA9A0 , 32'hFBB0B718 , 32'h12B75480 , 32'h022F94EC , 32'hF39A3080 , 32'hFFB24234 , 32'h09DB9C90 , 32'h0D183210 , 32'h00CE33D0 , 32'hF3DE0EC0 , 32'hF6FE4690 , 32'hF3A8C7B0 , 32'hF49062B0 , 32'h049F4348 , 32'h00127164 , 32'hFE672820 , 32'hFEC5120C , 32'h01F4F40C , 32'hF8CC1BE8 , 32'h05CBDBD0 , 32'hFB3635F0 , 32'h049FBDB8 , 32'h06164F60 , 32'h06B64C88 , 32'hF5CD4FF0 , 32'h0283EEEC , 32'hFD314000 , 32'h038BB334 , 32'hF6B2DB90 , 32'h0DD16F80 , 32'hF89DF2B0 , 32'hFB205A70 , 32'h098C8AA0 , 32'h01470F14 , 32'hED52C040 , 32'hFF52645E , 32'hFD45EBA0 , 32'hFB894E20 , 32'hFC347368 , 32'hFB6E7020 , 32'hF9DAAEE0 , 32'hFD54BE38 , 32'hFB681AB8 , 32'hFB1D7A68 , 32'h04A3E308 , 32'hFC05E234 , 32'h03179694 , 32'hF891D408 , 32'h02EBF994 , 32'hFE6B411C , 32'hFD37A9FC , 32'hFA36EC28 , 32'hFB4B27E8 , 32'hF97E5518 , 32'hFFF965D9 , 32'hFEA2D9C8 , 32'hFEF59314 , 32'h010A60D4 , 32'hFAA3F3A0 , 32'hFF127B3B , 32'h0A274070 , 32'hFDA63924 , 32'h038B42DC , 32'h0225D798 , 32'hFB6CD748 , 32'hF8707928 , 32'hFC4239B0 , 32'hFCEBB668 , 32'hFFE6A8BE , 32'h022C4110 , 32'hFE237160 , 32'hFF2F8BE5 , 32'hFFFC77AB , 32'hFFFDF7D2 , 32'hFFFF43CF , 32'hFFFFC423 , 32'h0000DA20 , 32'h00025544 , 32'hFFFF869E , 32'h0002E828 , 32'h00007A60 , 32'h00052912 , 32'h0000C55B} , 
{32'hDB105E00 , 32'h2DA7D4C0 , 32'hF747EEB0 , 32'hEF71C360 , 32'h13286620 , 32'hDB0ABCC0 , 32'h2CFC2640 , 32'h2ABD1880 , 32'hE3A6FA80 , 32'hFCCDBC5C , 32'hEA410E00 , 32'h18DCD1E0 , 32'h16BA2C80 , 32'hF194E7D0 , 32'h04154970 , 32'h174F4D60 , 32'h12DF5C80 , 32'h11450580 , 32'h08B785A0 , 32'hE9462720 , 32'h0D95D590 , 32'h0A786610 , 32'h03DF3FF8 , 32'h1C1848A0 , 32'h08843CA0 , 32'hF6D33620 , 32'h08A030C0 , 32'hEA5885E0 , 32'h0082FBEA , 32'hF52B1740 , 32'hEC9241A0 , 32'hFF30CEB8 , 32'h0158BE48 , 32'hFC86D21C , 32'h025EECE4 , 32'h0506A450 , 32'hFBB972A0 , 32'h0131C8FC , 32'h03DA17BC , 32'h0BD14200 , 32'h0D554470 , 32'h007A9E10 , 32'h0014DEC0 , 32'hF71A3B00 , 32'hF5E56490 , 32'hFFF52C4F , 32'h0C72EB20 , 32'h0941FD30 , 32'hF7B677A0 , 32'h086F4EC0 , 32'hFCE7C32C , 32'h0752A650 , 32'hFA64E1E0 , 32'hFF9A5F36 , 32'hFBEBE390 , 32'hFE618174 , 32'hF76CFE30 , 32'h0224B674 , 32'hFF5D6931 , 32'hFF7F55F2 , 32'h08A39550 , 32'hF2E8DB90 , 32'hFA1058F0 , 32'h0D494720 , 32'hFD913644 , 32'h0059F548 , 32'h0263B5A4 , 32'hFD49D2D4 , 32'hFFE17499 , 32'hFA134650 , 32'h00AF2A7C , 32'hFEC48754 , 32'hF61A8EB0 , 32'hFCCC9F14 , 32'h012BBD58 , 32'hFC6CFDC0 , 32'h028A765C , 32'h00C097B3 , 32'h00571CA5 , 32'hFE5F8760 , 32'hFC44DB48 , 32'hFFBEB70A , 32'hFBC6D518 , 32'hFF115A39 , 32'h00ABC74E , 32'hFC602C2C , 32'hFEE516C0 , 32'h024100F4 , 32'hFFF51ED8 , 32'h007F95CC , 32'h0000B6E1 , 32'hFFFFCBC7 , 32'h0001937E , 32'hFFFF82B2 , 32'hFFFFCB08 , 32'hFFFE86FB , 32'hFFFFBFC5 , 32'hFFFE90F3 , 32'h00002932 , 32'h0000E269} , 
{32'hF3373250 , 32'h0050EA33 , 32'hF3BA69B0 , 32'h114EFDE0 , 32'h05D2EFB0 , 32'h115FC640 , 32'hFCC65BB0 , 32'hFD779624 , 32'hF549BD00 , 32'h06EBC498 , 32'h01157B30 , 32'h072DFEC0 , 32'hFAC45300 , 32'hF8054488 , 32'hEEC010C0 , 32'h03C15384 , 32'hF33852A0 , 32'hFB908680 , 32'h015E8A80 , 32'h025C1C38 , 32'hFA9791F8 , 32'h0629FE38 , 32'hFE24AE98 , 32'hFD38EC8C , 32'h08546840 , 32'h01ACF52C , 32'hF687CD50 , 32'hFFC052BB , 32'hF80AC070 , 32'hEE225EA0 , 32'h0B72BD80 , 32'h0C5B4B70 , 32'hFF9C50E2 , 32'hFE78007C , 32'hFB59B3F0 , 32'hFF8A76D5 , 32'h06EF9E08 , 32'h030DA30C , 32'hFF4B790A , 32'h060FAC28 , 32'h00187CDC , 32'h0427CE68 , 32'h071278A8 , 32'hFE0DF924 , 32'hFE886F4C , 32'hFA46DA78 , 32'hFD546F0C , 32'h02BE30B8 , 32'h018F2040 , 32'hFDB5602C , 32'hF817C850 , 32'hF3D77FB0 , 32'hF925D0E0 , 32'hF7B81930 , 32'hFC5D246C , 32'hF7BB91C0 , 32'hFD9D9BEC , 32'h085B7840 , 32'h0211E470 , 32'hFDD01C4C , 32'h02D13FD4 , 32'hFDE5CAA0 , 32'hFD317C94 , 32'hFE60350C , 32'hFF87D1B1 , 32'hFF844DB4 , 32'h033081F0 , 32'h06F8FF18 , 32'h0372E1C0 , 32'hF9DB8F80 , 32'hFC202680 , 32'h02478780 , 32'hF998B8F8 , 32'h00162039 , 32'h008A0723 , 32'h02EE0664 , 32'h002A7263 , 32'h0018ADCD , 32'hFBDB4538 , 32'hFDA027CC , 32'h069FDA68 , 32'hFE2B0E08 , 32'hFF35B642 , 32'hFE1DA174 , 32'h00FFF6E7 , 32'h0197B090 , 32'h033138A4 , 32'hFE0E8114 , 32'h00E6501B , 32'hFFD7DD5A , 32'hFFFDAC47 , 32'h00042EA4 , 32'h000227B6 , 32'h00017DE4 , 32'h0000703E , 32'h0000D763 , 32'hFFFDD505 , 32'h00001BE9 , 32'hFFFD7794 , 32'h000029A8} , 
{32'hF9F35AF8 , 32'h0537D568 , 32'h01838574 , 32'h0843F780 , 32'h01BEBC78 , 32'hFF433FDF , 32'hFAFC10B8 , 32'h040914F0 , 32'hFDA083D4 , 32'hFB4726E0 , 32'hF89084C8 , 32'hFEE21FBC , 32'h0504BD10 , 32'hF9F34F10 , 32'h01405594 , 32'hFFE02810 , 32'hF6FE0180 , 32'h05C75488 , 32'hFF2B29C8 , 32'h012E8318 , 32'hFA74F198 , 32'hF922EA70 , 32'hFFEC9BA9 , 32'h0703F2D8 , 32'h01D57E70 , 32'hFDD28FA4 , 32'h05A996B8 , 32'hFCD7D17C , 32'hF8D61458 , 32'h05984680 , 32'hF76D4FC0 , 32'hF6FDD200 , 32'hFCB5B210 , 32'h002D7464 , 32'hF8C9D638 , 32'h02D0F2C0 , 32'h051C34E0 , 32'h0946B820 , 32'h054A7AF8 , 32'h001A8853 , 32'h0402E7B0 , 32'h03A58B00 , 32'hFE99F4D8 , 32'h03272300 , 32'hF8DC65F0 , 32'h032BA584 , 32'hFBDE9298 , 32'h02F7A964 , 32'hFDA90CFC , 32'hFF585435 , 32'hFF364247 , 32'h0289F728 , 32'hFA9F1EF0 , 32'h02D58BBC , 32'h03EC5D9C , 32'h0466FAD0 , 32'hFFAB273C , 32'hFD218298 , 32'h02FCC8F4 , 32'h063D1EA0 , 32'h053E00B8 , 32'hFB4F0AC8 , 32'h03735040 , 32'hFF65033F , 32'hFDEFA25C , 32'hFD240968 , 32'h01D030E8 , 32'h004B811D , 32'hFE10B040 , 32'h007A2F6C , 32'hFC8D2304 , 32'hFF42A08C , 32'h029777E0 , 32'hFFEBEE1F , 32'h0233F7E4 , 32'hFEFC7A10 , 32'h095AD3E0 , 32'hFEA3BA14 , 32'hFEEA96AC , 32'hFF7F56E2 , 32'h001280F3 , 32'h02B88EEC , 32'hFFBAA6C3 , 32'hFC37FFDC , 32'hFC832D84 , 32'h014436D4 , 32'h00E3F4AC , 32'hFF065511 , 32'h01229A94 , 32'h0050A378 , 32'hFFFDA82B , 32'hFFFB182E , 32'h0000ED36 , 32'hFFFF396E , 32'h0001BB18 , 32'h00028F77 , 32'h0000AF40 , 32'h00016533 , 32'h0004C1F4 , 32'h00000038} , 
{32'h076CF3C8 , 32'hEF920AA0 , 32'h05F7A148 , 32'hEF1214A0 , 32'h09697450 , 32'hEE9BBDE0 , 32'hF379E9A0 , 32'hE6AF9760 , 32'hE29BA400 , 32'h0EE08130 , 32'h14D4CD20 , 32'hF9FB7170 , 32'hEFA60D00 , 32'hF05D3D90 , 32'hF4198610 , 32'hE9B70940 , 32'hFC4EEC24 , 32'h11D818A0 , 32'hEF1C2F40 , 32'hF60CD340 , 32'hFF7C9990 , 32'h06D07D00 , 32'hFA70C8A8 , 32'hFBEE56C8 , 32'h06C96F60 , 32'hF5BE13D0 , 32'hFC313C8C , 32'h075DD718 , 32'hEB3D4480 , 32'hEDC4AB00 , 32'h00401834 , 32'hF7D7CA90 , 32'hFD3E11C0 , 32'hFB0F1F48 , 32'h029CAB20 , 32'hFC187BD8 , 32'hF10D2D10 , 32'h120EA4A0 , 32'hFDC4BB3C , 32'hF2DF5580 , 32'h0DBF4280 , 32'h011F0448 , 32'h122F7920 , 32'hFFCB2BA7 , 32'hF3A6D5B0 , 32'h02F52398 , 32'h02BDA8B0 , 32'hFD170044 , 32'h06C31D40 , 32'h0A663B40 , 32'h03CC7484 , 32'h045103B8 , 32'h0B143CB0 , 32'h02F68388 , 32'hFD1EB5D4 , 32'h03AAEDD0 , 32'hED4E4EE0 , 32'hFBE7FF00 , 32'hFA6291C0 , 32'h060213B0 , 32'h028F6174 , 32'hFF66BC56 , 32'hF23E63B0 , 32'hFF8DB09F , 32'hFD973B58 , 32'hFED82324 , 32'hF8B1B778 , 32'hFFC9F888 , 32'h03647DD0 , 32'h05183518 , 32'hFDA2E960 , 32'h0360CA2C , 32'h0A458480 , 32'hFBA71FC8 , 32'hFD83E22C , 32'h030A6580 , 32'h01607020 , 32'hFEF15828 , 32'h00720019 , 32'h03A01E54 , 32'hFC6DE830 , 32'h0541A7C0 , 32'h012306A4 , 32'hF9D044B8 , 32'h00D12B2A , 32'hFED78F2C , 32'hFF43DFA4 , 32'h014DFCA0 , 32'hFEA25F18 , 32'hFF319E78 , 32'hFFFEE3E3 , 32'hFFFFB2DF , 32'h0001A29C , 32'hFFFE595A , 32'h0001277E , 32'h00000AC2 , 32'hFFFBCFFC , 32'hFFFEC745 , 32'h00009622 , 32'hFFFECC7E} , 
{32'h0DFA7D60 , 32'h03B6F490 , 32'hFEAC5548 , 32'h06CDAAC0 , 32'h10C857A0 , 32'h05930548 , 32'hEFCF6560 , 32'h0A448470 , 32'h1EDF4880 , 32'hEFB4D6C0 , 32'h0615C608 , 32'hFF6F6856 , 32'hFBBA1CD0 , 32'hF2B6E560 , 32'h0367F8AC , 32'hEDAC6AC0 , 32'h05D78EC0 , 32'h0801D460 , 32'h0FD45620 , 32'hFAEDDAE0 , 32'h0C4FBA70 , 32'hFF71B0FD , 32'hFF749BA5 , 32'h038C52C8 , 32'hF8F49BE8 , 32'hFE28E0F4 , 32'h171155E0 , 32'h088CEF10 , 32'h03CFF350 , 32'h058EF8C0 , 32'hFCCB7C5C , 32'h067A22F8 , 32'hFC675554 , 32'h0520D408 , 32'hF4061120 , 32'h0B641690 , 32'hFDE3D824 , 32'hFD86B450 , 32'h0CF99C30 , 32'h061FC330 , 32'hF4D19640 , 32'h15A340C0 , 32'hFC30E484 , 32'h02945BF4 , 32'hF342CA60 , 32'h0943C620 , 32'h078FDAB8 , 32'h035D0A70 , 32'hFD8D02B4 , 32'hF5318520 , 32'hFF10434C , 32'h09BD7D20 , 32'hF77FD200 , 32'h01C2FF6C , 32'hF732AE10 , 32'hFD913AA8 , 32'hFAE8FFA0 , 32'hF57CB4B0 , 32'hFFB5540B , 32'hFF758DAF , 32'h02783838 , 32'h038AB290 , 32'h0087B419 , 32'hFA303F30 , 32'h00C1C139 , 32'h01DBCA78 , 32'hFB99A260 , 32'hF8CB0A70 , 32'hFC9A11A8 , 32'hFFB0071F , 32'h00B0EFC3 , 32'hF9C7D3F8 , 32'hFB8C38C0 , 32'h02D34328 , 32'h038D87BC , 32'h02A7B55C , 32'h059CA0A8 , 32'h05E1E038 , 32'hFF4BCE3D , 32'h02F382B8 , 32'hFB2356E0 , 32'h00F541DF , 32'hFE59C438 , 32'hFFF76B74 , 32'hFD73B438 , 32'hFF2A2258 , 32'hFFC1BBA0 , 32'hFB05A6B0 , 32'hFF6CD123 , 32'h00443749 , 32'h000101F9 , 32'hFFFE8DDF , 32'h00007678 , 32'h0003472D , 32'h000179A8 , 32'hFFFE2E4E , 32'h00028A68 , 32'h0001C0F2 , 32'hFFFFA9F1 , 32'h0003099D} , 
{32'hFFFD6F9E , 32'h000257D3 , 32'hFFFE2D93 , 32'hFFFC715F , 32'h0004BE93 , 32'h00083361 , 32'hFFFD7D0D , 32'hFFFD514A , 32'hFFFF419D , 32'hFFFDE87B , 32'hFFFF99C6 , 32'hFFF8D882 , 32'hFFFFFC1C , 32'hFFFF8BB9 , 32'h0003E969 , 32'h00008E6E , 32'h000183B2 , 32'hFFFD315F , 32'h0002929B , 32'hFFFD178C , 32'h00006D1A , 32'hFFFBEC1A , 32'h0006E2DA , 32'h00011F40 , 32'hFFFFDEA6 , 32'h0000B3D4 , 32'hFFFEFDD6 , 32'h0004729D , 32'h0007039D , 32'hFFFEC44B , 32'h0001480D , 32'hFFFF0655 , 32'hFFFCFB88 , 32'hFFFCE3C9 , 32'h0004F2E8 , 32'h00022672 , 32'hFFFBFB47 , 32'h0007A05E , 32'h0002CD6C , 32'hFFFDF55B , 32'hFFFC7A10 , 32'h00008315 , 32'h0004A9D1 , 32'h00030AEC , 32'hFFFB4D60 , 32'hFFFBEA25 , 32'h0001B782 , 32'hFFF9643A , 32'h000300DE , 32'hFFFF76A3 , 32'h000433C5 , 32'h000113BE , 32'h00013DB2 , 32'hFFFEE518 , 32'hFFFFE5EF , 32'h0000B7DE , 32'hFFFBA2C8 , 32'h0000B57C , 32'hFFFFCACE , 32'h0002C15D , 32'h00030C48 , 32'hFFFFA48C , 32'hFFFFCA95 , 32'h000023D9 , 32'h00009476 , 32'hFFFBED3D , 32'h0003A6DF , 32'h00006A9A , 32'h000290C3 , 32'h00014205 , 32'h00003E87 , 32'hFFFF2543 , 32'hFFFD6D9D , 32'h00020AE1 , 32'hFFFF7F22 , 32'hFFFEACBA , 32'hFFF796A0 , 32'h0001D6F7 , 32'h000177C9 , 32'h000487C8 , 32'hFFFD4A9A , 32'h0003D918 , 32'hFFFFB296 , 32'hFFFC4BD7 , 32'h0004E71B , 32'h00005558 , 32'hFFFB406E , 32'h0002BFC8 , 32'hFFFFA827 , 32'h00051787 , 32'hFFFFD455 , 32'h0005089A , 32'h00042D5D , 32'hFFF9083B , 32'hFFFFAC14 , 32'hFFFE9153 , 32'hFFFD6F75 , 32'h0002C27B , 32'h0006C7FF , 32'h000305B7} , 
{32'h0EC9FB40 , 32'h32182040 , 32'h1AAB47A0 , 32'h13D1A260 , 32'h3120DB00 , 32'hF4F90B80 , 32'h0875F5F0 , 32'h0EF737A0 , 32'hFCFFD110 , 32'h19683840 , 32'hDE203240 , 32'h0C054AA0 , 32'h09F80A30 , 32'hFCD07D44 , 32'h08D60010 , 32'h19B7AF60 , 32'h080A95D0 , 32'hFDE908D0 , 32'hEE202760 , 32'h00BA05B9 , 32'h092C4240 , 32'h124D7800 , 32'h02C5B2D0 , 32'hEABD2320 , 32'h00B5268B , 32'h0BF3ACE0 , 32'hFA85FFA8 , 32'h09BB78C0 , 32'hF5FADBA0 , 32'h03DBAEEC , 32'hFE253474 , 32'h028426E8 , 32'hFA93E900 , 32'hFA2DF3A8 , 32'hEE64B820 , 32'h025C08E4 , 32'h0B19ABA0 , 32'hEE7F1B60 , 32'hFE495214 , 32'hF6080F10 , 32'hFAE411F8 , 32'h046132A8 , 32'h036B2FCC , 32'hFCB9C498 , 32'h0B00C5D0 , 32'h021CED80 , 32'h0391BD5C , 32'hFC357764 , 32'hF7EC5B50 , 32'hFC5ACDBC , 32'h032F9C68 , 32'hFF58AF74 , 32'hFC47FED0 , 32'h024C69F4 , 32'hFC691A0C , 32'h0775DD18 , 32'hF58E0080 , 32'hFD2EB494 , 32'hFC814318 , 32'hED57E4E0 , 32'h0116E158 , 32'h060A4CB0 , 32'h0283161C , 32'h03023D40 , 32'h053DA0D0 , 32'h032B6700 , 32'hFEA60090 , 32'hFFF96AD9 , 32'h03B8C21C , 32'h0922B7F0 , 32'hF62C1A70 , 32'hF6D31DA0 , 32'h00419EEB , 32'hF50CF230 , 32'h02909BE0 , 32'h075E4760 , 32'h02A9BEE0 , 32'h01E6EADC , 32'h00F28F7B , 32'h03A70134 , 32'hFE5937E4 , 32'hFBE15380 , 32'h0393821C , 32'hFF1BF8EB , 32'h00863452 , 32'hFE911800 , 32'h04271B70 , 32'hFF3EBACD , 32'hFF4DCD12 , 32'hFFC6CAC4 , 32'hFFFD4DD0 , 32'hFFFEE22F , 32'h00006D4D , 32'hFFFD73BF , 32'hFFFF0A1C , 32'h0001AAA0 , 32'hFFFEE95C , 32'h000047BA , 32'hFFFF4695 , 32'h00002969} , 
{32'hF8A59300 , 32'hFF3BE4AB , 32'h13251040 , 32'hD93ECFC0 , 32'hE623DAA0 , 32'hE3BB4CE0 , 32'hF4716660 , 32'h02D24B14 , 32'h2EA84700 , 32'h06CF2270 , 32'hFC89FAFC , 32'hFFF88D84 , 32'h089B6C80 , 32'h094CE3B0 , 32'h044FA780 , 32'hF7628960 , 32'hFEE42C28 , 32'h20576A00 , 32'h08612E30 , 32'h0FC045A0 , 32'hE72C5A00 , 32'hFC1B4540 , 32'hFE810578 , 32'hF5C39310 , 32'h081A4340 , 32'hFA42EEA8 , 32'h0315A3D0 , 32'h090EB120 , 32'hFA001388 , 32'hF6D89870 , 32'h104C3F80 , 32'hF424C440 , 32'hEC2EB020 , 32'hED5DB0A0 , 32'h042CEA68 , 32'hFBB4B340 , 32'hF7FA02A0 , 32'hFA9010C8 , 32'hFAC13BF0 , 32'h02BFD978 , 32'h04AB1C50 , 32'h0633AD00 , 32'hF010E8E0 , 32'h0B4875C0 , 32'h05DAEE18 , 32'hFC88DD98 , 32'hF5A4F5C0 , 32'h00158D99 , 32'hFEF493F0 , 32'hFA903E68 , 32'h03AF4328 , 32'hF766FE20 , 32'h04786D80 , 32'hFCBEEEF4 , 32'h053B64E0 , 32'hF4B85190 , 32'h047A5390 , 32'hFE3E6B38 , 32'h04345638 , 32'hFA317F90 , 32'hF8C08940 , 32'hFC914A98 , 32'h028D5A20 , 32'h0E0C75E0 , 32'h039878C0 , 32'h008966A0 , 32'h02119C3C , 32'h00F1D101 , 32'h051256D8 , 32'hFF02F631 , 32'hFA1260C0 , 32'h08B911E0 , 32'hF9D26498 , 32'hFDBA3840 , 32'h04280D68 , 32'h007B1DDC , 32'h013A8704 , 32'hFFEC31D5 , 32'hFFA6E206 , 32'hFCC6C894 , 32'hFAC65960 , 32'hFEEB76B0 , 32'hFC271BBC , 32'hFDDFBA50 , 32'h0125A5F4 , 32'h0369023C , 32'hFDDEF99C , 32'h05DF94B0 , 32'h026E73C0 , 32'h002D485A , 32'hFFFEF4E5 , 32'hFFFD9A9C , 32'hFFFF98D2 , 32'hFFFF4284 , 32'hFFFF77F2 , 32'h00000E91 , 32'h0001DE26 , 32'h0001D8DA , 32'h00004EE6 , 32'h00024628} , 
{32'h00023A8B , 32'h0000E54D , 32'hFFFDCAF3 , 32'h00038549 , 32'h00059698 , 32'h0002979B , 32'hFFFFB536 , 32'hFFFD0F0E , 32'hFFFE8FCB , 32'h000171DD , 32'h00003549 , 32'hFFFD46F0 , 32'hFFFEC65B , 32'h0001B91D , 32'h00062ACC , 32'h00044D4E , 32'h0001D46E , 32'hFFFF74A3 , 32'h000213C8 , 32'hFFFF8CC0 , 32'h00027763 , 32'hFFFE46DB , 32'h0000AF86 , 32'hFFFAF760 , 32'hFFFDD5C3 , 32'h00046A64 , 32'h000039AF , 32'h00039BC6 , 32'h0001A24E , 32'h0002CAA0 , 32'hFFFE8844 , 32'hFFFD760D , 32'hFFFE559B , 32'h0000C2AE , 32'hFFFD6CE3 , 32'hFFFF217A , 32'hFFFEACFB , 32'hFFFFB477 , 32'h00019F93 , 32'h0000C093 , 32'h000008EE , 32'hFFFDC1FB , 32'h000018A3 , 32'hFFFE921C , 32'h0001A7BD , 32'hFFFC409B , 32'h0002EBD3 , 32'h00021C16 , 32'hFFFF5BF8 , 32'h000064EB , 32'hFFFFDA64 , 32'hFFFFB160 , 32'h000221C5 , 32'hFFFE2982 , 32'h00010A2E , 32'h0001E003 , 32'hFFFBEB09 , 32'hFFFFEB28 , 32'hFFFDF032 , 32'hFFFF7066 , 32'h00023F14 , 32'h000195F8 , 32'h00006AF9 , 32'hFFFCDD10 , 32'h00008C4E , 32'h00044317 , 32'h00037EF6 , 32'hFFF8678E , 32'hFFFF21E1 , 32'hFFFCF6FF , 32'hFFFCC096 , 32'hFFFF6AA9 , 32'hFFFEED33 , 32'h0000757B , 32'h00037607 , 32'hFFFB9598 , 32'h0000528F , 32'h00016D83 , 32'h0001B9CE , 32'hFFF6DC61 , 32'hFFFFF7BA , 32'hFFFD0738 , 32'hFFFF42D4 , 32'h00012CF4 , 32'h0001014E , 32'hFFFFA85E , 32'h0004B02C , 32'hFFFB44AE , 32'hFFFB4A9B , 32'h000781F2 , 32'hFFFE0176 , 32'h0000200D , 32'h000129FB , 32'h0002A613 , 32'h0000F74E , 32'h0001318D , 32'h000318AE , 32'hFFFFCD96 , 32'h000215FF , 32'hFFFF5B28} , 
{32'h9FDE6000 , 32'h1F9D39E0 , 32'h24F53100 , 32'hEF1C7820 , 32'h05990168 , 32'h1EE389C0 , 32'hDD3D5180 , 32'h0F374D20 , 32'hEAE2C940 , 32'h1430BC60 , 32'hE6D43640 , 32'hFC2C8E4C , 32'hF26C79D0 , 32'h01A9FDE4 , 32'h0BE30610 , 32'h10059340 , 32'hFFF7131A , 32'h03C4CC30 , 32'hFEC2DF20 , 32'hFA816CC0 , 32'h091432B0 , 32'hF46D35E0 , 32'h046DCFD8 , 32'h0DC89E00 , 32'h04319240 , 32'h03B9FC9C , 32'hF983DE30 , 32'hF519FA70 , 32'hFDF17A40 , 32'h11B233A0 , 32'hFC279288 , 32'h1B9CCB40 , 32'hF6C3F120 , 32'h0CF87570 , 32'hFFD3BB12 , 32'hE7DA8320 , 32'hFC849568 , 32'hF42C5440 , 32'h0F362500 , 32'hFCB2F8BC , 32'h0C875BC0 , 32'hE5CBA760 , 32'h02A9B8D4 , 32'h09FB3F70 , 32'h007BB0A1 , 32'h02F5979C , 32'hF9EF2D48 , 32'hFB601D80 , 32'hF6B18E60 , 32'h03EE74F4 , 32'hF25D0C60 , 32'h00A49FCF , 32'hFC5C8A30 , 32'h0072690F , 32'hFBA1E120 , 32'hFA318260 , 32'h045225D8 , 32'h00A5BC2D , 32'h07A913E8 , 32'h089A0680 , 32'hFF99FB37 , 32'h0284AC64 , 32'h038D1788 , 32'h0153B150 , 32'h067F94F8 , 32'hFAB052D8 , 32'hFBD21A80 , 32'h05507258 , 32'hFD7AE928 , 32'h08335C10 , 32'h051D5D50 , 32'hFF9CCEDE , 32'hFEA6F5D4 , 32'h0285D2C0 , 32'hFD788938 , 32'hFDADB8F8 , 32'h05DFB648 , 32'h0648E898 , 32'h00478F36 , 32'h013E1E80 , 32'h0235CDA4 , 32'h030F7930 , 32'h002231E3 , 32'hFF2B9D19 , 32'h01902DAC , 32'h00E74147 , 32'hFD45CF88 , 32'hFE4EA150 , 32'hFF00CB25 , 32'hFFFC2045 , 32'hFFFFA1B1 , 32'hFFFFC0BB , 32'h000291FE , 32'hFFFF0075 , 32'hFFFFE7A1 , 32'hFFFF81A5 , 32'hFFFEA9A2 , 32'h000160AF , 32'hFFFFE325 , 32'hFFFFD774} , 
{32'hFFFD931C , 32'h00004687 , 32'h0000CA49 , 32'hFFFF2BA6 , 32'h0001B760 , 32'h00019679 , 32'hFFFE9DFE , 32'hFFFBB491 , 32'h00003986 , 32'h0002A89E , 32'hFFFEB6BC , 32'hFFFDCF3F , 32'h000097E7 , 32'h0002D53D , 32'hFFFFE2D4 , 32'h0004FD39 , 32'h0001C3BB , 32'h0001E024 , 32'hFFFFC1A8 , 32'hFFFD5D55 , 32'h0002C862 , 32'h0001FAD4 , 32'h000059D7 , 32'h00056051 , 32'hFFFE480E , 32'h00021213 , 32'h0000B74B , 32'h0000DB42 , 32'hFFFFE97D , 32'h0003C822 , 32'h00017F78 , 32'h0003649A , 32'h0001C98C , 32'h00008287 , 32'h0002B584 , 32'h0001F19B , 32'hFFFBBDA1 , 32'hFFFD13B2 , 32'h00001EA3 , 32'h00054019 , 32'h000092CF , 32'hFFFDAEF1 , 32'h00048035 , 32'h0002750E , 32'hFFFF23A0 , 32'h0003191F , 32'hFFFD219B , 32'h00034886 , 32'hFFFE83EA , 32'h0001FE9C , 32'hFFFABD8C , 32'hFFFFA55B , 32'h00015995 , 32'h0001A24F , 32'hFFFF5327 , 32'h00029573 , 32'h00008D6B , 32'h0005B81F , 32'hFFFF0BBD , 32'hFFFF5022 , 32'h00003052 , 32'hFFFC41AE , 32'h00022907 , 32'h000046F8 , 32'h000052AF , 32'h000160D9 , 32'h0003AD11 , 32'hFFFBDD1E , 32'hFFFC5B34 , 32'h00037D4D , 32'hFFFD0630 , 32'hFFFCE7A5 , 32'h0004CC9E , 32'h0001EFE7 , 32'h000229D8 , 32'h0000B93B , 32'h0001C3E0 , 32'h000238A6 , 32'h000060BC , 32'hFFFB81E2 , 32'h00026EEC , 32'h00017CD4 , 32'hFFFCA71D , 32'hFFFDEBBA , 32'h0004176C , 32'hFFFFDE08 , 32'hFFFC4ACD , 32'h000341BA , 32'h0003E3DE , 32'h00023789 , 32'hFFFFB674 , 32'h00034D89 , 32'hFFFFB430 , 32'hFFFDF80A , 32'hFFFC92E2 , 32'hFFFFC706 , 32'hFFFE9B8D , 32'h0003A99B , 32'hFFFDC303 , 32'hFFFED7AA} , 
{32'h1430D6E0 , 32'hEFC40820 , 32'hE99FB6C0 , 32'hD6D537C0 , 32'hF7989470 , 32'hE50951E0 , 32'h09F9AF30 , 32'hFA310FE0 , 32'hF4680BD0 , 32'h0783D988 , 32'h0B851150 , 32'h1168FB80 , 32'hFFCAE9A4 , 32'hE48092A0 , 32'h05176AB8 , 32'h1B7D2680 , 32'h0292F1FC , 32'hFF04CDAE , 32'hFF8C319F , 32'hFBE7AD68 , 32'hF3C1B0E0 , 32'h072BF070 , 32'hF2CBE330 , 32'h0144F914 , 32'hFEADA130 , 32'h150A9B40 , 32'hF3D111F0 , 32'hFDD8F060 , 32'hEDF0F240 , 32'h0770BBC8 , 32'h0A2E1550 , 32'hFC1DC0F0 , 32'hFF1B3BC4 , 32'h096D8AB0 , 32'h10B2F160 , 32'h01010BA8 , 32'h0C6781A0 , 32'hF985E148 , 32'hF458D520 , 32'h05CD7320 , 32'hFBA2A008 , 32'h0D6A30B0 , 32'hF8EA2350 , 32'h06EE9188 , 32'hFD164A78 , 32'h03D6BE38 , 32'hF8C54410 , 32'hF86ADEA0 , 32'hF6B8AB10 , 32'hF61722B0 , 32'hFBBDE2D0 , 32'h02ACDC94 , 32'h00A4055E , 32'hFBD25B00 , 32'hF760CE20 , 32'h05E94338 , 32'h02AA2590 , 32'hFF4110F1 , 32'h09395E70 , 32'hF6AD5990 , 32'h001F6BAF , 32'hFCD2686C , 32'h03E59804 , 32'hF4334400 , 32'hF3A4F5D0 , 32'hFDCC8728 , 32'hFCB25934 , 32'h02CA3274 , 32'hFE19C458 , 32'hFFE87F99 , 32'hFF6F300A , 32'hFFEBF2D0 , 32'hF8B09208 , 32'h02118D34 , 32'hFDEBB4D8 , 32'h01E95FDC , 32'h00895808 , 32'hFF292014 , 32'h082B5680 , 32'h03E9B4EC , 32'h006ABF75 , 32'h02812B54 , 32'h013E57EC , 32'hFC129EE8 , 32'hFBF6F590 , 32'h0091C904 , 32'h0087B938 , 32'h02505694 , 32'h015C7E28 , 32'hFFD78EEE , 32'hFFFFAA37 , 32'h0000CC3A , 32'hFFFDE71E , 32'h0002CA89 , 32'h0000D5B4 , 32'hFFFE2C18 , 32'hFFFE603C , 32'h0001A67E , 32'hFFFF700F , 32'h00016A9C} , 
{32'h201DE480 , 32'hD70FCE80 , 32'h036D02D4 , 32'h1B9B7640 , 32'hDCAA0940 , 32'h2EFFF140 , 32'h28F54140 , 32'h0570AF50 , 32'hEC614080 , 32'hE4DF90E0 , 32'h0FF300B0 , 32'h130419A0 , 32'hFFF0D22C , 32'h1A4FF4E0 , 32'hDE256EC0 , 32'h113C0B00 , 32'h0CA65880 , 32'h21EA2F00 , 32'h095A09C0 , 32'hE5416F80 , 32'hFF32A344 , 32'hFF40EE73 , 32'h0AA620B0 , 32'hEBDCE800 , 32'hF4EDCD80 , 32'h0878C8F0 , 32'hF4ABC960 , 32'hED03DD60 , 32'hFCCCD484 , 32'hEF674340 , 32'hFCC37DE8 , 32'hEFFDB220 , 32'hF24CD1B0 , 32'h0010D92B , 32'hF9244BD8 , 32'hFFA235C8 , 32'h04FFA798 , 32'hF5F9A050 , 32'h03F30C7C , 32'h096B47A0 , 32'hF63FC900 , 32'hF6F2DF70 , 32'h09B1F7A0 , 32'h06E02C98 , 32'h1AB353E0 , 32'h00DB6794 , 32'h007F4687 , 32'h040B1898 , 32'hF9806610 , 32'hFE69DDCC , 32'h037B3CA0 , 32'hFB178670 , 32'hFEFA41F8 , 32'hF9AEF928 , 32'h011FE1C4 , 32'h03CACB24 , 32'hFA5814F0 , 32'hF7D320D0 , 32'hFE6328F4 , 32'hFC97CE94 , 32'h04935C20 , 32'hFD993A7C , 32'hF8380DE0 , 32'hFC5838B8 , 32'h07836838 , 32'hFA7B0E20 , 32'hFE61A330 , 32'hFBA49168 , 32'h02A7B4AC , 32'hFCC54200 , 32'h07AFF3B8 , 32'h04965728 , 32'hFFBC37D4 , 32'h006EDDD3 , 32'h0042F62E , 32'hFEC23958 , 32'h0305A268 , 32'h0083C26B , 32'h021AA0D8 , 32'hFCFB2FA4 , 32'hFC492448 , 32'hFDBF1CFC , 32'hFFABD84A , 32'hFE96A674 , 32'h00D44659 , 32'h005903D7 , 32'h024F4130 , 32'hFEDD041C , 32'h01BAC8B4 , 32'hFF5FBB1C , 32'hFFFEC483 , 32'h0001FD87 , 32'h0000D400 , 32'h00019087 , 32'hFFFFC21A , 32'h0000757D , 32'h00011067 , 32'h000230A6 , 32'h00048043 , 32'hFFFFAB88} , 
{32'h00022489 , 32'hFFFCE01C , 32'hFFFF43EA , 32'hFFFF75C3 , 32'hFFFF53E1 , 32'h00007EC4 , 32'hFFFD0005 , 32'hFFFBFBF9 , 32'hFFFC7C37 , 32'h00069E3A , 32'hFFFB2C4A , 32'h0001AAD5 , 32'h0002D67D , 32'hFFFE68C3 , 32'h000681F9 , 32'h00007BD7 , 32'h00008184 , 32'h00006E0D , 32'h0004F62A , 32'h0000C52A , 32'h00009D3F , 32'hFFFB3FBC , 32'h000206C5 , 32'h0004BC67 , 32'hFFFFAE0E , 32'hFFFEB476 , 32'hFFFFD359 , 32'hFFFF2419 , 32'h000173B3 , 32'h00041BFC , 32'hFFFFFF88 , 32'hFFF9FAC6 , 32'hFFFFFF35 , 32'hFFFE018E , 32'h00016FFE , 32'hFFFE14FD , 32'h00019003 , 32'h00011ADF , 32'h0000ECA4 , 32'h0002B5FE , 32'h00002E47 , 32'hFFFD6D03 , 32'hFFFC2611 , 32'hFFFD7CEC , 32'h00030F34 , 32'hFFFB25C3 , 32'h000014CC , 32'hFFFFFFEA , 32'h00039989 , 32'h0001DA93 , 32'h00031FA6 , 32'h00009EFA , 32'hFFFBC23A , 32'h00035457 , 32'hFFFD55B6 , 32'hFFFE2D8D , 32'h00039CA1 , 32'h00019070 , 32'hFFFF780A , 32'h000124FE , 32'h0001DE55 , 32'hFFFEB0A6 , 32'h00014C00 , 32'hFFFF16A5 , 32'h00016ADA , 32'h00010039 , 32'h0001131A , 32'h00011124 , 32'hFFFE1420 , 32'hFFFE0D1D , 32'h0002D074 , 32'h00014AFF , 32'hFFFE14A3 , 32'h0001B827 , 32'h000525C6 , 32'h000125A3 , 32'h0000CCDE , 32'hFFFA6FEB , 32'hFFFFE503 , 32'hFFFF79D4 , 32'hFFFB69AB , 32'h000102FA , 32'h0000B68F , 32'h000172CE , 32'hFFFFC50C , 32'hFFFE2716 , 32'h00034B64 , 32'h0002DA4D , 32'h00033DA0 , 32'h00010962 , 32'h00021E99 , 32'h00013B1C , 32'h00015BB3 , 32'h00024E11 , 32'h00029692 , 32'h00021044 , 32'hFFFDE7EA , 32'h0000065C , 32'h0000D297 , 32'hFFFFF413} , 
{32'hFFFAE0A0 , 32'h00006C2C , 32'hFFFF1E97 , 32'hFFFDE59C , 32'h00019531 , 32'hFFFF9F06 , 32'h000014C8 , 32'h00026057 , 32'hFFFC6D28 , 32'h0000D690 , 32'hFFFEC374 , 32'h00000DE7 , 32'h0001ABF0 , 32'hFFFE5783 , 32'h0003C9C3 , 32'hFFFE3D6F , 32'h0003BA31 , 32'hFFFEEA4C , 32'h00021047 , 32'hFFFD02B4 , 32'h0002DCA1 , 32'h000346FD , 32'hFFFD2A57 , 32'h000138F4 , 32'h00011766 , 32'hFFFC458F , 32'hFFFECE00 , 32'hFFFCA02E , 32'hFFFF9956 , 32'h00010578 , 32'hFFFCEDB7 , 32'hFFFB8095 , 32'h00008B11 , 32'hFFFCA588 , 32'h0000C20B , 32'hFFFF6964 , 32'h0001EFD8 , 32'hFFFD4448 , 32'hFFFFFD4A , 32'hFFFF2127 , 32'h00045EEF , 32'hFFFCFE22 , 32'h0000BFB1 , 32'hFFFEBC0B , 32'hFFFDADC7 , 32'hFFFED9AF , 32'h00005CEE , 32'hFFFC446C , 32'h00043390 , 32'hFFFE0C6E , 32'hFFFC0AA0 , 32'hFFFF689A , 32'h00039295 , 32'h0003E659 , 32'h0000BCDC , 32'h00002E99 , 32'h0003B960 , 32'h0002E2A4 , 32'hFFFBE5E0 , 32'h0001534B , 32'hFFFBA6D2 , 32'hFFFEB59F , 32'hFFFF9389 , 32'h00009F7B , 32'h0002BA04 , 32'h00039AEB , 32'h0003DF3C , 32'h0002AD1A , 32'hFFFBD3A9 , 32'h0000E24D , 32'h00049ADB , 32'h0001DED7 , 32'h000004CD , 32'h0001B362 , 32'hFFFC0BFC , 32'h00051361 , 32'h0000D587 , 32'h00030992 , 32'h00012556 , 32'hFFFEC6DC , 32'h00043361 , 32'hFFFE0298 , 32'h0002045F , 32'hFFFFBFFF , 32'hFFFDB9D0 , 32'h00041EBD , 32'hFFFD1FA8 , 32'h00035F67 , 32'h000299AA , 32'h0000EFA8 , 32'hFFFCC782 , 32'hFFFEB757 , 32'h0001E23B , 32'h00007D55 , 32'h0002A514 , 32'h00022122 , 32'h00021C8B , 32'h0001537B , 32'h00031B14 , 32'h00031F44} , 
{32'hFFFD77B0 , 32'h0000DCD6 , 32'h000012A5 , 32'hFFFCCC2C , 32'hFFFF9E7A , 32'h00029C68 , 32'hFFFD0B26 , 32'h0004B138 , 32'hFFFF9197 , 32'h00004789 , 32'h00010CD6 , 32'h0000CB35 , 32'h0003789B , 32'h00042236 , 32'h00018A3A , 32'h0001D89B , 32'hFFFFF7A5 , 32'h0000843B , 32'h00028422 , 32'hFFFEFB10 , 32'hFFFCED68 , 32'hFFFD9103 , 32'hFFFF2590 , 32'hFFFF8D3E , 32'hFFFDD72D , 32'h000133EE , 32'h00011FB9 , 32'h0001B16B , 32'h000085C0 , 32'hFFFE755F , 32'h00004E7D , 32'hFFFDEBCF , 32'h0004FA0A , 32'hFFFA7789 , 32'hFFFF8209 , 32'h00051216 , 32'hFFFF083E , 32'h00025E11 , 32'hFFFCD562 , 32'h00013EA6 , 32'h0003C952 , 32'hFFFF7255 , 32'hFFFEEE51 , 32'hFFFDAF73 , 32'h000304B5 , 32'h0002C1A6 , 32'h00014A29 , 32'hFFFF8A6D , 32'hFFFF5376 , 32'hFFFFC2A2 , 32'hFFFF5E22 , 32'h00023F59 , 32'hFFFE28EE , 32'h00011AAB , 32'h0002EDFE , 32'h00004CA1 , 32'h00038251 , 32'h0000757F , 32'h000235DA , 32'h0001CA6D , 32'hFFFAD657 , 32'h0003C8AD , 32'h00013074 , 32'h00019722 , 32'hFFFC63F2 , 32'h0004ADB6 , 32'hFFFF2464 , 32'h0000589D , 32'h0000A522 , 32'h0002E070 , 32'hFFFEE6D5 , 32'hFFFE2EA2 , 32'h000191A7 , 32'hFFFE4B12 , 32'hFFF9F899 , 32'hFFFF9AC3 , 32'h00006FB0 , 32'h0000151D , 32'h0001A3B1 , 32'h0000A5F7 , 32'hFFFFE747 , 32'hFFFC4E1D , 32'hFFFE4A59 , 32'h0003B706 , 32'hFFFF5A7F , 32'h00044843 , 32'hFFFA9FE1 , 32'hFFFEB12F , 32'h0001FB3A , 32'hFFFFF2F4 , 32'hFFFE6DB4 , 32'h00010DD5 , 32'hFFFF570D , 32'hFFFED9DF , 32'hFFFECECC , 32'hFFF67C73 , 32'h0003257D , 32'hFFFDB085 , 32'hFFFDFAAE , 32'hFFFEAFC5} , 
{32'hFFFBB54E , 32'hFFFF79A7 , 32'h00002941 , 32'h0000104F , 32'hFFFD21DA , 32'h00024676 , 32'hFFFF5750 , 32'h0001AB45 , 32'hFFFEA568 , 32'hFFFE30BA , 32'h00002A20 , 32'h0000CE40 , 32'h0003705C , 32'h00009BD2 , 32'hFFFF9C2B , 32'hFFFFFC57 , 32'hFFFAFC6F , 32'h0003064D , 32'h00016DA9 , 32'h0003CEF5 , 32'hFFFE0AFB , 32'hFFFE3B2B , 32'hFFFD4CC6 , 32'h0000B10E , 32'hFFFFCCC3 , 32'hFFFEB448 , 32'hFFFE24DB , 32'hFFFDD6A3 , 32'hFFFE3070 , 32'h0002B509 , 32'h00026813 , 32'hFFFDDF5B , 32'hFFFEF613 , 32'h00067FDF , 32'h00014B06 , 32'h00001AFC , 32'hFFFE1507 , 32'hFFFE6F5C , 32'hFFFA6A70 , 32'hFFFFE14A , 32'h0000DFE9 , 32'h00039148 , 32'h00014248 , 32'h00027660 , 32'h00009515 , 32'h00057687 , 32'hFFFD4323 , 32'hFFFE8728 , 32'h00036360 , 32'h00012AA5 , 32'hFFFD84F6 , 32'hFFFCCED9 , 32'hFFFDC667 , 32'hFFFF37DB , 32'hFFFA3911 , 32'h00005B25 , 32'hFFFE5242 , 32'h0006DD3C , 32'hFFFC4381 , 32'hFFFF0B6A , 32'hFFF85A73 , 32'h00003D70 , 32'hFFFDA227 , 32'hFFFD9524 , 32'h000043BC , 32'hFFFE7EFD , 32'h0002C9C9 , 32'hFFFCC7EB , 32'hFFFF9D66 , 32'hFFFC1CA9 , 32'hFFFBC2DE , 32'hFFFD7B89 , 32'h0002DE8F , 32'h00027D6A , 32'h0003BE66 , 32'hFFFFF737 , 32'hFFFC4BAF , 32'hFFFF52EE , 32'hFFFCBCCC , 32'h00013687 , 32'h00054EBA , 32'hFFFCED07 , 32'hFFFD87D0 , 32'hFFFFB592 , 32'hFFF7C2C6 , 32'h00026B8E , 32'h000059EA , 32'h000463B5 , 32'h00018D71 , 32'h0001CF7F , 32'hFFFE78BC , 32'h00045186 , 32'hFFFE9254 , 32'hFFFF5B19 , 32'hFFFDCEE5 , 32'h00016024 , 32'h00019E72 , 32'hFFFE0405 , 32'h0003AA20 , 32'h00015413} , 
{32'hFFFB9CB2 , 32'hFFFFAE95 , 32'h0001525A , 32'hFFFEC286 , 32'hFFFEFD6F , 32'h000167E9 , 32'hFFFECCC9 , 32'hFFFE553E , 32'hFFFE946D , 32'h00007F39 , 32'hFFFE8B7D , 32'h0000174D , 32'hFFFC6055 , 32'h000184E3 , 32'h0000DE50 , 32'hFFFE5115 , 32'h00004948 , 32'hFFFB3F34 , 32'hFFFD6E30 , 32'h00073070 , 32'hFFFE9E79 , 32'hFFFD0524 , 32'hFFFE144B , 32'hFFFE8187 , 32'h00003007 , 32'h0000F2AF , 32'hFFFF487B , 32'hFFFE914F , 32'hFFFC8856 , 32'hFFFC815A , 32'hFFFF413E , 32'h000005C2 , 32'h00004E67 , 32'h0000EB2A , 32'h00021AF1 , 32'h00005EE2 , 32'h00001365 , 32'hFFF92C35 , 32'hFFFBCEE5 , 32'h00018735 , 32'hFFFD656C , 32'hFFFF9D72 , 32'hFFFF9E62 , 32'h00007CC8 , 32'hFFFF2BD6 , 32'h0004F2F8 , 32'h00015292 , 32'h000148DA , 32'h0000AC5A , 32'hFFFF7841 , 32'h00023549 , 32'h00022C77 , 32'h0002DC1B , 32'hFFFED3A1 , 32'h00024028 , 32'h000284C5 , 32'hFFFEB766 , 32'hFFFEE0AE , 32'hFFFDFA40 , 32'hFFFCE7BC , 32'hFFFF89B8 , 32'hFFFF79F2 , 32'hFFFEC6E0 , 32'hFFFCAB8E , 32'h00026B64 , 32'h0003C152 , 32'hFFFF4B83 , 32'hFFFED622 , 32'h0002B998 , 32'hFFFC58F2 , 32'hFFFEA538 , 32'hFFFD36F6 , 32'h0000F869 , 32'hFFFFBE19 , 32'h0001F531 , 32'hFFFDFDB5 , 32'h0001149D , 32'h0001D75A , 32'hFFFD7081 , 32'hFFFD4EE3 , 32'hFFFDC0C3 , 32'hFFFF1C60 , 32'h0001DA06 , 32'h0005EB82 , 32'h0000DADE , 32'h0000A19C , 32'hFFFF8F1A , 32'hFFFEE041 , 32'h00037C94 , 32'hFFFFBD53 , 32'h0004FBEE , 32'h00017DF0 , 32'h00026337 , 32'h000181A5 , 32'h0002B52B , 32'hFFFCDACE , 32'hFFFEEB85 , 32'hFFFBFB3C , 32'hFFFFCAFD , 32'h0000008F} , 
{32'h00015DD8 , 32'h0002D12D , 32'h000293D8 , 32'h00030267 , 32'hFFFFCD00 , 32'h000073E3 , 32'h0002AAD9 , 32'hFFFDAA0E , 32'h0001960E , 32'h00016A97 , 32'hFFFC5A9B , 32'h00030CC2 , 32'hFFFFE1A4 , 32'hFFFD3942 , 32'hFFFBCD24 , 32'h00012CA6 , 32'h0002EEF3 , 32'h000563C2 , 32'h00009551 , 32'hFFFEAB4F , 32'hFFFD133A , 32'h000185B1 , 32'h00018D8C , 32'hFFFD2221 , 32'hFFF9A7B9 , 32'hFFFE9C8B , 32'h0001123F , 32'h00030517 , 32'h0003A429 , 32'h0002FC38 , 32'hFFFE628D , 32'hFFFA1F0F , 32'h00020BA6 , 32'h00019304 , 32'hFFFC0DA5 , 32'hFFFF6B90 , 32'hFFFE47DD , 32'hFFFF4756 , 32'h0002C25F , 32'hFFFEA6F7 , 32'hFFFF1052 , 32'h000261A6 , 32'h0000FC85 , 32'h00037A9C , 32'hFFFD9071 , 32'h0003D21F , 32'hFFFB20FC , 32'h0000614E , 32'h0000B756 , 32'hFFFCE39E , 32'hFFFFB6B9 , 32'hFFFC2C3B , 32'h0001519C , 32'hFFFAE6D0 , 32'hFFFC8C19 , 32'h00019A0C , 32'hFFFEEE0D , 32'hFFFFD022 , 32'h000129D0 , 32'h00027E2B , 32'h00019EFB , 32'h00010896 , 32'h00015BB7 , 32'h00014E81 , 32'h0001DA7F , 32'hFFFE67AE , 32'h0003C06F , 32'hFFFEE039 , 32'h00014E9A , 32'h0002049B , 32'hFFFC05E0 , 32'hFFFED3BE , 32'h000028FA , 32'hFFFF62FA , 32'h00016256 , 32'h0001C1F9 , 32'h000311E9 , 32'hFFFF81D7 , 32'hFFFE622B , 32'hFFFC4D28 , 32'hFFFDC3EC , 32'h00004DD1 , 32'hFFFCFBDB , 32'hFFFFA0D4 , 32'hFFFEF71C , 32'h0002591E , 32'h00042F3C , 32'h0000C1EA , 32'h0004A45B , 32'hFFFC7443 , 32'hFFFFC8BE , 32'h000409E1 , 32'h00009A47 , 32'h000226CA , 32'hFFFEB542 , 32'hFFFD0D79 , 32'hFFFD46B0 , 32'hFFFE93D1 , 32'hFFFC1D53 , 32'h00003104} , 
{32'h032AC040 , 32'hE1F091C0 , 32'h00D2E975 , 32'h12749A40 , 32'hF7D31370 , 32'hFD9FC408 , 32'h0B122430 , 32'hED01AA00 , 32'hF01C4F80 , 32'hF820D6D0 , 32'h07857F00 , 32'h0A352710 , 32'h0D495190 , 32'h07E08FA8 , 32'h0FBFF270 , 32'hF0D0C3F0 , 32'h01394DF8 , 32'h13351CA0 , 32'hF144FD80 , 32'h0F141F10 , 32'h0EF27A60 , 32'hFB4ACF70 , 32'hFBB0A620 , 32'hF3DFFEA0 , 32'h0B8233A0 , 32'h0173DF08 , 32'h02E3600C , 32'h077E4FA0 , 32'h0361B778 , 32'hFD1B8FC4 , 32'hFDE06A98 , 32'hF674F060 , 32'hF95B5858 , 32'h0522E648 , 32'h00165DC0 , 32'h03489ACC , 32'h0217E200 , 32'hFC654C4C , 32'hFC8F4E30 , 32'h0387C1D0 , 32'h01A760E8 , 32'h086741D0 , 32'hFA0AD190 , 32'hFE352E70 , 32'hF60AD430 , 32'hFCF82424 , 32'h0327BE24 , 32'hFD546B10 , 32'hF85CD150 , 32'h076B03B8 , 32'hF8DEF5C8 , 32'hF503FEE0 , 32'hFE3098C0 , 32'hF8139C18 , 32'hF4F50780 , 32'h0867FB90 , 32'h04452E90 , 32'h0038CAEC , 32'hFC3DA328 , 32'h04CE05A8 , 32'hFF8789E5 , 32'h00EAF6FE , 32'hFA4D3348 , 32'hFF620B94 , 32'hF8E05130 , 32'h02EF4A00 , 32'hFAD01118 , 32'h09EC4D90 , 32'hFCAA6498 , 32'hFEFCEAC0 , 32'h03C075F4 , 32'hFB6DEC98 , 32'h0334C4FC , 32'h0344A124 , 32'hFDAE73BC , 32'h01ED7B2C , 32'h04319270 , 32'hFBD6C8A8 , 32'hFAF7DEE8 , 32'hFDE6C414 , 32'h01F33B08 , 32'h02ADF2A8 , 32'hFF324704 , 32'hFEE9DEC0 , 32'h03ADDECC , 32'hFD6B5234 , 32'hFE8F2B98 , 32'h02E303B0 , 32'h03173470 , 32'hFFE881C1 , 32'hFFFC4AA1 , 32'hFFFFDA14 , 32'h00022D0C , 32'hFFFC260A , 32'hFFFECCB9 , 32'hFFFFF208 , 32'h000034D5 , 32'h0000CE0B , 32'hFFFF510C , 32'h00022804} , 
{32'hF0B34A00 , 32'hA9D16900 , 32'h10A3BAA0 , 32'h0A423E80 , 32'hFE69C0A8 , 32'hF9F675A8 , 32'h225CF7C0 , 32'h1FF9AB20 , 32'hFC533E18 , 32'hE40CD460 , 32'hEC16C9E0 , 32'h064A9760 , 32'hF70A77D0 , 32'hF88A68B8 , 32'h14628C80 , 32'hFB14B990 , 32'hFF21724B , 32'h037A5134 , 32'h02120734 , 32'h07323010 , 32'h016802B4 , 32'hFD05C6E4 , 32'hF4709A80 , 32'h0955FAB0 , 32'hF3A0F550 , 32'hFFE392CA , 32'hFDF9FF78 , 32'h02F2EFDC , 32'hFA0B5CC0 , 32'h039D24C8 , 32'hEFF45BE0 , 32'hFA7F12F0 , 32'h0E238860 , 32'hFC3AE108 , 32'hF9ABFDD8 , 32'hFFAA3417 , 32'hEF116EE0 , 32'h18ECD7C0 , 32'hED0171C0 , 32'hFE538640 , 32'hF721EA50 , 32'hFDA6B0BC , 32'h0DC89600 , 32'hF906F520 , 32'h0077155A , 32'hFD34CBC0 , 32'hFC4FB394 , 32'hF1173E50 , 32'h000C3288 , 32'hFA4D0A60 , 32'hF8364340 , 32'h057902F0 , 32'h0179D5D8 , 32'hF0D7A2F0 , 32'h0AA25BE0 , 32'hFAF57A80 , 32'h0B16B9E0 , 32'hF8143178 , 32'hFDC429C8 , 32'hF55ED6A0 , 32'h0B10A590 , 32'h015883F0 , 32'hFF6C68C0 , 32'h04CAF540 , 32'hFF814C24 , 32'h02197744 , 32'h06B34320 , 32'hFD4411C4 , 32'h0A3928D0 , 32'hFC0FAD24 , 32'hFC7C355C , 32'h0393C620 , 32'h05A7ABD8 , 32'hFF3D8EB3 , 32'h075D3950 , 32'h04C2C708 , 32'h048DB640 , 32'hFD23B4BC , 32'hFEBCEFD0 , 32'h00B1F909 , 32'h02D45504 , 32'hFEAB3128 , 32'hFF1D0195 , 32'h017C3FD4 , 32'hFFD250A7 , 32'h022FA86C , 32'h054D09E8 , 32'h010120AC , 32'hFDE0FB78 , 32'hFF341FD0 , 32'h0002123E , 32'h000095E4 , 32'h00026427 , 32'hFFFDF6F4 , 32'hFFFDED3E , 32'hFFFC197B , 32'h000111E9 , 32'h00010C2D , 32'hFFFF52CE , 32'h000071BB} , 
{32'h3603C5C0 , 32'hFA375308 , 32'hCD7B80C0 , 32'h30EB1B00 , 32'hE8AE73A0 , 32'hF4E5E2B0 , 32'hF9278488 , 32'h19BDEAE0 , 32'h2A819740 , 32'hEA04E480 , 32'hF0149710 , 32'h0134E320 , 32'hD69E2DC0 , 32'h0CA68F00 , 32'h0573A2A0 , 32'hFFDFBDF3 , 32'h0E7A2830 , 32'h1D7A2F40 , 32'h044152C0 , 32'h0F928960 , 32'h01087BB0 , 32'hEEACB480 , 32'hF48F24F0 , 32'h14B66680 , 32'h150990C0 , 32'hFC940974 , 32'h03EB4AC4 , 32'hF9A87888 , 32'h028E9E40 , 32'hFD6D9C34 , 32'h08E632D0 , 32'h07EF9D18 , 32'h08B69A50 , 32'hF838FBC0 , 32'hFA950020 , 32'hFE8C59F8 , 32'h00CAD26B , 32'h036C88C8 , 32'hEB074420 , 32'h0CC0A010 , 32'hF9EE38A8 , 32'h01F4401C , 32'h08FFE000 , 32'hF27B15E0 , 32'hF8FDA840 , 32'h026807FC , 32'h0A04BEA0 , 32'hF8BDDB40 , 32'h043FB458 , 32'h0F1C76A0 , 32'hE74E1900 , 32'h064DD5B0 , 32'h03DBBE34 , 32'h0035A73B , 32'h07EAAC40 , 32'h0D0175C0 , 32'h0388D7F0 , 32'hF62A4360 , 32'hFC444B60 , 32'h026A34B0 , 32'hFDD3BE90 , 32'h062B6508 , 32'hFEC8CC68 , 32'h003182AB , 32'hFA848518 , 32'h05EE4148 , 32'h00D056C0 , 32'hFE8763A8 , 32'hFEB20C20 , 32'hFFEA4194 , 32'h011E375C , 32'h00D877D5 , 32'h03B2EA28 , 32'h008F4B41 , 32'h037624FC , 32'h037FB3D0 , 32'hFB81E318 , 32'h068B1B98 , 32'h0300F61C , 32'hFB07C5B0 , 32'hFE541150 , 32'hFD6A1E30 , 32'h0162BEC4 , 32'hFDCA8498 , 32'h01568EC4 , 32'hFFB13616 , 32'h01019E60 , 32'h001304B0 , 32'hFDB49B04 , 32'h00C37CDF , 32'hFFFF0752 , 32'hFFFEC764 , 32'hFFFDBA15 , 32'h0002B995 , 32'h0000D299 , 32'h00037517 , 32'hFFFF42A4 , 32'hFFFED448 , 32'h00008506 , 32'h00005D2E} , 
{32'h0F782B60 , 32'hFC8411B8 , 32'hFEF668F0 , 32'h06F4E328 , 32'hDF8CDF80 , 32'hEFCB19A0 , 32'hEF935E80 , 32'h064A4B90 , 32'h13D79FC0 , 32'hE5B4F580 , 32'hFEE3A884 , 32'hFF10314C , 32'h00641CF8 , 32'hF1BCAAA0 , 32'h0A842230 , 32'h13FAF220 , 32'h0C761B10 , 32'h0657EDB8 , 32'hF5B8E7E0 , 32'hF80A18A8 , 32'hFA25E808 , 32'hF1853730 , 32'hF89AAB60 , 32'h07B65620 , 32'h03F9EE8C , 32'hF18EC8C0 , 32'h113E6520 , 32'h0172C560 , 32'hF95767F8 , 32'h11842540 , 32'hE7B98280 , 32'h0215ADC8 , 32'hF4974300 , 32'h10065640 , 32'hFBECB540 , 32'hF8E49698 , 32'hFE44324C , 32'hF3109610 , 32'h04260C58 , 32'h0E569CE0 , 32'h04978AD8 , 32'h0264A004 , 32'h067121D8 , 32'h01D87670 , 32'hFF937822 , 32'h0CA77DA0 , 32'hFE43F758 , 32'hF49F6650 , 32'h123DB9A0 , 32'hFF03BF11 , 32'h05A684D0 , 32'hEE61E2C0 , 32'hFAFA7C30 , 32'h05EC70C8 , 32'h01AC500C , 32'h04CBA028 , 32'hF8CDDDA8 , 32'h052C5250 , 32'hFAC41858 , 32'h04238F38 , 32'hFE7EE8BC , 32'hF85F5808 , 32'hFCB3CF84 , 32'hFB586CF0 , 32'h06607218 , 32'hFEABED40 , 32'hF8B3E2E0 , 32'hFFA7CBD3 , 32'h053E1120 , 32'h03136410 , 32'hF7A4C4F0 , 32'h06922C08 , 32'h04016A70 , 32'h0413E110 , 32'hFE5BAD04 , 32'hFE4517FC , 32'h04177700 , 32'h00300D97 , 32'hFE294380 , 32'hFF0FBAC2 , 32'hFD2CCD38 , 32'h00EE6A18 , 32'h0117A720 , 32'h03523C18 , 32'hFF7D467C , 32'hFDD7AD34 , 32'hFFF80675 , 32'hFF82F8C8 , 32'hFF6E6EEC , 32'hFFDA728A , 32'h0000E641 , 32'hFFFEF87A , 32'hFFFE2B19 , 32'hFFFE460D , 32'hFFFD8462 , 32'hFFFFB6F5 , 32'h0002018A , 32'hFFFE4EE3 , 32'hFFFEC225 , 32'h00007319} , 
{32'h136DCEA0 , 32'hE7EF2B80 , 32'hFEAEEF90 , 32'h06D68AA0 , 32'hDBED9340 , 32'hE85550E0 , 32'hF6F44DD0 , 32'h0927C360 , 32'h157450E0 , 32'hE8145C20 , 32'h04B43C50 , 32'hF8D3ACF8 , 32'h09940850 , 32'hF9585EB0 , 32'hF4B17DF0 , 32'h15818B80 , 32'h101075C0 , 32'hF6E15BD0 , 32'hFE051360 , 32'h08F49A20 , 32'h003B9654 , 32'hF30D7F40 , 32'h08EDF880 , 32'h0D960740 , 32'h082B0DB0 , 32'h021E96E8 , 32'hFD43CE1C , 32'hFD41A7A4 , 32'hF7C96F30 , 32'hEFFC6EC0 , 32'hF9457EC8 , 32'h0195A080 , 32'hF2C74C70 , 32'h0824AE90 , 32'hFFD2E209 , 32'h03741A8C , 32'hF1A315F0 , 32'hFF2DDCEB , 32'h07484780 , 32'hF4B2C110 , 32'hFF92206C , 32'h026BE5E8 , 32'h03453AF4 , 32'hF8A14CD8 , 32'h027C63B4 , 32'hFD83DFB0 , 32'hF252FB90 , 32'hEF1FC1E0 , 32'hF34810F0 , 32'h104206C0 , 32'hFD91DC18 , 32'hFD14970C , 32'hEB2EC460 , 32'h058DBBA0 , 32'hFD608894 , 32'h03E32628 , 32'hFDD1F574 , 32'h0462C988 , 32'h00941DEC , 32'h0166F848 , 32'hF434BE20 , 32'h065E9388 , 32'h025DED04 , 32'h03EE57BC , 32'h015CEEA0 , 32'h00E33428 , 32'h00BD3C22 , 32'h0546A290 , 32'h05BDCAF0 , 32'hF49BF700 , 32'h01543764 , 32'h019E3808 , 32'h00769307 , 32'hFE90AEC0 , 32'hFEFE23AC , 32'hFFC44407 , 32'hFF752BDA , 32'hFE93AF74 , 32'h009CE43C , 32'h04A56D30 , 32'hFE93F10C , 32'h0131CD8C , 32'h05CF7F70 , 32'hFD950B98 , 32'hFEEA4B18 , 32'h0240ED4C , 32'hFF9D590D , 32'h015CC76C , 32'h04D08760 , 32'h002743D6 , 32'h000469F7 , 32'hFFFE96C9 , 32'hFFFE79F1 , 32'h000020B7 , 32'h0000ACB9 , 32'hFFFFB68A , 32'hFFFF5F91 , 32'h0001DE39 , 32'h0000205E , 32'hFFFDF871} , 
{32'h02CD7D2C , 32'hFDA3D55C , 32'hE92F6520 , 32'h137B5280 , 32'h0B281560 , 32'hE0D4DDA0 , 32'hDF965B00 , 32'hEA21F440 , 32'hF15CCCA0 , 32'h04A77D00 , 32'h014481C4 , 32'h07D803B0 , 32'h08BAA570 , 32'h021316A4 , 32'hF2C86670 , 32'h1940C800 , 32'h0520E078 , 32'h09CC6F80 , 32'hFAF74C78 , 32'hF31AEA30 , 32'hF425AB20 , 32'hFD693D60 , 32'h14E81920 , 32'h10F3C360 , 32'h0150FDB4 , 32'h0CA64660 , 32'h06BD2FF0 , 32'hF9F15A50 , 32'hF1505430 , 32'hED534040 , 32'hFDE0313C , 32'h09E04040 , 32'h02CA2FC8 , 32'hFCD26D5C , 32'h00429EEC , 32'hFF7CF95D , 32'hEBB97D80 , 32'h063DF278 , 32'hFC668050 , 32'hF977A528 , 32'hFD8D88E8 , 32'h01BA5408 , 32'h0D224440 , 32'hEF6520C0 , 32'h080AE690 , 32'h02AA1430 , 32'hFF2D09B0 , 32'h0659DAE8 , 32'h00053FE6 , 32'hF4E09760 , 32'hFC6AF760 , 32'h0C75F440 , 32'h05C66D78 , 32'hFF159941 , 32'hED238BE0 , 32'hF31099B0 , 32'hFF76BDE1 , 32'hFC8E1184 , 32'hFC600C54 , 32'h000EDD5D , 32'hFDD85008 , 32'hFDA1BBE4 , 32'hFC8012D8 , 32'h03FF5894 , 32'hFDB6D84C , 32'h043EA9A8 , 32'hF4AE0560 , 32'hFE9537D0 , 32'hF81BF4C0 , 32'hFC53252C , 32'hFF61CD57 , 32'hFDE438A0 , 32'h00BDF72E , 32'h02FCE6E4 , 32'hFD2459EC , 32'h025EA77C , 32'hFF59D313 , 32'hFFB3B9FF , 32'h02B9AB7C , 32'hFDC58D50 , 32'h005BBEA6 , 32'hFDEAADE8 , 32'h032C3D50 , 32'h02A73CD8 , 32'h03FED49C , 32'h03E23820 , 32'hFF506B5F , 32'hFF7B2AB0 , 32'hFF573207 , 32'hFFA17A46 , 32'hFFFED544 , 32'hFFFE5BFE , 32'hFFFFB25E , 32'hFFFE5C54 , 32'h00011232 , 32'hFFFEC0CA , 32'h0000F92D , 32'h000132C3 , 32'h00000A79 , 32'h00001AF9} , 
{32'h0004C639 , 32'h0001B66D , 32'hFFFFEC33 , 32'h0000BE3A , 32'h0004479E , 32'h00000C17 , 32'h00010FB5 , 32'hFFFFD5D9 , 32'hFFFC6F74 , 32'hFFFDE03A , 32'hFFFC3FD9 , 32'h00034198 , 32'h000157DE , 32'h0002F2F1 , 32'h0001A63A , 32'hFFFE0165 , 32'hFFFBBDD1 , 32'hFFFDF530 , 32'hFFFB278A , 32'hFFFEF092 , 32'hFFFFC06D , 32'hFFFF8C9F , 32'hFFFD843E , 32'h0001C7D7 , 32'h00040542 , 32'h000206FC , 32'h0000BFFB , 32'h00013736 , 32'hFFFF3AF0 , 32'h0000F964 , 32'hFFFDF07F , 32'h00014197 , 32'hFFFD5EE7 , 32'hFFFF8C58 , 32'h0004A230 , 32'hFFFD00BD , 32'hFFFF0F66 , 32'h00054469 , 32'h0001549E , 32'hFFFE2C3B , 32'h0004DA0F , 32'hFFF8D683 , 32'h0000AA63 , 32'h0000F420 , 32'h0004BD04 , 32'hFFFD7DBA , 32'h00011D1A , 32'hFFFDC72A , 32'hFFFFAC01 , 32'hFFFCCCDD , 32'h0003DF8C , 32'h0001A88C , 32'hFFFE3C1B , 32'hFFFC0D2F , 32'hFFFC5F7B , 32'hFFFDE548 , 32'hFFFFF706 , 32'hFFFF0964 , 32'h0000E744 , 32'h000144FA , 32'h00024BCE , 32'h000159D5 , 32'h00020A4A , 32'h0000D891 , 32'hFFF964B0 , 32'h0004A5A1 , 32'hFFFF3B7A , 32'h0000BA18 , 32'h00062BAC , 32'h00012FEF , 32'h0004B0B3 , 32'h0000C40E , 32'hFFFE17D1 , 32'hFFFCE7BD , 32'h000210BA , 32'h0003A012 , 32'hFFFFEA89 , 32'hFFFE7FDD , 32'hFFFF88B1 , 32'hFFFD3FE8 , 32'h0001EDA0 , 32'h0003B8E8 , 32'h000163F8 , 32'hFFFF52B7 , 32'h0001051A , 32'hFFFE4821 , 32'h00023361 , 32'hFFFF0099 , 32'h00007275 , 32'h00024F0C , 32'hFFFF5A08 , 32'h0004F95A , 32'hFFFEAAE8 , 32'hFFFDFCFE , 32'hFFFC8DE1 , 32'hFFFC87A4 , 32'h00033AB1 , 32'h00001A00 , 32'h00024DD4 , 32'h000021C1} , 
{32'h0001D333 , 32'h000748CD , 32'hFFFEE684 , 32'h00013EA6 , 32'h0000835B , 32'h0001E450 , 32'hFFFE3F38 , 32'h00009513 , 32'h00023C87 , 32'hFFFD6A63 , 32'hFFFE67DC , 32'hFFFBEF7C , 32'hFFFBFD61 , 32'hFFFE87CD , 32'h00038CA4 , 32'h0001D6EC , 32'h00056540 , 32'h00021937 , 32'hFFFB1C7C , 32'h0004A755 , 32'h00015B20 , 32'hFFFEC40B , 32'h0000830D , 32'hFFFC7A28 , 32'hFFFDF15E , 32'hFFFDE1FA , 32'h0001D72D , 32'h0001AE42 , 32'h000276D9 , 32'hFFFF9A35 , 32'hFFFAD7BB , 32'h000317EC , 32'h00038F30 , 32'hFFFC7F19 , 32'hFFFFCDED , 32'hFFFC24DC , 32'h000418D0 , 32'h0002E234 , 32'h0000186B , 32'h00028E9C , 32'hFFFD7986 , 32'h000296C0 , 32'hFFFD56B4 , 32'hFFFEACB8 , 32'hFFFF05A4 , 32'h000621A1 , 32'h00010E8A , 32'hFFFDE0AC , 32'hFFFC34EC , 32'hFFFF9F71 , 32'h00013D3D , 32'hFFFF89D5 , 32'hFFFEEBB9 , 32'h0007ED8A , 32'h00032E17 , 32'h0002133E , 32'h000042F9 , 32'h0000E582 , 32'h00049193 , 32'hFFFDB353 , 32'hFFFCF31F , 32'hFFFEFCDF , 32'hFFFCA33E , 32'hFFFD7876 , 32'h0002CBDC , 32'hFFFD401E , 32'h0003A8DE , 32'hFFFEC1E6 , 32'hFFFE7C4C , 32'hFFFEB616 , 32'hFFFE147B , 32'hFFFEE456 , 32'h0001DF82 , 32'hFFFDA160 , 32'hFFFEC89B , 32'h0001ACCB , 32'h0003368B , 32'h000403E1 , 32'hFFFEBE6C , 32'h0001EA8D , 32'h0000714E , 32'h0000C843 , 32'h0001696B , 32'h0002310D , 32'hFFFF4795 , 32'h00035B89 , 32'hFFFE8EC9 , 32'h00049B9F , 32'hFFFF023C , 32'h00031C71 , 32'h00021DC7 , 32'hFFFC931E , 32'hFFFDFD34 , 32'hFFFBE9D1 , 32'hFFFD3FB5 , 32'hFFFEADC5 , 32'h0001318A , 32'h00006A6E , 32'h000247EE , 32'hFFFE6EBD} , 
{32'hFFFEB2F1 , 32'hFFFBBE24 , 32'hFFFE0EA9 , 32'h00010F00 , 32'hFFFEF3E9 , 32'hFFFDE467 , 32'h0001FC67 , 32'hFFFD0E11 , 32'h00021E80 , 32'hFFFCE1CC , 32'h0001133A , 32'hFFFBC595 , 32'hFFFEFC18 , 32'hFFFFB527 , 32'h0001CFDA , 32'h0005A64C , 32'h0004017F , 32'hFFFFB045 , 32'hFFFCE496 , 32'hFFFE31C4 , 32'hFFFF240A , 32'h00020CC3 , 32'hFFFDF106 , 32'h0001763E , 32'hFFFF388C , 32'hFFFF0DA8 , 32'hFFFD8EE8 , 32'h00009956 , 32'hFFFE7F5B , 32'h00035589 , 32'h00019EDF , 32'h0002C60F , 32'h00028981 , 32'hFFFF3164 , 32'hFFFC2681 , 32'hFFFD9C95 , 32'hFFFDDA71 , 32'hFFFF79D2 , 32'hFFFC0224 , 32'h000448E0 , 32'h000043DB , 32'h00007EDA , 32'h0001CCB7 , 32'h0000F72E , 32'h0000BA8A , 32'hFFFE7B28 , 32'hFFFEE932 , 32'hFFFE7256 , 32'h0001E100 , 32'h000019EE , 32'h0000BC18 , 32'h0001B0C6 , 32'h0006A858 , 32'h0000DAA1 , 32'h00037ACC , 32'hFFFD3266 , 32'hFFFE3E46 , 32'h0000B495 , 32'h00033341 , 32'hFFFEF493 , 32'h00028B1E , 32'h00024EC5 , 32'hFFFEBBDC , 32'hFFFFE3B1 , 32'h0001F5E5 , 32'h0001FD4C , 32'hFFFDDEAC , 32'hFFFFD042 , 32'hFFFDC856 , 32'hFFFFB6E3 , 32'hFFFD5E7A , 32'h0001B37C , 32'h0001CAD5 , 32'h0000A67C , 32'h000016E7 , 32'hFFFEB637 , 32'h00020463 , 32'h0000427B , 32'hFFFD8FD7 , 32'h000076CB , 32'hFFFFD54B , 32'h000133DC , 32'h00003BB9 , 32'hFFFE0E2B , 32'hFFFF6906 , 32'h0001B69E , 32'h00031256 , 32'h0000F143 , 32'h00027A5C , 32'hFFFFDC18 , 32'hFFFF2340 , 32'hFFFF4AF6 , 32'h0004920A , 32'h0001B33F , 32'hFFFF5531 , 32'hFFFF8F8E , 32'h0001A78C , 32'h0001B62A , 32'hFFFF8D3A , 32'hFFFFF930} , 
{32'hFFFCCC92 , 32'h0003BA3A , 32'h0000C113 , 32'hFFFDD6F5 , 32'hFFFEC262 , 32'hFFFCA988 , 32'hFFFED244 , 32'h00018522 , 32'hFFFE6481 , 32'hFFFF3298 , 32'hFFFD2161 , 32'h00024030 , 32'hFFFEBC46 , 32'hFFFD780F , 32'h00065803 , 32'h000009AC , 32'hFFFE4070 , 32'hFFFBBE97 , 32'hFFFEB43F , 32'h0003C143 , 32'hFFFB3461 , 32'hFFFEA199 , 32'h000044AF , 32'hFFFD4108 , 32'hFFFBDD3C , 32'hFFFD05B9 , 32'h0000F87D , 32'hFFFF99D0 , 32'hFFFB821B , 32'hFFFBF606 , 32'h00033920 , 32'h0001E33A , 32'hFFFE3361 , 32'hFFFF4549 , 32'h0000B8CF , 32'hFFFFCF35 , 32'h00010F81 , 32'hFFFCA635 , 32'hFFFDB23A , 32'hFFFDCF46 , 32'h000275F0 , 32'hFFFC3AF0 , 32'hFFFCD64E , 32'hFFFFB34A , 32'hFFFF37E3 , 32'hFFFEC09F , 32'h00013994 , 32'hFFFD72B5 , 32'hFFFE951B , 32'hFFFEB5EA , 32'h00042260 , 32'hFFFECE72 , 32'h00051F18 , 32'hFFFE434F , 32'hFFFF4714 , 32'hFFFBF363 , 32'h000212BD , 32'hFFFE0999 , 32'h00020B67 , 32'hFFFFC507 , 32'h0000DC85 , 32'h00066437 , 32'hFFFFC885 , 32'hFFFC1B1E , 32'hFFFBC49C , 32'hFFFFCA89 , 32'h0001492A , 32'h00057790 , 32'h000516A3 , 32'hFFFED4B4 , 32'h00002C50 , 32'hFFFE1753 , 32'hFFFF5AF9 , 32'hFFFE771F , 32'hFFFD2D1B , 32'hFFFD6621 , 32'h0002EDEF , 32'hFFFDDF76 , 32'hFFFF613E , 32'hFFFE117C , 32'h0000242B , 32'h00022DD9 , 32'hFFFBF4F5 , 32'hFFFCFA1F , 32'h00011551 , 32'h0003FFE6 , 32'hFFFE12FE , 32'hFFFF258B , 32'hFFFFD6FE , 32'hFFFBF141 , 32'hFFFD9CEA , 32'hFFFED1A8 , 32'h00054A31 , 32'hFFFE78E0 , 32'h00011B95 , 32'hFFFD9913 , 32'hFFFE2D2A , 32'h0006FB1F , 32'hFFFEBC1F , 32'hFFFEEEE0} , 
{32'hFFFF21BF , 32'hFFFF6C00 , 32'hFFFDF99E , 32'hFFFFD42B , 32'h00072F9E , 32'h0000942F , 32'h000135AB , 32'h000285EF , 32'h0000B281 , 32'h00035DF3 , 32'hFFFB6E4F , 32'h00038933 , 32'h0000D28F , 32'hFFFCB25F , 32'h00022CF0 , 32'h0002BCD4 , 32'hFFFC6D8F , 32'h000207F2 , 32'hFFFF046A , 32'hFFFD209C , 32'hFFFFE862 , 32'h00044462 , 32'h00010AC1 , 32'h0008900D , 32'hFFFE7ECE , 32'hFFF90E43 , 32'hFFFC294E , 32'hFFFD2425 , 32'hFFFD7119 , 32'h0004A842 , 32'hFFFFCD51 , 32'hFFF73B43 , 32'h00063ED7 , 32'h00022A08 , 32'h0002087C , 32'h000131F9 , 32'hFFFE99C5 , 32'hFFFDADC6 , 32'hFFFAE025 , 32'hFFFF58F2 , 32'h0000AFFF , 32'hFFFFE7E6 , 32'hFFFD2803 , 32'h0003D8D0 , 32'hFFFE1B88 , 32'h00018CAB , 32'hFFFE9A0D , 32'h00050DA6 , 32'hFFFDC18D , 32'hFFF7C63F , 32'h00039A4E , 32'hFFFA2754 , 32'h000242B2 , 32'hFFFDC6FE , 32'h0000FF35 , 32'hFFFCF346 , 32'hFFFFD879 , 32'hFFFA50A3 , 32'h00003E0A , 32'hFFFE94A8 , 32'hFFFE7B24 , 32'hFFFC23F6 , 32'h0000B66C , 32'h00004358 , 32'hFFFF2280 , 32'h00026016 , 32'h00008DE8 , 32'h0002B590 , 32'h00055308 , 32'hFFFEB0B1 , 32'hFFFF04A9 , 32'h00004845 , 32'h0001E892 , 32'hFFFAF9FE , 32'h000022BF , 32'h0001CADF , 32'hFFFFA84C , 32'h0004A1DC , 32'h00024BCA , 32'h0005892B , 32'hFFFE1504 , 32'h0003F52F , 32'h00020588 , 32'h0000FBF3 , 32'h0001CE55 , 32'hFFFBB8B7 , 32'h000085AD , 32'hFFFF4167 , 32'hFFFC952B , 32'h00000269 , 32'h0000D974 , 32'h00027F74 , 32'hFFFCC836 , 32'h0001BC2A , 32'hFFFF0603 , 32'hFFFCCBF9 , 32'hFFFD9A5F , 32'h0001465D , 32'h00044A88 , 32'hFFFE42B1} , 
{32'h05C2FF80 , 32'h0A208530 , 32'h04DB36F8 , 32'hF816B518 , 32'h03930360 , 32'h06C931B8 , 32'hF9EF0DF0 , 32'h06987630 , 32'h19903540 , 32'hF62837C0 , 32'hF895AD48 , 32'hFB8E1338 , 32'h0959E9D0 , 32'h05DD7678 , 32'hFD1E434C , 32'hF8434228 , 32'hFB53BC90 , 32'hF8495E38 , 32'h152BBA80 , 32'hFECC8670 , 32'h06170698 , 32'hFD1484E0 , 32'hE428A700 , 32'hFC2ED73C , 32'h160A5EC0 , 32'hF808FA40 , 32'hFCB1FFE0 , 32'h021E5C04 , 32'hF57EDB90 , 32'hFE96D974 , 32'hF4CCB470 , 32'hF11FE080 , 32'h039C34D0 , 32'hFCD60984 , 32'hFEAF0650 , 32'hFF4914D6 , 32'h0E322800 , 32'hF555F7D0 , 32'hF238B690 , 32'hFD17219C , 32'hF6F24590 , 32'hFCEEDCE8 , 32'hF4F05860 , 32'h05BC2380 , 32'h039C4DCC , 32'hFBFB3DF0 , 32'h168DBA60 , 32'hF4FFAFB0 , 32'h02BD0DEC , 32'hFFA314A1 , 32'h0E9D6030 , 32'hFB07FD40 , 32'hFF4DAA5B , 32'h0951BE90 , 32'h04174CE8 , 32'h01C6FFF0 , 32'hFDA57538 , 32'h034EA068 , 32'h07A044E0 , 32'h01444B0C , 32'h006DC979 , 32'h0653E888 , 32'hF9F645A8 , 32'h03355C78 , 32'h0115D884 , 32'h019648EC , 32'hFBC0ABC0 , 32'hFBDBFBD8 , 32'hFEB3C550 , 32'hF63ECE50 , 32'hFFBA8943 , 32'hF9D31D10 , 32'hFCE55504 , 32'h03FF2DB8 , 32'hFCA7C3A0 , 32'h00D5ABE6 , 32'hFE0C25D0 , 32'hFC563200 , 32'hF9A23750 , 32'hFED20DC8 , 32'hF9F04F18 , 32'hFE38FB14 , 32'h006029C9 , 32'hFE32ABBC , 32'hFEC128D0 , 32'h01DEC2E4 , 32'hFD57E648 , 32'h00EAAE86 , 32'hFAE5E0E0 , 32'hFF7B97C8 , 32'h0000A2EC , 32'h0000E344 , 32'h0000A53C , 32'hFFFE7926 , 32'h00012AB5 , 32'hFFFD7152 , 32'hFFFCF7F5 , 32'h00011177 , 32'h00002BEF , 32'hFFFEB0A3} , 
{32'h006123BD , 32'h2F4CCE00 , 32'hFC996AB0 , 32'hF7379A20 , 32'hF7027E00 , 32'hFE687784 , 32'hFF2C2165 , 32'h05E3B190 , 32'hF6769F80 , 32'hE997CD00 , 32'hF8F62798 , 32'h121BB780 , 32'hF2BA5C60 , 32'h08694F10 , 32'hF0EE7030 , 32'h11A5E040 , 32'h0C86E440 , 32'h039B541C , 32'h081BF840 , 32'h04575F98 , 32'hF432F630 , 32'h0A9C8C30 , 32'h04DF4D60 , 32'h02609704 , 32'hF3B04910 , 32'h0212BD28 , 32'h090337A0 , 32'hEB20DD20 , 32'h1674C460 , 32'hF928AFC8 , 32'h029B1A54 , 32'hFAADAB20 , 32'h0DC5F940 , 32'h074B2BB8 , 32'h02D0C580 , 32'hE4BFC6A0 , 32'h02AF02B8 , 32'h0FF61990 , 32'h0551A4B8 , 32'hF49AED40 , 32'hFDB46DA4 , 32'h0927ADC0 , 32'hFE1A746C , 32'h03F54D7C , 32'h0FFBEC10 , 32'h04522ED8 , 32'h057C9538 , 32'hF95B8078 , 32'h0074540D , 32'hFF8AAB87 , 32'h0E368690 , 32'hF434A140 , 32'h04BFCFF8 , 32'h0899A7A0 , 32'hF3118690 , 32'hFE810D80 , 32'hFC34750C , 32'hF77BE330 , 32'h098F1600 , 32'h028B32D4 , 32'h04A30B50 , 32'h03735470 , 32'h05572A40 , 32'hFBDF1288 , 32'hFEF06EF4 , 32'hFA9321E0 , 32'h09275CB0 , 32'hFF0E94A7 , 32'hFFB20C0D , 32'h001144C3 , 32'hF93BA920 , 32'hFEA41584 , 32'h030D0350 , 32'h05F08A18 , 32'hFF09A49C , 32'h06E34B10 , 32'hFFC01A5F , 32'hFD64EFF4 , 32'hFAE1E2C0 , 32'hFD49FC00 , 32'h04209168 , 32'h057EA740 , 32'hFCEB6330 , 32'hFFB619A4 , 32'hFD370914 , 32'h04C3B370 , 32'h01B0AD08 , 32'h00A2AFA0 , 32'hFC783F38 , 32'h000B6317 , 32'hFFFFD6D9 , 32'hFFFFF74C , 32'hFFFFB75F , 32'hFFFFAFC2 , 32'hFFFEFD6A , 32'h00007238 , 32'hFFFF8257 , 32'hFFFEB2C8 , 32'h0000395B , 32'h0000E384} , 
{32'h17D01680 , 32'hFD49F710 , 32'hFC2454D0 , 32'h11E43C40 , 32'hD5962A80 , 32'hF3069010 , 32'hD6EA1100 , 32'hEF852E40 , 32'h1349A840 , 32'hF23BDB00 , 32'hD21BD240 , 32'h0B5BB610 , 32'h26946580 , 32'hFC7AC9B0 , 32'h04C72CF0 , 32'h07C6E7B0 , 32'h06ACAA00 , 32'hFA0E0978 , 32'hF16A4C40 , 32'h1074D760 , 32'h1AB4D5E0 , 32'h0CD12300 , 32'h034C8724 , 32'hEB15F9C0 , 32'h095BD940 , 32'hF52FC320 , 32'h02A07170 , 32'hFF6D31B0 , 32'h008D695A , 32'hF94BF230 , 32'h0E3372C0 , 32'h03778DA8 , 32'h08423860 , 32'hFE3E5074 , 32'hF9562E90 , 32'hFECC0FC0 , 32'hF90EDF88 , 32'h05001168 , 32'h1652C660 , 32'h1744D4A0 , 32'hF77E1630 , 32'hFA3C3540 , 32'h0DED1BC0 , 32'hF7FF67C0 , 32'h02972E38 , 32'h0C5031D0 , 32'hF612A1C0 , 32'hF53F6C00 , 32'h02111E40 , 32'hFCB6F8A4 , 32'h02FFD268 , 32'h0738FF70 , 32'hFE87C9F8 , 32'hEFA1EFA0 , 32'hFFEAE89B , 32'hF9BBE750 , 32'h04F795C0 , 32'h065D8318 , 32'h0AE45530 , 32'h02293D40 , 32'hF8FE44A0 , 32'hFE9C8CE8 , 32'hF666C9C0 , 32'hFD19B284 , 32'hFEE4B644 , 32'hFBDFFCA0 , 32'h0301EFB8 , 32'h0181CBBC , 32'hFE1A02F0 , 32'hFCEF8134 , 32'hF8C22878 , 32'hF8E57DF0 , 32'h0233A38C , 32'h015D2268 , 32'hFDD58AAC , 32'h02C764C0 , 32'hFBF13050 , 32'hFBF5FF68 , 32'h049CE3F8 , 32'h06B3C3D8 , 32'hFB4A5650 , 32'h03190990 , 32'hFE09CBF0 , 32'hFD60B5AC , 32'h00F6BD1E , 32'hFCD83C54 , 32'h00CF9868 , 32'h0469D690 , 32'hFD296D88 , 32'h00F9B948 , 32'hFFFF1731 , 32'hFFFFE425 , 32'h000151A5 , 32'h00020E67 , 32'h00010DFC , 32'hFFFF146E , 32'hFFFE708A , 32'hFFFF2BF4 , 32'h00011A06 , 32'h00018BBB} , 
{32'h0002C800 , 32'hFFFFB276 , 32'hFFFED710 , 32'hFFFBB4AB , 32'hFFFF5322 , 32'hFFFDE81E , 32'h0003994D , 32'h0002B0DE , 32'hFFFFAE23 , 32'hFFFF43C8 , 32'h0003CCFD , 32'h000176B7 , 32'h00030CB7 , 32'h0005BF92 , 32'h0003B988 , 32'hFFFF5182 , 32'h0000F3C5 , 32'h00041869 , 32'hFFFF018F , 32'hFFFC572E , 32'h0004D93E , 32'hFFFD032D , 32'hFFFCE5D1 , 32'hFFFE3287 , 32'hFFFEB044 , 32'h00026F11 , 32'hFFFE25A0 , 32'h000142BE , 32'h0004C060 , 32'h0001FCF4 , 32'h0001989F , 32'hFFFD338B , 32'hFFFCFC13 , 32'hFFFBBBAA , 32'hFFFBFB84 , 32'h0002AF34 , 32'hFFFF05F3 , 32'h0001F1EA , 32'h00019AC0 , 32'h00006956 , 32'hFFFF06C1 , 32'h00037934 , 32'h0002D454 , 32'h000109BA , 32'h0000DDCC , 32'hFFFD74F4 , 32'hFFFDD412 , 32'h00001BC5 , 32'hFFFE60B3 , 32'h00030C69 , 32'hFFFF48A8 , 32'hFFFF9F49 , 32'h00013303 , 32'h00000267 , 32'h0004F07D , 32'h000088E5 , 32'hFFFF1C9E , 32'h00004EAD , 32'hFFFE4DE2 , 32'hFFFFA4D9 , 32'hFFFE17F1 , 32'hFFFDC655 , 32'h0003377D , 32'h00019DD5 , 32'hFFFEC532 , 32'hFFFD3592 , 32'h000125C0 , 32'hFFFFDFE8 , 32'hFFFC38B2 , 32'hFFFF4ED6 , 32'hFFFE3911 , 32'hFFFAEB51 , 32'hFFFE3ADD , 32'h00016867 , 32'hFFFED28C , 32'h00008587 , 32'hFFFCD609 , 32'hFFFD86A4 , 32'hFFFB06DC , 32'h00031D0A , 32'h0000B53F , 32'hFFFF0E5C , 32'h0001FD3F , 32'h0002C482 , 32'hFFFC50A0 , 32'hFFFDC26B , 32'hFFFCF73F , 32'h00000357 , 32'h000682F9 , 32'h000382D5 , 32'h0008EAED , 32'hFFF9C70C , 32'hFFFD3900 , 32'h0003B583 , 32'hFFFE0730 , 32'h00008ABA , 32'h00012D73 , 32'h00023925 , 32'hFFFC7035 , 32'hFFFF0371} , 
{32'hFFFE0271 , 32'hFFFD1D20 , 32'hFFFB4C2B , 32'hFFFDB8E0 , 32'h0001882E , 32'h00026D44 , 32'h0000DFB1 , 32'h000043E6 , 32'hFFFD6E9B , 32'h00004918 , 32'h0004DF34 , 32'hFFFD3553 , 32'h0000A798 , 32'hFFFE52EE , 32'hFFFE867C , 32'h00001128 , 32'hFFF6C7D7 , 32'h00043341 , 32'h00047044 , 32'h000168AE , 32'hFFFFFA45 , 32'h000348EE , 32'hFFFF9DD7 , 32'hFFFD1206 , 32'h000192F9 , 32'hFFFEFAD0 , 32'hFFFDEB49 , 32'h00029FCB , 32'h0004B925 , 32'h000179DE , 32'h00027B7C , 32'h00000830 , 32'hFFFFA1AE , 32'hFFFD9EC1 , 32'hFFFDF0B8 , 32'h00017B27 , 32'hFFFD9E9A , 32'h0003F47E , 32'hFFFA73F7 , 32'h000374EF , 32'h0003BAE2 , 32'hFFFD01ED , 32'hFFFF9B43 , 32'h0003F60C , 32'h000207CB , 32'h00039664 , 32'h0001127B , 32'h0002CE0C , 32'hFFFCCB61 , 32'h00014DF7 , 32'hFFFE6FD2 , 32'hFFFF066C , 32'h00009DA0 , 32'hFFFFD214 , 32'hFFFDF3E6 , 32'hFFFFA799 , 32'hFFFEC72D , 32'h00045172 , 32'hFFFBE12F , 32'h0002974D , 32'hFFFE215A , 32'h0000BD9A , 32'h0000EE12 , 32'hFFFF0183 , 32'hFFFD47E7 , 32'hFFFEC8A8 , 32'hFFFFDC90 , 32'h000347B9 , 32'h0003FDA1 , 32'h000044A9 , 32'h00051043 , 32'h0004ACE8 , 32'h00019F2E , 32'hFFFE0F2B , 32'hFFFD29AC , 32'hFFF88776 , 32'hFFFDA553 , 32'h00001BAE , 32'h000468F4 , 32'h0002B6E1 , 32'h0000610C , 32'h0003C30F , 32'hFFFF30A4 , 32'hFFFDEC51 , 32'h00021D2A , 32'h0001CA8C , 32'hFFFFCBE2 , 32'h000141B8 , 32'hFFFE5AF9 , 32'h0000E22F , 32'h0007ABE2 , 32'h00031BD1 , 32'hFFFE9BBD , 32'h00014033 , 32'hFFFD3CD6 , 32'h0002257F , 32'hFFFF0337 , 32'hFFFBB9F0 , 32'h00060C73 , 32'hFFFBB7A8} , 
{32'hFFFF3E94 , 32'h00014F1D , 32'hFFFF7AEA , 32'h00012A4B , 32'h000021C7 , 32'hFFFE2AE9 , 32'hFFFDC66B , 32'hFFFE17C3 , 32'h0000C2C6 , 32'hFFFE7A3C , 32'h000051CB , 32'hFFFEE159 , 32'hFFFD1243 , 32'hFFFD6154 , 32'hFFFF8C2F , 32'hFFFB65D5 , 32'h0000EAF8 , 32'hFFFD1756 , 32'h000088D9 , 32'h0005149A , 32'h0002044B , 32'h000233D4 , 32'hFFFF6223 , 32'h00006921 , 32'h00023DE2 , 32'h0001DD67 , 32'hFFFE3F3E , 32'h00011CCA , 32'h0003CFFC , 32'hFFFE6B85 , 32'hFFFF5CB8 , 32'hFFFD51BF , 32'hFFFF4CBB , 32'hFFFCD0D0 , 32'hFFFAF00F , 32'hFFFFBC08 , 32'hFFFD5A01 , 32'h00012B4E , 32'hFFFD5FBA , 32'h0003B7CE , 32'h00020A96 , 32'h000138FF , 32'h00006883 , 32'hFFFD3DDA , 32'hFFFF5005 , 32'hFFFCF724 , 32'h00066B5F , 32'h00011816 , 32'h00006133 , 32'hFFFDBAEB , 32'hFFFDFDA4 , 32'hFFFDECD3 , 32'h00010E77 , 32'hFFFCFD43 , 32'hFFFDFE6B , 32'hFFFE500D , 32'hFFFE2334 , 32'hFFFC7482 , 32'hFFFD20AD , 32'h0000A457 , 32'hFFFA75EA , 32'h00005F14 , 32'hFFFA72A4 , 32'hFFFC2A05 , 32'hFFFEC025 , 32'h0001D4E5 , 32'h00040086 , 32'hFFFF4792 , 32'hFFFE2CC7 , 32'hFFFFAC48 , 32'h00029DF0 , 32'hFFFEFADF , 32'hFFFC522B , 32'h0000AE86 , 32'hFFFC4D1E , 32'h0001C631 , 32'hFFFE39FC , 32'h00030706 , 32'h0002A0FF , 32'h00017400 , 32'h0002FADD , 32'hFFFDF171 , 32'hFFFE0045 , 32'h0001FF41 , 32'h00019441 , 32'h000154AA , 32'hFFFE6FB1 , 32'h0001A8A0 , 32'h00007F90 , 32'h000431C4 , 32'h00042F8D , 32'h000191B1 , 32'h00025CA6 , 32'h000200D1 , 32'h00020D5E , 32'hFFFC8F7B , 32'hFFFE935E , 32'hFFFD39C7 , 32'h0001DED6 , 32'h0000DC9F} , 
{32'h0004FE81 , 32'hFFFC34D4 , 32'hFFFE9006 , 32'h00013B0C , 32'hFFF8775A , 32'hFFFD9976 , 32'hFFFFF5DD , 32'hFFFED1C8 , 32'hFFFDB495 , 32'hFFFE10B4 , 32'hFFFFDB7A , 32'hFFFF694B , 32'hFFFCEEC5 , 32'hFFFCA5C8 , 32'h0000146B , 32'h0004702E , 32'h0001CB47 , 32'hFFFDC535 , 32'hFFFEF17A , 32'h00011A7D , 32'hFFFFD3CC , 32'h000354E4 , 32'hFFFE843F , 32'hFFFEB8F9 , 32'h00012338 , 32'h000265F8 , 32'h0000E3F3 , 32'h0003D204 , 32'hFFFE42A7 , 32'hFFFEB39D , 32'h00009769 , 32'h00037BB0 , 32'hFFFEE24D , 32'hFFFFEBCA , 32'hFFFFE460 , 32'hFFFF2EEC , 32'hFFFCCD5E , 32'hFFFEE834 , 32'hFFF94D5D , 32'h0004F1BA , 32'hFFFF9FA3 , 32'h0001EE3C , 32'h0004D038 , 32'h00022848 , 32'hFFFC124D , 32'hFFFEA519 , 32'h00037B51 , 32'hFFFD11C2 , 32'hFFFE4119 , 32'hFFFC3DA3 , 32'h0006DC83 , 32'h00065DA8 , 32'hFFFDA8A0 , 32'hFFFF5E4D , 32'hFFFA6057 , 32'hFFFF1B6B , 32'hFFFE3968 , 32'hFFFDF360 , 32'h00034D51 , 32'h00031728 , 32'hFFFB9197 , 32'hFFFE51DC , 32'h0002F2BA , 32'h00009700 , 32'hFFFE1EDB , 32'hFFFEB6E1 , 32'hFFFD3DA4 , 32'h000746C5 , 32'h0000014D , 32'hFFFDD4CD , 32'h00027BE1 , 32'hFFFDD75F , 32'hFFFBAC73 , 32'h0000FD0A , 32'h0000E6BA , 32'h00009DEA , 32'hFFFD8752 , 32'h000383FD , 32'h000021AC , 32'hFFFF1232 , 32'h000128F1 , 32'h0004416B , 32'h00028ABF , 32'h00006599 , 32'h00015F12 , 32'h000115EE , 32'hFFFEA74C , 32'hFFFDE844 , 32'hFFFAFBD4 , 32'h0000CABE , 32'h00017422 , 32'h0002EB1B , 32'hFFFB0074 , 32'hFFFEE9B5 , 32'h000547F9 , 32'h0003B959 , 32'h000350D7 , 32'hFFFCDAD9 , 32'h00033A47 , 32'hFFFF861E} , 
{32'hF3398A10 , 32'hFB4D15D8 , 32'hF23B34B0 , 32'h06BA73E8 , 32'h1488B980 , 32'h18AFD3A0 , 32'h0A152940 , 32'h01BCEF88 , 32'h042636B8 , 32'h064F1DA8 , 32'h09EC6920 , 32'h052A1640 , 32'hF075ED80 , 32'hF7CD5E10 , 32'h02182638 , 32'hFB800F50 , 32'hFF3F8252 , 32'h06DD6D38 , 32'h04BD0278 , 32'h11C03D40 , 32'hF1865400 , 32'h085AD5D0 , 32'h04000620 , 32'hF3402630 , 32'h0A9579F0 , 32'hEDEE5100 , 32'hF85A6BA8 , 32'h03D24FD8 , 32'hFDCB67DC , 32'hFB9390E8 , 32'h062C27B8 , 32'h073C06C8 , 32'hFC0E3FBC , 32'hFE97142C , 32'h047084B8 , 32'hF69A4230 , 32'h075695D0 , 32'h09293BF0 , 32'h00F85D0B , 32'h0D262C30 , 32'h05810410 , 32'hFE66AA74 , 32'h04BA7C88 , 32'h0DCBE270 , 32'hFE59B900 , 32'h05561418 , 32'h02EE5008 , 32'h00AD92A8 , 32'hFB6BD908 , 32'h00ACEA6D , 32'hF66980A0 , 32'hFFB5510C , 32'hFDFE422C , 32'h0013702B , 32'hF6FB8020 , 32'h0DA20C20 , 32'hFDB8EA5C , 32'h03FE4874 , 32'h04683878 , 32'h012DEAA0 , 32'h069FF280 , 32'hF80275B0 , 32'hFC8CE8E4 , 32'h0140D438 , 32'h0037DE84 , 32'h081AA2A0 , 32'h0144E480 , 32'hFFE0F30F , 32'hFEC10D9C , 32'h0072A9BE , 32'h013E1500 , 32'h084FE9F0 , 32'hFA8961E8 , 32'h05575208 , 32'h01B725D8 , 32'h0277C6D4 , 32'hFB58C0B8 , 32'hF9C4CE28 , 32'hFF1E72B4 , 32'h024C0C10 , 32'h0666D530 , 32'hF7364940 , 32'hFFCD068C , 32'hFC93E05C , 32'hFD18B930 , 32'hFF667200 , 32'h0262D374 , 32'h00F07BF3 , 32'hFE1202DC , 32'h00660699 , 32'h000096F6 , 32'hFFFD5C5D , 32'hFFFF16FB , 32'hFFFCA8F2 , 32'hFFFE5794 , 32'hFFFC63FF , 32'h0003A915 , 32'h00017424 , 32'hFFFDFCB5 , 32'hFFFEB9B7} , 
{32'hB8C71980 , 32'hC0925D00 , 32'hF7E340A0 , 32'hEECB9140 , 32'h0FDE7140 , 32'hE23D5020 , 32'h279A61C0 , 32'h14F3DF80 , 32'h1E09DEA0 , 32'hE62FAAA0 , 32'h154D5F00 , 32'hE69174E0 , 32'hE7773F00 , 32'hEE087440 , 32'h2E943B00 , 32'h03D94E4C , 32'h319AAA40 , 32'hFAF87EC8 , 32'hF4E2D1B0 , 32'h06A6DDB8 , 32'h01F83B54 , 32'h09D76B00 , 32'h13B457E0 , 32'hF4D1FF20 , 32'h0CDB9870 , 32'hF5C5F6B0 , 32'hE261E0C0 , 32'hF693B690 , 32'hFB30E118 , 32'hFC2F3C9C , 32'h001BBEA7 , 32'h009E0FA0 , 32'h1D2B10A0 , 32'hFE70E7C8 , 32'hE7A5C4E0 , 32'hFB2DE188 , 32'h0917E480 , 32'hFD7B2570 , 32'h0B9983A0 , 32'hF13D2B20 , 32'hF68027D0 , 32'h04934288 , 32'h045F6208 , 32'h0DC03900 , 32'h048E4CD0 , 32'h00EE9783 , 32'hF3423810 , 32'h0720A400 , 32'hF8926DD0 , 32'hF76C09C0 , 32'hFD737470 , 32'hFDD625F8 , 32'h066D1FB0 , 32'h038E11BC , 32'h02C6D2B8 , 32'h019E8800 , 32'hF9C7D068 , 32'h0AAD4020 , 32'h0281099C , 32'h03469E48 , 32'h05E0E138 , 32'h0733CF78 , 32'h01D712EC , 32'hFE06B0D0 , 32'hFBE31658 , 32'h0321E674 , 32'hFB4E44E0 , 32'h017BF930 , 32'hFABC08B8 , 32'hFD7D1D8C , 32'hFBFF64F8 , 32'h041A98A0 , 32'h02246CE0 , 32'h0561EBC8 , 32'h00C40A3D , 32'h03EBBF6C , 32'h032D5F80 , 32'h0019769F , 32'hFCE94BFC , 32'hFED465B4 , 32'hFDCBEF60 , 32'hFDFA355C , 32'hFFF57733 , 32'hFE53EDAC , 32'h03268B04 , 32'h02F6C610 , 32'hFDB88DD8 , 32'h0058E2D9 , 32'h021DF0F0 , 32'h0071F641 , 32'hFFFFC2F4 , 32'h0001347F , 32'h00024983 , 32'h00007E6B , 32'h00013E32 , 32'h00014998 , 32'hFFFE9BC4 , 32'h00009896 , 32'h000257D2 , 32'h00001E8C} , 
{32'h0001319E , 32'h000444FF , 32'h000002C2 , 32'h000035FE , 32'hFFFCF031 , 32'h0000A350 , 32'h0003DEC1 , 32'hFFFF3ADE , 32'h000241F0 , 32'hFFFB7931 , 32'h00002F96 , 32'h000238A9 , 32'h00044A10 , 32'h000123D9 , 32'hFFFF6C77 , 32'hFFFD8C6C , 32'h00049A2A , 32'h0002027C , 32'h00015C65 , 32'hFFFEC16F , 32'hFFFFC3F7 , 32'hFFFFCF05 , 32'h00018EBA , 32'hFFFE7E2C , 32'hFFFF6812 , 32'h0000E2C8 , 32'h0002C514 , 32'h00006741 , 32'hFFFFC8DC , 32'h0000D28D , 32'h0001F2D5 , 32'hFFFAB6F5 , 32'h0000B8B5 , 32'h0001662B , 32'hFFFF3E37 , 32'hFFFFDE07 , 32'h000162C2 , 32'h00006E94 , 32'hFFFE96CC , 32'hFFFCD580 , 32'hFFFFE2F9 , 32'h0000B3FE , 32'h00010FEB , 32'h00033386 , 32'h00002423 , 32'hFFFF8088 , 32'hFFFC7D95 , 32'h00006E6C , 32'h0004009E , 32'hFFFE0EC8 , 32'h000043D2 , 32'h0004498E , 32'hFFFFD4FA , 32'hFFFFBF0C , 32'hFFFB2186 , 32'hFFFDEA96 , 32'h00026724 , 32'h0003BDC1 , 32'h000205DB , 32'hFFFF0F45 , 32'hFFFBD247 , 32'h00004982 , 32'hFFFE94F2 , 32'h00018627 , 32'hFFFF7F44 , 32'hFFFE1427 , 32'hFFFF1457 , 32'hFFFD9935 , 32'h00055200 , 32'hFFFC3185 , 32'h0000A25D , 32'h0004F51B , 32'h000177E5 , 32'hFFFD3703 , 32'hFFFEBE98 , 32'h0000E41C , 32'hFFFE01B0 , 32'hFFFF4CE0 , 32'hFFFD8882 , 32'hFFFC1542 , 32'h0004ADDB , 32'hFFFD07E4 , 32'hFFFE69C2 , 32'hFFFEBD2E , 32'h0002FDE4 , 32'h000086E4 , 32'h00020D95 , 32'h000024FA , 32'h0003BCFC , 32'hFFFF0165 , 32'h0001A142 , 32'hFFFA977C , 32'hFFFB4CCD , 32'hFFFD4143 , 32'hFFFD9931 , 32'hFFFFB6D9 , 32'hFFFBBB18 , 32'h000172DD , 32'h0001BEC8 , 32'h0001AD25} , 
{32'h00055FC7 , 32'h0003419E , 32'h000159E4 , 32'hFFFE3B98 , 32'hFFFD509A , 32'h000298C0 , 32'hFFFAB7EC , 32'h00013C4A , 32'hFFFAD244 , 32'hFFFEEEF1 , 32'h000154D7 , 32'hFFFAA659 , 32'hFFFE8D4B , 32'hFFFD5717 , 32'h00020094 , 32'hFFFF9A03 , 32'hFFFD9BC4 , 32'hFFFF05B6 , 32'hFFFFB2F4 , 32'hFFFCDCD1 , 32'hFFFE766C , 32'h0001CFE5 , 32'h000074A6 , 32'hFFFEEFC4 , 32'h0001C869 , 32'hFFFEF9B6 , 32'h0001B7CF , 32'hFFFB1243 , 32'h0003B035 , 32'h0000FCC1 , 32'h00019A6A , 32'hFFFF5B75 , 32'h0001EFCE , 32'hFFFF7151 , 32'h0001EC4F , 32'hFFFFB0F4 , 32'hFFFDCA8D , 32'hFFFF6DED , 32'h00024E2A , 32'h00011CF0 , 32'hFFFDB474 , 32'h000283F3 , 32'hFFFF679F , 32'hFFFF43BA , 32'h0001DC8D , 32'h0001373C , 32'hFFFEE539 , 32'hFFFF8955 , 32'h0000D1C6 , 32'h000139E5 , 32'h0000F2CE , 32'hFFFD9EDB , 32'h00042B5E , 32'h0000C3C7 , 32'h0000370D , 32'hFFFEBE3E , 32'h00026C63 , 32'h00015465 , 32'h0001759D , 32'hFFFBBAE4 , 32'hFFFE631D , 32'hFFFC928E , 32'hFFFD272F , 32'h00016D31 , 32'hFFFE8BB7 , 32'hFFFC7193 , 32'hFFFFC493 , 32'hFFFD7AE6 , 32'hFFFCED80 , 32'h00054BF4 , 32'h0001A7D1 , 32'hFFFD23D7 , 32'hFFFF90F1 , 32'hFFFF6C3A , 32'hFFFD90DB , 32'h00004D43 , 32'h00037F60 , 32'h000271B2 , 32'h000069D2 , 32'h000252B1 , 32'hFFFE46F0 , 32'h0000F8B6 , 32'hFFFF3AAC , 32'hFFFD90DF , 32'h0001FD32 , 32'hFFFED56B , 32'hFFFFA2D2 , 32'h0004D7B2 , 32'hFFFD6A88 , 32'h00030396 , 32'hFFFEE775 , 32'hFFF89F52 , 32'h00007885 , 32'hFFFFE3F7 , 32'h0002688C , 32'hFFFCAB32 , 32'h000060B7 , 32'hFFFD1FAD , 32'hFFFFBAD9 , 32'hFFFFF6C3} , 
{32'h00001E30 , 32'hFFFBFFE9 , 32'hFFFD2266 , 32'hFFFF6E75 , 32'hFFFF1273 , 32'h0004E6B6 , 32'hFFFFF87B , 32'hFFFFDC70 , 32'h00047EB3 , 32'hFFFCDA01 , 32'h0002CF78 , 32'h0003B9D8 , 32'hFFFE05C4 , 32'h0001C5B3 , 32'hFFFD3805 , 32'h000034BE , 32'h00026519 , 32'h000195CC , 32'hFFFDDA95 , 32'hFFFDD5E6 , 32'h000195B1 , 32'h0000E802 , 32'h000151CF , 32'h0002C483 , 32'hFFFE5052 , 32'h00018F7B , 32'hFFFAB487 , 32'h00009D5B , 32'h0001CC1B , 32'hFFFE4194 , 32'h00003B92 , 32'h0000426A , 32'h0000D98E , 32'hFFFF0B6C , 32'h00021A2A , 32'hFFFFCD8A , 32'h00007689 , 32'hFFFD3CB9 , 32'hFFFD8E1E , 32'hFFFC5D15 , 32'h000311D6 , 32'hFFFCD99A , 32'hFFFBFD13 , 32'h00013563 , 32'h000868B4 , 32'h0000C531 , 32'hFFFF3EE7 , 32'hFFFDECA1 , 32'h00078008 , 32'hFFFDCA53 , 32'h00039BCE , 32'hFFFF370C , 32'h0001295B , 32'hFFF94232 , 32'hFFFDE092 , 32'h0001D8FA , 32'h00022C28 , 32'h0001C599 , 32'hFFFC1386 , 32'hFFFBB77D , 32'h00029AB4 , 32'hFFFE0175 , 32'hFFFE5AF4 , 32'hFFFE19FF , 32'hFFFEF761 , 32'hFFFD7BC7 , 32'hFFFEECB2 , 32'hFFFC258F , 32'h000152C4 , 32'hFFFE8482 , 32'h00029B12 , 32'h0000713F , 32'hFFFECB49 , 32'hFFFEC57A , 32'hFFFDF05C , 32'h0004E2BF , 32'h00039E0C , 32'h0005524A , 32'h0000A702 , 32'h00015175 , 32'hFFF9EAC2 , 32'hFFFF5551 , 32'hFFFD7ED4 , 32'hFFFE9298 , 32'hFFFAF54B , 32'h00003442 , 32'h00052543 , 32'hFFFE4E2C , 32'hFFFF9BDE , 32'hFFFF1FDA , 32'hFFFDBBB4 , 32'hFFFFEF00 , 32'hFFFE0729 , 32'hFFFF171D , 32'hFFFE6243 , 32'hFFFE5684 , 32'h00006ABB , 32'hFFFDA715 , 32'h0000108C , 32'h0001325D} , 
{32'h24DF0C00 , 32'hD3C73B00 , 32'h14ACE260 , 32'hC93D1600 , 32'hCBF0F780 , 32'hFF5B01A7 , 32'h29FF8DC0 , 32'hF415AE20 , 32'hD0F2A600 , 32'hFF76FBB3 , 32'h0DFB92C0 , 32'hF60ED030 , 32'hF6443790 , 32'h11C12E20 , 32'hFE8A9FBC , 32'hD81DCD80 , 32'h07B37078 , 32'h10C2E720 , 32'h046FB3D8 , 32'h0EE51C60 , 32'h0BFAC6F0 , 32'h09F53560 , 32'hF67A50B0 , 32'h0E59BD40 , 32'h1D4931E0 , 32'h0BB9E120 , 32'hFF054079 , 32'hF6A1A980 , 32'h080A8B00 , 32'hF88E3148 , 32'h0F711740 , 32'h048CAE98 , 32'hF706F6C0 , 32'hF83A4750 , 32'hF5E53D30 , 32'hF8CD0D80 , 32'h05E03E00 , 32'hFE1276D8 , 32'h0B0B3750 , 32'hFB594260 , 32'hF98BA3F8 , 32'h03AC4E54 , 32'hF81051A0 , 32'hF6D250C0 , 32'hFED73B5C , 32'h139955A0 , 32'hE8161A80 , 32'hFDC1AFD4 , 32'h063E77B8 , 32'h0372CDDC , 32'h0894EF70 , 32'hFCEECA64 , 32'hF6B851D0 , 32'h02F5A5CC , 32'hFE22FE78 , 32'h00C29F54 , 32'hFA04FBC0 , 32'h00D3C04E , 32'h0232CEC0 , 32'hF8761CD0 , 32'hFFB0F9D3 , 32'hFF02EC2E , 32'hF7A23EB0 , 32'h02FA9158 , 32'hF5D0F4B0 , 32'hF9FFBB30 , 32'h02B9AFEC , 32'h036667DC , 32'hFF973696 , 32'h05417B00 , 32'h01A68748 , 32'hF920CE38 , 32'h0133316C , 32'h03EA5460 , 32'h04FB0B18 , 32'hFB41D1D0 , 32'h02E6B264 , 32'hFD816D58 , 32'hFE82A6E0 , 32'hFF4B7FCD , 32'h047097B0 , 32'hFE73DC68 , 32'hFF836093 , 32'hFFAD6EB8 , 32'hFE3F9C70 , 32'h03557B48 , 32'hFDFFF784 , 32'hFE1A6D48 , 32'hFBE42818 , 32'hFFE8EFA4 , 32'hFFFD8BF4 , 32'hFFFFE9BE , 32'h000096E9 , 32'hFFFF533E , 32'hFFFEAE4B , 32'hFFFE7F64 , 32'h0001EB7E , 32'hFFFED360 , 32'hFFFE37C6 , 32'hFFFFC62E} , 
{32'h05748360 , 32'hD5328F00 , 32'h0B0AEC30 , 32'h0D489D50 , 32'hF2AFD890 , 32'h551A3700 , 32'hDD5369C0 , 32'h06B6BDB0 , 32'h251F9240 , 32'hDC9B7F80 , 32'h107DA780 , 32'h256C5380 , 32'h025F72C0 , 32'hED8AF5E0 , 32'h07105E98 , 32'h23AE0500 , 32'h04B4A748 , 32'h10969340 , 32'hEFE24520 , 32'hFF30F087 , 32'h0551F900 , 32'h1203A040 , 32'hF7A3F290 , 32'hF316F990 , 32'h105173A0 , 32'h0E3926A0 , 32'hF4855ED0 , 32'h0289CAD8 , 32'h0BD20D00 , 32'h00310DC3 , 32'h0234489C , 32'h0FA44040 , 32'h01FEDD34 , 32'hFC15367C , 32'h05623600 , 32'h0D588040 , 32'hF47251C0 , 32'h06D3F0B0 , 32'hF2A65DE0 , 32'hFF01DFCD , 32'h0CDD6390 , 32'h09201D50 , 32'h04EE19B0 , 32'h06538640 , 32'hFF94EE7E , 32'h01A57930 , 32'h083EE350 , 32'h030A6EB8 , 32'hFA46E5A8 , 32'hFD4DF72C , 32'h028F1A7C , 32'hFBF10990 , 32'hFFBDAF6C , 32'h05774468 , 32'h074DDC50 , 32'hFFA9B896 , 32'hEFC30FA0 , 32'h05609668 , 32'h000E26C4 , 32'hFF0B0C8C , 32'hFCF49188 , 32'hF527F5C0 , 32'h02410828 , 32'hFE2E723C , 32'h00797FB5 , 32'hF547E120 , 32'h020DE374 , 32'hFF2DB3AE , 32'h012E5EDC , 32'h04709220 , 32'hFFDB8877 , 32'hFD350E58 , 32'h01C41500 , 32'hFB8F1648 , 32'hFEA6B4A0 , 32'hFFD1284C , 32'h030EC61C , 32'h03E2AD34 , 32'hFEB2B734 , 32'h00560B81 , 32'h02DEE7B0 , 32'hFE852E40 , 32'hFF785088 , 32'h01405360 , 32'h0129E054 , 32'h04211F88 , 32'hFE35A9CC , 32'h026F85E4 , 32'hFFEA9369 , 32'hFF8CF43E , 32'h0003CD8E , 32'hFFFFF95B , 32'hFFFFD932 , 32'hFFFEBC1A , 32'h000062CA , 32'hFFFC585D , 32'h00016793 , 32'hFFFE1FA1 , 32'hFFFF641E , 32'h0000352D} , 
{32'hCB431680 , 32'hC7F5B7C0 , 32'h0906B360 , 32'h0C206510 , 32'hE1F3B980 , 32'hCA1A2780 , 32'hE53940A0 , 32'h087AD960 , 32'h0F6F68A0 , 32'h16228A60 , 32'h10242640 , 32'h15A66680 , 32'h12AA30A0 , 32'hF8535B58 , 32'hDD850F40 , 32'h08ABD600 , 32'h003A446B , 32'h04166C08 , 32'hECF8B4C0 , 32'h00E27334 , 32'h01A1F614 , 32'h0C44A1A0 , 32'h0BA3C820 , 32'h1040A780 , 32'hE9CD8040 , 32'hDF87F180 , 32'hFF7215F8 , 32'hFEEFC178 , 32'h1D6C5660 , 32'hFB6EFFA8 , 32'h070CA668 , 32'h00F6E3E4 , 32'h0D4693E0 , 32'hFBFC12A0 , 32'h0871BCA0 , 32'h044C3F20 , 32'hFFDCB097 , 32'hFA228F70 , 32'h04500BC0 , 32'h05A0C6B8 , 32'hF6DC02D0 , 32'hFB20DB68 , 32'hF847CC60 , 32'h093C49E0 , 32'h004166E6 , 32'hFABA7778 , 32'hF8A33F28 , 32'h014FB314 , 32'h0D5CDAE0 , 32'hFB9ECB98 , 32'hF6663D30 , 32'hF949A480 , 32'hF9B872F0 , 32'h04F14078 , 32'h0CA60210 , 32'h0371DC1C , 32'hFA0D29C8 , 32'hF38B6560 , 32'h064740F0 , 32'hFECDB27C , 32'h08278E10 , 32'h04ED2FB0 , 32'h014204A8 , 32'h05A0EC58 , 32'hF54A35F0 , 32'h07F33080 , 32'h0090DAB5 , 32'h08E152C0 , 32'hFADE9628 , 32'h04320180 , 32'hFE22DD48 , 32'hFD029DCC , 32'hFF1C1789 , 32'hFDBF6094 , 32'hF9A32478 , 32'hFEE5D944 , 32'h03211B44 , 32'h04D9DD90 , 32'h029BB31C , 32'h0049E35D , 32'hFC6AFA5C , 32'hFED9826C , 32'h016E4F84 , 32'hFFD6732D , 32'h01639E48 , 32'hFE63C380 , 32'h01FB10A0 , 32'h0138EEB8 , 32'hFEC274D4 , 32'hFCB87390 , 32'h00017DBA , 32'hFFFF4BB2 , 32'hFFFEE56E , 32'hFFFFF174 , 32'h00018352 , 32'h00004F26 , 32'h0000216E , 32'h0000F4BC , 32'hFFFF6A65 , 32'hFFFF3FE2} , 
{32'hFFFC102B , 32'hFFFF5FCE , 32'hFFFEEB22 , 32'h00019287 , 32'h00017AC9 , 32'h0000A04D , 32'hFFFE0EA8 , 32'hFFFF7DBD , 32'hFFFCA2E6 , 32'hFFFF4A9B , 32'hFFFFE887 , 32'h0000017A , 32'hFFFF10EF , 32'hFFFEE319 , 32'hFFFD556A , 32'h0000FD71 , 32'hFFFD3E17 , 32'hFFFEBE40 , 32'h0002DE12 , 32'h00010746 , 32'h0001447E , 32'h00066C15 , 32'hFFFCEA72 , 32'h000442E0 , 32'hFFFE0F57 , 32'hFFFDFB81 , 32'h000086E3 , 32'hFFFF23E8 , 32'h0008942C , 32'hFFFEF063 , 32'hFFFF31F9 , 32'hFFFC915C , 32'h00016A10 , 32'h0002B9E2 , 32'hFFFDD743 , 32'hFFFD4342 , 32'hFFFEEFF9 , 32'hFFFF0984 , 32'h00007C0A , 32'hFFFE53B5 , 32'h00025A2D , 32'h00003CA5 , 32'h00029D4F , 32'h00014A44 , 32'hFFFDB4F8 , 32'h0002F95A , 32'hFFFEA9E7 , 32'h0003687A , 32'h00069D44 , 32'h0001F877 , 32'hFFFF2B8F , 32'h00025175 , 32'hFFFF7537 , 32'h0000E752 , 32'h00023C54 , 32'h00031DDD , 32'h0000C157 , 32'h00014843 , 32'hFFFF32B0 , 32'h0001890F , 32'hFFFE563D , 32'h0000BDD2 , 32'h00002BF6 , 32'h0005AA49 , 32'h0002A7E9 , 32'h0002411B , 32'hFFFEFCB5 , 32'hFFFAE08F , 32'h00004CFB , 32'h0000F113 , 32'h0005728C , 32'h00002E12 , 32'hFFFEA6EC , 32'h0001CC2A , 32'hFFFBBAF1 , 32'hFFFFEF33 , 32'hFFFFC57B , 32'hFFFC20BE , 32'hFFFE751A , 32'hFFFF2F76 , 32'hFFFE9375 , 32'hFFFBA79F , 32'hFFFDD9E0 , 32'hFFFE4C00 , 32'h0001CA34 , 32'h00023368 , 32'h000134DC , 32'hFFFCC4A1 , 32'hFFFD6577 , 32'h00025292 , 32'hFFFEE252 , 32'hFFFA0AA7 , 32'h0000FDAB , 32'h000280A6 , 32'hFFFD6BBF , 32'h00080CF3 , 32'hFFFF2EAE , 32'hFFFEDA6C , 32'hFFFFCC6F , 32'h00016CC6} , 
{32'h0001CB22 , 32'h0001B08C , 32'hFFFCD076 , 32'hFFFF71F2 , 32'hFFFD80CE , 32'h00020A55 , 32'hFFFB0848 , 32'hFFFCE193 , 32'hFFFE8400 , 32'h0000A0E9 , 32'hFFF769E2 , 32'h000211CE , 32'h0000E35C , 32'h0000A769 , 32'hFFFB61B8 , 32'h0004EED6 , 32'h00011F81 , 32'hFFFD02B8 , 32'hFFFC2EDD , 32'hFFFF27C5 , 32'h0004184E , 32'h0000EC07 , 32'h00006735 , 32'h0003827A , 32'h0006EFED , 32'h0002D4CC , 32'h000060EA , 32'hFFFE507D , 32'h00042EAE , 32'hFFFD7F58 , 32'h00024BFD , 32'h0000570A , 32'h0005397C , 32'h0003BFB6 , 32'h0000868A , 32'h00032A98 , 32'hFFFA9CFC , 32'h0004B24C , 32'h00008709 , 32'hFFFD302F , 32'h00008365 , 32'hFFFEAD20 , 32'h0004E706 , 32'h0000A98C , 32'h000070EF , 32'h0004444E , 32'h00062500 , 32'h0006B97B , 32'hFFFBD546 , 32'h000134A9 , 32'h00001050 , 32'h0000EF00 , 32'hFFFD9F56 , 32'h0003F136 , 32'hFFFFE37A , 32'hFFFFB66E , 32'h0000F259 , 32'h0003BA24 , 32'h0004F86B , 32'hFFFD3DC0 , 32'hFFFC6A1F , 32'h0000E71D , 32'hFFFE2CB3 , 32'hFFFC0442 , 32'hFFFEB102 , 32'hFFFE2B88 , 32'hFFFB82C4 , 32'hFFFDB89C , 32'hFFFF5BCA , 32'h00001103 , 32'hFFFE0644 , 32'h000172C8 , 32'h00057A61 , 32'h00039F1F , 32'hFFFD2A0D , 32'hFFFC8282 , 32'h00028AB4 , 32'h000470FF , 32'h00023421 , 32'hFFFE7750 , 32'hFFFE8015 , 32'h00045667 , 32'h0000AB95 , 32'h00011492 , 32'hFFFC825D , 32'h00020C4D , 32'hFFFBC95A , 32'hFFFF757D , 32'h000680FA , 32'hFFFCECD1 , 32'hFFF8161A , 32'hFFFCC50F , 32'h0005B1D1 , 32'h00032351 , 32'hFFFEAA95 , 32'hFFFD1626 , 32'h000188FE , 32'h00014130 , 32'hFFFDBAB3 , 32'hFFFD4B1F} , 
{32'h0003DC22 , 32'hFFFEBCD7 , 32'hFFFEEA4C , 32'h0003119E , 32'h000199D2 , 32'hFFFFCC52 , 32'h00028266 , 32'hFFFE0CDF , 32'h0001D832 , 32'hFFFB44A5 , 32'h00013247 , 32'hFFFE0E6E , 32'h000209C1 , 32'h00016F1F , 32'h0000B669 , 32'hFFFD4C9A , 32'h00051AFF , 32'h00049E82 , 32'hFFFDDAFF , 32'hFFFF7B2A , 32'h0001EC97 , 32'hFFFD7ACD , 32'h00038329 , 32'hFFFEA148 , 32'hFFFFFCB2 , 32'hFFFF3ECC , 32'h00036B5F , 32'hFFFB457A , 32'hFFFEECF4 , 32'hFFFF75E6 , 32'h000408E7 , 32'hFFFFCB1D , 32'h000066E1 , 32'h0001204C , 32'h0003B56D , 32'hFFFED822 , 32'hFFFEDC48 , 32'h00003075 , 32'h000019B8 , 32'h00021711 , 32'h0001D727 , 32'h0001380E , 32'hFFFC1BBB , 32'hFFFFFE25 , 32'h0004D57C , 32'hFFFE15D1 , 32'hFFFEDC74 , 32'h000325E8 , 32'h000184BF , 32'hFFFC8F26 , 32'hFFFEDAA4 , 32'h00034B7E , 32'hFFFE7C57 , 32'hFFFE44BE , 32'h000041A4 , 32'h00007508 , 32'h00002572 , 32'hFFFEDB98 , 32'h00048CC0 , 32'hFFFD458F , 32'hFFFFE27D , 32'h0000313F , 32'h00022A02 , 32'h0002F54C , 32'h000109B6 , 32'h0003D407 , 32'hFFFF00DA , 32'h00004377 , 32'h00014EEC , 32'h0000F969 , 32'h00009ABD , 32'h0007A01D , 32'hFFFF389A , 32'h00040F1C , 32'h00010012 , 32'h000774D8 , 32'h00003A9C , 32'h00022207 , 32'h000206C9 , 32'hFFFB1F88 , 32'h0000DFA0 , 32'h000203D3 , 32'h0002DF0A , 32'hFFFDA1E9 , 32'hFFFF45AE , 32'hFFFC8AC2 , 32'hFFFF9B3F , 32'h00006568 , 32'hFFFFCE08 , 32'h0000AEA4 , 32'h0004E947 , 32'hFFFEB446 , 32'hFFFE1A37 , 32'hFFFF1ACC , 32'h00036109 , 32'hFFFC59F1 , 32'hFFFE6CFC , 32'hFFFECD44 , 32'hFFFA7A38 , 32'h0001A9CF} , 
{32'h05F2D2C0 , 32'hF7F18EF0 , 32'h08C40BC0 , 32'hEF2F7D00 , 32'h00FBAEB9 , 32'hF0DBBD80 , 32'h0B4DFD90 , 32'hF38C8DE0 , 32'hFD95D034 , 32'hFED63A60 , 32'h09C8C7D0 , 32'h008E95F4 , 32'h05E24880 , 32'hFA3C38C0 , 32'hF1B30150 , 32'hF075DCD0 , 32'h0ECF3C80 , 32'hFEED7CAC , 32'hFC1E1D64 , 32'h0F180440 , 32'h0F2E39D0 , 32'hF75CC470 , 32'h06314C78 , 32'h0584E690 , 32'h09E63130 , 32'hF946DFE8 , 32'hFC754944 , 32'hFDA2EF10 , 32'hFDDAA860 , 32'hFF86A5C3 , 32'hFA25B950 , 32'hF7495F50 , 32'hFF3047F0 , 32'h03094324 , 32'h044A6630 , 32'h013FE294 , 32'hFB2652A0 , 32'h05B7E6F8 , 32'h0280A51C , 32'hF88AEBE0 , 32'h0B3D13C0 , 32'h05BC2778 , 32'hFBC14288 , 32'hF6204F00 , 32'h09DCFE60 , 32'h08F0A8C0 , 32'h0B44BDD0 , 32'hF8D6E5A0 , 32'hF92A9CB0 , 32'h01EC2F18 , 32'hFDD49170 , 32'h027666C4 , 32'h086DD140 , 32'h02486A20 , 32'hFB3CA670 , 32'h024802B8 , 32'h09D932F0 , 32'hF86197E8 , 32'hFDB2E854 , 32'hFBEB8F58 , 32'h035ED828 , 32'h0499E9B0 , 32'h067BF378 , 32'hFC0901C0 , 32'h00D89852 , 32'h013C0B8C , 32'hFE9E7A18 , 32'h04E89AC0 , 32'hFF68C27B , 32'h0A935400 , 32'hFFBC8F6C , 32'h08EBCC30 , 32'hFB40BC70 , 32'h01427EFC , 32'hFE541170 , 32'hFD8D1E38 , 32'h05C86008 , 32'hFB9418E8 , 32'hFD07206C , 32'hFE9EA250 , 32'hF8E4EB08 , 32'h03E09C78 , 32'hFFC2968F , 32'hFEC78470 , 32'h00D72A15 , 32'h0080D532 , 32'h0231B484 , 32'h00055674 , 32'hFF44D6CA , 32'h005BEE0A , 32'hFFFFB4C5 , 32'h00039864 , 32'h0000EC65 , 32'hFFF9B8AE , 32'h00019589 , 32'hFFFF8AB2 , 32'h00007A59 , 32'h000078DF , 32'hFFFF1776 , 32'hFFFE7159} , 
{32'h03B1B1AC , 32'h039554F4 , 32'h0DA2D290 , 32'hFBD638D8 , 32'h083E1110 , 32'h0F8D0790 , 32'hFD4B2ACC , 32'hF434C750 , 32'hFE399EC8 , 32'hF5A27140 , 32'hF9518A40 , 32'hF8DDF270 , 32'hF6EF4010 , 32'hF68C0F70 , 32'h09A83990 , 32'h0A3DF7F0 , 32'hF1AB4260 , 32'hF5EB8120 , 32'hFD55058C , 32'h05F4B168 , 32'hF83D6C78 , 32'hF73D5F10 , 32'hFBC52000 , 32'hF8C3CF78 , 32'hFF6FFA1C , 32'h0261B38C , 32'h01CE4B68 , 32'h098A60E0 , 32'hFCC3FBC8 , 32'hFFAD76A6 , 32'hFD87CA30 , 32'hF4F40BA0 , 32'h0A8897C0 , 32'hF65A1E80 , 32'h004F0A08 , 32'hF21A1120 , 32'hFE1B4AFC , 32'hF5248670 , 32'h00FFEEB4 , 32'hFA649F18 , 32'hF85AC5C0 , 32'h022DF470 , 32'h09A2E080 , 32'hF2F78BA0 , 32'hF9FCC3B0 , 32'h012F4710 , 32'hFDAFD88C , 32'h096C15D0 , 32'hFBE874B8 , 32'hFE05FD98 , 32'h01449E80 , 32'hFDD1303C , 32'hFFEE05D2 , 32'h0328470C , 32'h0737B5F8 , 32'h0191F5B4 , 32'hFABD16F8 , 32'hF7E1E570 , 32'hFC80353C , 32'hFECC8C84 , 32'hFC753148 , 32'hF83362D0 , 32'h03FB7654 , 32'h002CD96C , 32'h01BD5BF4 , 32'hFE4E13F0 , 32'hFFECF246 , 32'h03696068 , 32'hFCAAEE1C , 32'hF5BC1D40 , 32'h069DCB78 , 32'h08819FD0 , 32'hFAED61A8 , 32'h0028DACA , 32'hFE086DF0 , 32'h00B21062 , 32'h039D3B20 , 32'h00506F5F , 32'h05D928F0 , 32'h01B2BFA8 , 32'hFE1EA8DC , 32'hFE11AE58 , 32'h01EBF398 , 32'hFC790474 , 32'hFCB23120 , 32'hFD578BA8 , 32'hFDEE0274 , 32'hFD680414 , 32'hFFC9BDEF , 32'hFFCAAB77 , 32'hFFFE08BB , 32'h000204A7 , 32'hFFFECBAD , 32'h000097B9 , 32'h0000EEFF , 32'hFFFD0287 , 32'hFFFEDD98 , 32'hFFFF5ABE , 32'hFFFE2DE2 , 32'h00010A34} , 
{32'h34BB59C0 , 32'hE0F5B580 , 32'hDF0CF640 , 32'h1831FD20 , 32'hE20AC0E0 , 32'hBA761A00 , 32'h1B7ABD00 , 32'hDDD38780 , 32'hFF41EE0C , 32'h35E6E0C0 , 32'hF1865E30 , 32'h01F2FDA8 , 32'hE9EEAF60 , 32'h144F74A0 , 32'h215FC900 , 32'h14E5E560 , 32'h12819D40 , 32'hFF22CE7C , 32'h0794BF60 , 32'h00D8EAF1 , 32'h12E4FBA0 , 32'hE6C22E40 , 32'hF77D1900 , 32'hFADE4470 , 32'h007AA526 , 32'h0683F2F0 , 32'hF878CC10 , 32'h067C2BB0 , 32'h03048FB4 , 32'hFA602F58 , 32'h024DF890 , 32'hF0E2DAB0 , 32'hFB7D7108 , 32'h0C8C8FB0 , 32'hFAEF6C78 , 32'hFE2D7E88 , 32'hFEA78B68 , 32'h09DDB040 , 32'h0602E848 , 32'h07052D08 , 32'h0AF73290 , 32'h01D05C8C , 32'h036B21B8 , 32'h072D6EC0 , 32'h08A5DB60 , 32'hDEF84A80 , 32'h040F2338 , 32'h08E4A140 , 32'h07991DA0 , 32'hFCCB5C08 , 32'hFE2F3CCC , 32'hFB9D4420 , 32'h0BC41AB0 , 32'hFA7CB2C0 , 32'h00C240F9 , 32'h004893C4 , 32'h0014EB7F , 32'h021E5D20 , 32'h00AFFED9 , 32'hFC2E7FC0 , 32'h02A29D58 , 32'hFDFF3F88 , 32'h0586F290 , 32'hFE6F3B30 , 32'h006B0DC0 , 32'hFAE7A798 , 32'h04FF7B28 , 32'h02621464 , 32'h02359A9C , 32'hFBF8FE98 , 32'h07B8E940 , 32'hFDB7C608 , 32'h03F5499C , 32'hFD2B5330 , 32'hFE1BF120 , 32'h02253CD0 , 32'h0414A838 , 32'h0153CF98 , 32'h02555268 , 32'h02B87E34 , 32'h005DC0D8 , 32'h03C2B2FC , 32'hFE75F2E4 , 32'h0296EDDC , 32'hFD84405C , 32'h01774524 , 32'hFC13DD24 , 32'hFCF21DCC , 32'hFF1EDA11 , 32'hFF4F4A5B , 32'h00001907 , 32'hFFFF6FA9 , 32'hFFFFAE2D , 32'h00012811 , 32'hFFFEF8EA , 32'h00008009 , 32'h00015D6B , 32'hFFFE14AD , 32'hFFFE9405 , 32'h00002B88} , 
{32'h00016B79 , 32'hFFFD78AC , 32'hFFFE81BF , 32'hFFFE6DE2 , 32'hFFFD9CCD , 32'h0001C620 , 32'h00009D9A , 32'hFFFE59F7 , 32'h0002243A , 32'h0001BF80 , 32'h0003B64C , 32'hFFFFF941 , 32'h000447B5 , 32'h0000F4A6 , 32'hFFFF9EEC , 32'h0000FDCE , 32'h00014B7D , 32'hFFFA5A96 , 32'hFFFDEE5F , 32'hFFFF41EC , 32'h00036601 , 32'hFFFF7424 , 32'hFFFD369F , 32'hFFFCCA0B , 32'hFFFF4E67 , 32'hFFFE7E24 , 32'hFFFF3583 , 32'hFFFFC7A8 , 32'h00016F07 , 32'h00053499 , 32'h0002AD00 , 32'hFFFD12D8 , 32'h0000D048 , 32'hFFFEB564 , 32'h00003E7C , 32'hFFF8DCA6 , 32'h00023790 , 32'h00019BB8 , 32'hFFFECD9A , 32'hFFFEE140 , 32'h0001FE2F , 32'h0002C066 , 32'hFFFD218B , 32'hFFFECF21 , 32'h0004D18C , 32'h00006B62 , 32'h00005707 , 32'h0002C1D1 , 32'hFFFF7C8D , 32'h0000DC00 , 32'h00000147 , 32'h0000E917 , 32'h0001519B , 32'hFFFC6B59 , 32'hFFFF2923 , 32'hFFFF72EB , 32'hFFFF8AD2 , 32'hFFFB6BAD , 32'hFFFCBF80 , 32'hFFFEECDE , 32'h00003684 , 32'h0000F87B , 32'hFFFFA5B1 , 32'h00064813 , 32'hFFFF1E8E , 32'hFFFE5DD3 , 32'hFFFA61F8 , 32'hFFFF5EFF , 32'hFFFFDE8B , 32'hFFFFEC12 , 32'h0000D78F , 32'h0000B789 , 32'hFFFB3506 , 32'hFFFE5B1F , 32'hFFFAA7C7 , 32'h0001F785 , 32'hFFFE7319 , 32'h0001681D , 32'hFFFEA9E3 , 32'h000331FB , 32'hFFFDD926 , 32'hFFFF20F6 , 32'h0005AD13 , 32'hFFFAF5F2 , 32'h0002A678 , 32'hFFFE0AA1 , 32'hFFFC37A4 , 32'h000395C0 , 32'h0001CA71 , 32'h0001DDD1 , 32'h0002FADB , 32'hFFFD9976 , 32'hFFF9A2EA , 32'hFFFBAD4F , 32'h0003B3A3 , 32'hFFFBACA1 , 32'hFFFF5F72 , 32'h00000AF1 , 32'h00040C33 , 32'h00005205} , 
{32'h0086E77A , 32'h03712610 , 32'hFC853A38 , 32'hFC5065E4 , 32'hFD833DAC , 32'h0131F498 , 32'hF9638A28 , 32'h001C60A7 , 32'h00E83B67 , 32'hFD0D0A84 , 32'h00F3A57C , 32'hFF34C4D9 , 32'h00E6D036 , 32'h0194A864 , 32'h02498E6C , 32'h040FDE48 , 32'hFD8E82F4 , 32'hFECA0EE0 , 32'hFF894686 , 32'hFE985348 , 32'hFA4F6930 , 32'hFE6F0724 , 32'hFAD19610 , 32'hFA7D1820 , 32'hFFEB3731 , 32'h02697C64 , 32'hFD0636A0 , 32'h0461B880 , 32'hFCAE5EEC , 32'h00FB6107 , 32'h02D24E50 , 32'hFF293FBE , 32'hFCA5DE58 , 32'hFDCBA2D0 , 32'h01A34AF0 , 32'hFFFBDEBD , 32'hFE2DCFF8 , 32'hFEBF3AB4 , 32'h0039A19B , 32'hFB173908 , 32'hFFE5C199 , 32'h02456258 , 32'hFF5C2AC4 , 32'h02D44E68 , 32'hFF155D23 , 32'hFD3B6E44 , 32'h00B9982D , 32'h015DD55C , 32'hFC4D68EC , 32'hFBAAAD10 , 32'hFDABE834 , 32'h020AAF40 , 32'h0080A86B , 32'hFF156ED9 , 32'hFFD11FB4 , 32'h00A81AD5 , 32'hFEF5B0C4 , 32'hFE00517C , 32'h0245F028 , 32'hFE8A227C , 32'h01A2F0DC , 32'hFF77450D , 32'hFF1B25F4 , 32'h00046526 , 32'h013FFAA0 , 32'h02DF2720 , 32'hFE2FAAF8 , 32'hFDF31284 , 32'h000FC5A4 , 32'hFF99DE89 , 32'h005E3524 , 32'h015E8534 , 32'h00AE0963 , 32'h028BFEB4 , 32'hFE91C5B8 , 32'hFEBF1550 , 32'hFF3F10A1 , 32'h0213E120 , 32'hFE2B1D7C , 32'hFE51DAE0 , 32'hFF778942 , 32'h00211FF5 , 32'hFE940ED4 , 32'hFF943D5A , 32'h0059D4A0 , 32'hFFD67492 , 32'hFDEB7D54 , 32'h03AC64D4 , 32'h00B3A4C9 , 32'hFFF1DEE1 , 32'hFFFECC05 , 32'h00046314 , 32'hFFF9F1FE , 32'h0001A4DA , 32'hFFFBEE36 , 32'h000240B1 , 32'h00071B3E , 32'hFFFE2D70 , 32'hFFFF803A , 32'h00005A1C} , 
{32'hFFFCDE7C , 32'hFFFAE1AA , 32'hFFFF324B , 32'hFFFB0E63 , 32'h00021984 , 32'hFFF9FE2A , 32'hFFFD468A , 32'hFFFCD3C9 , 32'h0005C93A , 32'h0001023B , 32'h000118FA , 32'h0002D615 , 32'hFFFCF3D0 , 32'h000065FE , 32'h0009456F , 32'h0004D4E5 , 32'hFFFCDB0E , 32'h00038CDD , 32'h0000B79D , 32'h00039733 , 32'hFFF86632 , 32'hFFF7BF4B , 32'hFFFDA8C8 , 32'h0004F659 , 32'hFFFB378C , 32'hFFFD1768 , 32'h00028AB8 , 32'hFFFF3F5A , 32'h00030DBF , 32'h000164F0 , 32'hFFFB8124 , 32'hFFFECCAA , 32'h000325A8 , 32'h00027250 , 32'h0001ABC3 , 32'h00007243 , 32'hFFFDB004 , 32'hFFFB1817 , 32'h000074F1 , 32'hFFFFA417 , 32'hFFFD0D48 , 32'h00024C9C , 32'hFFFCC823 , 32'hFFFD99AE , 32'h00046F39 , 32'hFFF83D75 , 32'h00007BC9 , 32'h000126AF , 32'hFFFEDE64 , 32'h0002448A , 32'h000397D4 , 32'hFFFFCD77 , 32'hFFFEC700 , 32'hFFF8B198 , 32'hFFFD7D34 , 32'h00024237 , 32'h00014523 , 32'h00001CEC , 32'hFFFFA6FB , 32'h0004866B , 32'h0003AFA0 , 32'h000172E4 , 32'hFFFF10F5 , 32'hFFFEF976 , 32'hFFFB5DED , 32'hFFFFA80F , 32'hFFFF3E7E , 32'hFFFFFEC9 , 32'hFFFF0596 , 32'hFFFD876D , 32'hFFFDCD13 , 32'h000779BF , 32'h0001CA7A , 32'h0003766F , 32'hFFF91C08 , 32'h0000221C , 32'h0001611C , 32'h0004834A , 32'hFFFC73DD , 32'hFFFCDA5A , 32'h00006181 , 32'hFFFF38F2 , 32'hFFFC8261 , 32'hFFF853F7 , 32'hFFFCD88E , 32'h0001B6CD , 32'h000137C8 , 32'hFFFC424B , 32'hFFFFEA16 , 32'hFFFF961C , 32'hFFFE6528 , 32'h0001C5ED , 32'h0001D5F2 , 32'h0000F740 , 32'h00010192 , 32'h00003D19 , 32'hFFFFAD21 , 32'h0001934A , 32'hFFFEF134 , 32'hFFFB3C69} , 
{32'hFAB95D50 , 32'hF6F22C40 , 32'h13138B20 , 32'hEE8B05A0 , 32'h136C34E0 , 32'h1676D240 , 32'h2ED31100 , 32'hF8026ED0 , 32'hEC543780 , 32'h3693C500 , 32'h05812E60 , 32'h03BF6E84 , 32'hF5133DF0 , 32'hF7FFC590 , 32'hE5934700 , 32'hE7278B40 , 32'h03246C44 , 32'h00F4F30A , 32'h0524E140 , 32'h027FB6BC , 32'h16EFD8E0 , 32'h069F0070 , 32'h1C6023C0 , 32'hF5004FC0 , 32'hF7203BB0 , 32'hF2786CE0 , 32'hFCD9D0E4 , 32'h10F124E0 , 32'hFB5AA2F8 , 32'h03C090B8 , 32'h027D635C , 32'h0A769FD0 , 32'h107EB6E0 , 32'h00A0D02B , 32'h0BA87850 , 32'h0B1DA0D0 , 32'hFD84CCA8 , 32'h00BE3E60 , 32'hE57DA5C0 , 32'h0C4C4480 , 32'hF9DDE660 , 32'h021111EC , 32'h0A7BD170 , 32'hF1EEB570 , 32'hFEAE62C4 , 32'hFCFB6104 , 32'h00254ADE , 32'h00B5A3C4 , 32'hF7176EB0 , 32'h07CBFD60 , 32'h00B96B8E , 32'hFED8CFE0 , 32'hFA7CB700 , 32'hF8E48FE0 , 32'hFEB4EC40 , 32'h0AF06F00 , 32'h02F54214 , 32'h07AD9CD0 , 32'h02026950 , 32'h01BF18E8 , 32'hFD66C8DC , 32'h00FD371F , 32'hFC4428B0 , 32'hFE0263C4 , 32'h042720B0 , 32'hFE6BFE7C , 32'h023DDBCC , 32'hFC4B12D4 , 32'hFE0DE324 , 32'h04F420B0 , 32'hF9F8C9F8 , 32'h00A85BD5 , 32'hFF5C5BD0 , 32'h01FEBEB4 , 32'h07AE06C0 , 32'hFE665948 , 32'h00FDB44A , 32'hFDA4E960 , 32'h01D91A78 , 32'h01850F48 , 32'hFA731108 , 32'h018DBF20 , 32'hFDD4CB74 , 32'hFDD063DC , 32'hFCFD2BC4 , 32'h01C57A48 , 32'hFCCE0AB0 , 32'hFD8DFDA8 , 32'h020456E0 , 32'hFFD8F69C , 32'h0002F4D1 , 32'h00016AB0 , 32'h0000037B , 32'hFFFFB97D , 32'h0000C9E0 , 32'h00004CC8 , 32'h0001B5F2 , 32'hFFFF5E1E , 32'h0000CE01 , 32'hFFFFB87A} , 
{32'h0002ADD4 , 32'hFFF7055E , 32'h0007FFF9 , 32'hFFFF70C8 , 32'h0003AC87 , 32'hFFFCC075 , 32'hFFFFC761 , 32'hFFFE28A1 , 32'h000007D9 , 32'h00038C42 , 32'hFFFD87EE , 32'hFFFFC7CB , 32'h00010269 , 32'h000396EA , 32'hFFFE8E8E , 32'hFFFA3F73 , 32'h000009CF , 32'h0001E469 , 32'hFFFDB118 , 32'hFFFBD80D , 32'h00018A65 , 32'h0004E64B , 32'hFFF9D9B0 , 32'hFFFB5CA7 , 32'h00072401 , 32'h00026E3C , 32'hFFFF81E1 , 32'h00006C7D , 32'hFFFDE74B , 32'hFFFFD6A8 , 32'hFFFBD0AB , 32'h0003A3F6 , 32'h000193C8 , 32'hFFFBBF60 , 32'hFFFEFFEE , 32'hFFFDE9FA , 32'h0001E1DF , 32'h000272D1 , 32'h000189C6 , 32'hFFFDC989 , 32'h000172A3 , 32'hFFFC4894 , 32'hFFFB4658 , 32'hFFFB0FD2 , 32'hFFF86CAA , 32'h00006BC7 , 32'h0000B091 , 32'hFFFC117B , 32'h00059385 , 32'h00027830 , 32'hFFFF6624 , 32'hFFFEF5F1 , 32'h0003AC18 , 32'h00047EAD , 32'h0006C1AF , 32'hFFFE05DC , 32'hFFFF35F6 , 32'h0004DB63 , 32'h0002F5B8 , 32'h0003EC6E , 32'hFFFE57C9 , 32'hFFFA895C , 32'h00025950 , 32'h0001BFBF , 32'hFFFFC437 , 32'hFFFD962B , 32'hFFFC5B01 , 32'h00064BA5 , 32'hFFFE982F , 32'hFFFE8080 , 32'h00051548 , 32'hFFF98B4A , 32'h0001A3FB , 32'h000379EB , 32'h0005A815 , 32'h0001692D , 32'h0000EDAB , 32'h0001E552 , 32'hFFFDCBCB , 32'hFFFB9DE5 , 32'h000181A4 , 32'hFFFFA4B0 , 32'h0003883D , 32'h00039D85 , 32'hFFFA75A4 , 32'h000717A3 , 32'hFFFEB21C , 32'hFFFD154C , 32'h0001F8DF , 32'hFFFF38A5 , 32'h00006335 , 32'h0000F350 , 32'h000268DD , 32'h00036F9F , 32'hFFFF782A , 32'h00017FCE , 32'hFFFCD469 , 32'hFFFF0136 , 32'hFFFF14A8 , 32'h000118CA} , 
{32'h175E7B60 , 32'hCE837C00 , 32'h2C6EF540 , 32'h01BEB808 , 32'h3BF77500 , 32'h4C691180 , 32'hD85FC3C0 , 32'hF4A2C720 , 32'hEC228AC0 , 32'h201CDD40 , 32'h0C035E60 , 32'hEA4B4B80 , 32'h191231E0 , 32'h08870260 , 32'hF0CF27C0 , 32'hFCC38878 , 32'h21903B80 , 32'h087B1530 , 32'hE4B9A100 , 32'h23868900 , 32'hFF4296D3 , 32'h0355A4E8 , 32'h0D9B1D30 , 32'h10C1D9A0 , 32'h0E5DD530 , 32'hEA1B1E40 , 32'hFDF37304 , 32'h00AD1FC4 , 32'hF343D490 , 32'h0E775040 , 32'hFF6765D4 , 32'hED24C5E0 , 32'hFFE81A9C , 32'h04FAA528 , 32'h0CD90160 , 32'hFBEADB10 , 32'h000626CF , 32'h1F039D60 , 32'h0BD123F0 , 32'h02E8A2EC , 32'hFC4BAAFC , 32'hFF07B67F , 32'hFAC53A20 , 32'h043C5058 , 32'hFAA6DC90 , 32'hFB1A98A0 , 32'hF9D7D7A8 , 32'h04944FD8 , 32'h03FA8E20 , 32'hF3518700 , 32'h07A96D58 , 32'h07999338 , 32'h05531F98 , 32'hF5057FA0 , 32'hFC34C56C , 32'hFB381948 , 32'hF4889150 , 32'h03E43C0C , 32'hFBF21698 , 32'h00FA5F62 , 32'h005B3736 , 32'h041BD408 , 32'h03162ED8 , 32'hFED80178 , 32'h06B76678 , 32'hFE9519C4 , 32'h04104B90 , 32'hFE426810 , 32'h03AE62D8 , 32'hF8A69CD8 , 32'h021AB078 , 32'hFE10D268 , 32'hFC3D9F48 , 32'h02FA7970 , 32'hFFB83FC2 , 32'h001FBF5D , 32'hFA6C1CA0 , 32'h0462D248 , 32'hFFBCE214 , 32'hFA7B5298 , 32'h003A10E6 , 32'hFDF35468 , 32'h052E23C8 , 32'h00053257 , 32'hFE808C8C , 32'hFE743F64 , 32'h004E222D , 32'hFEE36FF4 , 32'hFF419424 , 32'hFF79C1EB , 32'h000038F5 , 32'hFFFE77EA , 32'hFFFDAF0A , 32'h000136B6 , 32'hFFFEB53B , 32'h000064A0 , 32'h00010705 , 32'h000135B9 , 32'h0001A616 , 32'hFFFFE9F6} , 
{32'hFFFE3517 , 32'h00010E11 , 32'h00025FCC , 32'hFFFF4687 , 32'h00004C2A , 32'hFFFE1857 , 32'h0001B8C9 , 32'h000318A1 , 32'hFFFDC25B , 32'hFFFDDB49 , 32'h00024011 , 32'h0002EAA1 , 32'h00000CA3 , 32'hFFFCD449 , 32'h0001AEAA , 32'hFFFD46CC , 32'hFFFF7B79 , 32'h00020516 , 32'h00001C85 , 32'hFFFDEE03 , 32'hFFFE5D40 , 32'h000338BC , 32'h00025F0A , 32'hFFFBE235 , 32'hFFFEB867 , 32'h0000A933 , 32'hFFFCECEF , 32'h0004C827 , 32'hFFFC4C3F , 32'h0002BD7A , 32'h0000D2DD , 32'hFFFD4303 , 32'hFFFD9E2F , 32'hFFFF728B , 32'h00003FBF , 32'h0000618D , 32'h000423F1 , 32'h00070188 , 32'hFFFC0089 , 32'h0000121F , 32'hFFFC228E , 32'h0000B5EB , 32'hFFFCE3B3 , 32'h0003CCF3 , 32'h0001F377 , 32'hFFFD29F7 , 32'hFFFE25A2 , 32'hFFFFE7F6 , 32'h00001759 , 32'h000837D5 , 32'hFFFDEBD4 , 32'hFFFED326 , 32'hFFFD5CD2 , 32'hFFFBD765 , 32'h0000C777 , 32'h0001EDDC , 32'h0001096F , 32'h00018F51 , 32'h000520ED , 32'hFFFDCB4D , 32'hFFFB0613 , 32'h00001A7C , 32'hFFFFA1F2 , 32'h00017594 , 32'h00005FFF , 32'h0002B78D , 32'hFFFC56C5 , 32'h0004E7ED , 32'h000442FD , 32'hFFFF6009 , 32'h00042255 , 32'h0002D34A , 32'hFFFB0458 , 32'hFFFF400B , 32'h00059A30 , 32'hFFFC6155 , 32'hFFFAA018 , 32'hFFFC2F93 , 32'hFFFE7A6E , 32'hFFFC0F33 , 32'h0001423B , 32'h00025D20 , 32'hFFFF541E , 32'hFFFEDEF4 , 32'hFFFF4A7B , 32'h0002919D , 32'hFFFDE2AE , 32'hFFFE5486 , 32'hFFFBB53F , 32'hFFFCD061 , 32'h0004C2A0 , 32'hFFFBD03F , 32'hFFFF668C , 32'h0001BCDF , 32'hFFFF7DFC , 32'hFFFD8105 , 32'h0000D156 , 32'hFFFD881A , 32'h00005DD0 , 32'h00027988} , 
{32'h06E11380 , 32'h4AF03580 , 32'h21A7E840 , 32'h1A873A20 , 32'h1F82CDE0 , 32'h0B863550 , 32'h3E1DA980 , 32'h35306B00 , 32'h19110AA0 , 32'h1D6713A0 , 32'hECF93980 , 32'h061BCF90 , 32'h06C74B88 , 32'h058E26A0 , 32'hF79E2610 , 32'hFCA0ECD4 , 32'h1B17ACA0 , 32'hF1A90600 , 32'hED991A20 , 32'hFF51EA1C , 32'hF351A710 , 32'hF7640390 , 32'hF521C6F0 , 32'h11420A00 , 32'hF43E86F0 , 32'hF81294B0 , 32'hF87D2BE8 , 32'h116C4160 , 32'h03F3EE98 , 32'hEDF72780 , 32'hF6616BC0 , 32'hE214EB20 , 32'hFEEB24C8 , 32'hF3E72E60 , 32'h009B3390 , 32'hF90E0038 , 32'hFD5D95B4 , 32'h04AE92E0 , 32'h0F768970 , 32'hFC49C518 , 32'hE4E23520 , 32'hFAD95980 , 32'h0891D2B0 , 32'hF93D1C48 , 32'hF4767B60 , 32'h0DAACB30 , 32'h04F6C418 , 32'h00BB5768 , 32'h0A44BFA0 , 32'h01F91648 , 32'hF8CDE908 , 32'hF984AE10 , 32'h01B25E3C , 32'hFDF9F4FC , 32'h05641DD0 , 32'hFCB7E210 , 32'hFA7A9C80 , 32'h00FE14B2 , 32'h03B27CBC , 32'h00737E4A , 32'hF8F44968 , 32'hF6B58DB0 , 32'h028A437C , 32'hFB5234A8 , 32'hFC2A0C78 , 32'h04202978 , 32'hFE4949FC , 32'h0411B930 , 32'h023FA8C4 , 32'h06A5FC40 , 32'h02B34400 , 32'h00FFB7C9 , 32'h035FEBE8 , 32'hFCA7B640 , 32'hF9F11A08 , 32'hFBF11628 , 32'hFB26A0C8 , 32'hFE0352F8 , 32'hFE7B494C , 32'h007855EE , 32'h068FCD10 , 32'h006270CE , 32'hFDAC8CEC , 32'h006025C5 , 32'hFFC8E52F , 32'h02FF69D0 , 32'hFE1F8CB0 , 32'h00243C35 , 32'h02A08608 , 32'h0095205B , 32'h00003444 , 32'hFFFFC526 , 32'h00006518 , 32'h0001B7CE , 32'h000158DB , 32'hFFFF1608 , 32'h00008D57 , 32'h0001728E , 32'h00005D34 , 32'hFFFF9C6A} , 
{32'h228D9340 , 32'hF838EEB0 , 32'hF6530D20 , 32'h24346100 , 32'hFF5E2CC9 , 32'hEF59F700 , 32'hF7471E80 , 32'hFAE49770 , 32'hFAE2C428 , 32'hD93F4580 , 32'hF7186C00 , 32'h18A69980 , 32'hF43EBF70 , 32'h0D655130 , 32'hE64C8440 , 32'hED646C00 , 32'h12798A00 , 32'h01338910 , 32'h0614C430 , 32'hFAD422F0 , 32'hF1EEDA50 , 32'hF319EC30 , 32'h0E33B090 , 32'h01C388B8 , 32'hF9FBF968 , 32'h03424020 , 32'h05E32618 , 32'hF87E0CE0 , 32'hD5EF1A40 , 32'hFB5FDA28 , 32'hF52D6560 , 32'hEFFB4620 , 32'hFB0B5160 , 32'h00C60896 , 32'h07260428 , 32'hF6781AF0 , 32'h086237F0 , 32'hFC9C1B44 , 32'h0485C1A0 , 32'hF66A8750 , 32'h02BA6ED8 , 32'hFA253720 , 32'hFC9A8F70 , 32'h0438B720 , 32'hEF4EE660 , 32'h04E0CDE8 , 32'hF97F00C0 , 32'hFED3BB08 , 32'h020D1368 , 32'hFD5E3000 , 32'hFF70FCC2 , 32'h0B503BE0 , 32'hFB0F76C8 , 32'h00BB4677 , 32'hFD86F8E0 , 32'h048A0000 , 32'hFF8C7C5D , 32'hF84984E0 , 32'h05145CC0 , 32'h02A8BAC4 , 32'hFDB27CF0 , 32'h07203638 , 32'hFF2225A3 , 32'hFCB4C7DC , 32'h053B2710 , 32'hFBAA4228 , 32'hFF6F4494 , 32'h07398CB0 , 32'h05BD88D0 , 32'hFB978C20 , 32'hF9F4B8C8 , 32'hFE1C657C , 32'hFE55E17C , 32'hFF53A80B , 32'hFDE6216C , 32'h006F020C , 32'h0223CE70 , 32'hFFD5F3CC , 32'hFC42235C , 32'h021F2788 , 32'hFF0C4C0C , 32'hFA868E08 , 32'hFA64C4E0 , 32'h093EF480 , 32'h039E0294 , 32'hFE3A7430 , 32'hFC09C54C , 32'hFE479CF0 , 32'hFFE290BF , 32'hFF3175E1 , 32'h000177A0 , 32'hFFFF41EC , 32'h0000B0C0 , 32'h0000CFD7 , 32'hFFFEFD6F , 32'hFFFBE8D7 , 32'hFFFFAC78 , 32'hFFFF727C , 32'hFFFE662E , 32'h00017300} , 
{32'hA9020C00 , 32'h172217C0 , 32'h41753D80 , 32'hC7D5B580 , 32'hD6501B00 , 32'h06D973C8 , 32'h048F8A30 , 32'hF21EC5E0 , 32'h02A264CC , 32'hF2045CC0 , 32'hDBD26FC0 , 32'h07478D30 , 32'h080E13C0 , 32'h1BEDF520 , 32'hF064A7B0 , 32'h05AF1E50 , 32'h1BFADA40 , 32'hFF07B3FE , 32'h0DD0F9B0 , 32'h0E270F30 , 32'hF93D8320 , 32'hE6797260 , 32'h10DC3B80 , 32'hFF51A976 , 32'hFE1DFF84 , 32'h1DB8B280 , 32'h186C7D00 , 32'h04976C60 , 32'h0075EBC4 , 32'h0806D410 , 32'h0DC60190 , 32'hE8FC08A0 , 32'h1082E580 , 32'h02882360 , 32'hFE7CCE10 , 32'h08A7B710 , 32'hF912D880 , 32'hFA760720 , 32'h00D8153F , 32'h0406F980 , 32'h0116D048 , 32'h0EBAEEF0 , 32'hF88448F0 , 32'hFFF73FED , 32'h024F823C , 32'hFBA4FE50 , 32'h020EAB9C , 32'h09FEB640 , 32'hF861D6A8 , 32'hFCC04228 , 32'hF8A1AA00 , 32'h02C664BC , 32'hF9077E78 , 32'hF77DFF70 , 32'h07A945B0 , 32'h012B1E58 , 32'hF52BE090 , 32'h077D7670 , 32'hF35908E0 , 32'h05791430 , 32'h016DA890 , 32'h04FABEC0 , 32'hF89611B0 , 32'hF7877880 , 32'hFE329EF0 , 32'h05311C20 , 32'hFD6FA170 , 32'hFB233E68 , 32'hFF4B06CF , 32'h0038E26F , 32'hFBD8D668 , 32'hFCE81BA4 , 32'h02C39F64 , 32'hFA50A770 , 32'hFF34C736 , 32'hFFFCC8C1 , 32'hFB7ACB88 , 32'hFC9F8900 , 32'h0095DE68 , 32'hFFC8CB26 , 32'h064F6E30 , 32'h028A79E0 , 32'hFD7FA38C , 32'h01BA3E3C , 32'hFE8913DC , 32'hFDCBDD8C , 32'h018EC178 , 32'h01353140 , 32'hFD1C4F8C , 32'hFFECEAD3 , 32'h00030250 , 32'h000041BA , 32'hFFFF08F3 , 32'hFFFE0E1D , 32'h0000F63B , 32'hFFFF3D94 , 32'h000051C6 , 32'h00008F95 , 32'hFFFF9FC8 , 32'hFFFE67E2} , 
{32'h0E4D9870 , 32'hD4F55C40 , 32'hF83BA0F8 , 32'h54E59700 , 32'h099282D0 , 32'h269D44C0 , 32'h0DE0B6F0 , 32'hC4B04940 , 32'h2BE9D300 , 32'h081F81E0 , 32'h0C0D71A0 , 32'h1FC50AE0 , 32'hEC5FD520 , 32'h1EE63E00 , 32'hEB49FC40 , 32'h03E4F9E8 , 32'h142C19E0 , 32'hE9949E80 , 32'h120DDAE0 , 32'h07CF1BE8 , 32'hF507CC70 , 32'h1675CA60 , 32'hFBD09F68 , 32'h15059AE0 , 32'hF7614B70 , 32'h03554000 , 32'h155F22E0 , 32'h192567A0 , 32'h02541C1C , 32'hEFF94080 , 32'hEEA72360 , 32'hF41F1610 , 32'h003AD5DB , 32'h0A302010 , 32'hF5F7DD60 , 32'hF18B3690 , 32'hF492FFF0 , 32'hF4738290 , 32'h0865DEE0 , 32'hFC830330 , 32'h11B345E0 , 32'hF9C03CC0 , 32'hF99F9D68 , 32'h03DEBF38 , 32'h018CB820 , 32'hF9CAD870 , 32'hF96CDB40 , 32'h02C804CC , 32'hF307FC50 , 32'h08DA4BF0 , 32'h044D5640 , 32'h06A6D1A8 , 32'hFD777DBC , 32'h000AEAF5 , 32'hF91975A8 , 32'h04B8D768 , 32'h0B145170 , 32'h0AB9A550 , 32'h040900E8 , 32'h055CF978 , 32'hFEC71F18 , 32'hFF2868D9 , 32'hFFF1375C , 32'h0347F320 , 32'hF639F9B0 , 32'h041AB608 , 32'h0330C12C , 32'hFA2B4AA0 , 32'hFEC69964 , 32'h0583F7E0 , 32'hFFF84E42 , 32'h00AD8B3C , 32'hFFBFE08E , 32'hFDA7F138 , 32'h0081629B , 32'h0104D7E4 , 32'h02D813F8 , 32'h053BFB68 , 32'hFE28CDA0 , 32'h01CD3A08 , 32'hFFCC0E11 , 32'h0123DB98 , 32'hFFFAF78D , 32'hFCD47CA8 , 32'hFE504A44 , 32'h01A65BF4 , 32'h02A654C8 , 32'h00E1C134 , 32'hFFD7D362 , 32'h00696319 , 32'h00006F22 , 32'h00025C11 , 32'hFFFFFC3B , 32'h00003786 , 32'h0000BAF4 , 32'hFFFF2221 , 32'hFFFFB32D , 32'hFFFF445C , 32'hFFFFB32E , 32'h00000ADF} , 
{32'h00024761 , 32'h00012E04 , 32'hFFFD2966 , 32'h00043CE8 , 32'h0001BBD9 , 32'hFFFB8152 , 32'h00011D17 , 32'hFFFE63A6 , 32'h00038D4A , 32'h00025FCA , 32'hFFFAA8BB , 32'hFFFACED7 , 32'hFFFA478F , 32'h00011F3B , 32'h0002B42C , 32'hFFFF3BAE , 32'hFFFFCB33 , 32'h00014B31 , 32'hFFFF662E , 32'hFFFE8865 , 32'hFFFC45E9 , 32'h0001CD69 , 32'hFFFD0968 , 32'h00018DFF , 32'hFFFFE591 , 32'h0000820D , 32'h00034B04 , 32'hFFFDB269 , 32'hFFFAFCDB , 32'h00017241 , 32'h00009A3D , 32'hFFFED327 , 32'hFFFAEA80 , 32'h0003F900 , 32'h000426D5 , 32'hFFFD4585 , 32'h0000C548 , 32'h00024694 , 32'h00005BB0 , 32'hFFFD74B9 , 32'hFFFF2C7D , 32'hFFFD6BE7 , 32'h0000246C , 32'h0000068F , 32'hFFFF63BE , 32'h0001BF9F , 32'hFFFE9074 , 32'hFFFFDC9D , 32'hFFFB9E05 , 32'h000063DF , 32'hFFFF258B , 32'h0001238A , 32'hFFFECEDD , 32'hFFFCC782 , 32'h00002DB1 , 32'h0001955B , 32'h000067AC , 32'hFFFE8A7D , 32'h000018CB , 32'h0003A03A , 32'h0001A36F , 32'h00020BB6 , 32'hFFFF7A0B , 32'h0001E622 , 32'h00016D5F , 32'h000428D0 , 32'hFFFF55CD , 32'hFFFE89CD , 32'hFFFD6619 , 32'h00030F13 , 32'hFFFD9936 , 32'h0002C335 , 32'h0001F95C , 32'h0002C662 , 32'h0001ABC5 , 32'hFFFCC206 , 32'h000202B3 , 32'hFFFC6BB9 , 32'hFFFC5C52 , 32'h000378A6 , 32'hFFFED43E , 32'h00037DB3 , 32'hFFFF4538 , 32'h000084CB , 32'hFFF9F22C , 32'h0000E89C , 32'hFFFD41E3 , 32'hFFFD4F94 , 32'h000532EA , 32'hFFFCE848 , 32'h000457A2 , 32'h0000B80D , 32'hFFFFF741 , 32'h00008BE1 , 32'h000064FE , 32'h0000C26F , 32'h0000F63B , 32'hFFFE8234 , 32'h00006F1C , 32'h0000BAF0} , 
{32'h04F6AE28 , 32'h02CD8508 , 32'h1C629460 , 32'hEB2867A0 , 32'hFCE99754 , 32'hDD71A940 , 32'h06B88238 , 32'hEFCC1D60 , 32'hF47005E0 , 32'hF911DA78 , 32'hF20F4A70 , 32'hE9A4B580 , 32'h00533913 , 32'h00E9A0C5 , 32'h033A1728 , 32'h04C3F728 , 32'hF9DE2D10 , 32'h01C67B78 , 32'hFCB53E9C , 32'hFB5EB4A0 , 32'h09C04F80 , 32'hF0190410 , 32'hF8704CE0 , 32'h0BDBC210 , 32'hE81615E0 , 32'h1144BE20 , 32'hEE47B2A0 , 32'h08545E90 , 32'h05C0C840 , 32'h056CD830 , 32'hF93EA538 , 32'hE52806A0 , 32'h0393904C , 32'hF8A1C5E0 , 32'h08775540 , 32'h12E0FB60 , 32'hFBE4E2B0 , 32'hFBA48040 , 32'hF5D067A0 , 32'hFAF96900 , 32'h03842AE8 , 32'hF7ED6590 , 32'h03B53548 , 32'hFF218A1E , 32'hFD043F30 , 32'h069FB810 , 32'hF7FF81B0 , 32'hF8029C28 , 32'hF7A49A80 , 32'h0B60BD50 , 32'h11CC9A20 , 32'h00001FA3 , 32'h057434C0 , 32'h08EC2960 , 32'h03A83FC4 , 32'hFCF32F90 , 32'hFAA01598 , 32'hF83FA5F0 , 32'hF95B8DE8 , 32'h04ECF0B0 , 32'hFF765111 , 32'hFE7BD2EC , 32'hFF8C9907 , 32'hFE93BDE0 , 32'hFE63DDBC , 32'h06E62838 , 32'h0522E3B8 , 32'h0346974C , 32'hFC8DFB18 , 32'hFFDDE15A , 32'hFF6FF5FC , 32'hFABE93B0 , 32'hFA92BE88 , 32'h07EEABA0 , 32'h01BCE924 , 32'h00F1D1D1 , 32'h007671D2 , 32'h03788AD4 , 32'h04B9B5A8 , 32'h01321158 , 32'h00758182 , 32'hFFB0634C , 32'hFF656561 , 32'hFCE66040 , 32'h04105020 , 32'hFE50CE90 , 32'hFED928EC , 32'h00656E8E , 32'h00D5566F , 32'hFF36143F , 32'h00017E70 , 32'h000219A2 , 32'h00015DDE , 32'h000070F5 , 32'hFFFD9281 , 32'hFFFEB6E7 , 32'hFFFF7B2D , 32'h00016652 , 32'hFFFDDD4C , 32'hFFFFD44E} , 
{32'hF93F84A0 , 32'hFF1FF05A , 32'h04033BC0 , 32'hFDD338D0 , 32'hFF6B78BD , 32'hFCC5E2AC , 32'h00109A08 , 32'h012456BC , 32'h053BC480 , 32'h0149F9E4 , 32'hFB73E640 , 32'h06786498 , 32'h05861030 , 32'hFACDA6B8 , 32'hFFE99F22 , 32'hFC87B0C8 , 32'hFB201080 , 32'h1080D520 , 32'hFAA2AD98 , 32'h05F40B70 , 32'hFAD9E480 , 32'hFEB03EEC , 32'hFEB99E9C , 32'hFD9C6E44 , 32'hFFBAD308 , 32'h02F46220 , 32'h03CD48A8 , 32'h000E4FFA , 32'h01B53A70 , 32'hFD4D4228 , 32'h04E03D68 , 32'hFE6B1278 , 32'h02D022B0 , 32'hFE7CB49C , 32'h02A771C8 , 32'h009BB9C2 , 32'hFEE3A1E0 , 32'hFFE63A4B , 32'hFAD0DDE0 , 32'hFEF4C4DC , 32'hFCB22884 , 32'h054A7610 , 32'hF86F3F70 , 32'hFC31C9EC , 32'hFF3B1C52 , 32'h041861A8 , 32'hFB68B040 , 32'hF94459C0 , 32'h042AA6E8 , 32'hFDAAA294 , 32'hFCA55B7C , 32'hFD8907C4 , 32'h00405EC3 , 32'h0242029C , 32'h08979BF0 , 32'hFD5F96CC , 32'hFE193A1C , 32'h011ECB48 , 32'h03B32BD0 , 32'h02B96C68 , 32'hFC965EB4 , 32'hFEFC81F0 , 32'h07E86990 , 32'hFF15D833 , 32'hFC888508 , 32'hFF88AA1B , 32'hFD538C90 , 32'hF996AC78 , 32'h04DA0AF8 , 32'h0179AC10 , 32'hFFA888B6 , 32'hFDA1FB0C , 32'hFF2214D9 , 32'h012082E4 , 32'hFB6F4500 , 32'hFFF73491 , 32'h03826D08 , 32'hFFFEA9A4 , 32'hFEF3ED00 , 32'hFDACB96C , 32'h00F82C50 , 32'hFDABFA40 , 32'h02308C4C , 32'h0129114C , 32'hFD580C88 , 32'h00C45F9D , 32'hFDC6FE5C , 32'hFDF3A3A0 , 32'hFF6AAF3E , 32'h005A59B1 , 32'hFFFD8940 , 32'hFFFF761F , 32'h0002D1B8 , 32'hFFFCFC9A , 32'h00046CCA , 32'h00010E8F , 32'hFFFE8363 , 32'hFFFDCA42 , 32'h00028AD2 , 32'hFFFC57FE} , 
{32'hFFFF1833 , 32'h000345AC , 32'hFFFC03C9 , 32'hFFFF0A59 , 32'hFFFDB891 , 32'hFFFFD419 , 32'h00005418 , 32'h0004FC97 , 32'h0001CF99 , 32'hFFFCA88E , 32'h00011438 , 32'hFFFD8AE6 , 32'hFFFC2B2F , 32'h00011F29 , 32'h0001425C , 32'hFFFDE1D4 , 32'h000097E0 , 32'hFFFC2785 , 32'h0000833F , 32'hFFFDDD11 , 32'hFFFB70D6 , 32'hFFFE0BD8 , 32'h000392DC , 32'h000110B6 , 32'hFFFAC083 , 32'hFFFE84DE , 32'h0000315B , 32'hFFFE3AD6 , 32'hFFFD7CE4 , 32'h0002FDF5 , 32'h00005E0F , 32'h00015016 , 32'h0003ADF4 , 32'hFFFE0CD4 , 32'hFFFF0A8C , 32'hFFFE2FB0 , 32'hFFFEEF23 , 32'hFFFDF6BB , 32'hFFFE5017 , 32'h0001D68A , 32'h00039024 , 32'h000094EE , 32'hFFFECEE1 , 32'hFFFF2C9F , 32'h00048CEA , 32'h00025536 , 32'h00000234 , 32'hFFFC3D25 , 32'h00003211 , 32'h0002D910 , 32'hFFFEFC78 , 32'h000154FF , 32'h00019CB5 , 32'hFFF97D25 , 32'hFFFD0388 , 32'h0000E3A8 , 32'hFFFF3A54 , 32'h000012E1 , 32'h00004688 , 32'hFFFC0EDE , 32'h0004824F , 32'hFFFBD5ED , 32'hFFFD4FC5 , 32'hFFFFBA38 , 32'h0005EA8A , 32'h00014A03 , 32'h00013752 , 32'h00005391 , 32'hFFFFC045 , 32'hFFFDAC06 , 32'hFFFC99C9 , 32'h00016AB9 , 32'hFFFD229C , 32'h00021157 , 32'hFFFFF537 , 32'h00023BF1 , 32'h0000EB37 , 32'hFFFBD8C8 , 32'h00020313 , 32'h00012716 , 32'h000353FF , 32'hFFFBC9C4 , 32'hFFFF585B , 32'hFFFDDADB , 32'h0001D415 , 32'hFFFE7AC3 , 32'h0000E327 , 32'hFFF9A8B9 , 32'hFFFE9D46 , 32'h00050C86 , 32'h0002D4B3 , 32'hFFFF518F , 32'hFFFDC2D0 , 32'hFFFF2E38 , 32'hFFFF19F7 , 32'h00002169 , 32'h000064DD , 32'h0002210B , 32'hFFFDD46C , 32'hFFFF5F87} , 
{32'h0B001720 , 32'hF25CB240 , 32'h0BBCF970 , 32'hF7A94F90 , 32'h1CFDC6C0 , 32'h0333A9A8 , 32'hEFDBCD20 , 32'h1CDC5240 , 32'hFBC020C8 , 32'hFDC3F754 , 32'h04D46AF8 , 32'hF3C08FD0 , 32'hFF6D0492 , 32'h060C2B78 , 32'hFC42EDFC , 32'hEE5E00C0 , 32'h02C71A00 , 32'h10211EA0 , 32'h022FABC8 , 32'h0231A26C , 32'h059C6A58 , 32'hF01297A0 , 32'h06A195A0 , 32'hFEA7A7A8 , 32'hFCAF8D60 , 32'hF21136D0 , 32'hEE3215A0 , 32'h1DE4E3C0 , 32'h02417AC4 , 32'hEF3616E0 , 32'h02F5EFEC , 32'h00395C7E , 32'h0177BBA4 , 32'h0A922830 , 32'hFF6970CC , 32'h090BC390 , 32'h0E435CA0 , 32'h056D27E8 , 32'h047310E0 , 32'hFB74AD80 , 32'h00078860 , 32'hFD285318 , 32'hFF4A7EE5 , 32'h035616E0 , 32'h02031390 , 32'h0242FB3C , 32'hFE18F5B0 , 32'hF8844388 , 32'h02453D70 , 32'hF4DD3790 , 32'hFCA00754 , 32'hF61E8A40 , 32'h07B0D3F8 , 32'h077F6760 , 32'h03768A2C , 32'hF6AE44C0 , 32'h06EC50C0 , 32'hFB2C12F0 , 32'h01E31A10 , 32'hFC98C07C , 32'h009B0CC9 , 32'hEFA35100 , 32'hFBD738E0 , 32'hFFE9280D , 32'h0A4F46B0 , 32'hFF891F59 , 32'h0185239C , 32'hFF5B5D41 , 32'hFB7BBD38 , 32'hF9E38000 , 32'h041DECD0 , 32'hFF127A0F , 32'hFC844578 , 32'hFDCABC18 , 32'h076DE978 , 32'hFC81680C , 32'h030A70D0 , 32'hFF345D28 , 32'h04259900 , 32'h022834FC , 32'hFDA21D40 , 32'h0639E220 , 32'hFCFA7B7C , 32'h0556E640 , 32'hFE4B1A04 , 32'h001C83DF , 32'h010BF320 , 32'h01F6066C , 32'h0036BE03 , 32'h007FFDB6 , 32'hFFFE8DC0 , 32'h00011CBA , 32'h000062FB , 32'h0001736C , 32'h000087AA , 32'hFFFE32C1 , 32'hFFFE7BF7 , 32'hFFFEA335 , 32'hFFFFD715 , 32'hFFFECCF4} , 
{32'hFFFF62D9 , 32'h000132EE , 32'hFFFD7B44 , 32'h00019113 , 32'h0000DECA , 32'hFFFFD13F , 32'h00004D32 , 32'hFFFCC501 , 32'hFFF9EB81 , 32'h000044B2 , 32'hFFFECFE4 , 32'hFFFCF11D , 32'h000002E2 , 32'hFFFBFAD9 , 32'h00019F4D , 32'h00018259 , 32'h00026C2E , 32'hFFFDCDBA , 32'h00012C05 , 32'hFFFFE66F , 32'h00014155 , 32'hFFFFB027 , 32'hFFFEA1B6 , 32'hFFFF7815 , 32'hFFFC936B , 32'hFFFDD72F , 32'hFFFF45C4 , 32'hFFFFCA65 , 32'hFFFDDC5D , 32'hFFFD6EF2 , 32'h0005CFA4 , 32'hFFFF741D , 32'h0002F181 , 32'hFFFE8D83 , 32'hFFFDF16C , 32'hFFFD5DD7 , 32'h000149E7 , 32'h0000AC9F , 32'hFFFEE725 , 32'h0002723A , 32'h00022637 , 32'hFFFE3ECE , 32'h0000CFA8 , 32'hFFFE9B35 , 32'hFFFF4AF0 , 32'hFFFE5054 , 32'h00036765 , 32'h0000B140 , 32'hFFFF32CC , 32'hFFF95215 , 32'h00003F06 , 32'hFFFFAF50 , 32'hFFFBC484 , 32'hFFFFBCFE , 32'h00015C0E , 32'hFFFA241F , 32'hFFFA866A , 32'hFFFF7E3F , 32'h0000EEFE , 32'hFFFECB08 , 32'h0002F16E , 32'h0007812B , 32'h0003A02D , 32'h0002D2BE , 32'hFFFE4B3F , 32'h0001A1C0 , 32'h0000F88D , 32'hFFFBDEAE , 32'h0000B99D , 32'hFFFF3CE5 , 32'hFFFF2A9F , 32'h000393B1 , 32'hFFFF8AC9 , 32'h00011B37 , 32'h0001DAAC , 32'h0000DF40 , 32'hFFFF1F68 , 32'hFFFD700E , 32'hFFF920EA , 32'hFFFFB1F0 , 32'hFFFF4D93 , 32'h0000EF06 , 32'hFFFADBAF , 32'hFFFF4A8C , 32'h00028202 , 32'hFFFC3F88 , 32'h0003CA17 , 32'h0005A8BF , 32'h0001C4DD , 32'hFFFDA54A , 32'h0000F36C , 32'hFFFECD20 , 32'hFFFBF034 , 32'h0000BF9D , 32'hFFFD96A1 , 32'hFFFFD81B , 32'hFFFE49E8 , 32'hFFFAE7FE , 32'h000160D7 , 32'hFFFFBFCB} , 
{32'h01F3FB00 , 32'hFC26BABC , 32'h07CBC400 , 32'hFBAAE050 , 32'hFEF1C3E8 , 32'h08368520 , 32'h0129BED4 , 32'hFED07B70 , 32'h02354CD8 , 32'hFF52F149 , 32'hF51DC830 , 32'h01B2D11C , 32'hFA7E6580 , 32'hF7B57880 , 32'hF6A065B0 , 32'h00E723AD , 32'hFFBB0D51 , 32'hFF03D60A , 32'hFCA40570 , 32'hFEFE2DD4 , 32'hFBBB2010 , 32'hFAF98E28 , 32'hFDB69460 , 32'h049271B0 , 32'hF9C16010 , 32'h027C87C0 , 32'hFD662420 , 32'hF95CFD60 , 32'h026A3108 , 32'hFA9E0DF8 , 32'h01C029A4 , 32'h02A61450 , 32'h024A6E1C , 32'h01D2DECC , 32'h07F57660 , 32'hFA6ED5A0 , 32'hFC249B98 , 32'h024D2CE0 , 32'hFE01F324 , 32'hFE79A5F8 , 32'hFEDEBCB4 , 32'h032790EC , 32'h03FF79F4 , 32'h095DF170 , 32'hFEBFD000 , 32'h01056718 , 32'h02138718 , 32'h0038B284 , 32'h019ED524 , 32'hFE9236E8 , 32'hFEED877C , 32'h05E13608 , 32'hFFF62CEF , 32'hFF0F5DD1 , 32'hFEA6BA30 , 32'hFCDEF858 , 32'h0894A5B0 , 32'hFA4C9BC8 , 32'hFD148FC4 , 32'h055CA1C8 , 32'h04A66268 , 32'h02664090 , 32'hFCAD9264 , 32'h07E49898 , 32'h0235FFB4 , 32'hF8E98948 , 32'hFE3271C8 , 32'hF9291200 , 32'hFA7D1100 , 32'hFF09FBBE , 32'h012B0BE0 , 32'hFACEE188 , 32'h012AB4AC , 32'hFBA324F8 , 32'hFE9B40F0 , 32'hFDE609E0 , 32'hFD79A1BC , 32'hFE439A24 , 32'hFDC0C780 , 32'h00AB5790 , 32'hFB386A90 , 32'hFCF9026C , 32'h00818B37 , 32'hFC5E46FC , 32'hFEFC6D9C , 32'h042A97E0 , 32'h00499ECC , 32'h04104C80 , 32'hFF703D85 , 32'h008E8684 , 32'hFFFDA9AB , 32'hFFFD2DDE , 32'hFFFEC515 , 32'h0003DDCF , 32'h00009F2E , 32'hFFFE5167 , 32'h00006B1B , 32'hFFFE4533 , 32'hFFFE573A , 32'hFFFFFB2F} , 
{32'h2D431B80 , 32'hEA642A80 , 32'h3E130E80 , 32'h02B4EFD0 , 32'h15B17380 , 32'h25831D40 , 32'h159E3B40 , 32'h015ECBBC , 32'h0BFF7A20 , 32'h0FEFC260 , 32'hCC56C400 , 32'h14BC7440 , 32'hFD98A134 , 32'h110EE6C0 , 32'h13259800 , 32'h0937EA80 , 32'hF1DEC120 , 32'hEEB40200 , 32'hEBC80B20 , 32'h0EEBD7D0 , 32'hF751B3C0 , 32'hF743DF70 , 32'h06B07A00 , 32'hF3FE2BB0 , 32'h1A913C60 , 32'hF74419C0 , 32'h05DBCC78 , 32'hF39B8590 , 32'hE7705160 , 32'hFB9ACD60 , 32'hF2EF8F30 , 32'hFD3F733C , 32'h0CBDCD90 , 32'h07ECE830 , 32'h08550C30 , 32'h0D8123D0 , 32'h03E38DC8 , 32'hEEEAC800 , 32'hFD509828 , 32'h01595464 , 32'hFBF54120 , 32'h080A7C70 , 32'h054E4BC0 , 32'h01F46190 , 32'hF71F0B30 , 32'h00B2637D , 32'hF9FA5518 , 32'h0BD7EE80 , 32'h08D82600 , 32'h08D08420 , 32'hF8E16BA0 , 32'hFF877250 , 32'h039079E0 , 32'h07CD1E50 , 32'hF93ABC20 , 32'hF3EC0830 , 32'h0C8B1A30 , 32'hF0CFAF30 , 32'hFD2D4870 , 32'hFF9FFA7F , 32'h014618B4 , 32'hF9F6E088 , 32'h0CD42190 , 32'h03C38CC0 , 32'hFDB35E54 , 32'hFD0CC680 , 32'hFBCEEE20 , 32'hFC251D7C , 32'h01666C7C , 32'h02B770C0 , 32'hFF826F18 , 32'hFC0D8F4C , 32'h01B4B50C , 32'h05BCEC08 , 32'hFEF3D5F0 , 32'hFC15CAB8 , 32'h00A07749 , 32'hFE1B3C40 , 32'hFCE132C0 , 32'h0433B9E8 , 32'hFF7C1DAA , 32'hFBF8D450 , 32'h02549D98 , 32'hFB920DB8 , 32'h0200A5C4 , 32'h030209AC , 32'hFEC38A7C , 32'hFE6B341C , 32'hFE6A5790 , 32'hFF983B77 , 32'h000133E6 , 32'h0000B749 , 32'h0000D3DE , 32'hFFFDFD0D , 32'h00002FB4 , 32'h0000EBC4 , 32'h00014145 , 32'hFFFE6540 , 32'hFFFFD77E , 32'hFFFF879C} , 
{32'h416B9D00 , 32'h1652B1E0 , 32'h0FAC5DE0 , 32'h082DAB90 , 32'h072E4130 , 32'h1F40E3A0 , 32'hE82A86E0 , 32'hF67FB5F0 , 32'h0E5714D0 , 32'h066A1460 , 32'h02AFAA64 , 32'hF51DFE70 , 32'hFCF779D8 , 32'hF4A76420 , 32'h05065AB0 , 32'h09616A30 , 32'h0E8B3750 , 32'hFE807F24 , 32'h19FC7600 , 32'h05449CD8 , 32'h0DEF1DA0 , 32'h038B67B0 , 32'h01DFE344 , 32'h08725F30 , 32'h06509830 , 32'hF1363600 , 32'h0A9A9AA0 , 32'hED2E78E0 , 32'h07872D78 , 32'h06D4AB58 , 32'hEE4E90E0 , 32'hF2086260 , 32'hF8D6EE80 , 32'hF7CD4760 , 32'hEEA07060 , 32'hFDB33F10 , 32'hFC77D438 , 32'h03CCAB34 , 32'hF68C43F0 , 32'hF3327060 , 32'hFF3B3575 , 32'hFC83B5C0 , 32'h037CE454 , 32'hF6582900 , 32'hFBB76568 , 32'h02A4718C , 32'hFC290448 , 32'h0D1F0D60 , 32'hF45E7110 , 32'hFB0F1048 , 32'h0272F284 , 32'hFC37BBCC , 32'hF7492A00 , 32'hF727A090 , 32'h012A4A88 , 32'h0B10FB70 , 32'h063128B8 , 32'hFF9DB7E8 , 32'h078CBDA8 , 32'hF7773710 , 32'h0D6B5210 , 32'hF8BFD188 , 32'h02A13494 , 32'h001B797C , 32'h0762B950 , 32'hFF0EBBC3 , 32'hFED52928 , 32'h039C789C , 32'hFC1788C0 , 32'h020C4200 , 32'h032EC2C4 , 32'h01B4F654 , 32'h0426CE20 , 32'h0365E2AC , 32'h031E3928 , 32'h06655B88 , 32'hFE2CC9C4 , 32'h03551224 , 32'h01E8327C , 32'h037D1758 , 32'hFD8995E4 , 32'h008403A0 , 32'hFF234300 , 32'hFFB13948 , 32'hFD26F410 , 32'hFDFC4654 , 32'hFA613D10 , 32'h031CEFF8 , 32'hFF6948EF , 32'hFF316956 , 32'hFFFEA066 , 32'hFFFF5577 , 32'h00012ED0 , 32'hFFFFF1BC , 32'hFFFEA633 , 32'h00009D6E , 32'hFFFF3CCF , 32'hFFFE39AF , 32'h0001A849 , 32'hFFFEB294} , 
{32'hFFFCAFB4 , 32'h00028691 , 32'hFFFDD2F2 , 32'h00015921 , 32'hFFFD0B72 , 32'hFFFF9B4F , 32'h00001EE9 , 32'h0001C953 , 32'h00027B2C , 32'h0004D1A5 , 32'h00000A9E , 32'h00023AA7 , 32'hFFFEAB4E , 32'h0004F81B , 32'h0003718C , 32'hFFFFA133 , 32'h000078BB , 32'hFFFD6297 , 32'hFFFEEF62 , 32'h0004B5B6 , 32'hFFFEE01B , 32'h00031D8E , 32'hFFFEBCE7 , 32'hFFFDB5C3 , 32'h0000423C , 32'hFFFBAB07 , 32'hFFFCC3F8 , 32'hFFFC20A2 , 32'hFFFCEF8C , 32'h00022A5B , 32'hFFFBDE19 , 32'hFFFF6949 , 32'hFFFB0C41 , 32'h00015A77 , 32'hFFFDA90A , 32'h00008E8B , 32'hFFFEC8C3 , 32'h00009076 , 32'hFFFDBF7B , 32'h00004F1D , 32'h00023B15 , 32'h00007814 , 32'hFFFCBCF4 , 32'h0002E424 , 32'hFFFE83F5 , 32'hFFFDE52C , 32'h00018DED , 32'h00041326 , 32'h0000EEF7 , 32'h0005B482 , 32'h0002B1F4 , 32'hFFF7DAFE , 32'hFFFF30D9 , 32'hFFF9489C , 32'hFFFD5294 , 32'h000517F5 , 32'hFFFF255E , 32'h000242F4 , 32'hFFFC7976 , 32'h00013EB0 , 32'hFFFF5BA5 , 32'hFFFDF2F5 , 32'h00038202 , 32'hFFFF0F7C , 32'hFFFE4131 , 32'hFFFD7649 , 32'hFFFBFB91 , 32'h000200A7 , 32'hFFFFA562 , 32'h0002B00D , 32'h0002D7E1 , 32'h00048842 , 32'h0000C53C , 32'hFFFDD673 , 32'hFFFE8454 , 32'hFFFB4118 , 32'h000196CE , 32'hFFFFDF33 , 32'hFFFDCF6E , 32'hFFFD476A , 32'hFFFC50E9 , 32'h00032223 , 32'h00055E9A , 32'hFFFF5047 , 32'h00013468 , 32'hFFFF214E , 32'hFFFD6EE8 , 32'hFFFFDF91 , 32'hFFFD312A , 32'hFFFC0B6F , 32'hFFFE6592 , 32'h00035E1C , 32'hFFFA66DC , 32'hFFFD41CD , 32'h00018803 , 32'h000131C9 , 32'h00018F20 , 32'h0001201F , 32'h00002F27 , 32'hFFFCC587} , 
{32'h0002C0E8 , 32'h00027BA9 , 32'hFFFC0B91 , 32'hFFFE649A , 32'hFFFA2B56 , 32'hFFFF92DF , 32'h000135D2 , 32'hFFFB2004 , 32'h00019142 , 32'h0002FDC9 , 32'hFFFDDFFB , 32'h0005B103 , 32'h00037CB6 , 32'hFFFF04CF , 32'hFFFD7926 , 32'hFFFDE1BC , 32'h0001E0EA , 32'hFFFEF176 , 32'h0001E207 , 32'h0001C02C , 32'hFFFE0147 , 32'hFFFEE4BE , 32'hFFFF1D98 , 32'hFFF978D8 , 32'hFFFF16E5 , 32'hFFFE594A , 32'hFFFBC8EE , 32'hFFFFA063 , 32'h0003A9FA , 32'hFFFF7D8F , 32'h0002ADD0 , 32'h00036E26 , 32'hFFFDAB50 , 32'h0004BBFF , 32'hFFFC983D , 32'hFFFB5B42 , 32'h0000A5DE , 32'hFFFFA355 , 32'h0002D8F0 , 32'h00028CDD , 32'h00005C47 , 32'h00022900 , 32'hFFFFEAD6 , 32'h00055505 , 32'h00027EEF , 32'h00017E7C , 32'h0000884D , 32'h0000E656 , 32'hFFFA9B4E , 32'h0000C054 , 32'hFFFD0ADF , 32'h00021744 , 32'h0001535D , 32'hFFFC56C9 , 32'hFFFE29A0 , 32'h000242C6 , 32'h0002E681 , 32'h00011596 , 32'h00041A88 , 32'hFFFD2350 , 32'hFFFD4101 , 32'hFFFFE4A8 , 32'h00007BA6 , 32'hFFFE9017 , 32'hFFFF4ED5 , 32'hFFFFAB8B , 32'hFFFD981B , 32'hFFFEC0AD , 32'h0001040A , 32'hFFFFBC8E , 32'hFFFD1EB0 , 32'hFFFFBA81 , 32'h00076EDA , 32'h000084E0 , 32'h0002D341 , 32'h000012DE , 32'hFFFDEE50 , 32'hFFFCB8F1 , 32'hFFFEE52E , 32'hFFFE2A47 , 32'h00018B81 , 32'h0002C41D , 32'h0002B5BC , 32'h00024B98 , 32'hFFFCA473 , 32'h00014CB9 , 32'hFFFFDB6F , 32'h0001445B , 32'hFFFFB598 , 32'hFFFCD95F , 32'hFFFF011E , 32'h0000870B , 32'hFFFD6F1C , 32'h0000D210 , 32'hFFFEBC4C , 32'hFFFDA977 , 32'hFFFC95E4 , 32'h000008AB , 32'h0000C3D6 , 32'hFFFDC551} , 
{32'hCE684180 , 32'h13AA4B80 , 32'h19647620 , 32'hFF63DE8C , 32'h06404BA0 , 32'h13219960 , 32'hF83A2DB0 , 32'hF5489930 , 32'hDDC81940 , 32'h02716928 , 32'hEE930240 , 32'hE7FAF5A0 , 32'h0724D540 , 32'h22C3C540 , 32'h00F0870E , 32'h03C3C8D8 , 32'hF997A990 , 32'hFDEF6DC4 , 32'hFA148DB8 , 32'h0FD196D0 , 32'h0C5D53A0 , 32'h051CD3B8 , 32'hFF1310BC , 32'h0A4FAA80 , 32'h03B73448 , 32'hE99E6BC0 , 32'hF00DE050 , 32'hF4B92B80 , 32'h0266CEB0 , 32'h02F2D6A8 , 32'hFA2BB808 , 32'hF0D928D0 , 32'hEE939960 , 32'h043B90D8 , 32'hF18F36F0 , 32'h0A6F4030 , 32'h0B610510 , 32'hF0118070 , 32'hF77DB950 , 32'hF291D9B0 , 32'h06857D40 , 32'h0EF1A850 , 32'h07AE0B88 , 32'h065C4540 , 32'h06B11320 , 32'hF73E7D80 , 32'h0266E23C , 32'hF09A0370 , 32'h046019F0 , 32'h088A2860 , 32'h00B55068 , 32'h0FAD2780 , 32'hFEA29124 , 32'h02F488D4 , 32'h026B9DFC , 32'hFDF40EB4 , 32'hFFF16267 , 32'h015C500C , 32'h076166A8 , 32'hFCB6DCBC , 32'hFCB54AB8 , 32'hFCAD1C70 , 32'hF83A0E60 , 32'hF9E22E68 , 32'hF993F488 , 32'h0389B018 , 32'h0045267D , 32'hFE15EAE0 , 32'hFA07BE80 , 32'h03936544 , 32'hF743BC60 , 32'h04CD15F8 , 32'h07CF7700 , 32'hFF4F3F72 , 32'hFDAE3410 , 32'h04D30430 , 32'h065EE958 , 32'h0518EF60 , 32'h0626EC68 , 32'hFF52595D , 32'h01411970 , 32'hF902A858 , 32'h00A369E7 , 32'h031DFE58 , 32'hFBE64AF8 , 32'h00A02D8C , 32'h002E31BF , 32'h03A01C6C , 32'h005B9F7B , 32'h00E2F0DA , 32'h0001A0BC , 32'hFFFF96D2 , 32'hFFFF4F17 , 32'h00035DE1 , 32'hFFFFFCC1 , 32'hFFFFA4D8 , 32'h0000FEED , 32'h0001F257 , 32'hFFFDDDDA , 32'h000056A1} , 
{32'h000351CC , 32'h0001CBD8 , 32'h0000A7F3 , 32'hFFFE2D97 , 32'hFFFD0D7A , 32'h00040471 , 32'h0001E2C0 , 32'h0001E845 , 32'hFFFE37AD , 32'hFFFD0F18 , 32'h0003818B , 32'hFFFF86A9 , 32'hFFFFA593 , 32'h000157FE , 32'hFFFF732C , 32'h0003EADB , 32'h00024E3E , 32'hFFFFB7E7 , 32'hFFFDFCC4 , 32'hFFFCCFE3 , 32'h00014427 , 32'h00011C48 , 32'h00025E89 , 32'h000161A7 , 32'h000043AC , 32'h00051A4F , 32'h0003EDB9 , 32'h0004304E , 32'hFFFD41E1 , 32'h000485E2 , 32'hFFF90E00 , 32'h0001DC0B , 32'h0000F740 , 32'hFFFF4350 , 32'hFFFE8A48 , 32'h000446DC , 32'hFFFE2A4C , 32'hFFFD7540 , 32'hFFFF2CE0 , 32'h00014243 , 32'hFFFEBAAB , 32'hFFFCDD9D , 32'h00009472 , 32'h0003C8AE , 32'hFFFE7153 , 32'hFFFECC6C , 32'hFFFEE562 , 32'hFFFD48A6 , 32'h000187AD , 32'hFFFFEA80 , 32'h00033D26 , 32'h0001DE09 , 32'h0004D558 , 32'h0001F306 , 32'h00012FF4 , 32'hFFFD2EC2 , 32'hFFFD2969 , 32'h0005D55E , 32'hFFFE7E00 , 32'hFFFEA0D0 , 32'h00012ECE , 32'hFFFE3207 , 32'h000290EC , 32'hFFFC4CCF , 32'hFFFDA431 , 32'hFFFD9E6F , 32'hFFFCC499 , 32'hFFFDEAB9 , 32'h0002E049 , 32'h0005972A , 32'hFFFF1A6F , 32'h00011D59 , 32'h000051DD , 32'h000044B1 , 32'hFFFF430F , 32'hFFFE5771 , 32'hFFFC92BF , 32'h00000075 , 32'h0001F6E3 , 32'h00012049 , 32'h000434E4 , 32'hFFFEDE74 , 32'h00006905 , 32'h00013711 , 32'h00051B09 , 32'hFFFE70CC , 32'hFFFC3B94 , 32'hFFFCCBB5 , 32'h0003077A , 32'hFFFCDC31 , 32'h00009B89 , 32'h000309E1 , 32'h00045108 , 32'hFFFFD1DE , 32'hFFFE2DA4 , 32'h0000B86D , 32'hFFFC2980 , 32'hFFFD3444 , 32'h0003229C , 32'h0002DB9B} , 
{32'h33CAEB00 , 32'h04319538 , 32'hF7687B20 , 32'h1C5805C0 , 32'h193E2DC0 , 32'h093AB510 , 32'hF82826C0 , 32'hEDE557E0 , 32'hEC3974A0 , 32'h068F4710 , 32'hF09CFED0 , 32'h14663AE0 , 32'h1AA7DDA0 , 32'h09A11280 , 32'h11B52520 , 32'hFEB2701C , 32'h06106810 , 32'hFF89AF8A , 32'hF11B6890 , 32'h0B350920 , 32'hFF9571F3 , 32'hF4D15C40 , 32'hEB76F840 , 32'hEB7EBAA0 , 32'hF9BC7A98 , 32'hF0307000 , 32'hFE068DC0 , 32'hEB018EA0 , 32'h1EFA4560 , 32'hFBECAD28 , 32'h1AD56460 , 32'h0B276A20 , 32'h0C03C530 , 32'hFEFDCF6C , 32'hE7A28AE0 , 32'hF0586730 , 32'hEC7D8FE0 , 32'hFB3D19F8 , 32'hF3C0D4E0 , 32'h01807790 , 32'h0047137D , 32'hFC7E34AC , 32'hF43B43B0 , 32'hFC02E80C , 32'hEC4395A0 , 32'h0562EEC0 , 32'h0317D260 , 32'hF6B7FD00 , 32'hF6916D50 , 32'h0029900F , 32'h04E6B860 , 32'h0218AE24 , 32'h08109AD0 , 32'h07695970 , 32'hFA0C3958 , 32'h05F35CD0 , 32'hF8671380 , 32'h043FB938 , 32'hFF75E8DE , 32'hFEB5ECD8 , 32'hF6A231E0 , 32'hFD1AF32C , 32'hFC996554 , 32'h078F6420 , 32'h081AA430 , 32'h07740E58 , 32'hFFE1105E , 32'h07A1D858 , 32'h01D750FC , 32'h02584E68 , 32'h0889E850 , 32'h083C6520 , 32'hFEE9FD0C , 32'hFD4E4424 , 32'h00053634 , 32'hFFA568B9 , 32'hFFF08051 , 32'h00A54B90 , 32'h00739322 , 32'h0339A004 , 32'hFBD50A80 , 32'hFFFC6147 , 32'hFC913434 , 32'h04A28688 , 32'h013AF258 , 32'h00ACFC53 , 32'hFEB5420C , 32'hFE1825E0 , 32'hFE2CC5BC , 32'hFFFDFD7E , 32'h0003249B , 32'hFFFF06BD , 32'hFFFF4B83 , 32'h00019974 , 32'h0000FF61 , 32'h00005764 , 32'h00008C15 , 32'h0002A53F , 32'h000046E3 , 32'hFFFF979D} , 
{32'h000316C3 , 32'hFFFE4785 , 32'h00005425 , 32'hFFFF7C49 , 32'h00002C6F , 32'hFFFD5082 , 32'h0000C5E7 , 32'hFFFF7D77 , 32'h000011E7 , 32'h00011A5B , 32'hFFFF5CE3 , 32'h0000EE5D , 32'hFFFDFC0E , 32'h00044F50 , 32'h0001CDF7 , 32'h00051EB5 , 32'hFFFDE956 , 32'h000321AD , 32'h0003212D , 32'hFFFF4986 , 32'h000127E2 , 32'hFFFED035 , 32'h000182B0 , 32'h000362C2 , 32'hFFFA9F79 , 32'h0000B080 , 32'h000026A3 , 32'h00039274 , 32'h00010950 , 32'hFFFC294D , 32'h00014C98 , 32'hFFFA623C , 32'h0003669C , 32'h00014200 , 32'h0000788F , 32'h0007CB57 , 32'h000196D9 , 32'h00031EC8 , 32'hFFFC15A2 , 32'hFFFE3243 , 32'h00033040 , 32'hFFFF5C8D , 32'h0000058C , 32'hFFFCE22D , 32'hFFFD29E1 , 32'h0004CF70 , 32'h000366EC , 32'h00013871 , 32'hFFFC9D0B , 32'h0000634E , 32'h000023A7 , 32'hFFFB6509 , 32'h00003274 , 32'hFFFFCBCB , 32'hFFFCC4AC , 32'hFFFFD9EF , 32'h000424DA , 32'hFFFF728D , 32'h0002811F , 32'hFFFB345A , 32'hFFFACA40 , 32'h0001D406 , 32'hFFFD3474 , 32'hFFFD0AB3 , 32'h0000E2C8 , 32'h0004A7BE , 32'h0001A755 , 32'hFFF7B51B , 32'h00042E50 , 32'h0003FBEC , 32'h000174B8 , 32'h0000350F , 32'hFFFEB057 , 32'hFFFDCD3F , 32'hFFFECF6E , 32'h00001AC3 , 32'h0003824E , 32'hFFFFCC67 , 32'hFFFED4D4 , 32'hFFF8F2DB , 32'h00025F7D , 32'h0000C5D6 , 32'hFFFF6410 , 32'h0001B24B , 32'h0003BC0C , 32'hFFFD9E44 , 32'h0005413A , 32'h00006283 , 32'h0000B161 , 32'hFFFF8BD1 , 32'h000088FC , 32'h0001841C , 32'hFFFD4697 , 32'h0000C6AE , 32'hFFFEBB5C , 32'h0004DFC8 , 32'h00040BDF , 32'h000053D5 , 32'h0005C005 , 32'h00005713} , 
{32'hFF761237 , 32'h0317A6B8 , 32'hFFD8845A , 32'h025E0E50 , 32'hFE35AE18 , 32'h062DE460 , 32'hFE9A6148 , 32'h04BB3970 , 32'h00DADEE3 , 32'hFDA2BA24 , 32'h05D61308 , 32'h0302BD78 , 32'h066E1010 , 32'h039790A0 , 32'hFFADAC09 , 32'h03B5708C , 32'h02D4FBFC , 32'hFE08F7AC , 32'hFD620700 , 32'h03E4F1C4 , 32'hFE4FCC44 , 32'h02310E24 , 32'h0399F6C4 , 32'h01D4884C , 32'h05E58248 , 32'hFCE9AEB8 , 32'h02D23C2C , 32'h050074C0 , 32'hFF7ECAC9 , 32'hFE1D67BC , 32'hFCB91EBC , 32'h01D3D44C , 32'h016782BC , 32'hF8F1A258 , 32'hFECF41A4 , 32'h014E16FC , 32'h02F1BBD8 , 32'h00D94ED1 , 32'h03B18DB4 , 32'h02803044 , 32'h00F17E8B , 32'hFEA99218 , 32'hFF246119 , 32'hFC9B4CC0 , 32'h005C41E7 , 32'h0285E25C , 32'hFFE0737B , 32'h02A293F4 , 32'hFF9F1CD8 , 32'h023B8580 , 32'hFD008250 , 32'hFE93ABD8 , 32'h0291ED1C , 32'h01D8F9BC , 32'hFE1D345C , 32'h04366F20 , 32'hFEF85FE8 , 32'h00BA9283 , 32'h00803B4F , 32'hFBE14F10 , 32'hFBEA7120 , 32'h021A2748 , 32'h01EF27CC , 32'h02F2C098 , 32'h03ACA604 , 32'h01E306A8 , 32'hFF72AEDA , 32'hFD49ECBC , 32'h03B481DC , 32'h01789ECC , 32'hFE9B0D34 , 32'h016CCA24 , 32'hFF6B7DBF , 32'hFB1FB4B8 , 32'hFE405360 , 32'hFFC36E63 , 32'h01A244C0 , 32'h00266B67 , 32'hFF58711B , 32'hFF29E895 , 32'h0251EBB8 , 32'hFC69EEB8 , 32'h0285AA10 , 32'h002BC6CC , 32'h03684630 , 32'hFF18BD6B , 32'hFFCF1AA4 , 32'hFF12C5F1 , 32'h00523991 , 32'h004E087C , 32'hFFFDA856 , 32'hFFFEF9FC , 32'hFFFF6AA8 , 32'hFFFEACAB , 32'h0000BF93 , 32'h00036902 , 32'hFFFCEAD3 , 32'h0002CF25 , 32'hFFFFE437 , 32'hFFFDF8A7} , 
{32'h00007910 , 32'hFFFBF49D , 32'hFFFBBF00 , 32'h00033676 , 32'h0001C890 , 32'hFFFE1746 , 32'h00045599 , 32'h00003744 , 32'h00009F44 , 32'hFFFDF9EC , 32'h000040A6 , 32'h00053E33 , 32'hFFFF73FD , 32'h00012EE9 , 32'hFFFF37E1 , 32'h0000FCD6 , 32'h0002EB02 , 32'hFFFF097E , 32'hFFFD9327 , 32'h000158D8 , 32'h00004865 , 32'h000112F2 , 32'h0001B5D3 , 32'hFFFF9909 , 32'h00028E19 , 32'hFFFDE4A0 , 32'hFFFF9658 , 32'h000380B0 , 32'h00032E66 , 32'h000234FF , 32'h00012381 , 32'hFFFC6FC4 , 32'hFFFC0A5E , 32'h00030351 , 32'hFFFB7511 , 32'h00018FA8 , 32'hFFFF808C , 32'hFFFC169E , 32'hFFFFE5F9 , 32'h0001A86A , 32'hFFFA84A8 , 32'h00025180 , 32'hFFFDBE9F , 32'h000404DE , 32'hFFFE4E53 , 32'hFFFDF54D , 32'hFFFCBDBC , 32'hFFFDB9CB , 32'hFFFDE14F , 32'h0000BE1F , 32'hFFFFB9ED , 32'h000435EC , 32'hFFFFE76D , 32'h00062D91 , 32'hFFFEBA24 , 32'hFFFEA673 , 32'h0002776D , 32'hFFFF7DE4 , 32'hFFFE93A9 , 32'hFFFFCF34 , 32'hFFFF9DED , 32'h00035814 , 32'hFFFF14A7 , 32'hFFFFC6A0 , 32'h000330CB , 32'hFFFEE312 , 32'hFFFF7D70 , 32'hFFFF36D6 , 32'hFFFE3C3A , 32'h0002D46D , 32'h0000090C , 32'hFFFCD165 , 32'h0000E842 , 32'hFFFFD711 , 32'hFFFCA817 , 32'h00019B21 , 32'hFFFC9D42 , 32'h0001315E , 32'h00025102 , 32'h0005C832 , 32'hFFFB1355 , 32'h0001AEE3 , 32'h0001D496 , 32'hFFFF8E74 , 32'h0005CE44 , 32'h000296C6 , 32'h0000B143 , 32'hFFF9CEA0 , 32'hFFF9CC7F , 32'hFFFCC55A , 32'hFFFF423A , 32'h00057E7D , 32'hFFFE2A5A , 32'h00011E24 , 32'h0001DAEF , 32'hFFFF0B4E , 32'h00002121 , 32'h0001BEAE , 32'h00020D0E , 32'hFFFEBA4F} , 
{32'h21A8AE80 , 32'h3474E100 , 32'hE52B4820 , 32'hED246DE0 , 32'hFDAAF748 , 32'hFD59011C , 32'hFF280205 , 32'h0B25E670 , 32'h1418C620 , 32'hFBCA99D8 , 32'hF756BB90 , 32'h087CC200 , 32'hEE90E4C0 , 32'hED373A20 , 32'hE51685E0 , 32'hF1C2FD90 , 32'h039A87E0 , 32'hF2F70CA0 , 32'h05C5B748 , 32'hF98B2E28 , 32'h06FC7E58 , 32'h10CE6980 , 32'hF56134E0 , 32'h0562F270 , 32'hF95F3910 , 32'h06297938 , 32'hEC499B00 , 32'hFEC18F90 , 32'h00D4AFCD , 32'hFBC9DFC0 , 32'h0558EAC0 , 32'hF3B7B480 , 32'h00489D3E , 32'hF24E1CC0 , 32'h00EFEFD4 , 32'hFA355AB8 , 32'hF2BF8780 , 32'hF00EB9A0 , 32'h08363D70 , 32'hFBE971A0 , 32'hF70F4DD0 , 32'h07A8EEB0 , 32'hFFF748BA , 32'h149B4160 , 32'h02C28D28 , 32'h0621FFA8 , 32'hFD250A08 , 32'h04F95FE0 , 32'hFDB0B348 , 32'h059094D8 , 32'hF9D80EB0 , 32'h0BE603A0 , 32'h00FB2485 , 32'hF7C01D10 , 32'h0563B3D0 , 32'hFE35C2A8 , 32'hFBAC73A8 , 32'hFBFC3068 , 32'hFEA0C310 , 32'hFFB5C552 , 32'hFE2D0604 , 32'hF743A590 , 32'h025F077C , 32'h0B85CDD0 , 32'h049EDF28 , 32'h01AB87C8 , 32'hF9144A10 , 32'h01FDD7B4 , 32'hFE8FB138 , 32'hFEB758F8 , 32'hFF80A280 , 32'hFD4CAC54 , 32'hFB8DED80 , 32'h01282374 , 32'h0244DFE8 , 32'h07A208C8 , 32'h01F0D31C , 32'h008E142D , 32'h02F09C4C , 32'hFB75EC78 , 32'hFFA6C2EE , 32'h0519E270 , 32'h01712E88 , 32'h037DD498 , 32'hFDCF7C9C , 32'h022E9E74 , 32'h048A79D0 , 32'hFE753214 , 32'h010491B0 , 32'h000FDA6D , 32'hFFFEB580 , 32'hFFFFEBFC , 32'h00010905 , 32'hFFFD05E5 , 32'hFFFF40E5 , 32'h0001726E , 32'hFFFFAA28 , 32'hFFFCD315 , 32'h00016406 , 32'hFFFEFC7A} , 
{32'h000029BD , 32'h00007042 , 32'h0002DA46 , 32'h00016435 , 32'hFFFD31F9 , 32'h0001F9F3 , 32'hFFFF13DF , 32'hFFFE8E67 , 32'h00023E39 , 32'h0004F5D9 , 32'hFFFEA746 , 32'hFFFD3D8A , 32'hFFFEC1C2 , 32'hFFFDE566 , 32'hFFFFB17F , 32'h00002EC9 , 32'h0003DB47 , 32'hFFFF2948 , 32'hFFFFD524 , 32'h0001E2A0 , 32'hFFFF62C9 , 32'h00001ABB , 32'hFFFF1155 , 32'h0003D7D7 , 32'hFFFD59C4 , 32'hFFFF8462 , 32'hFFF99692 , 32'h0002715A , 32'hFFFF25D2 , 32'h00027BB3 , 32'h000197B5 , 32'hFFFE6C89 , 32'h0002F543 , 32'h0003E4EB , 32'h00042761 , 32'hFFFEAD90 , 32'h000497AF , 32'h00036B0E , 32'hFFFD7F0C , 32'h0000C139 , 32'hFFFDBFFD , 32'hFFFF04CC , 32'hFFFCDEE5 , 32'hFFFF763C , 32'h000027E6 , 32'h0001B18C , 32'h00032307 , 32'hFFFECBA2 , 32'hFFFE5E46 , 32'h0004937D , 32'hFFFF0C4C , 32'h0002343B , 32'hFFFE3D7B , 32'hFFFEEFFE , 32'h000175C3 , 32'hFFFC0830 , 32'h0003FF18 , 32'hFFFD0167 , 32'h0004E244 , 32'hFFFF84E2 , 32'hFFFFBFF4 , 32'hFFFD9EB2 , 32'h000389EC , 32'hFFFB3460 , 32'h00008B95 , 32'hFFFD9947 , 32'hFFFF5950 , 32'h0000422F , 32'hFFFFDA8B , 32'h00044294 , 32'hFFFEA512 , 32'h00017866 , 32'h000079B4 , 32'hFFFCDB29 , 32'h00040FF6 , 32'hFFFB286F , 32'hFFFE3762 , 32'h0000A9ED , 32'h00004DFB , 32'h00016342 , 32'hFFFB27E1 , 32'hFFFE23EE , 32'h00052B51 , 32'hFFFB79E7 , 32'h0003110E , 32'hFFFC61A3 , 32'h0004705B , 32'h0000F6B6 , 32'h00008881 , 32'h0000D575 , 32'hFFFE1F3E , 32'hFFFE27D4 , 32'h00024492 , 32'hFFFF0260 , 32'h0000CE56 , 32'h00050C5A , 32'hFFFDBBC9 , 32'hFFFDBAC7 , 32'h0000618C , 32'hFFFC66BC} , 
{32'h0001B8EF , 32'hFFFDF52D , 32'hFFFE4E7E , 32'hFFFB56F8 , 32'hFFFD7326 , 32'h0001DDDF , 32'h0001C2EC , 32'hFFFC56E5 , 32'hFFFD6FCC , 32'hFFFDB361 , 32'hFFFB68DD , 32'hFFFDD158 , 32'hFFFFEC83 , 32'h00008117 , 32'hFFFD74BE , 32'h0000EB3A , 32'h000060A2 , 32'hFFFECABE , 32'hFFF7CFFD , 32'h000116D8 , 32'h00044B64 , 32'h0001738F , 32'h0002AD49 , 32'hFFFC254A , 32'hFFFE9AE8 , 32'h0000E107 , 32'hFFFC00ED , 32'h0000603B , 32'hFFFC5751 , 32'h0004572C , 32'h0003B825 , 32'hFFFD3A5E , 32'h00011AC4 , 32'hFFFFEEC1 , 32'hFFFC6FA5 , 32'h00017491 , 32'h000469C0 , 32'h0001C550 , 32'h0001D550 , 32'hFFFFB791 , 32'hFFFEFD55 , 32'hFFFDE24B , 32'h0002A1AA , 32'h00023713 , 32'hFFFED050 , 32'hFFFF5BE3 , 32'hFFFECE11 , 32'hFFFD810F , 32'h00001380 , 32'hFFFEDB99 , 32'hFFFCCD08 , 32'hFFFF13D3 , 32'hFFFE5657 , 32'hFFFC9609 , 32'h00029475 , 32'h0001D564 , 32'hFFFE637A , 32'h00051333 , 32'hFFFEE51F , 32'hFFFD5808 , 32'hFFFB46DA , 32'h000265C7 , 32'hFFFF75D7 , 32'h0000EBC1 , 32'hFFFD7FDD , 32'hFFFE7100 , 32'h000192A2 , 32'h0002215E , 32'h000359F6 , 32'hFFFAAFA5 , 32'hFFFF2CBA , 32'h00001934 , 32'hFFFB2D95 , 32'hFFF9D07C , 32'h00028B1D , 32'h00013D84 , 32'h000363E3 , 32'hFFFA4CDB , 32'hFFFF07EE , 32'h0001F5A5 , 32'h000324F5 , 32'hFFFFCC45 , 32'h0001EA98 , 32'hFFFE55DA , 32'hFFFCE01A , 32'hFFFEDE51 , 32'hFFFE5779 , 32'h0001F1AD , 32'hFFFE6583 , 32'hFFFC2DD3 , 32'h0002D13F , 32'h00039322 , 32'hFFFABD87 , 32'hFFFEDE7D , 32'h00066EEA , 32'hFFFEACE5 , 32'h0002C284 , 32'hFFFD7632 , 32'h00004A4D , 32'h00016F01} , 
{32'hFFFD285D , 32'hFFFFD6AB , 32'h000181F7 , 32'hFFFF2A44 , 32'h0001E8A1 , 32'hFFFE15AD , 32'h00005C05 , 32'h0001321F , 32'hFFFE5995 , 32'h00006689 , 32'h00020F6D , 32'hFFFFF916 , 32'h00033D06 , 32'h0001682B , 32'h00009505 , 32'h00024231 , 32'h00011227 , 32'hFFFE06C6 , 32'h0005DD04 , 32'hFFFF7D7A , 32'h00000587 , 32'hFFFE110C , 32'h0000689E , 32'hFFFFF804 , 32'hFFFD6939 , 32'h0000C34A , 32'hFFFE62B3 , 32'hFFFCF850 , 32'h00063262 , 32'h0001B4C2 , 32'hFFFDF82F , 32'h0003B172 , 32'h00005103 , 32'hFFFECC8B , 32'h00020629 , 32'h0002410B , 32'h00059924 , 32'hFFFBF3F2 , 32'h0005C946 , 32'hFFFF2B61 , 32'hFFFDDC00 , 32'hFFFE5B56 , 32'h0002121D , 32'h0004F480 , 32'h000235A4 , 32'hFFFEF81E , 32'h00019D02 , 32'h0001B8A9 , 32'h0002293D , 32'hFFFB38F2 , 32'h00024EA8 , 32'hFFFE1233 , 32'hFFFF6000 , 32'hFFF9BD7E , 32'h0003067A , 32'h0003255B , 32'h00009599 , 32'hFFFB7EA4 , 32'hFFFBDA2B , 32'hFFFCC80B , 32'h0001D028 , 32'hFFFD3ACC , 32'hFFFFB19D , 32'h0004ADB9 , 32'hFFFEED4D , 32'h000257DB , 32'hFFFD868A , 32'h00003D07 , 32'h0000A480 , 32'hFFFF8407 , 32'hFFFB7D1A , 32'h0000401E , 32'h0001DC69 , 32'hFFFFF82B , 32'h00004C4B , 32'hFFFFD672 , 32'h0002CB87 , 32'h0000CEDC , 32'h0002BDBD , 32'h000191BC , 32'h00038301 , 32'hFFFFDEAF , 32'h00016F40 , 32'h0003E4BE , 32'h0001D0B7 , 32'hFFFDFA51 , 32'hFFFD6B1B , 32'hFFFF0845 , 32'h0000A0F8 , 32'h0000EC11 , 32'hFFFB002B , 32'hFFFB8B58 , 32'hFFFD2A03 , 32'hFFFBB886 , 32'hFFFFB45A , 32'h0003ECDA , 32'h00000859 , 32'h00021A44 , 32'hFFFCDB98 , 32'h0001178D} , 
{32'hF9166250 , 32'hFDAA5EDC , 32'hE0D12940 , 32'hE4A812E0 , 32'hD1C5D680 , 32'hF1B5C9E0 , 32'h090DBB10 , 32'h0050F27B , 32'hE3497DC0 , 32'h18D7F640 , 32'h07B11E20 , 32'h06B72F28 , 32'h06A20228 , 32'hF8D5AD98 , 32'hF2EBB890 , 32'h227B4CC0 , 32'h0BC7B500 , 32'h09CABA90 , 32'hE6535DC0 , 32'h19443EA0 , 32'hEA77B9C0 , 32'hFD790F1C , 32'h05DBC9E0 , 32'hF231D7B0 , 32'hF6FE7820 , 32'hF9E35A60 , 32'hF13D81D0 , 32'h07E1BAF8 , 32'hFDC777CC , 32'h021381A8 , 32'hEE69D800 , 32'h0235A414 , 32'h02817ABC , 32'h0C214D50 , 32'h06515F90 , 32'hE70EC4C0 , 32'hF7046940 , 32'hFBF7EA88 , 32'h015FACB4 , 32'hFB583DF0 , 32'h0374C7F0 , 32'h129D2560 , 32'hFE53CED8 , 32'hF5B9FC80 , 32'hFFC098A3 , 32'hFEC0549C , 32'h0B24D4C0 , 32'hF90296B0 , 32'h02048908 , 32'h0176BF7C , 32'hF67F5CC0 , 32'hFF4E2B4E , 32'h000CA055 , 32'h07C0D280 , 32'h028A5F48 , 32'hFE42D6D8 , 32'h04641320 , 32'hFBCD2128 , 32'h000894C1 , 32'hFF094B55 , 32'hFB3B04D0 , 32'hFAD047C8 , 32'h03DD2FAC , 32'h014EC7B4 , 32'h04BF3278 , 32'hFD7C54B0 , 32'hFF5832D1 , 32'h002BEF38 , 32'hFCB941C8 , 32'hFD636D58 , 32'hFC995E78 , 32'hFB9E95F0 , 32'hFFC141AB , 32'hFA85CF78 , 32'h05C2B070 , 32'h0622DBC8 , 32'hFE4E79A8 , 32'hFA1B4AE8 , 32'h02E95CAC , 32'hFBA01978 , 32'hFE50A768 , 32'h003BA698 , 32'hFBD98178 , 32'h015E9ED4 , 32'hF9C739F8 , 32'hFEF0C634 , 32'hFBBB85D0 , 32'hFDC3C3CC , 32'hFD5CE5CC , 32'h00C38606 , 32'h000045B9 , 32'hFFFF710B , 32'h00014CC2 , 32'hFFFE217C , 32'h00001BDC , 32'hFFFF7949 , 32'hFFFE26CB , 32'h00018636 , 32'hFFFF3626 , 32'hFFFFF432} , 
{32'hDF980D80 , 32'h080BF720 , 32'hF68234E0 , 32'h29C25AC0 , 32'h19DA4F00 , 32'hE57B6560 , 32'h13F668A0 , 32'hCD924AC0 , 32'h07893400 , 32'hFB1A9C50 , 32'h004A44CA , 32'hE74924E0 , 32'hD54AA640 , 32'hFE94B2FC , 32'h07A6EFE0 , 32'h0C961EB0 , 32'h0225AF60 , 32'h29764A80 , 32'hFD6C1F08 , 32'h202A4500 , 32'hFFB0890A , 32'h21617A00 , 32'hFF53B0CB , 32'hEDAE92E0 , 32'hF4B1BFE0 , 32'hF3B9A690 , 32'hF55485B0 , 32'h0191A93C , 32'h0C7AB250 , 32'hFA650BA0 , 32'hED5CD520 , 32'h000AD503 , 32'h0136627C , 32'hFB0E2020 , 32'h08B03550 , 32'hFF6AE12D , 32'hF96290F0 , 32'hFB897258 , 32'h01748390 , 32'h095558D0 , 32'h00314BEC , 32'h00B85293 , 32'hF7FBCC40 , 32'h04A0A780 , 32'hFBC670A8 , 32'h028DACE0 , 32'h0899BD90 , 32'hFC616280 , 32'hF9FBB020 , 32'h03C5FCA0 , 32'hFD06C79C , 32'h0B2043E0 , 32'hF652D400 , 32'h04370A18 , 32'h020DBFBC , 32'hF93CCF70 , 32'hFBE097D8 , 32'hF9D62D38 , 32'hFDD167D8 , 32'h01A410FC , 32'h036080F8 , 32'hFAD4F810 , 32'h04690960 , 32'hFA7AD3E0 , 32'hFCAF0074 , 32'hFB9D5B68 , 32'h03F36838 , 32'hF909E7A8 , 32'h061C3A00 , 32'h062B3778 , 32'hFF9C3E19 , 32'hF9584CA8 , 32'hFC2F1920 , 32'h05979D90 , 32'hF7E6B5B0 , 32'hFA308CB8 , 32'hFBB61278 , 32'hFA19BEC0 , 32'hFFE8452E , 32'h027E891C , 32'hFC32EB4C , 32'h0191295C , 32'hFF0BAEC4 , 32'h0548E388 , 32'h008DDFD6 , 32'hFE6F9D54 , 32'h00BDBE53 , 32'hFE778230 , 32'h0156C1D4 , 32'h00052EF1 , 32'h00001646 , 32'hFFFFB30A , 32'hFFFD9727 , 32'h0000CB3F , 32'hFFFCC017 , 32'h00007613 , 32'h00005325 , 32'h00013A6E , 32'h0001EFB9 , 32'h0001FEEB} , 
{32'hFFFF1203 , 32'h0004FAC7 , 32'h00001BD3 , 32'h0000868B , 32'h0007A9D6 , 32'h00022464 , 32'h00000B2C , 32'h00014629 , 32'h0000CDA9 , 32'h00025ED1 , 32'h000201CC , 32'hFFFE3525 , 32'hFFFF4BF6 , 32'hFFFFC861 , 32'h0003F235 , 32'h00008D4B , 32'h00039920 , 32'h000320E4 , 32'h0003AC29 , 32'hFFFB2F51 , 32'h000107FB , 32'hFFF70B32 , 32'hFFFD1089 , 32'h00029140 , 32'hFFFEFE77 , 32'hFFFBB52F , 32'h00032F97 , 32'h0000F995 , 32'hFFFC191F , 32'hFFFE5E8A , 32'hFFFBEE39 , 32'h000774A9 , 32'h000511B3 , 32'hFFFFAC01 , 32'hFFFBF68A , 32'hFFFFF6EF , 32'h0002272B , 32'h000200A0 , 32'hFFFF8786 , 32'h00024644 , 32'hFFFFE66C , 32'hFFFDE476 , 32'hFFFF6772 , 32'hFFFFC117 , 32'h00025DA4 , 32'h000144E0 , 32'hFFFE1EFF , 32'h0000C455 , 32'hFFFEE17B , 32'h00041124 , 32'hFFFAEA58 , 32'h0000E28C , 32'hFFFEC410 , 32'hFFFE6D7A , 32'h00053EF8 , 32'h0000566B , 32'h0000586D , 32'hFFFD8E57 , 32'h0000C13D , 32'hFFFCA9AF , 32'hFFFEA54F , 32'h0002FFF2 , 32'hFFFC03C6 , 32'h0001F8C8 , 32'hFFFEAA3E , 32'hFFF9591C , 32'hFFFF53CE , 32'h00022463 , 32'h00014604 , 32'h0003F797 , 32'hFFFD677F , 32'h0001C23B , 32'hFFFD68AA , 32'h000122BE , 32'h0000BC91 , 32'hFFFF5F2A , 32'h00051865 , 32'h00059342 , 32'hFFFF69F6 , 32'hFFFAB728 , 32'hFFFDC4D8 , 32'h000364B4 , 32'h00007025 , 32'h0002D8F0 , 32'hFFFEDB31 , 32'h00028B71 , 32'hFFFFF069 , 32'h0004432D , 32'h000209D3 , 32'h0003BB16 , 32'h000076DD , 32'h00001A23 , 32'h000075B2 , 32'hFFFE6BEA , 32'hFFFAF600 , 32'hFFFE16DB , 32'hFFFD8AAA , 32'h0001CB8B , 32'hFFFCB669 , 32'hFFFCBED9} , 
{32'hFFFC2C40 , 32'hFFFAFAD7 , 32'h0000737A , 32'hFFFFE884 , 32'h00015961 , 32'hFFFFB6C3 , 32'hFFFF82FB , 32'h00010473 , 32'hFFFE9771 , 32'hFFFC4AF7 , 32'hFFFD14E8 , 32'h000555FC , 32'hFFFDE9A7 , 32'h000074D1 , 32'hFFFEA8C1 , 32'h00034E6A , 32'hFFFFFFB7 , 32'h000251B8 , 32'hFFFDD278 , 32'h000191CA , 32'hFFFF3F57 , 32'hFFFB4518 , 32'h00001539 , 32'hFFFF33CB , 32'h0008FBDB , 32'hFFFE38EF , 32'h00000FD6 , 32'hFFFFFBC4 , 32'h000174E5 , 32'h0000DCB8 , 32'h00017164 , 32'h00021926 , 32'h00010486 , 32'hFFFF78E6 , 32'hFFFC2ACF , 32'h00018D2C , 32'h00030268 , 32'hFFFE38BE , 32'hFFFDE703 , 32'hFFFCB365 , 32'hFFFEF64C , 32'hFFFBA27D , 32'h000085F1 , 32'h0003CE03 , 32'h000728C8 , 32'h00011BF9 , 32'hFFFEE9A6 , 32'h00005ABC , 32'hFFFA9CD7 , 32'hFFFC0B18 , 32'hFFFA1642 , 32'h000015DC , 32'hFFFF6469 , 32'h0004BAB3 , 32'hFFFC6877 , 32'hFFFC578D , 32'h0000CF96 , 32'hFFFC3469 , 32'h0005B088 , 32'hFFFCFC6B , 32'hFFFD7232 , 32'hFFFFA5B5 , 32'hFFFFBDA8 , 32'h0001694C , 32'hFFFDAC7B , 32'hFFFC7682 , 32'hFFFBE6E4 , 32'hFFFEA279 , 32'h0002CBB7 , 32'h00017555 , 32'h00009371 , 32'hFFFFC006 , 32'h00024690 , 32'hFFFF00FB , 32'h0002F6BB , 32'hFFFE80B6 , 32'hFFFD82E4 , 32'hFFF6FEAE , 32'h00022254 , 32'h00014474 , 32'h0001B560 , 32'hFFFE83FE , 32'hFFFA76A6 , 32'h00040E9D , 32'hFFFE1958 , 32'hFFFD2BA5 , 32'h0001F084 , 32'hFFFB17FD , 32'hFFFE36E1 , 32'hFFFF3DE0 , 32'hFFFD0F44 , 32'hFFFAB83F , 32'hFFFB4937 , 32'hFFFD142C , 32'hFFFE9E68 , 32'h00005927 , 32'hFFFD1F09 , 32'h0001E635 , 32'hFFFEF75C , 32'hFFFF1754} , 
{32'h0001DB8D , 32'hFFFF5DFB , 32'h00055E9E , 32'h00005041 , 32'hFFFBE56E , 32'h0002039F , 32'h00003A38 , 32'h0001BDBF , 32'hFFFE7847 , 32'hFFFF9DEA , 32'h0002A474 , 32'h0003F274 , 32'h00017AF8 , 32'h00049884 , 32'h00040641 , 32'hFFFA3CDE , 32'hFFFD692F , 32'hFFFC7B45 , 32'h0000650D , 32'hFFFF884F , 32'h00002A4B , 32'hFFFFFF43 , 32'h00042FA7 , 32'hFFFF878D , 32'hFFFEFD2B , 32'hFFFEC6FA , 32'h00059A51 , 32'h0000398B , 32'h00002ADA , 32'h00027F06 , 32'hFFFF4909 , 32'hFFFECD61 , 32'hFFFF0BBA , 32'h00027A58 , 32'h0005D896 , 32'hFFFB98BD , 32'hFFFAF46B , 32'h0001C5A6 , 32'hFFFD2770 , 32'hFFFDD7C1 , 32'hFFFDCF8E , 32'h0000E2A3 , 32'h0000B86D , 32'hFFFF0A91 , 32'hFFFF414C , 32'h00032F40 , 32'h00020C21 , 32'hFFFA9C81 , 32'hFFFCFCE0 , 32'h0002E422 , 32'hFFFA2BAB , 32'hFFFE0AB5 , 32'h0002C43F , 32'hFFFE7AB3 , 32'h000298F1 , 32'h00063872 , 32'h00010233 , 32'hFFFF9F7F , 32'h0000E9FA , 32'h00020F27 , 32'hFFFDFEDB , 32'hFFFF8BF9 , 32'h0002A6C4 , 32'hFFFFA343 , 32'h0005A117 , 32'hFFFFB3CC , 32'h0001FFD3 , 32'hFFFCB252 , 32'h00001D61 , 32'h00061107 , 32'hFFFFA520 , 32'hFFFB0B9D , 32'h0000AEF5 , 32'h0001A63D , 32'hFFFF2B12 , 32'hFFFF74CD , 32'hFFFF1A17 , 32'h0001B615 , 32'h0000F8DD , 32'hFFFDA97D , 32'hFFFD3D95 , 32'hFFFA303F , 32'hFFFEF89E , 32'hFFFF4DCA , 32'hFFFDDF3D , 32'h00027108 , 32'hFFFF695C , 32'h000256E5 , 32'hFFFFCA7F , 32'hFFFD9DAB , 32'hFFFD3F16 , 32'h0005D2FB , 32'hFFFD38BC , 32'h000416E7 , 32'h0000723B , 32'h0003D7C1 , 32'hFFFD9948 , 32'h00013114 , 32'hFFFF2B5B , 32'h000332CC} , 
{32'hFFFF60BF , 32'hFFFFC745 , 32'h0001ABF5 , 32'hFFFE7636 , 32'hFFFEE063 , 32'hFFFF4AAD , 32'h0004752C , 32'h0002F0C5 , 32'h0000B73E , 32'h00001B6B , 32'h00000C0F , 32'h0000D927 , 32'h0000972E , 32'h00003453 , 32'h00004326 , 32'h00045120 , 32'hFFFD3AB2 , 32'h000221B3 , 32'hFFFE805F , 32'h0001460D , 32'hFFFCEB5A , 32'hFFFDA983 , 32'hFFFE0A08 , 32'h0000FF9E , 32'hFFFD22A4 , 32'h00051873 , 32'h00012DF9 , 32'h0001AD38 , 32'hFFFE8686 , 32'h00024777 , 32'hFFFF1773 , 32'h00028FAB , 32'h00021FDE , 32'hFFFDD84E , 32'hFFFD41E3 , 32'hFFFD3F98 , 32'h00006AD7 , 32'h00006F3F , 32'h000133DC , 32'hFFFA8357 , 32'h0001AAA5 , 32'h000037BC , 32'hFFFEF2FE , 32'h0006CE0F , 32'h0001F495 , 32'hFFFDE4D8 , 32'h00000825 , 32'hFFFDC161 , 32'h0000F712 , 32'hFFFFA223 , 32'h00008D86 , 32'h0001C3D8 , 32'h00043A2C , 32'h000011A4 , 32'hFFFE3A0B , 32'h000207EA , 32'h00023075 , 32'h0003E3C5 , 32'h0000D21B , 32'h00007DBF , 32'hFFFEDAFE , 32'hFFFC96A2 , 32'h00011047 , 32'hFFFF76A5 , 32'hFFFBA776 , 32'hFFFF1B74 , 32'hFFFD4587 , 32'h00005E39 , 32'hFFFF7376 , 32'h0001B84E , 32'h0000ED19 , 32'h00015CCE , 32'hFFFF6718 , 32'hFFFE95B8 , 32'hFFFFA1E5 , 32'hFFFA6A29 , 32'h00003FC2 , 32'h0001099A , 32'h00006245 , 32'h00045297 , 32'hFFFF340B , 32'h0001A705 , 32'hFFFEBA03 , 32'hFFFFFF64 , 32'h00021322 , 32'hFFFEA4D7 , 32'h0003C888 , 32'h00040F3C , 32'h0002E670 , 32'h0001CBCB , 32'hFFFFC2E3 , 32'hFFFF18F8 , 32'h000093B9 , 32'hFFFE7719 , 32'h00024F01 , 32'hFFFCE875 , 32'h00031D22 , 32'hFFFC5A86 , 32'h0000E304 , 32'h00000045} , 
{32'hEA97EC40 , 32'hED691E60 , 32'h225A93C0 , 32'h1DF22160 , 32'h244E57C0 , 32'h24C68040 , 32'h1A3FEEE0 , 32'hF555DF90 , 32'h0ADC6270 , 32'h0CC71870 , 32'hD6989EC0 , 32'hFE63D948 , 32'hFC674D44 , 32'hFD928940 , 32'hE63C0740 , 32'h0568FFE0 , 32'hE5626B40 , 32'hF190B730 , 32'hF82CF1B0 , 32'h129A75E0 , 32'hFD929FA4 , 32'h07330540 , 32'hE4AE7640 , 32'hF4AB3E50 , 32'hF5E237D0 , 32'hFE1C21A0 , 32'hFF6E4F19 , 32'hEAABB340 , 32'hFCFF7498 , 32'h04643438 , 32'h00252128 , 32'hFA85DB58 , 32'hFB708BB8 , 32'h0598EAA0 , 32'h0BE62F50 , 32'h0D5FBE40 , 32'hF940CE30 , 32'h0AF62C90 , 32'h0286DDD0 , 32'h116371A0 , 32'h0E152D60 , 32'hF9E1AF18 , 32'h02565E24 , 32'h090A0D60 , 32'h144B4340 , 32'h02B17BE8 , 32'h0051F374 , 32'hFBC7ADB0 , 32'hFDD80694 , 32'hF44A4DC0 , 32'hF8193CE0 , 32'h003CFB3C , 32'hFB2ADA80 , 32'h0DCBCCD0 , 32'h037427F4 , 32'h004D53C1 , 32'hF94A7CF0 , 32'hFAA6B988 , 32'h049CFC00 , 32'hF7AFCD00 , 32'hF9517A20 , 32'h0BF446A0 , 32'hFDC41AEC , 32'h042BBDE0 , 32'hFB12B630 , 32'h058C8850 , 32'hFE620FA4 , 32'h06555670 , 32'hFE484E80 , 32'hFB60BD48 , 32'h06196380 , 32'hFFAAADAE , 32'h08396E70 , 32'h03F983D8 , 32'h08365AD0 , 32'h043DD738 , 32'hFEFF1298 , 32'hFD38C054 , 32'hFB6D3EA0 , 32'h007B4BFF , 32'hFF21D707 , 32'h03FCF964 , 32'hFDCA6398 , 32'h01E659B8 , 32'h04124298 , 32'h01F85024 , 32'hFDD7C238 , 32'hFDD24D58 , 32'h016D4B74 , 32'h004BCB5B , 32'hFFFD659F , 32'hFFFF28BF , 32'h00016250 , 32'h00008DF7 , 32'h000093FF , 32'hFFFF871B , 32'hFFFD7394 , 32'hFFFF03CB , 32'h000188A0 , 32'h0000C70C} , 
{32'h116AD100 , 32'h0E0C1740 , 32'h24D84200 , 32'h1361E6C0 , 32'hE5FB7460 , 32'hED9F02E0 , 32'hFA54CB18 , 32'hF097EFC0 , 32'hEABC6CE0 , 32'h07DB0D80 , 32'h08C79CA0 , 32'h130812A0 , 32'hEC72F320 , 32'hFB6EB7F8 , 32'hF1FAB150 , 32'hFA8B0E10 , 32'hFD97F288 , 32'hFBD739C8 , 32'hEBEA52E0 , 32'hF9E9D4B0 , 32'h067082E0 , 32'hFD4D6EE4 , 32'h060002B0 , 32'hFB869DF8 , 32'h18F0A1E0 , 32'hFFA58698 , 32'h0514D9C0 , 32'h08AB73D0 , 32'hFB5C9DA0 , 32'h130D9420 , 32'h0B3CD4A0 , 32'h096737A0 , 32'hF7AAB5F0 , 32'h03ED7760 , 32'hF84F6B20 , 32'h0A2E3E00 , 32'hFFA64271 , 32'hF763E040 , 32'h08A2F070 , 32'h024D2F14 , 32'hE5768DC0 , 32'hFF7C6BEC , 32'hFFFBD8FC , 32'hFA794BC8 , 32'h023CD38C , 32'hF91B1F58 , 32'h032A48E0 , 32'hF892A178 , 32'hFB27A410 , 32'hF78167B0 , 32'h05E43450 , 32'h0C4105E0 , 32'h04C66F98 , 32'h125693A0 , 32'hFD170664 , 32'h006DD994 , 32'h03BC702C , 32'hFEA092D4 , 32'hFD067768 , 32'h02BAA0F8 , 32'h1247C0C0 , 32'hFD1A11B8 , 32'h00305CB7 , 32'h06432B50 , 32'hFDD0BD84 , 32'h02C1EF84 , 32'hFAD69CC0 , 32'hFD430E38 , 32'h11C16EE0 , 32'h0477F558 , 32'h0650EAE8 , 32'h00174DDA , 32'hFCBB51EC , 32'hFF49865F , 32'hFBEAECB8 , 32'h04320A38 , 32'hFE7986C4 , 32'hFDB4B818 , 32'h02B30838 , 32'hFD2AEB6C , 32'h02CD5850 , 32'h0435D9C0 , 32'hFCF90C00 , 32'hFE3E1F50 , 32'h0188DBCC , 32'h04809420 , 32'h01F36530 , 32'h03273EA8 , 32'h01A81248 , 32'h00064EC5 , 32'h00004977 , 32'hFFFDDC3F , 32'hFFFFE3EC , 32'h0004582D , 32'h0002D172 , 32'hFFFE8283 , 32'h00006A5F , 32'h000114AD , 32'h00008A79 , 32'hFFFFE4A8} , 
{32'h239EC080 , 32'h0AEFB720 , 32'h2F34E3C0 , 32'hEE11A1A0 , 32'h08E66DB0 , 32'hD6931580 , 32'hD7AF5140 , 32'h03939FB0 , 32'hDFBC8600 , 32'hF80DF688 , 32'h0190F9E8 , 32'hF5B3AC80 , 32'h06509140 , 32'h17A3D300 , 32'hFF885379 , 32'h0A1428C0 , 32'hF3773750 , 32'h025878D4 , 32'h04E649F0 , 32'h053BD300 , 32'hFE4EC6BC , 32'hFDDB7088 , 32'hECCED3C0 , 32'h02458188 , 32'h04D944B8 , 32'hEFC00620 , 32'h0A5C55B0 , 32'h0EC81690 , 32'hE71AD760 , 32'hF8491CE0 , 32'hF6DE4CC0 , 32'h0E40F5E0 , 32'h162DDFE0 , 32'hFD673C18 , 32'h022B4F4C , 32'hF9ADD498 , 32'hED66A7E0 , 32'h01965F00 , 32'hF9BDAEB0 , 32'h037F6250 , 32'hFCBDF39C , 32'h06444E40 , 32'hF1FA4A60 , 32'h157A17E0 , 32'hFECBFE2C , 32'hF9079708 , 32'h045BDE00 , 32'h01FAE7A8 , 32'hF9108098 , 32'hFBB926E0 , 32'h0191546C , 32'h0C1C2CF0 , 32'hFF972009 , 32'hFBBA9AA0 , 32'hF7F55C10 , 32'h070FE5B0 , 32'hFE19AAC8 , 32'h05B820C8 , 32'h06EDA0E0 , 32'h02DE640C , 32'h0BA39210 , 32'hFE59E760 , 32'h01B3FE34 , 32'hFF30B5AC , 32'hFE1F0584 , 32'h023807C4 , 32'hFC0003B8 , 32'hFFC222B4 , 32'h00FB5255 , 32'hFCB43768 , 32'hFF039AE6 , 32'hFE57EFDC , 32'h0278D9C4 , 32'hFAA20FF8 , 32'h06A32260 , 32'hFDABDDC0 , 32'h0172C388 , 32'hFE3954A0 , 32'hFCDA139C , 32'hFE2A0998 , 32'h01C6BB40 , 32'h02BD1890 , 32'hFE5093D8 , 32'h02D7A338 , 32'h011D8F24 , 32'h00BBAD06 , 32'hFF44C1B3 , 32'hFF6EEF8B , 32'h02DE3E6C , 32'hFFDEFCFB , 32'hFFFF30C7 , 32'h0003AB96 , 32'hFFFFE571 , 32'hFFFF7CCA , 32'h000355A3 , 32'h000210A8 , 32'hFFFEE4FA , 32'hFFFEFC2A , 32'h000015E5 , 32'hFFFE7427} , 
{32'hF23D9D40 , 32'hEEEA0C60 , 32'hDE34BB40 , 32'hFEA1D66C , 32'hBEAE6D80 , 32'hF28DB330 , 32'hE663EE20 , 32'hEDE24800 , 32'hE53AA4C0 , 32'hFEE7A474 , 32'hE9495440 , 32'h1DDF29C0 , 32'hEF6089A0 , 32'hEED2BE20 , 32'h0065B7D0 , 32'h0B9206B0 , 32'h10177000 , 32'hF3D2CAA0 , 32'h0DCF9F90 , 32'hEA178260 , 32'hF56EF160 , 32'hE83F3DE0 , 32'h01BE26B0 , 32'hE19571E0 , 32'h0916ED50 , 32'hDD1E1640 , 32'hEDC61500 , 32'h03161948 , 32'hF4287120 , 32'hFBBA1570 , 32'h040DC1F0 , 32'hE8C0BF40 , 32'hFD8798AC , 32'h096FA920 , 32'hFC0C5190 , 32'hF7E8E3F0 , 32'hF9FAAFD8 , 32'hFF42F1A8 , 32'hE9A84C40 , 32'hF377D790 , 32'hFCD34404 , 32'hFA56DEB0 , 32'hEF6EDEA0 , 32'hFCCBE13C , 32'hFD2177EC , 32'h0AFE9410 , 32'hFCF54148 , 32'h038B0608 , 32'h0345540C , 32'hF49BE710 , 32'hFBF4CA80 , 32'h01581E0C , 32'hFFC2EBFA , 32'hFDA8A968 , 32'h00AD51F0 , 32'hFE4EA3D4 , 32'h050A99F0 , 32'h04420E58 , 32'h00D2C2B9 , 32'hFB13BBC0 , 32'hFF4F1ECE , 32'hFF96906D , 32'hF5282E80 , 32'h03F8A8C0 , 32'hFD36C5A8 , 32'h0037EA6C , 32'h03CEFC28 , 32'hFBA8F138 , 32'hF6708000 , 32'h08677320 , 32'hFD4C73DC , 32'hF84E9758 , 32'hFF2D5AB1 , 32'hFF33B832 , 32'h0370F6F8 , 32'hF999FBA0 , 32'hFB5FB228 , 32'h0330FF84 , 32'hFCBE66F0 , 32'h00376E48 , 32'h04ECD888 , 32'h02A825D8 , 32'h05E14088 , 32'hFDCC5518 , 32'h03205F7C , 32'hFF2369C0 , 32'h0267B3D0 , 32'hFAC87728 , 32'h02D3E204 , 32'h00BB6BAC , 32'hFFFF50DC , 32'hFFFC3B73 , 32'h0001412D , 32'h00014954 , 32'hFFFF09BE , 32'hFFFF5F42 , 32'h000000A1 , 32'hFFFFE6ED , 32'h00029CE4 , 32'h0000A854} , 
{32'hE71FFEC0 , 32'hDE4BBD80 , 32'h19C88400 , 32'h05BA6D98 , 32'hE3D86E40 , 32'hEFACA3E0 , 32'h09200B70 , 32'h0F5B6470 , 32'h11F572A0 , 32'hF2D4DAA0 , 32'h05ABA410 , 32'hF6879A80 , 32'h02B26D28 , 32'hEE3ECCA0 , 32'hEABAF280 , 32'h11185860 , 32'hFB10C990 , 32'h0ED48730 , 32'hFE809BB8 , 32'h188A3B40 , 32'h16C4E220 , 32'h085F2520 , 32'h033F98F4 , 32'hFE94D9C8 , 32'hF70A3B10 , 32'hF5A50FD0 , 32'h05D8B7E8 , 32'hF04C7EE0 , 32'hF8B0C8D0 , 32'hF5BD3ED0 , 32'h06FE64A0 , 32'hFC308B74 , 32'h0057CAD9 , 32'hFEEF4A94 , 32'h09B97870 , 32'hFC441340 , 32'h0E8D83F0 , 32'hF8D40CB8 , 32'hF773B800 , 32'h00356114 , 32'hFC3B1EC4 , 32'h004EE064 , 32'hF8A71F38 , 32'hF98B36B8 , 32'hF0067810 , 32'hEFDE50C0 , 32'hF46BEFF0 , 32'hF127EEE0 , 32'hFEBE6734 , 32'hFBC263D0 , 32'h077B3B48 , 32'h07F45918 , 32'hFCF5B914 , 32'hFFCE0CDF , 32'hFDAC95F0 , 32'hFA968DF8 , 32'h05A3DA20 , 32'h0B9C3650 , 32'hF762FC20 , 32'hFC45812C , 32'hFE9F4C14 , 32'h04BF4BD8 , 32'h03EBEAD0 , 32'h01D62120 , 32'h0D95B040 , 32'h017EA9F0 , 32'h08BFF220 , 32'hFB91E6D8 , 32'h050B06A8 , 32'h010D1458 , 32'hFB64CF60 , 32'h03D5634C , 32'h01CD5FDC , 32'hFA41A1F0 , 32'hF822D3A8 , 32'h002229AA , 32'hFF2B3207 , 32'h06C55278 , 32'hFE9D36FC , 32'hFE75B640 , 32'h01FE69C0 , 32'h05D36608 , 32'h003610B8 , 32'h00CE0304 , 32'h03B4AA1C , 32'hFF6581A9 , 32'hFFAF03EF , 32'hFE132AE8 , 32'hFE36F21C , 32'h014C2570 , 32'hFFFA1F45 , 32'h00017FD5 , 32'h00033F6B , 32'hFFFEEA8A , 32'h0000930B , 32'h00007F7E , 32'h0002E2C9 , 32'hFFFD10DA , 32'hFFFF7AB2 , 32'h00005CEE} , 
{32'hFFFE8431 , 32'hFFFD4FE5 , 32'h00043738 , 32'hFFFF09B2 , 32'hFFFE8F2B , 32'h0000F421 , 32'h00005A3E , 32'hFFFE2A99 , 32'hFFFDF234 , 32'hFFFEE311 , 32'h00033466 , 32'hFFFC0127 , 32'hFFFD32CB , 32'hFFFD746E , 32'hFFFC1AAE , 32'h000356B1 , 32'hFFFF5DA3 , 32'h00039119 , 32'h000038D9 , 32'hFFFFA766 , 32'hFFFE8EE3 , 32'h00033C31 , 32'h00044F66 , 32'hFFFF5877 , 32'hFFFC5FC4 , 32'h00028A96 , 32'hFFFC6AAB , 32'hFFFB525F , 32'h00008577 , 32'hFFFF4BC9 , 32'hFFFDF5B5 , 32'hFFFE6200 , 32'hFFFD012E , 32'h00006DF6 , 32'hFFFE7B16 , 32'hFFFF62F8 , 32'hFFFFA66F , 32'hFFFF1547 , 32'hFFFE2183 , 32'h0005D2BA , 32'hFFFF28F7 , 32'hFFFFB084 , 32'h0000C843 , 32'h0001FD66 , 32'hFFFE61FF , 32'hFFFDC8EC , 32'h00002195 , 32'h0002A9B6 , 32'hFFFCD0BE , 32'hFFFD8832 , 32'hFFFF3181 , 32'hFFFD925B , 32'h000147E5 , 32'hFFFE53C3 , 32'hFFFE9695 , 32'hFFFEA79E , 32'hFFFFF74C , 32'h00016283 , 32'hFFFD7140 , 32'h0001DBCE , 32'hFFFCD962 , 32'h0002B8FA , 32'hFFFE320F , 32'hFFFFADBB , 32'hFFFCCB0C , 32'hFFFED1D9 , 32'hFFFDFEDD , 32'hFFFC211C , 32'h00009954 , 32'h00064F4C , 32'hFFFD01C3 , 32'h00006F64 , 32'hFFFFA3F9 , 32'hFFFD724B , 32'hFFFEF9C3 , 32'hFFFEBCB0 , 32'h0000A599 , 32'h00001817 , 32'h00009569 , 32'hFFFFAF6C , 32'hFFFF80E5 , 32'h000352D5 , 32'h00003494 , 32'hFFFFAFC4 , 32'h000274A7 , 32'h000055F0 , 32'hFFFD544C , 32'hFFFF52DD , 32'h000237B0 , 32'h00044F07 , 32'h0000366D , 32'hFFFE2D3C , 32'hFFFC6703 , 32'h00050008 , 32'h000199D8 , 32'hFFFFE230 , 32'hFFFE1284 , 32'h000406ED , 32'h0001353C , 32'hFFFFB6FC} , 
{32'h0001B908 , 32'hFFFDBA16 , 32'h0002AFAD , 32'hFFFED4B0 , 32'hFFFEC1BA , 32'hFFFE799E , 32'hFFFC800A , 32'h0001D0F2 , 32'h0003C073 , 32'h00007C70 , 32'h0002B608 , 32'hFFFEEB54 , 32'h00016E67 , 32'hFFFCCA70 , 32'h000331BF , 32'hFFFF0BBF , 32'h0004862A , 32'hFFFD3031 , 32'h000254AE , 32'h0000241E , 32'h0000A12E , 32'h00030306 , 32'h00021BEB , 32'hFFFCC610 , 32'hFFFD82AD , 32'hFFFE4EF2 , 32'hFFF8F7FE , 32'h00030A0B , 32'h00002894 , 32'h00018702 , 32'h0005EFF4 , 32'hFFFD7161 , 32'hFFFC7923 , 32'hFFFFB6E6 , 32'h00005AF8 , 32'hFFFC4AB4 , 32'h0001143C , 32'h00017A61 , 32'h00017257 , 32'hFFFE912F , 32'h000377C3 , 32'hFFFE1F55 , 32'hFFFFB5DC , 32'hFFFF365B , 32'h0003C68C , 32'h000861E6 , 32'h00053FD4 , 32'hFFFB4FF5 , 32'hFFF7D204 , 32'hFFFD01F0 , 32'h00016BC1 , 32'hFFFDE53A , 32'h00004D6F , 32'hFFFA5CF5 , 32'h0000C9B3 , 32'hFFFC3C24 , 32'hFFFE4742 , 32'hFFFF3EF8 , 32'h00032D73 , 32'h000221A8 , 32'h0002C680 , 32'hFFFF343E , 32'hFFFF8A99 , 32'hFFFFD6F2 , 32'hFFFEF63C , 32'hFFFFA919 , 32'h00015AB3 , 32'hFFFF6958 , 32'hFFFEA99F , 32'hFFFC60B1 , 32'h00041031 , 32'hFFFD3DE9 , 32'hFFFC3BA8 , 32'hFFFC7D39 , 32'h00007862 , 32'h00035ABB , 32'h0000B67F , 32'hFFFD8DCD , 32'h00021A4B , 32'h0001BF52 , 32'hFFFF3F25 , 32'h000074C1 , 32'h000248DD , 32'hFFFD0283 , 32'h00008B97 , 32'h0005B633 , 32'h00011CFC , 32'h0005AF2C , 32'h0005D0B2 , 32'hFFFDBF2A , 32'hFFFE558F , 32'hFFFFCEFA , 32'h0000F632 , 32'hFFFE776E , 32'h00003274 , 32'h0001A52C , 32'h0003C588 , 32'hFFFFE6DC , 32'hFFFFBB12 , 32'hFFFC29CE} , 
{32'h0000AFF0 , 32'h00034B3C , 32'h0001D255 , 32'h0001B7A8 , 32'h0004C3EA , 32'hFFFFEF5F , 32'h00037077 , 32'hFFFF7825 , 32'h00028C55 , 32'hFFFFF596 , 32'h000303F6 , 32'hFFFFA116 , 32'h000161C9 , 32'hFFFE13E7 , 32'h00025FE6 , 32'hFFFF3A20 , 32'h00054186 , 32'hFFFDEC1C , 32'hFFFF67DA , 32'h000369C7 , 32'h00007C8A , 32'hFFFFC83C , 32'h00036348 , 32'hFFFD2989 , 32'h00025D36 , 32'h0000F86F , 32'hFFFAC15D , 32'h0000879F , 32'h0000CD8F , 32'h00023EDE , 32'h00002A00 , 32'hFFFEC31F , 32'h00042405 , 32'h00013336 , 32'h0001B920 , 32'hFFFB9EC1 , 32'h0004D4A0 , 32'h0001F954 , 32'h00034627 , 32'h000239A1 , 32'hFFFEB0B0 , 32'h00017FED , 32'hFFFF6829 , 32'h00052AE2 , 32'hFFFFAF0D , 32'h0002CFA6 , 32'hFFFECED2 , 32'h0000C256 , 32'h00027A86 , 32'hFFFE8B33 , 32'hFFFEA1D7 , 32'h00005E87 , 32'h0003B879 , 32'hFFFC4ECE , 32'h00023E2A , 32'hFFFF608D , 32'h0004A5B9 , 32'hFFFD85A8 , 32'hFFFEEFEC , 32'h00006B09 , 32'hFFFEA5E6 , 32'h0002A627 , 32'hFFFB3444 , 32'hFFFB4993 , 32'h0000E78D , 32'hFFFEB3A2 , 32'h0002CE42 , 32'h000249CA , 32'h00026A9D , 32'hFFFFDAB5 , 32'h00009DFB , 32'h0002539D , 32'hFFFD3761 , 32'hFFFFECB6 , 32'h000360EF , 32'hFFFECAA3 , 32'h00025C79 , 32'h0004AB85 , 32'hFFFAEB74 , 32'hFFFE768A , 32'h00023B3A , 32'h0005F72F , 32'hFFFAB17E , 32'h0002E665 , 32'hFFFA8C78 , 32'h0004490B , 32'hFFFD27ED , 32'hFFFED210 , 32'h000018DF , 32'hFFFF9647 , 32'h00029FB1 , 32'hFFFE9AF4 , 32'hFFFD7E1B , 32'h000078F5 , 32'h0000C107 , 32'hFFFF4E54 , 32'hFFFFE637 , 32'hFFFE7D9B , 32'h00008B13 , 32'hFFFE6C00} , 
{32'h04330460 , 32'h04F623E8 , 32'hF3DCBE50 , 32'h04EA1138 , 32'h0154E7C0 , 32'h032E1B50 , 32'hF6CBA670 , 32'h08BCE7C0 , 32'h02FD7D18 , 32'h08650A40 , 32'h0CCC6BE0 , 32'h00BCD005 , 32'h0B0CCEA0 , 32'hFF669771 , 32'h029897F8 , 32'hFDE2DC7C , 32'hFFC12E96 , 32'h063FFAA8 , 32'h05F5E700 , 32'h076DE460 , 32'h088FEFA0 , 32'hFE69DC24 , 32'hFE549C44 , 32'h023747A0 , 32'h00549CAE , 32'h04515CE0 , 32'h05B67D30 , 32'h01B373B8 , 32'hF7E56700 , 32'h02CED604 , 32'hFD2A62C0 , 32'hFA1E3640 , 32'h00F292F2 , 32'hED5A7920 , 32'hFA9AAD40 , 32'h001DC1E7 , 32'h06730D50 , 32'h0743CE68 , 32'hFD0FBEA8 , 32'hFF3B9B98 , 32'hFBFBF400 , 32'hFDF11690 , 32'hFA0E59D8 , 32'hF2FD0C60 , 32'hFFAB28C1 , 32'hFF166428 , 32'h0689BFC8 , 32'hFE34C844 , 32'hFF09E477 , 32'h05CFB2C0 , 32'h05CA4F80 , 32'hFDDB5E84 , 32'h00BE1445 , 32'hFE6304AC , 32'h02112E98 , 32'h087C06B0 , 32'hF8A67DE0 , 32'h0562B098 , 32'h03FF9AE4 , 32'h009C1FA0 , 32'hF6231B10 , 32'hFDB55A6C , 32'h00AF2154 , 32'h001DF58E , 32'h03993404 , 32'hFBF53CC0 , 32'hFE10C9B4 , 32'hFE6BA7D4 , 32'hFF5BB401 , 32'h0586D188 , 32'hFFFB1FCD , 32'h01B59E48 , 32'h023CA51C , 32'h01A4235C , 32'hFDB991BC , 32'h0252AC08 , 32'h0394E528 , 32'h00B6D853 , 32'hFD7B4E50 , 32'hFDD25810 , 32'hFFB9C174 , 32'hFD2521F0 , 32'hFB1D5290 , 32'h0041F91C , 32'h046574D8 , 32'h04245F40 , 32'h04B91AC8 , 32'hFDB8744C , 32'h033482E0 , 32'hFF37B1D2 , 32'hFFFEBADC , 32'h0002938B , 32'hFFFD97F3 , 32'h00004BE4 , 32'h00017A6C , 32'hFFFF4B3F , 32'h000149B5 , 32'hFFFDDAFE , 32'h0000C1BB , 32'hFFFF8AE2} , 
{32'h00042F06 , 32'hFFFC867B , 32'h00003C33 , 32'h000488A6 , 32'hFFFC70DB , 32'h00005B4C , 32'hFFFE2095 , 32'h00018C6D , 32'hFFFAF467 , 32'hFFFBACFA , 32'hFFFEFA75 , 32'h0000F640 , 32'h0005AAC8 , 32'h0000FAA6 , 32'h0002A682 , 32'h000464AB , 32'hFFFE7A19 , 32'hFFFFCBC2 , 32'hFFFF8BD8 , 32'hFFFFE0EB , 32'hFFFF2BA0 , 32'hFFFE35DD , 32'h000248D8 , 32'h00007B96 , 32'h000305A3 , 32'hFFFC45EE , 32'h00027E54 , 32'h000001DF , 32'h00028DAB , 32'h0003E7B7 , 32'hFFFE3395 , 32'h00024095 , 32'hFFFEBC43 , 32'hFFFEB7C1 , 32'h000050A8 , 32'h00032B25 , 32'hFFFFCE5E , 32'h0001CA1C , 32'h00013367 , 32'h0003207E , 32'h00020F48 , 32'hFFFC5100 , 32'h00007BC0 , 32'h00024E9B , 32'h0000C617 , 32'hFFFE8D43 , 32'h00051959 , 32'hFFFC2096 , 32'hFFFFD620 , 32'hFFFF0364 , 32'hFFFD5E2B , 32'h000065ED , 32'h00033476 , 32'hFFFD043A , 32'h00022A43 , 32'hFFFF7C7C , 32'hFFF8E870 , 32'hFFFB99FE , 32'hFFFFDD95 , 32'hFFF6F7E2 , 32'h00000045 , 32'h00025362 , 32'h0004D156 , 32'h00011C2B , 32'h00020E83 , 32'h000073A7 , 32'hFFFEFCD2 , 32'hFFFE8B6B , 32'h0000994F , 32'hFFFE7944 , 32'hFFFD46D4 , 32'h0002939E , 32'h000061A8 , 32'h00012E77 , 32'h00000B9C , 32'hFFFC39DF , 32'hFFFA6645 , 32'hFFFE8602 , 32'hFFFE955E , 32'h00023355 , 32'hFFFCF0ED , 32'h00012233 , 32'h0003958F , 32'h0001FEE9 , 32'h0000DA30 , 32'h00023A84 , 32'hFFFF6C71 , 32'hFFFBCF3F , 32'h00007B71 , 32'hFFFEC66E , 32'hFFFCA848 , 32'h00039D60 , 32'hFFFFE2E1 , 32'h00037D7A , 32'hFFFCA2B3 , 32'hFFFEB0A2 , 32'hFFFF7A60 , 32'h0001A2C9 , 32'h00026B33 , 32'hFFFB5FBB} , 
{32'h0000A208 , 32'hFFFAD54A , 32'hFFFD27A4 , 32'hFFFF4410 , 32'h0002796D , 32'hFFFE20EE , 32'h0000746E , 32'h0001B548 , 32'h0002F9EE , 32'hFFFE15FE , 32'hFFFFDAB7 , 32'hFFFEFDF7 , 32'hFFFDC9D9 , 32'hFFFBDBBC , 32'h000169AF , 32'h00004088 , 32'hFFFC508C , 32'h00025278 , 32'h00006AAB , 32'h0003DBF3 , 32'h00003144 , 32'h0001E80B , 32'h0000D061 , 32'hFFF9AF7A , 32'hFFFF1D35 , 32'h00030098 , 32'h000314EB , 32'hFFFD21A6 , 32'hFFFD407E , 32'h00005A61 , 32'h0001DF74 , 32'h00062DBB , 32'h00026FEA , 32'hFFFF435C , 32'h0002A7BC , 32'h000059E3 , 32'hFFFFF9EB , 32'hFFFD281E , 32'h0002B504 , 32'h0006BA9A , 32'hFFFEE5AB , 32'h0000CC06 , 32'hFFFFAEF4 , 32'h00005615 , 32'hFFFF35A3 , 32'hFFFE50B9 , 32'h0001FE3B , 32'hFFFE84A2 , 32'hFFFABB32 , 32'hFFFFE1F9 , 32'hFFFB14E2 , 32'h00030E52 , 32'hFFFD1415 , 32'hFFF9F66C , 32'hFFFB0EC5 , 32'hFFFE09AA , 32'h00004247 , 32'hFFFE66E0 , 32'h0000470E , 32'h000413A1 , 32'h00035A99 , 32'hFFFE3100 , 32'hFFFF0724 , 32'h00021E3E , 32'h0001C911 , 32'hFFFD20A0 , 32'hFFFD43CB , 32'hFFFF192E , 32'hFFFA228C , 32'hFFFC6EFE , 32'hFFFA0712 , 32'hFFFEEA5F , 32'h00009F95 , 32'hFFFC51D2 , 32'h0000F5B2 , 32'h0000418B , 32'h00045FF0 , 32'hFFFD5531 , 32'h0005C4D9 , 32'h00047D04 , 32'h0001358A , 32'hFFFFBCC9 , 32'h0000055A , 32'hFFFFC833 , 32'hFFFFB03C , 32'h0003A304 , 32'hFFFD6AE3 , 32'h000020AC , 32'hFFFF0DA6 , 32'h00012F6E , 32'h00062C1E , 32'hFFFDDED6 , 32'h0004D1F4 , 32'hFFFE384F , 32'hFFFAD4CC , 32'hFFFFF1FD , 32'h0005A093 , 32'h0004C810 , 32'hFFFEFA34 , 32'h0001F6D2} , 
{32'h09076F50 , 32'hF3B78020 , 32'hF88CC1D8 , 32'h0C7EC7C0 , 32'h05A640E8 , 32'hECEED040 , 32'hEF347EC0 , 32'hFC89A020 , 32'h072DE3D0 , 32'hF145C840 , 32'h05109DC0 , 32'hF8709E28 , 32'h0F7DC0D0 , 32'hF95A14F0 , 32'h0A19D790 , 32'h077028F8 , 32'hFDD12994 , 32'hFF1C75A5 , 32'h001A4B17 , 32'h02E38134 , 32'hF7230D30 , 32'hFE5EF910 , 32'hFC3B89E0 , 32'h084F3680 , 32'hFF9D3DE2 , 32'hFFA22AA3 , 32'h0600B400 , 32'hF21A64F0 , 32'hFE604D44 , 32'hEE217EE0 , 32'h020F4FA4 , 32'h08D2E890 , 32'hFB850698 , 32'h00BF4E9D , 32'hEFEF7960 , 32'hFD2748E4 , 32'h02B8A6F0 , 32'h05B9F338 , 32'h0661CA88 , 32'h0042E506 , 32'h091B72B0 , 32'hFF8E2086 , 32'hFD6E661C , 32'h02C08AE8 , 32'hFA29E788 , 32'hFF350EC3 , 32'hFF0EB054 , 32'hFD1EB074 , 32'h08E5EA90 , 32'hFD652A9C , 32'h0AB767D0 , 32'h0A537600 , 32'h03FE745C , 32'h03A298F4 , 32'hFD7D41B0 , 32'hF762E3C0 , 32'hFF235E91 , 32'hFA4D8BE0 , 32'hFBECA438 , 32'hF8B7D2B8 , 32'h01AA1A34 , 32'h05C7B000 , 32'h005DF7F4 , 32'h014F3878 , 32'hFEDFFDB4 , 32'hF9047AE0 , 32'hFF70CEB2 , 32'hFDB87AC4 , 32'h0143F7C0 , 32'h01BB6858 , 32'h0292FD7C , 32'hFE7D0F38 , 32'h067921A0 , 32'hFB56B400 , 32'h063046D0 , 32'hFE85C79C , 32'hFCF10524 , 32'hFB0B9130 , 32'h06DD7960 , 32'hF86AE390 , 32'h000C1155 , 32'hFE6C30E0 , 32'h00CE4541 , 32'hF8359230 , 32'hF9ECB4C0 , 32'hFF7C9261 , 32'hFFDC449C , 32'hFC4E9DC0 , 32'h03B39A94 , 32'hFF94086A , 32'h0001875C , 32'h00028D4B , 32'hFFFEEE02 , 32'h00010400 , 32'h00008743 , 32'hFFFF8C9C , 32'h0001CC53 , 32'hFFFFDE3F , 32'hFFFEE367 , 32'hFFFFBD07} , 
{32'hFF003ACA , 32'hE6AB18A0 , 32'hBC0C9D00 , 32'hD4E636C0 , 32'h1CDCDE80 , 32'hFE66507C , 32'hFAFBAB98 , 32'hF1C6B450 , 32'hF514A4B0 , 32'hF9056D78 , 32'hE1C56940 , 32'hF7A0E4D0 , 32'h0F1D4720 , 32'h045064E8 , 32'hFB919CD0 , 32'hF83DB898 , 32'h010179FC , 32'h09A2B890 , 32'h19E6F7A0 , 32'h0E1FF2D0 , 32'hE6DC2700 , 32'h059D0D10 , 32'h0A8379E0 , 32'h0483A720 , 32'hF1229700 , 32'h024BA978 , 32'hF42CB810 , 32'hFD5C4658 , 32'hDEE402C0 , 32'hFA309CD8 , 32'hF749D560 , 32'h005B28D0 , 32'h06528E40 , 32'hEBCB8EA0 , 32'hFA5D4408 , 32'h155FEF60 , 32'hFF4080C2 , 32'hF26535E0 , 32'h0EB151B0 , 32'hFEA2AFBC , 32'h0D674A20 , 32'hF1016C90 , 32'h00425C7C , 32'hFC72C070 , 32'h011DDC74 , 32'hFBD9F828 , 32'h04301D70 , 32'hF81BC6D8 , 32'h113C88C0 , 32'hF9BB7320 , 32'hFCB6BFC8 , 32'hFAF7CA18 , 32'h03270B60 , 32'h08629AE0 , 32'h08F93610 , 32'h15061DA0 , 32'hFE7B37AC , 32'h0B6A6120 , 32'hFA9467E8 , 32'hFD209E38 , 32'h04EE5008 , 32'hFFFCCB2B , 32'h043293F8 , 32'h04C20908 , 32'h073339E8 , 32'hF87B8930 , 32'h00C0DCDD , 32'h027B0CDC , 32'h00D4CD0B , 32'h0A15CF50 , 32'h07FB4BB0 , 32'hFD19D61C , 32'hFED04D84 , 32'hFC969114 , 32'hFE0296B4 , 32'h014C2A5C , 32'hFF165A78 , 32'h002E0958 , 32'h00AAEDC9 , 32'h00A2E2CC , 32'h00BCC695 , 32'hFE97722C , 32'h03960FC4 , 32'h012614EC , 32'hFCE0C838 , 32'h00145157 , 32'h02F526A8 , 32'h026496A4 , 32'hFE0F6A48 , 32'h00C7C809 , 32'hFFFF916C , 32'hFFFF2BB9 , 32'h0000AACB , 32'h000153F5 , 32'h0002142E , 32'hFFFEB976 , 32'h0001C548 , 32'hFFFF7A35 , 32'h00000D6A , 32'h00016677} , 
{32'h0001A75B , 32'hFFFDDB9E , 32'h00036CAE , 32'h00006F2D , 32'h0002A285 , 32'h00064D3A , 32'hFFFBF498 , 32'h00007F56 , 32'h0000E780 , 32'h0004D22A , 32'h00002E26 , 32'hFFFD0A9F , 32'hFFFE9E19 , 32'hFFFE91ED , 32'hFFFE55F1 , 32'h0003D64B , 32'h00005BA9 , 32'hFFFCA841 , 32'hFFFAE858 , 32'hFFFF9437 , 32'h00049642 , 32'hFFFFEB6E , 32'hFFFFBDBD , 32'h0000DF30 , 32'h00020DC8 , 32'hFFFF2858 , 32'hFFFAE573 , 32'hFFFBD086 , 32'h0000FB20 , 32'h0000666D , 32'hFFFB47C9 , 32'hFFFD5183 , 32'h00030598 , 32'hFFFE9608 , 32'h0000CCCC , 32'h000002B9 , 32'h0000BA9D , 32'h0000CCBD , 32'hFFFDF7BF , 32'h00043F80 , 32'hFFFE6914 , 32'hFFFD9C12 , 32'h00001C6E , 32'h0003DDB2 , 32'h00017B39 , 32'hFFFDCF93 , 32'h000264FA , 32'h00011E74 , 32'hFFFD5240 , 32'hFFFF548A , 32'h0001724E , 32'hFFFE5588 , 32'h00012B3D , 32'h0001876B , 32'hFFFF465C , 32'h0002106D , 32'h0001C498 , 32'h000162EF , 32'h0001D30C , 32'hFFFF8A42 , 32'h0000382E , 32'hFFFFE9AF , 32'hFFFAE789 , 32'hFFFEE138 , 32'hFFFED6BB , 32'hFFFF0450 , 32'h000106B3 , 32'hFFFCAC20 , 32'h0000875E , 32'h0006B3B4 , 32'hFFFE3CB0 , 32'h0001A488 , 32'h0002F255 , 32'hFFFE11F5 , 32'hFFFFA89E , 32'h00026F17 , 32'hFFFE6FEA , 32'hFFFCB1A6 , 32'hFFFD5886 , 32'h000018E1 , 32'hFFFFE02C , 32'h000271B0 , 32'hFFFD7652 , 32'hFFFDB7DD , 32'h00022346 , 32'h0001F59C , 32'hFFFF9E0D , 32'hFFFE0D61 , 32'h00002C5A , 32'h000297FC , 32'hFFFE7806 , 32'h0003CC05 , 32'h000425D8 , 32'hFFFE48D4 , 32'hFFFE88F1 , 32'h0002AF8D , 32'hFFF922A4 , 32'hFFFD300F , 32'hFFFD99C8 , 32'hFFFF5F5C} , 
{32'hC8DCBAC0 , 32'h80000800 , 32'h07CE5A20 , 32'h045BDA70 , 32'h00E9BA4B , 32'hFAF4ECF8 , 32'h23EEE800 , 32'hF8CE1598 , 32'h115F4980 , 32'hE8E00CE0 , 32'hE5296CA0 , 32'hF0D15570 , 32'hEB1902E0 , 32'h1D669560 , 32'h15C67F60 , 32'h021B5FF0 , 32'hDE9B7D00 , 32'hFCE91594 , 32'h054F8A68 , 32'hE5391660 , 32'hFA6027F0 , 32'h0573A878 , 32'h0CF0D8C0 , 32'h12C4EE80 , 32'h1E1EC680 , 32'h03ED63B8 , 32'hFAF3E190 , 32'hFB4D13F8 , 32'hF3566600 , 32'h0993BAD0 , 32'h015FF950 , 32'hFC644FA4 , 32'h048DAD18 , 32'h00A91F0C , 32'h0F60A260 , 32'hF4D2B0D0 , 32'hFB8C2A60 , 32'h0DDBA0A0 , 32'h0258C00C , 32'h0600BC48 , 32'hF94DB510 , 32'h04524E20 , 32'h0401BEF8 , 32'hFE456C7C , 32'h02AB5954 , 32'h0C73E5D0 , 32'h02E19728 , 32'hFB8D8608 , 32'hFAECB6E8 , 32'hFDCEB380 , 32'h042CEC18 , 32'h04872050 , 32'h018DBA00 , 32'h00C56DBB , 32'hF76116C0 , 32'h08509290 , 32'hF74D9D90 , 32'hFE986898 , 32'h0281CBE8 , 32'hF2FD7A00 , 32'hF47EB050 , 32'hFC13BCBC , 32'h00E1BB96 , 32'hFB829A48 , 32'h04BC6D30 , 32'h05A11B70 , 32'h01F75EF8 , 32'h00879122 , 32'h01A7F0D0 , 32'h0454FF40 , 32'h04A94980 , 32'hFC5093B4 , 32'hF9500400 , 32'hF9B8FFF8 , 32'hFBA78E58 , 32'h00FEF8B2 , 32'hFFF65648 , 32'h05982F68 , 32'h0179124C , 32'hFFCC01DD , 32'hFBC4D6C8 , 32'h06A4BAA8 , 32'hFDE58250 , 32'h011E3CD0 , 32'h000477BE , 32'h009E08DC , 32'hFF8A8C49 , 32'h00A301BE , 32'hFF34071A , 32'h008A7081 , 32'hFFFE62ED , 32'h00001BEB , 32'hFFFE641D , 32'hFFFFCEAB , 32'h00001C60 , 32'h0001ABE9 , 32'hFFFEEB3A , 32'h0000F066 , 32'hFFFFA8D4 , 32'hFFFDC5C0} , 
{32'hF770E240 , 32'h136BA4E0 , 32'hFBD23148 , 32'h05494298 , 32'h0863D620 , 32'h07F7DA38 , 32'h07543E48 , 32'hFA52DD90 , 32'hFD3CA49C , 32'h06343A18 , 32'hFDDE0444 , 32'h00008630 , 32'hE7C40EC0 , 32'h0045AC87 , 32'h04A5D390 , 32'h0663CD10 , 32'hFEC86748 , 32'h0AB6FC10 , 32'h074239A0 , 32'hF74F9BB0 , 32'hF9493DA8 , 32'h031D1454 , 32'h0A1B83F0 , 32'hF816B498 , 32'hFD9DB400 , 32'hF63E92D0 , 32'hFB993ED0 , 32'h078D3638 , 32'hFE7F8F4C , 32'h09210700 , 32'h08A2D0D0 , 32'hFCFF1890 , 32'hFE9C3FFC , 32'hF91D1298 , 32'hFE6E7830 , 32'h0C7908C0 , 32'h0516D758 , 32'h0552A158 , 32'hFE0E80FC , 32'h0A7DDA70 , 32'h0137A97C , 32'hFD9EED8C , 32'h015AB2D4 , 32'h04807168 , 32'hFDEAAF98 , 32'h0023ACE0 , 32'hF92DC9A8 , 32'h029FA364 , 32'h007157E3 , 32'h03C109E4 , 32'hFDFD3A60 , 32'hF73DAC50 , 32'hFE4D165C , 32'hF47ADE00 , 32'hFA3ABB78 , 32'h02799B50 , 32'h003C6593 , 32'h04E7D268 , 32'hFE2FC5B4 , 32'hFA4D4088 , 32'hF6053D70 , 32'h013C956C , 32'hF61F8FB0 , 32'hFB32ADA8 , 32'h08403B20 , 32'h036096E8 , 32'hF9E47EC0 , 32'hF83BEEE8 , 32'h03F21B50 , 32'h01F9F964 , 32'hFCA9E89C , 32'hFA30ABB8 , 32'hFB22C608 , 32'h01BCFAB0 , 32'hFC46677C , 32'h0191CC68 , 32'h07842490 , 32'h0141AB3C , 32'h031F314C , 32'h00E70814 , 32'h034BC304 , 32'h01D9F7E4 , 32'hFF53DF58 , 32'h04248398 , 32'hFCD02514 , 32'h04C845E0 , 32'hFAC16650 , 32'h0126A5F4 , 32'hFF225815 , 32'hFF4E1D6B , 32'h00025C1E , 32'hFFFD564A , 32'h00013CC3 , 32'hFFFFA1B9 , 32'h00037012 , 32'h0001B98C , 32'hFFFC8EE2 , 32'hFFFF9B4B , 32'h0000852F , 32'h0000BFC1} , 
{32'h04F77890 , 32'hFE97C4B4 , 32'hECBA2060 , 32'hF1737A70 , 32'h013BE0B0 , 32'h027566F4 , 32'h12A8C7C0 , 32'hEC8CFF80 , 32'hF390B450 , 32'hF901E370 , 32'h0A7AECF0 , 32'h0E5AAE30 , 32'hF0675770 , 32'h0AB36950 , 32'hFC2A2160 , 32'hFD7FCDC8 , 32'h0E36A7B0 , 32'hF31A5990 , 32'h025EC008 , 32'hFE86A914 , 32'h144CE460 , 32'h0900ABA0 , 32'hFE9A9C8C , 32'h0ED7ACF0 , 32'h0F31BCE0 , 32'h01FD08CC , 32'h0338EED4 , 32'h1B5DEAA0 , 32'h08F73230 , 32'h019A9BE0 , 32'hFD5C8588 , 32'hFE71CF84 , 32'hFD1AC6D8 , 32'hFEA4FAF0 , 32'h07A9BD60 , 32'h01069CDC , 32'h02247550 , 32'hECE36040 , 32'hFA24C3A8 , 32'hFB907C60 , 32'hFE1B3E4C , 32'h00DF6EAA , 32'h05CB2BE0 , 32'h19C93900 , 32'hF442C6A0 , 32'h02F2CD54 , 32'hFE58D078 , 32'hFBF24A10 , 32'h081CA990 , 32'hF7E53410 , 32'hF8F961A8 , 32'h02C26C08 , 32'hFC097030 , 32'hFF55082A , 32'hF9AE7AD0 , 32'hF4C40040 , 32'hFF528667 , 32'hFACC6C88 , 32'h027416C8 , 32'hFCF2B5B4 , 32'h01C6814C , 32'hFE5A8308 , 32'hFB66A6A8 , 32'h04080BD0 , 32'h039BDD18 , 32'hFE5CBD30 , 32'h047C3410 , 32'h03B5C7AC , 32'hFF6BD0BF , 32'hF97AC9B0 , 32'h07D42030 , 32'hFEFC8AEC , 32'h0AD323B0 , 32'hFE833E84 , 32'hFE50C6BC , 32'hFFD5F45A , 32'h01F042A4 , 32'h05F10740 , 32'h03A2E080 , 32'h00B08C33 , 32'hFF3ECDE3 , 32'hFDFAD074 , 32'h00F93BED , 32'hFE57B70C , 32'h0098CF48 , 32'hFD9F5E18 , 32'hFFA43B25 , 32'h00EA1604 , 32'hFD9B9678 , 32'h00CA7277 , 32'hFFFDF4E9 , 32'h00012FC6 , 32'hFFFFD68C , 32'hFFFDC5F0 , 32'hFFFEB200 , 32'h0001BC4D , 32'h00003160 , 32'hFFFFBC3F , 32'h00020F67 , 32'hFFFF4BC6} , 
{32'hE87A8060 , 32'h00BB0A40 , 32'hDC28DB40 , 32'h16C68140 , 32'hD5863600 , 32'h1775C900 , 32'hFD49A4D0 , 32'h17E7E560 , 32'hFB554A58 , 32'h05B04040 , 32'hFE6A2924 , 32'hFEEA7A7C , 32'hFA9E6D68 , 32'h11AC7020 , 32'hFD40BA94 , 32'hF71CB0D0 , 32'hEB9E96C0 , 32'hEDA5CB40 , 32'hFCC52AD8 , 32'h1073FFA0 , 32'hEF153BA0 , 32'hF406DEA0 , 32'h04312378 , 32'hF1831AE0 , 32'hF98177D8 , 32'h0089E9DE , 32'hFECFD05C , 32'hFA0AF9A8 , 32'hF9CA9020 , 32'h0197F320 , 32'hF81E5540 , 32'h0FE446B0 , 32'h03CB3638 , 32'h031327EC , 32'h010EC4F4 , 32'h0AFE5100 , 32'hF1209B90 , 32'h010A81FC , 32'h01FAB2B8 , 32'hF77A11A0 , 32'hEAFE4F80 , 32'hFE4FCE6C , 32'h03342184 , 32'h122BAC20 , 32'hF4108920 , 32'h05C3E4A8 , 32'h0D52D180 , 32'h076F6F98 , 32'hF9742A10 , 32'h05947A70 , 32'h04434470 , 32'hFF3F7E6B , 32'hF0E693A0 , 32'hFB88B568 , 32'h09145110 , 32'hFD204540 , 32'hF8FE0718 , 32'h00BD41CF , 32'h0180E22C , 32'hFDB90308 , 32'h006EDFB5 , 32'hFFCA5D6D , 32'hF849C168 , 32'hFE160038 , 32'hFBE0CEE8 , 32'hF6CF1570 , 32'h0ADD1EE0 , 32'h07F83658 , 32'hFE997A54 , 32'hFD9F297C , 32'h01905420 , 32'h016080D0 , 32'h00A02F39 , 32'hFAE18DF8 , 32'hFB5E9F70 , 32'h001D3B59 , 32'h031C0790 , 32'hFAE2D040 , 32'h04365CA8 , 32'hFD333574 , 32'hFC9D7F28 , 32'hFFCFE1AC , 32'h01E683FC , 32'hFF96B168 , 32'hFE842A04 , 32'h01154024 , 32'hFE81C330 , 32'hFF28B959 , 32'hFE61C308 , 32'h00BACAB8 , 32'h00003BB6 , 32'h0002B4D0 , 32'h00007523 , 32'hFFFED238 , 32'hFFFFFC01 , 32'h00012B76 , 32'h000192AE , 32'hFFFE0863 , 32'h000092DA , 32'hFFFF814F} , 
{32'hFFFDD2B7 , 32'hFFFC481C , 32'hFFFDDA40 , 32'h0002952C , 32'h00017E7F , 32'hFFFC6E7C , 32'hFFFF1FD7 , 32'h00019960 , 32'h0001E228 , 32'h00031203 , 32'h0003394A , 32'hFFF9F427 , 32'hFFFBC711 , 32'h00021A4A , 32'h00026EA9 , 32'h0003274C , 32'hFFFDF7C2 , 32'hFFFBFB22 , 32'hFFFF1ED3 , 32'h000083DD , 32'hFFFCEC33 , 32'h00037A83 , 32'hFFFCEC8F , 32'h00020412 , 32'h0002A4CD , 32'h0000DC9D , 32'h0002C8E5 , 32'hFFFFBE02 , 32'h0000972B , 32'h00029C32 , 32'h000262D3 , 32'h00007885 , 32'hFFFE8717 , 32'h00019E21 , 32'h0001479C , 32'h0001073A , 32'h00001C2C , 32'h0001391F , 32'hFFFD7171 , 32'hFFFEDC15 , 32'h0002A88D , 32'hFFFF5395 , 32'h00007C67 , 32'hFFFF3E73 , 32'hFFFDDFCC , 32'h0000FCFB , 32'h00007CF7 , 32'h00012BCE , 32'h000383F3 , 32'h000565E7 , 32'h0001546E , 32'h00035658 , 32'h0000B1E2 , 32'h000465C7 , 32'hFFFC9D0A , 32'hFFFD8DAB , 32'hFFFD4A5E , 32'h0005665D , 32'hFFFF512F , 32'h0000779E , 32'h00024772 , 32'hFFFF46F7 , 32'hFFFD7ABC , 32'hFFFB8811 , 32'hFFFF51C5 , 32'h0001ACCD , 32'h000128A9 , 32'hFFFCA080 , 32'hFFFED390 , 32'hFFFF4846 , 32'hFFFFAA42 , 32'hFFFE3A61 , 32'h0001F9BE , 32'h0002CDD0 , 32'h0004C775 , 32'hFFFCD3AB , 32'h000078B7 , 32'h0000F73F , 32'hFFFE4CB6 , 32'h000178A9 , 32'h00002F60 , 32'h00029BB3 , 32'hFFFBFD74 , 32'hFFFF11C4 , 32'h00013D53 , 32'hFFFFE0EB , 32'hFFFE1AB1 , 32'h00008669 , 32'h0003D9D6 , 32'h000043BC , 32'h000105CC , 32'h00042916 , 32'h0001E56E , 32'h0003348D , 32'hFFFEFE87 , 32'h00007F5A , 32'hFFFE2B7F , 32'h0003F289 , 32'h0001AA17 , 32'hFFFFEBA4} , 
{32'h0B0A70F0 , 32'hF8F1DD28 , 32'hF8B0DD08 , 32'h0E4DBE70 , 32'hE2727020 , 32'h0F0F3D50 , 32'h09841D90 , 32'h0704BF68 , 32'hFD682CD0 , 32'hFB7A37D0 , 32'h059BC8F8 , 32'hF9AFFCC8 , 32'h05FCCD00 , 32'hFF7ACC69 , 32'h07B77970 , 32'h106DE6C0 , 32'h080F2B40 , 32'hE84FB9A0 , 32'h07CD1028 , 32'h0C0063B0 , 32'h0B79B220 , 32'hFA2A6A18 , 32'hFF6D1391 , 32'h029296B8 , 32'hF8102E70 , 32'h035C1910 , 32'hF8A09198 , 32'hFD9D65F4 , 32'h001BBD2F , 32'hEF372240 , 32'hFE416960 , 32'hFFE293B4 , 32'h09707AD0 , 32'hF8769C10 , 32'h070825A8 , 32'hFE0E49A4 , 32'h0424AA90 , 32'h11B07BA0 , 32'h0FCD4150 , 32'h0427CCA8 , 32'h15C7A960 , 32'hFDDB3D0C , 32'h029AB534 , 32'h03D9C138 , 32'hFE207F38 , 32'h03786C20 , 32'hF76DC310 , 32'hFA7D1AF8 , 32'hFA342340 , 32'hF2D98ED0 , 32'hFE7AE814 , 32'hF691DD20 , 32'hFF57885A , 32'h0D5776E0 , 32'hFCB36900 , 32'h09FB42C0 , 32'h001855AF , 32'hFB2F74F8 , 32'h025A2538 , 32'hFC33D838 , 32'hFE699C40 , 32'hFAAB2468 , 32'h0258D0FC , 32'h03E17474 , 32'hFC81DA78 , 32'h10D134C0 , 32'hFBFBE820 , 32'hFA4FD388 , 32'h03B6468C , 32'h04578430 , 32'hFD09DEB0 , 32'hFC3EC804 , 32'hF80498B8 , 32'h01A77940 , 32'hFFEFB189 , 32'hFAB815C0 , 32'h02B2B4B0 , 32'hF8393B78 , 32'h06030A80 , 32'hFF310628 , 32'h01B69F98 , 32'hFE864408 , 32'h031E9B8C , 32'hFDB608D4 , 32'h00DDE2C3 , 32'hFACDBB88 , 32'h00DC1422 , 32'hFFDB1004 , 32'hFE239B88 , 32'h00B29F4D , 32'h00013900 , 32'h0003A120 , 32'h0000995B , 32'h00025EF6 , 32'hFFFF96AE , 32'h0000FAA4 , 32'h000195A2 , 32'hFFFC6F56 , 32'h0000B312 , 32'hFFFED65D} , 
{32'h16BDBDE0 , 32'h0CBF7250 , 32'h20788900 , 32'h0DD440E0 , 32'h13362880 , 32'hDBC8A9C0 , 32'h1089C920 , 32'h18614D00 , 32'hE6B0B160 , 32'hE75F1E20 , 32'hF81A0498 , 32'h126AA0C0 , 32'hF3582900 , 32'hF7924720 , 32'h081871E0 , 32'hF0856020 , 32'hFC88B9FC , 32'h0CD6FDD0 , 32'hFDC8ACEC , 32'h04C81D58 , 32'hF12B4550 , 32'h1A8EF5A0 , 32'h03226680 , 32'hF1505880 , 32'h09CC0F70 , 32'hF6FF13B0 , 32'h00F4DCA7 , 32'h19943E00 , 32'hF5CA7AC0 , 32'h0BADA3D0 , 32'hF5016720 , 32'h0E9D2BC0 , 32'hFDAF7E28 , 32'h0EF707A0 , 32'h0B7FF720 , 32'h0B73F230 , 32'hFEE9F448 , 32'h02979DF0 , 32'h14F2DE00 , 32'hEF25E920 , 32'h0730B5B0 , 32'h03A4D76C , 32'hEDE27640 , 32'hFA6681D0 , 32'h0635FFB8 , 32'hF36A3FB0 , 32'hF9FE1D40 , 32'h04285788 , 32'hF68118B0 , 32'h01CB923C , 32'hFF6DB3F6 , 32'hF6E4E630 , 32'hF97592F8 , 32'hF78A5F30 , 32'h0589C6F8 , 32'hFDE99868 , 32'h05B22620 , 32'h00875EA5 , 32'hF421D130 , 32'hFDF8B110 , 32'hF1137010 , 32'hF8A263E8 , 32'hFD8823A8 , 32'h02785288 , 32'hFE1E2EC4 , 32'h06581068 , 32'hFCA3B0F0 , 32'hFDB945B4 , 32'hF69FB480 , 32'hFD474DA8 , 32'h037595AC , 32'h075FEFA0 , 32'h05A592E8 , 32'h06705858 , 32'hF90F35E8 , 32'h07AAA2C8 , 32'hFA997080 , 32'hFF8E7E23 , 32'h006A8CBD , 32'hFCAF1004 , 32'hFB9FDF40 , 32'hFF99B186 , 32'h00DC899A , 32'hFFEC32DB , 32'h013E4E30 , 32'hFFD1631F , 32'h014578E4 , 32'hFEE628B0 , 32'hFDE9FCF8 , 32'hFFB21BD6 , 32'h00012B71 , 32'hFFFE35AC , 32'hFFFFD35C , 32'h00038F9B , 32'h0000A42F , 32'hFFFF04C5 , 32'h000148E6 , 32'hFFFF091B , 32'h0000D829 , 32'h0000BD02} , 
{32'hFA9DC0E0 , 32'hFDCEFAAC , 32'hF91E4980 , 32'h0EBEE4C0 , 32'hFC4094D4 , 32'h01861DD8 , 32'hF9E641D0 , 32'hF5F3A2C0 , 32'hF79E85A0 , 32'h033C7CCC , 32'hF4B334E0 , 32'hFDBEE898 , 32'h089BA840 , 32'h00232006 , 32'hF8B50000 , 32'hFADD0CC8 , 32'h047A41F0 , 32'h0ABB5C60 , 32'hF7554240 , 32'hFE252F14 , 32'hF9900F90 , 32'h000D3181 , 32'hFF9CA8B8 , 32'h08EF1410 , 32'h029B23A4 , 32'hFD03E258 , 32'hF9B629A8 , 32'h05DA3BB0 , 32'h0085B8EA , 32'h009C4AC3 , 32'hFD5324BC , 32'h01CD2834 , 32'hFDC5291C , 32'hFAF13548 , 32'hF5AB7E30 , 32'h020995CC , 32'hFC667754 , 32'h0DB389D0 , 32'hFA574320 , 32'hEDDDBC00 , 32'h08EA3DA0 , 32'hFD1BCA4C , 32'h041CBE58 , 32'hFC234E20 , 32'hFED79D34 , 32'hFD34919C , 32'hFF3544C9 , 32'hFD9A287C , 32'h02DA3984 , 32'h01427554 , 32'h06583878 , 32'hFB8A4788 , 32'hFFB22B05 , 32'hFEE57620 , 32'hFE51E800 , 32'h010885A0 , 32'h05A83E10 , 32'hFED9441C , 32'h06E090A8 , 32'h02442F18 , 32'h063439A8 , 32'hFAB21E30 , 32'hFF1B6098 , 32'hFCEB56FC , 32'hFCD0C5AC , 32'hFF7706BD , 32'hFF471010 , 32'hFB2B3EF8 , 32'hFE4228C0 , 32'hFCDE1208 , 32'hFCB00728 , 32'hFEA151E4 , 32'hFCF31C40 , 32'hFB7C3BD8 , 32'hF9620438 , 32'h06B0EDB8 , 32'h0075A29F , 32'h045A2248 , 32'hFE9F64E0 , 32'h01ACDEDC , 32'h00611CDE , 32'hFCDFAD68 , 32'hFC7EA67C , 32'h01DAC384 , 32'hFFBC87EE , 32'h00B1EDB3 , 32'h00972FCF , 32'hFC0E5D4C , 32'hFE64B01C , 32'h002A8D45 , 32'h0000BBE2 , 32'h000498F3 , 32'hFFFFCB64 , 32'h00007986 , 32'hFFFEFA86 , 32'h0001701B , 32'hFFFE7D44 , 32'h00004178 , 32'h00002520 , 32'h0000C21A} , 
{32'hFFFFD93E , 32'hFFFCB7BB , 32'h0000CA1C , 32'hFFFDA240 , 32'hFFFFA812 , 32'hFFFF8677 , 32'h0000C3F5 , 32'hFFF9BFD9 , 32'h0002668B , 32'hFFFD9CE6 , 32'hFFFF5EC9 , 32'hFFFF50CE , 32'hFFFD4E8D , 32'hFFFFCB2C , 32'hFFFE87C6 , 32'h000099AF , 32'hFFFE378F , 32'hFFFDA9A6 , 32'hFFFD4C7A , 32'h00018D8D , 32'hFFFDB03F , 32'h0001EEF0 , 32'h0001599B , 32'h000146CA , 32'hFFFDEC04 , 32'hFFFDCE94 , 32'h0001C261 , 32'h0003C979 , 32'hFFFCA3AE , 32'h0002AFA9 , 32'h00014718 , 32'hFFFCB371 , 32'hFFFFADC7 , 32'hFFFF7417 , 32'h0001026B , 32'hFFFE29B6 , 32'h0000501D , 32'hFFF9EF83 , 32'hFFFBF551 , 32'hFFFC0D2A , 32'h0001BF5D , 32'h00028706 , 32'h0003D1C8 , 32'h000117E0 , 32'hFFFC5CE9 , 32'h00015113 , 32'hFFFF8AE7 , 32'hFFFBC550 , 32'hFFFDEA06 , 32'hFFFDA4CA , 32'h00009A68 , 32'hFFFF47F9 , 32'h00001FD6 , 32'hFFFE7392 , 32'h00048AD4 , 32'h0001FEB4 , 32'h00009E47 , 32'hFFFBA2D3 , 32'hFFFEC9CD , 32'hFFFA1B5B , 32'hFFFE1655 , 32'hFFFFDB03 , 32'h000630EE , 32'h00007059 , 32'hFFFE5EF6 , 32'hFFFB5C6B , 32'h00008B06 , 32'hFFFECF4C , 32'h00054F01 , 32'h000092A5 , 32'hFFFF4092 , 32'hFFFB7195 , 32'hFFFDCDA3 , 32'hFFFF260F , 32'hFFFE625A , 32'h0000F5A1 , 32'hFFFFD579 , 32'hFFFD0E66 , 32'hFFFE8FBF , 32'h0000C268 , 32'hFFF94A70 , 32'h0004BE9F , 32'hFFFFB5CA , 32'h0002058F , 32'hFFFD7061 , 32'h00008536 , 32'hFFFFA374 , 32'hFFFEF449 , 32'h0001CD71 , 32'h0004B4FA , 32'h0001A9F8 , 32'hFFFF137B , 32'h000076E4 , 32'h00043F06 , 32'h00022BD8 , 32'h0002CEDA , 32'hFFFF3BE5 , 32'hFFFF02C1 , 32'hFFFEE401 , 32'hFFFEE682} , 
{32'h299F6B80 , 32'h04A9D8C8 , 32'hE9834360 , 32'hBD7C2D80 , 32'h0B5F6740 , 32'hE8A40C40 , 32'hC5A2E180 , 32'hF37E1AB0 , 32'hED9F3EA0 , 32'h036B8280 , 32'hFBC34FE0 , 32'h195310A0 , 32'hEBB64F00 , 32'h0151A33C , 32'h05F2A358 , 32'h0C0EEA30 , 32'hE8599920 , 32'hE7EDC940 , 32'h09B88FD0 , 32'h21CCF400 , 32'hFC7FC5CC , 32'h14701060 , 32'h01C5DC60 , 32'hF88CD9B0 , 32'hFBEA05B8 , 32'hF5D0C130 , 32'h08DA79C0 , 32'hFF969F06 , 32'hFD1AB1A0 , 32'h02788260 , 32'h0A61C390 , 32'hFB136AB0 , 32'h0569BCB0 , 32'h055EBC70 , 32'hFF61E659 , 32'hFEC30BB4 , 32'h09689E30 , 32'hFE8C205C , 32'h0534C048 , 32'hFD3FD578 , 32'hF9952FB0 , 32'hFD1CFD90 , 32'h16901AE0 , 32'hFF6F1BA4 , 32'hFDD3C58C , 32'h0E40BE20 , 32'hF223B600 , 32'hFEB92938 , 32'hF4EE2ED0 , 32'h0C557800 , 32'h05EE6AC8 , 32'hF2BF79F0 , 32'hFE10F824 , 32'hF9DC8178 , 32'h11611A60 , 32'h02850EBC , 32'h02F85C90 , 32'hF38DB700 , 32'hFEF83EF4 , 32'h063B42D8 , 32'h00D65B0E , 32'h09C20BD0 , 32'hFCD9FFF0 , 32'h052E8878 , 32'h052170E0 , 32'hFF6FC8BC , 32'hF9E1F2F8 , 32'hF3ED6860 , 32'h04A20540 , 32'hFD865B14 , 32'h05126F88 , 32'h01936C54 , 32'h00CD44E3 , 32'hFD309388 , 32'hFC0F7314 , 32'hFE63384C , 32'h047BCF50 , 32'h01B7F39C , 32'hFD06BC24 , 32'hFE67F3B0 , 32'h0192FC70 , 32'h03E5A350 , 32'hFDED6CA0 , 32'h00F03B05 , 32'hFE185D48 , 32'h00E2CD3A , 32'h012CF9B8 , 32'hFEA132F0 , 32'h019A6CAC , 32'hFFD95ED4 , 32'h00013AAB , 32'h00001013 , 32'h00008C9B , 32'hFFFF384D , 32'hFFFE3DCD , 32'h00010496 , 32'hFFFFD54A , 32'h00008200 , 32'hFFFF855B , 32'hFFFF604E} , 
{32'hDC48C540 , 32'h3AEEC340 , 32'hFAE37100 , 32'h53782080 , 32'h253B2F00 , 32'hE07C05E0 , 32'h26F43D80 , 32'hB8401C00 , 32'h08975AF0 , 32'hCA3CB580 , 32'h00DCF2AA , 32'hEC58E780 , 32'h1C6DDB20 , 32'hE60C1A20 , 32'hEE4E1760 , 32'h05E82E68 , 32'hF90EA828 , 32'h05804F38 , 32'h1CAB1900 , 32'hF38A55D0 , 32'hF3615540 , 32'h0FDB5B80 , 32'h011510D8 , 32'hED4435E0 , 32'h15EC5520 , 32'hE9993C40 , 32'h0087465B , 32'h0AF9B730 , 32'hFBF212F8 , 32'h0E072E60 , 32'h113D1FA0 , 32'hFCBE1A38 , 32'hFEB49418 , 32'hEF923800 , 32'h01B4978C , 32'hFF09045C , 32'hF44BF0E0 , 32'hFE693368 , 32'h0AE31440 , 32'hFFFB8900 , 32'hFEA0B9C0 , 32'hFC208504 , 32'h0DA06E40 , 32'hFB7DD720 , 32'h0294BBA8 , 32'hF778CDD0 , 32'hFBEEE628 , 32'hF90BD460 , 32'hFE40FAA0 , 32'hF96D9650 , 32'hFCC857B4 , 32'hFA1A45A8 , 32'h0385948C , 32'hFE6CF344 , 32'h05C85A40 , 32'hF4279430 , 32'h011DCD10 , 32'hFBD95B68 , 32'hFC1C3B10 , 32'h005C6C66 , 32'h07A0DD98 , 32'h01D0C218 , 32'h00185EFD , 32'hFED3BA0C , 32'h00434380 , 32'h031051C0 , 32'h003DD91C , 32'h04891888 , 32'hFDE11454 , 32'h04A6C2B8 , 32'h013062FC , 32'hFD628724 , 32'h03D05308 , 32'hFE708AE8 , 32'h01FE86C4 , 32'hFB6642C0 , 32'hFFBE8605 , 32'h0253588C , 32'hFE5340AC , 32'h01893530 , 32'h04F0F1A0 , 32'hFE694D14 , 32'hFCA860CC , 32'hFE57CADC , 32'hFEC40F88 , 32'h01017D40 , 32'hFD3DD7A0 , 32'hFED10EA4 , 32'hFFAE0C24 , 32'h0066AA70 , 32'h0002C9B8 , 32'h00010353 , 32'hFFFE4A15 , 32'hFFFDAF8D , 32'hFFFF4B12 , 32'hFFFF9F14 , 32'hFFFEE6A4 , 32'hFFFF461C , 32'hFFFD32E1 , 32'hFFFDAE97} , 
{32'h2EAFDD40 , 32'h0B628280 , 32'h1234F7E0 , 32'hED0AF6E0 , 32'h1C869540 , 32'hEDFF4BC0 , 32'hF9BBD328 , 32'hF1B182D0 , 32'h0446E030 , 32'h02CC402C , 32'h19CDAEC0 , 32'h2E6BBE40 , 32'hF8DD4450 , 32'h08C17A30 , 32'hF6BCA060 , 32'h01F0EF88 , 32'hF6E9E200 , 32'hF16CA2C0 , 32'h04A143C8 , 32'h026DC800 , 32'h02C0CEF4 , 32'hFC0646CC , 32'h05963480 , 32'h02B98D90 , 32'h036CC040 , 32'h099564B0 , 32'hF0DA38C0 , 32'hFAD54BF8 , 32'hFC093698 , 32'h0A081310 , 32'h03C005E0 , 32'hFFC1320D , 32'h0275E268 , 32'h0E3D34C0 , 32'hFB80ABF0 , 32'hF0ACA890 , 32'hFDD4E104 , 32'hF8F40D90 , 32'h06135A00 , 32'h05FCF1C8 , 32'h04FB5E40 , 32'h014D4EF4 , 32'hFEE28430 , 32'h072BD110 , 32'hFE2ED58C , 32'h031876AC , 32'h00B47FC3 , 32'hFF6D0E22 , 32'h0C37EF10 , 32'h0741F1C0 , 32'hF5EEB920 , 32'h02835458 , 32'hFE9929EC , 32'hF9C77F90 , 32'h00501015 , 32'hF78A68F0 , 32'hF2055670 , 32'h0C457920 , 32'hF2A68E60 , 32'hF3C06270 , 32'hFFE5F2E2 , 32'h022B4E54 , 32'h045E5530 , 32'h03726DAC , 32'h06AE7578 , 32'h0AFDEE00 , 32'h0616D3D0 , 32'hF93108B8 , 32'hF9017760 , 32'h0626F728 , 32'hFF49378E , 32'hFF9A6615 , 32'h0AA3EAA0 , 32'h063586A8 , 32'h03085C4C , 32'hFF634B8D , 32'h03DD134C , 32'hF99D9648 , 32'h03533750 , 32'hFA5F3178 , 32'hF95128E0 , 32'hFBDA3D90 , 32'hFE4B7560 , 32'h01D1C204 , 32'h02B87038 , 32'h000819DC , 32'h000B558A , 32'h033649FC , 32'h00143860 , 32'hFFE6670E , 32'hFFFECEE6 , 32'h0003BB58 , 32'h00026FA7 , 32'h0001109B , 32'hFFFFE458 , 32'hFFFF215E , 32'hFFFF6489 , 32'h00006CDC , 32'h00007BDA , 32'hFFFEAD04}
};

logic signed [31:0] US_3 [100][10] ='{
{32'hF4EEF580 , 32'hD30DD3C0 , 32'hC14D1640 , 32'hF4BF6F10 , 32'h44AA9900 , 32'h16E95AE0 , 32'h07986A40 , 32'hEC87F020 , 32'h1719EE60 , 32'hE380A2A0} , 
{32'h422E4A80 , 32'hD55E4000 , 32'h1C62E7E0 , 32'hF8372F50 , 32'hD012CA00 , 32'hF905D5D0 , 32'hFED427D0 , 32'h02C7A5A4 , 32'h16140760 , 32'h01E138C0} , 
{32'h1D82D8E0 , 32'h007F8A4E , 32'hD8448640 , 32'h33014140 , 32'h01165CE0 , 32'hD75132C0 , 32'h464B8280 , 32'hEA134BC0 , 32'h0881B1E0 , 32'h015B1EF8} , 
{32'h00016954 , 32'hFFFF66EE , 32'h00016B36 , 32'h0004B634 , 32'h000521E3 , 32'hFFF9FC69 , 32'h0003A13D , 32'hFFFFDD00 , 32'hFFFDE86D , 32'h00059EA9} , 
{32'hFFFBE89F , 32'h00057D13 , 32'hFFFE67E1 , 32'hFFFF86B6 , 32'hFFFFD67C , 32'hFFFEF224 , 32'hFFFB7D87 , 32'hFFFDE439 , 32'h000198E5 , 32'hFFFF59A2} , 
{32'h024EC018 , 32'h48387200 , 32'hBF958680 , 32'hF729D830 , 32'h176C3DA0 , 32'h1BA178A0 , 32'hD9721AC0 , 32'hEABAAC60 , 32'hE5A6F9E0 , 32'hF426B2D0} , 
{32'h36860440 , 32'h24A47BC0 , 32'h0B215FD0 , 32'hF8BDB310 , 32'h0726D6A8 , 32'h01E1E4E4 , 32'hFB1AB7F0 , 32'h20B4F640 , 32'hF84476C0 , 32'hF63CE460} , 
{32'hFAA8E5B8 , 32'h3A841D00 , 32'h23A24780 , 32'hFB2455B8 , 32'hB2A02C80 , 32'h1E0FB3A0 , 32'h14436620 , 32'h2201B600 , 32'h15A1F120 , 32'hE2C3F7A0} , 
{32'hFFFFD7A1 , 32'h0007F1FF , 32'hFFFF2410 , 32'hFFFCDF7A , 32'hFFFC316F , 32'h00011199 , 32'hFFFC1DE3 , 32'hFFFC8EBC , 32'hFFFCC96C , 32'h000559D1} , 
{32'hFFECAF05 , 32'hEF37F9E0 , 32'h567A5C80 , 32'h5204FB00 , 32'hE51EE660 , 32'h234C20C0 , 32'h0647CB30 , 32'hF9607478 , 32'h010A2458 , 32'hE5D2DC80} , 
{32'h0F4AD050 , 32'h1FBE31E0 , 32'hD35D7280 , 32'hD7C122C0 , 32'h0B58B6F0 , 32'h05404438 , 32'h13314340 , 32'hCE67EF40 , 32'hF5F11660 , 32'hFC81A1B4} , 
{32'hD619E0C0 , 32'h408E6100 , 32'hD0FDE6C0 , 32'hE8ABE5A0 , 32'hEF1DC4C0 , 32'hEA8C0920 , 32'h40CE1680 , 32'h0A5D26E0 , 32'hF38A8AD0 , 32'hF6FFBFE0} , 
{32'h01C1A1B8 , 32'hB4288100 , 32'h355AB340 , 32'h4D6ACC00 , 32'h38DE0D40 , 32'hE91B0640 , 32'h33E84B40 , 32'hECF09E80 , 32'hF5F25030 , 32'hEE349E80} , 
{32'h11B75DA0 , 32'h2881DC00 , 32'h2FB95900 , 32'h0401BB68 , 32'hDB929A80 , 32'hFCBB2284 , 32'h02315A34 , 32'hFCB8A6FC , 32'hEE252120 , 32'hDD35A780} , 
{32'hEC890820 , 32'hC666CB80 , 32'hE3796520 , 32'hF62E0930 , 32'h0629F7F8 , 32'hDC67FF00 , 32'hEBFF2BC0 , 32'h17DF1840 , 32'h2B8ABFC0 , 32'hE04D15E0} , 
{32'h067405D0 , 32'hE9441640 , 32'h13EE6260 , 32'hB0959B00 , 32'hDE10F7C0 , 32'h04ACCC88 , 32'hE8C49D60 , 32'h347CBB80 , 32'h0F0377D0 , 32'hF6334740} , 
{32'h5D2FE880 , 32'hFBC3B228 , 32'h097B2870 , 32'hE2629B80 , 32'hDAA624C0 , 32'hF95F4028 , 32'h276166C0 , 32'h26DDD900 , 32'h05FA0DA8 , 32'hEFF78040} , 
{32'h2DB426C0 , 32'hF7EEC530 , 32'hE30A7360 , 32'h2F43A380 , 32'hE5020180 , 32'hD4677580 , 32'h1033D280 , 32'h31166AC0 , 32'hFF2AB3E5 , 32'hEA7D4000} , 
{32'h3D7439C0 , 32'hD6BDF840 , 32'hFDE25478 , 32'hFC605614 , 32'hEAE9D980 , 32'hCE451F40 , 32'hC8508240 , 32'h0D52C4C0 , 32'hE2777D80 , 32'hE2C46E80} , 
{32'h0000A43B , 32'h0001EB4D , 32'h000209BA , 32'h0000B274 , 32'h00022EB1 , 32'hFFFE31D5 , 32'h0001C16C , 32'h00034754 , 32'h00001BD1 , 32'hFFFEB9B7} , 
{32'h3C5C0540 , 32'h44691880 , 32'h31C62C00 , 32'h16B1D5A0 , 32'h12413CE0 , 32'hF3F854C0 , 32'hFA381D88 , 32'hC1C36B00 , 32'h0F519970 , 32'hD60CA480} , 
{32'hE7774720 , 32'h0DEE1290 , 32'h3394F600 , 32'hD6959940 , 32'hFAEC55C8 , 32'hBBA33580 , 32'hF21E7090 , 32'hF2C516E0 , 32'h0F2D5620 , 32'hEACAF9E0} , 
{32'h22D4D540 , 32'hBED9D480 , 32'h10F48780 , 32'hC0317B40 , 32'hF6CE9460 , 32'h179DEF60 , 32'hFED027A8 , 32'hFBF7B0A0 , 32'h0198BBB8 , 32'hFD46E7A0} , 
{32'h00025E9C , 32'h0000BA33 , 32'h0000F41A , 32'h0001B00C , 32'hFFFE43BA , 32'hFFFB8B0B , 32'h0004A791 , 32'h00010411 , 32'h000418C3 , 32'hFFFE62AA} , 
{32'h7FFFF800 , 32'h14506EC0 , 32'hD662D380 , 32'hF9131F38 , 32'h07861328 , 32'h1E101DA0 , 32'hF443FCA0 , 32'hF5AD5020 , 32'h2E2D0540 , 32'hE918B0E0} , 
{32'h23ED7900 , 32'h4C266300 , 32'hF8810578 , 32'h0DE26AE0 , 32'h2D5FD500 , 32'h189389A0 , 32'hF7C33740 , 32'hFF2C5E54 , 32'h05CE2AC8 , 32'hF5778010} , 
{32'h170B2580 , 32'h1BBA6EE0 , 32'hFDA46F3C , 32'h05384BB8 , 32'h2A2BA900 , 32'hEA63B580 , 32'h0C66AC70 , 32'h0A4AB320 , 32'h23F33C40 , 32'hF2158610} , 
{32'h1ACE2E20 , 32'h15FC0F20 , 32'h12A62800 , 32'hEEF25560 , 32'h011D1F9C , 32'hF6FC6C10 , 32'hE79A3BA0 , 32'hEC10A520 , 32'hE583AD60 , 32'hF6F1D7D0} , 
{32'hF9964670 , 32'hE8FDBFA0 , 32'hEFC88C60 , 32'hDD0484C0 , 32'hF88F1F58 , 32'h18CEBA60 , 32'hE4611000 , 32'h2BF24000 , 32'hDF3AF540 , 32'h0EFAB140} , 
{32'hD4D83AC0 , 32'hEF824F20 , 32'hBB048F80 , 32'hF75B8BE0 , 32'h14357420 , 32'hFDE065A8 , 32'h1DDC9340 , 32'hCFA8A7C0 , 32'hD218C540 , 32'hE2E22C80} , 
{32'h54A3FE80 , 32'h210040C0 , 32'h3EA24D00 , 32'hEE9E2760 , 32'hF1170110 , 32'hEF8CE560 , 32'h2BC6C9C0 , 32'h0DD95530 , 32'hC0050D40 , 32'hD7448CC0} , 
{32'h34018800 , 32'hC27BC140 , 32'h341BAF40 , 32'hF8773D80 , 32'hEFB63CE0 , 32'h2429B000 , 32'h0DD8EE40 , 32'hE2937F80 , 32'hCCCF32C0 , 32'h00B88967} , 
{32'hA1B8A000 , 32'h1C2AD800 , 32'h1D349FC0 , 32'h1F3F6020 , 32'h15185D80 , 32'hE6AA34C0 , 32'h249F8880 , 32'h1BCE4E40 , 32'h164A2920 , 32'hF03E2790} , 
{32'hB4517D00 , 32'hFE643458 , 32'h358CAEC0 , 32'hD61F8780 , 32'h34371AC0 , 32'hC61B8A80 , 32'h4E617480 , 32'h38EC2080 , 32'h0315706C , 32'hF0FEC340} , 
{32'hFFFD4E0B , 32'h00020EA7 , 32'h00041E52 , 32'hFFFA3EC6 , 32'h0004B6DB , 32'hFFFFEC19 , 32'hFFFE264F , 32'hFFFA7A83 , 32'h0004AFC9 , 32'h0001EDBA} , 
{32'hFAD071B8 , 32'hC95EBC00 , 32'hEF0A3860 , 32'h13F011C0 , 32'h21F09840 , 32'hBAD59500 , 32'h0194E5B4 , 32'hFFC1EDB7 , 32'hF8CAF4C0 , 32'hF5214BA0} , 
{32'hF1743A90 , 32'hEE12A8C0 , 32'hD0261BC0 , 32'h0A7165D0 , 32'h1E5CF0E0 , 32'h122DBCE0 , 32'h1D058820 , 32'hECBA2640 , 32'h0530D220 , 32'hFF80D6A7} , 
{32'h02CA812C , 32'hC67EC0C0 , 32'h4589EA00 , 32'hC4A7BA40 , 32'hF54ECD20 , 32'h2F4C9B80 , 32'hF6550EB0 , 32'hEF0AE460 , 32'h0F886A00 , 32'hF0295250} , 
{32'h25D55AC0 , 32'hD4E33740 , 32'h092AFD40 , 32'hD2340B80 , 32'h156C2EC0 , 32'hF85C5B70 , 32'hE0A8F9A0 , 32'h0B702490 , 32'h2A4CA780 , 32'hF20C4EE0} , 
{32'h2CC45B80 , 32'hCFBA1C00 , 32'hFDEAE860 , 32'hD9A14AC0 , 32'h154B26E0 , 32'h2D52F680 , 32'hF98EFE38 , 32'h12EDFAA0 , 32'hE671C620 , 32'hF8B948C0} , 
{32'hD8A9D5C0 , 32'h20ED0C40 , 32'h3F7533C0 , 32'h0326527C , 32'hDDFE5BC0 , 32'h1964F6A0 , 32'h11045CE0 , 32'hC4F14CC0 , 32'h239AF8C0 , 32'hF7F67370} , 
{32'h011913D4 , 32'hFDEFB8B8 , 32'hFB1CEFB8 , 32'h04FE8470 , 32'h007EDBDF , 32'hFB04A150 , 32'hFFA6F778 , 32'h0265B180 , 32'hF9798E98 , 32'hFBD4A200} , 
{32'hF9A3A5F0 , 32'h0E5D8C30 , 32'h094361B0 , 32'h13ED3340 , 32'hFC071DD8 , 32'h050425E0 , 32'hF78BF3C0 , 32'h0B94D1D0 , 32'hE366F9A0 , 32'h01A568BC} , 
{32'hE30B8CA0 , 32'hEDBE2940 , 32'h37420BC0 , 32'hF482A3C0 , 32'h38BC7180 , 32'hDCFF4500 , 32'hE4E13B00 , 32'hEAF94280 , 32'h16897520 , 32'hEEEAC9A0} , 
{32'hF77FA5F0 , 32'h0B41B7F0 , 32'hA2E0B880 , 32'hFB98AD80 , 32'hB8F41980 , 32'hF57E2EB0 , 32'h0126CD60 , 32'h205D4180 , 32'h28102540 , 32'hF4463850} , 
{32'hE81F6D80 , 32'h16402740 , 32'hC72DD300 , 32'hE23F6900 , 32'hDC89FB40 , 32'h1CCD3BC0 , 32'h37234C00 , 32'h00B901E7 , 32'h12F18280 , 32'h00669950} , 
{32'h0329FBD8 , 32'h9E0F7780 , 32'hF9FA3D78 , 32'h0D9B5460 , 32'h19901860 , 32'hF71658C0 , 32'h24640B80 , 32'hEF5618A0 , 32'hC9A5CF00 , 32'hF1078EC0} , 
{32'h348BC680 , 32'hF5E05C70 , 32'hEE3CCD00 , 32'h46309A00 , 32'hDC579000 , 32'hE5E16120 , 32'hEA28E080 , 32'h0FB93360 , 32'hD8D28140 , 32'hEEC18D80} , 
{32'hF9DC95F0 , 32'h57C6C300 , 32'h07AFC930 , 32'hF19979F0 , 32'h0E214150 , 32'h1B431360 , 32'h2B1E8700 , 32'h2CB5B340 , 32'hF73B8E80 , 32'hEDC4F060} , 
{32'hC9B143C0 , 32'h3A429040 , 32'hF3A5B920 , 32'hDA4A1D80 , 32'hCF178080 , 32'h0F8FC920 , 32'h1AF504E0 , 32'hC8E77C00 , 32'h191AC2E0 , 32'hF1D0D320} , 
{32'hFD671554 , 32'h23B755C0 , 32'h1E07DF40 , 32'h03E941C0 , 32'h4FE10880 , 32'hF7AAA7B0 , 32'hF7BB6A10 , 32'hCA98C680 , 32'h0D4E3A00 , 32'hE7095660} , 
{32'hF517CFB0 , 32'hE5984C00 , 32'hDC711EC0 , 32'hEB6F0340 , 32'h3C65F800 , 32'h37AB1B80 , 32'h3B19C180 , 32'hF7C06B70 , 32'h21D1E300 , 32'hF32D10F0} , 
{32'h312BD380 , 32'hD8BD8140 , 32'hDAE020C0 , 32'h4EABF980 , 32'hD1F85F80 , 32'h0039BE91 , 32'h144B56C0 , 32'h133083E0 , 32'h181E8040 , 32'hFC270C80} , 
{32'hDAE36180 , 32'h0CE02150 , 32'h00BD8A3A , 32'h27391080 , 32'hFEBEAB34 , 32'h1F7C40C0 , 32'hF0A2F410 , 32'h35665EC0 , 32'hDD352100 , 32'hFC7A9C10} , 
{32'hF295C6B0 , 32'h09126760 , 32'h0640D6F0 , 32'hEEC96CC0 , 32'h2A387F00 , 32'hDE3C3740 , 32'hDDE6D500 , 32'h250F3080 , 32'hF91489C0 , 32'hF7F17DB0} , 
{32'hEB4517A0 , 32'h0F680110 , 32'hDA303480 , 32'hF63B8A90 , 32'hFB9BF770 , 32'h07F59788 , 32'hC9DC13C0 , 32'hF9125F20 , 32'h0736A088 , 32'hFA524280} , 
{32'hCF1B6880 , 32'hEDBD0BA0 , 32'hC71BBD40 , 32'hC84D5F80 , 32'hEC27C4E0 , 32'hCDD14700 , 32'hC49BF840 , 32'hF7EAED40 , 32'hE65EBF40 , 32'hDA64EDC0} , 
{32'h13722880 , 32'h02869C44 , 32'hB3D5C600 , 32'h3A96E300 , 32'hC21BAA80 , 32'h05215618 , 32'hFA37FB50 , 32'h06D53AA8 , 32'hF878D448 , 32'hF1A7C330} , 
{32'hDAA65FC0 , 32'h19074580 , 32'h259F17C0 , 32'h28CD58C0 , 32'hD83C74C0 , 32'h0BE7C940 , 32'h02FDF86C , 32'hF596DAD0 , 32'h0CE24250 , 32'hF2B06790} , 
{32'hC31B0600 , 32'h338B6240 , 32'hDE7C4180 , 32'hFF0F406D , 32'hD2D2E500 , 32'hCDD7B300 , 32'h1B0DC640 , 32'hE734D200 , 32'hD9070800 , 32'hEA5B3960} , 
{32'hF132A940 , 32'hB4AB7D80 , 32'hB6F02200 , 32'hDF545580 , 32'h10D91A40 , 32'h118FE9A0 , 32'hFBD56628 , 32'h214D7FC0 , 32'hF9B03478 , 32'hF34312B0} , 
{32'h04DF0EC0 , 32'hEFE99340 , 32'hE62B6900 , 32'h0268CD18 , 32'h360EAEC0 , 32'h2208DFC0 , 32'hF2389580 , 32'hDB160700 , 32'hF2D10C60 , 32'h0481A210} , 
{32'hFA6E5EE0 , 32'hFA0471A0 , 32'hFFB97694 , 32'hC8FB23C0 , 32'h03CD0A84 , 32'hF9F72E20 , 32'h62EC0800 , 32'h09ADFE00 , 32'h0760B1C0 , 32'hF185F9E0} , 
{32'hDE4A3B80 , 32'hE6DE73E0 , 32'hE21458E0 , 32'hE7CFA200 , 32'h0B3D3180 , 32'hF17E0C50 , 32'h05CE36A0 , 32'hED273480 , 32'hFBF13428 , 32'hF3D63970} , 
{32'h2B4DFC40 , 32'hEECC9220 , 32'hCA270400 , 32'h007D4651 , 32'h0B86B5B0 , 32'h320FA900 , 32'hE9D6BA80 , 32'hF0B3C1C0 , 32'h0C623480 , 32'hF4A6B7D0} , 
{32'hC1885880 , 32'hD0A97540 , 32'h053008D0 , 32'h009D1D21 , 32'hBC9A9580 , 32'h32FF6900 , 32'hF4FECCF0 , 32'hF17E1650 , 32'hF63DE060 , 32'hE57D9380} , 
{32'hFFFD7953 , 32'hFFFD7F4E , 32'h00030CB7 , 32'h000051A5 , 32'hFFFBE3A6 , 32'h00020842 , 32'hFFFC49F2 , 32'hFFFD9EE0 , 32'h000407C4 , 32'hFFFA1056} , 
{32'h20906F80 , 32'hFB405210 , 32'hEC8B3C80 , 32'h283F5DC0 , 32'h0DA28F80 , 32'hEBB322C0 , 32'h1D456680 , 32'h0AABE880 , 32'hD832D640 , 32'hE809B5E0} , 
{32'h027536E4 , 32'hEC751860 , 32'h06A2BCA0 , 32'hEDAAFD60 , 32'hEE6F5060 , 32'h0D0FF270 , 32'h1FC95C80 , 32'hF7E30C60 , 32'hF40C2B70 , 32'hF9293F58} , 
{32'h0917A680 , 32'hE011FA20 , 32'hC9FE0680 , 32'h266BA540 , 32'h034277C0 , 32'h1B02C080 , 32'h1824B360 , 32'h12AFE3A0 , 32'hF7725E60 , 32'hECA62CC0} , 
{32'hE9B98EC0 , 32'hFFBD915E , 32'h1A6EFF80 , 32'h071CB188 , 32'h28417200 , 32'h196D3CE0 , 32'h03A1C7C0 , 32'h32A64280 , 32'h00809090 , 32'hEB76DC80} , 
{32'h0A664510 , 32'h11B4A420 , 32'hF4D6EAE0 , 32'h358EF440 , 32'hECCB1820 , 32'h0C631A40 , 32'h14CCA880 , 32'h1B6C53A0 , 32'h0DCE0AA0 , 32'hF3F68B40} , 
{32'h0C671080 , 32'h31CCB540 , 32'h02B758D8 , 32'hFC385174 , 32'h30D6AC80 , 32'h32BCC0C0 , 32'hEEF2D5A0 , 32'hF3010060 , 32'hF08017D0 , 32'hEA7078C0} , 
{32'h06544F90 , 32'hEFEB2060 , 32'h04DCB428 , 32'hDEE4AB80 , 32'hF0BABFA0 , 32'hD4C6E100 , 32'h10091440 , 32'hEBB7B000 , 32'hF723A4E0 , 32'hFC664D70} , 
{32'h162926A0 , 32'hFEED9EAC , 32'h050082B8 , 32'h2A5701C0 , 32'h0F8BEBB0 , 32'h242DB6C0 , 32'h2229BFC0 , 32'h362BD240 , 32'h1B92FFC0 , 32'hE08CDAC0} , 
{32'h11106DE0 , 32'hF70BC250 , 32'h36D67780 , 32'hE3AB7A20 , 32'h0BB8B000 , 32'hE92A8D40 , 32'hE748C5A0 , 32'h0C3B0CC0 , 32'hEEE4E240 , 32'hFB236E08} , 
{32'hDD1C75C0 , 32'h1EF3C060 , 32'h3AE244C0 , 32'h0739F120 , 32'h037905AC , 32'h144DA3A0 , 32'h0E793A50 , 32'hFE59EE98 , 32'h07B7EBF0 , 32'hFF812C62} , 
{32'h211C2E80 , 32'h36FBDC80 , 32'hDD7BF640 , 32'h24CE73C0 , 32'h1625E0A0 , 32'h32653840 , 32'hC973FA00 , 32'h0479DBA0 , 32'h095B6930 , 32'hDD898A00} , 
{32'hA3D7F780 , 32'hD42FA340 , 32'hF47413F0 , 32'hF2FA2450 , 32'hE1143BE0 , 32'hF90960C8 , 32'hDAA72200 , 32'hEB8B3640 , 32'h092ED690 , 32'hCF8F3DC0} , 
{32'h2D6E2880 , 32'hCAD68A40 , 32'h3E9AA000 , 32'h0E02F1B0 , 32'hF93FC6C0 , 32'hF4545D30 , 32'h08249AB0 , 32'hD1705740 , 32'h308F0740 , 32'hF664FD90} , 
{32'hB8E93A00 , 32'h02329270 , 32'h1332D4A0 , 32'h32141600 , 32'hEF85DC40 , 32'h0D4AA620 , 32'hCE0E7840 , 32'hFAAEDCD8 , 32'h09BCB770 , 32'hE3FF7140} , 
{32'hFFCBF7EA , 32'h2C64BD40 , 32'h1104FCE0 , 32'h5963C500 , 32'hCC731DC0 , 32'hDF852E80 , 32'hF2ADE1B0 , 32'hCBC76700 , 32'h11007000 , 32'h05FA1B48} , 
{32'hEBBD7EC0 , 32'h228D0AC0 , 32'h331D2E40 , 32'hD6BFDD80 , 32'hE9E38620 , 32'h22C96800 , 32'hE1D9C980 , 32'h07837080 , 32'hFB6A12B8 , 32'hEAD71060} , 
{32'hFFFEABC7 , 32'h00048C21 , 32'hFFFEE11C , 32'hFFFDBB9B , 32'h00038246 , 32'hFFFED6D8 , 32'hFFFCE852 , 32'hFFFCC120 , 32'h00016478 , 32'h00051F47} , 
{32'h0783A510 , 32'h47F47580 , 32'h026EEF18 , 32'h05778B58 , 32'h31A13D00 , 32'h2C5D12C0 , 32'h03A97F10 , 32'h0F20D260 , 32'hDF122BC0 , 32'hFCD48F98} , 
{32'hD58FDCC0 , 32'h147681C0 , 32'h350CFE00 , 32'h005A23FA , 32'h2A1C5740 , 32'h13B8D360 , 32'hE8673AA0 , 32'h4A3EE980 , 32'h160111A0 , 32'hEC35CE60} , 
{32'h3732BE40 , 32'h1609AAA0 , 32'hD13C02C0 , 32'h020B7D34 , 32'h2D956740 , 32'hFEEF09C4 , 32'h068A9960 , 32'h12AE5600 , 32'h46E12F00 , 32'hEAF05000} , 
{32'h5B9EB600 , 32'hFD68E574 , 32'hF6B2E040 , 32'hB5642300 , 32'hE5EC4520 , 32'h23550B80 , 32'h34554680 , 32'hC4086A80 , 32'hFFA89BB2 , 32'hF6F3CEF0} , 
{32'hD53917C0 , 32'h024FD624 , 32'hE2F4F5C0 , 32'hC1E81C80 , 32'hC1A81CC0 , 32'hF3384E20 , 32'h13AEB5A0 , 32'hFAA4FBC8 , 32'hFFFC5E5F , 32'hE7C60620} , 
{32'h00005366 , 32'h00014E3A , 32'h00012CA8 , 32'h00034CFB , 32'h0000DCF0 , 32'h0000E864 , 32'h000204FC , 32'h0006558C , 32'h000058AE , 32'h0000EFB9} , 
{32'h31AC5400 , 32'h04C9C358 , 32'h0C78DD50 , 32'hEAE3D7A0 , 32'h1EA674A0 , 32'hB6BA5D00 , 32'hEC3249C0 , 32'hFCD8AD94 , 32'h0B759F90 , 32'hF7B66800} , 
{32'hFD3083AC , 32'h13C7D5A0 , 32'h0E6F49D0 , 32'h01301278 , 32'h08D04790 , 32'h012BA140 , 32'h046299C0 , 32'h1A2C3FE0 , 32'h110A3520 , 32'h0A0F9470} , 
{32'h16F783E0 , 32'h3E5F1140 , 32'h08323BD0 , 32'h0476A670 , 32'h033F6110 , 32'h121888A0 , 32'hFCCE3824 , 32'hF15869F0 , 32'hCEB76B80 , 32'hFD7C3B70} , 
{32'h42D1CF80 , 32'h32E90B00 , 32'h00986514 , 32'hC9C88680 , 32'hF5526F40 , 32'hC582BE80 , 32'hF1E85FF0 , 32'hF1B452B0 , 32'h0C4DCCC0 , 32'hE50B71E0} , 
{32'hFFFD9193 , 32'hFFFAFDB6 , 32'h0000C1E1 , 32'hFFFC6F4B , 32'h000305D2 , 32'h00026547 , 32'h0003AA28 , 32'hFFFBE813 , 32'h0003C707 , 32'hFFF969D6} , 
{32'hFAC124F8 , 32'hC7D62800 , 32'hDCABF6C0 , 32'h3884E540 , 32'h192FE5A0 , 32'hE1420100 , 32'hF33729C0 , 32'hECE3E260 , 32'hF9999700 , 32'hD325B1C0} , 
{32'hD421A2C0 , 32'hB7B80A00 , 32'h0921C6F0 , 32'h24A7B940 , 32'hECE3F740 , 32'h1CF316C0 , 32'h004A57CB , 32'hE367E340 , 32'h44E8A080 , 32'h05D5BDF8} , 
{32'hF2215C50 , 32'h9AED6980 , 32'h308C2080 , 32'hFDA54578 , 32'hE0E9BD40 , 32'h4C3D0500 , 32'h09B38A00 , 32'h0B94AFA0 , 32'hE234A6A0 , 32'hD7C4D480} , 
{32'hE30C8A60 , 32'h295D8FC0 , 32'hDEDF6AC0 , 32'hE850AAA0 , 32'hF5ACF150 , 32'h04B552B0 , 32'hE6541700 , 32'h0AEBFD80 , 32'h14CF6900 , 32'hE3ED57C0} , 
{32'h4B362580 , 32'hEF359F80 , 32'h0FB56400 , 32'hF40291F0 , 32'hD4C33BC0 , 32'hE2DF8480 , 32'hFF513F0D , 32'h1B6F8360 , 32'h23656C40 , 32'h1362AD40}
};
logic signed [31:0] bias_0[37] = '{32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000};
logic signed [31:0] bias_1[300] = '{32'hE1D84140 , 32'h0D158350 , 32'hFB98EC28 , 32'h25F12780 , 32'hF36849A0 , 32'hFA4EC5A8 , 32'hFE3B6F98 , 32'hF7138BB0 , 32'hFABEE7D0 , 32'hF0703490 , 32'hECCBC760 , 32'h0CBC0FC0 , 32'h20CA9400 , 32'hFE52B9C8 , 32'hF1488380 , 32'h01B4F764 , 32'hFE09B4CC , 32'h06099C20 , 32'hD9F73F00 , 32'hFEF0CCC8 , 32'hFE2F9B20 , 32'hF6780B80 , 32'h260CA540 , 32'h065972A8 , 32'h15ABC340 , 32'hFEDBDF34 , 32'hFC4B9158 , 32'h026CB170 , 32'hFEBDFEBC , 32'h2E8C74C0 , 32'hFDB1A0CC , 32'h0B318D10 , 32'hE8CACE20 , 32'hF7F9F890 , 32'hFF09E04F , 32'h02FDBE08 , 32'h161D8700 , 32'hE79BC8E0 , 32'hF78BC980 , 32'h009C932A , 32'hEAA079C0 , 32'hF80EAAC8 , 32'hFE2207A0 , 32'h0527E240 , 32'h23D1D380 , 32'h28D89500 , 32'hFF969002 , 32'hFF12B725 , 32'h09B85E20 , 32'hF8467D60 , 32'hFAC5D180 , 32'hFCC3D6AC , 32'hF4E069A0 , 32'h11D58160 , 32'hF8C53338 , 32'hFF333EBE , 32'hFC6272DC , 32'hFAF7D138 , 32'hFEF91280 , 32'hC72D5A80 , 32'hFC633068 , 32'hFD266B50 , 32'hFAE36B18 , 32'hFEA94B70 , 32'h11C67C40 , 32'hFB33BB38 , 32'hF3D00270 , 32'h03047E3C , 32'hFE360C38 , 32'hDE3FFCC0 , 32'hF6B182E0 , 32'hE41C8CA0 , 32'hFD0B5C34 , 32'hFEDEFF6C , 32'hFDF8C040 , 32'hDA886B80 , 32'hF568AFE0 , 32'hFE66AA44 , 32'h148CDE80 , 32'hEEEEB620 , 32'hF4BB59C0 , 32'h1C2DF920 , 32'hF7EDAD00 , 32'hFC31731C , 32'hDA00EE80 , 32'h14310500 , 32'hD2FDDA00 , 32'hEFF26B80 , 32'hEB1E1980 , 32'hE25E97A0 , 32'hFE6E5D10 , 32'h1B24F9A0 , 32'hFD8D0B28 , 32'hDF0D3880 , 32'hED62D2C0 , 32'hFE3A35AC , 32'hFED3E354 , 32'hFD42E1A4 , 32'hF61CDFA0 , 32'h08A79B80 , 32'h1F027CE0 , 32'hFDF49114 , 32'hD8372B00 , 32'h078E1AA0 , 32'h2EDCF380 , 32'hFE637ECC , 32'hE497AB20 , 32'hFEA86618 , 32'h10CD2940 , 32'h28B32800 , 32'hFC5BC694 , 32'h2F015F80 , 32'hF3E95EF0 , 32'hF9A7C030 , 32'hDA6BDDC0 , 32'h0C21F940 , 32'hE05E0400 , 32'hFEE1DB1C , 32'h0903B5A0 , 32'hFCC3E5F8 , 32'hEF25A7A0 , 32'hFA145CD0 , 32'hED411C80 , 32'hF0E71F30 , 32'h0F15F790 , 32'hF9BB25A0 , 32'hFCD180D8 , 32'hFDF3CDAC , 32'hFEFEF07C , 32'hFBE706F0 , 32'hFCE24DA4 , 32'hFD114A80 , 32'h0B219360 , 32'hF9873C78 , 32'hFD054E10 , 32'h2A785C40 , 32'h0D7BB040 , 32'hFE702028 , 32'hFE70241C , 32'hEC71A060 , 32'hF7901690 , 32'hFE1E0FBC , 32'hFB417C60 , 32'h187F6000 , 32'h1CCFA780 , 32'hF48885A0 , 32'hF1241280 , 32'hFF0B346B , 32'hEE44AAC0 , 32'hF9749428 , 32'hF7298700 , 32'hE97A3780 , 32'hFED120AC , 32'hF81B4E30 , 32'hF3B69130 , 32'hFDB6F870 , 32'h092B1B90 , 32'hD2D128C0 , 32'hEFF2B160 , 32'hF9EE6658 , 32'hFDECA728 , 32'hD65A5580 , 32'hF987AA78 , 32'h0D1D8150 , 32'h0EE9CEE0 , 32'hFE17C024 , 32'h124E9600 , 32'hFAA61C20 , 32'hFBBCD0D8 , 32'hF2AF72E0 , 32'hE8908380 , 32'hF4B87C80 , 32'hFEAFAA8C , 32'hF6CB5720 , 32'hED168000 , 32'hE9C3B700 , 32'h18EAEC40 , 32'hEEBE68C0 , 32'h069C4E18 , 32'hF09D3990 , 32'hE8663760 , 32'hFDB63BF4 , 32'hF9CD8398 , 32'hFE7F11DC , 32'hF48300E0 , 32'h1ABC3340 , 32'hEC9277C0 , 32'hF9580B70 , 32'h2B922540 , 32'h146C77A0 , 32'hFE2B86F4 , 32'hE96A53E0 , 32'h11301EC0 , 32'hF70E9A70 , 32'hFA994518 , 32'hFEB4D7D4 , 32'hE7E880A0 , 32'hEA3DA240 , 32'hE739FFC0 , 32'hFCE3ECBC , 32'hFBB1C918 , 32'hFF055385 , 32'hFE7C1CD0 , 32'hFE52D810 , 32'hF39FAB50 , 32'hEFDA1420 , 32'h05B1E018 , 32'hFFDAB13D , 32'hEEE7B500 , 32'h038A36B8 , 32'hFF1B0F46 , 32'hFE787364 , 32'hFEE8D37C , 32'hF85D7780 , 32'hFD5DEFBC , 32'hEC881880 , 32'h03207BF4 , 32'h0E16E2A0 , 32'hFD994D0C , 32'hFEE5F214 , 32'hFCD963B4 , 32'hFD0EB268 , 32'h0A17C570 , 32'hF45E1A60 , 32'hFC691870 , 32'hFBD56EF0 , 32'hFD24326C , 32'hF1AD71B0 , 32'h116688E0 , 32'hEE6E62A0 , 32'hFEB596C8 , 32'hFF2815CF , 32'hFF207C80 , 32'hE2F73D80 , 32'h0928F0B0 , 32'hFEB38244 , 32'hFE9643A4 , 32'hF49DE8F0 , 32'hFE09F0B8 , 32'hD101E300 , 32'hFD9777B4 , 32'h26CEDAC0 , 32'hFE6713E8 , 32'hFFCD908F , 32'hF2B68140 , 32'hF009C870 , 32'h2A746740 , 32'hF8C1BA08 , 32'hEF427840 , 32'hE552E780 , 32'hFEBF9030 , 32'h2E29BD40 , 32'hF52D0CA0 , 32'h018D4A3C , 32'h0B52AE40 , 32'h1B5E8C80 , 32'hF1D41B90 , 32'hFCDB93A0 , 32'hF9DC0AD8 , 32'hF45EF730 , 32'h1338DC20 , 32'hEA000300 , 32'hDFF11800 , 32'hFD2E0580 , 32'hFD37C3DC , 32'hFEB828F4 , 32'hF6493B40 , 32'hF9FA8130 , 32'hE1951A80 , 32'h0A34F180 , 32'hFD5009C4 , 32'hFD950F20 , 32'hFF37B7C3 , 32'hEFD6C7A0 , 32'h1FD0F740 , 32'h0167D424 , 32'hFC83E29C , 32'h006D4D08 , 32'hD41A0900 , 32'hFD4AC058 , 32'hFE0CB884 , 32'hF2914250 , 32'hFBCE8FF8 , 32'hF7ABD1D0 , 32'hFC932C78 , 32'hEE992480 , 32'hCA653580 , 32'hF7204B00 , 32'h06DF8780 , 32'hDF02C440 , 32'hDB859640 , 32'hFDF98EB8 , 32'hFE94DA18 , 32'hF4F73260 , 32'h1642E860 , 32'hE5A18760 , 32'hF5F73B50 , 32'h091D3490 , 32'hF7CFB110 , 32'hFB1E7C88};
logic signed [31:0] bias_2[100] = '{32'h074D40A0 , 32'hFD2DD604 , 32'h0470DE18 , 32'hFF218263 , 32'hDC706D40 , 32'h4EB3CB80 , 32'h1DC92A40 , 32'h2A191340 , 32'hFD6344D0 , 32'hDED5DF40 , 32'h1788AE80 , 32'h05D74C78 , 32'hD26E6B80 , 32'h3AD08380 , 32'h070AF5A0 , 32'h1845AE60 , 32'h04546920 , 32'h22FE9B00 , 32'h238AC380 , 32'hFC97830C , 32'h068CAEC0 , 32'h275B6700 , 32'hE96E16C0 , 32'hFCDDC7EC , 32'hF95E1A30 , 32'h19B8CA80 , 32'h0271EEE8 , 32'h2C4D6AC0 , 32'h0FAD1970 , 32'h152E0040 , 32'hF7C7D850 , 32'hED1FBC20 , 32'hE5BDFB20 , 32'h00D57DFA , 32'hFF20CA3D , 32'hE3F913A0 , 32'hE0F4FB00 , 32'hCFB61DC0 , 32'hEBFFA840 , 32'hE73ABD80 , 32'hFCB1D728 , 32'hD53F6280 , 32'h25143D40 , 32'hEF4D4580 , 32'h437F1800 , 32'h0D44F990 , 32'hDF538540 , 32'h2AE1C040 , 32'h20C23F00 , 32'h2859B5C0 , 32'hFB8EA450 , 32'hF21DAE60 , 32'h07534BC0 , 32'h2DE8C400 , 32'h15A17980 , 32'h47952F00 , 32'h3B64B100 , 32'h435D8600 , 32'h13B1B920 , 32'h40E7D780 , 32'hF0911DA0 , 32'hF5C277F0 , 32'hD37BE000 , 32'h04422AD8 , 32'h0F39AFA0 , 32'h02B76720 , 32'hECD9B060 , 32'h021B7A28 , 32'hEDF67A80 , 32'h0264D7C0 , 32'hD985E800 , 32'h0BDA9F90 , 32'hFC3565C0 , 32'h0801A2B0 , 32'hE61A9A20 , 32'h057A1568 , 32'hED870EA0 , 32'h0A0C7780 , 32'h0BA8A970 , 32'hF932AF38 , 32'h338B7100 , 32'h162733A0 , 32'h29411300 , 32'hF9473E10 , 32'h0FC7A470 , 32'h1699A500 , 32'hF36E4A70 , 32'h01F813B8 , 32'h07B80388 , 32'hFBF1C490 , 32'h274C2FC0 , 32'hFEAE4D70 , 32'h2ED46440 , 32'h3B08B6C0 , 32'hFDC03FA4 , 32'hFACC7B48 , 32'h0E416040 , 32'hE6043B80 , 32'h36EDBB80 , 32'h21B92D40};
logic signed [31:0] bias_3[10] = '{32'hFAB601C8 , 32'hDE7F0AC0 , 32'hFADF11A0 , 32'hFF50128A , 32'h05E4BB58 , 32'hE47F7B00 , 32'h03D3D510 , 32'hD9AAB740 , 32'h4827FF00 , 32'h099F4220};


endpackage
