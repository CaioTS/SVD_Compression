

library ieee;
use ieee.std_logic_1164.all;

library ieee_proposed;
use ieee_proposed.fixed_pkg.all;

use work.types.all;
package weights_constants is

    constant weight_n0_0 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(0.00020837431657128036)),(to_sfixed_a(-5.5579595937160775e-05)),(to_sfixed_a(0.00022957788314670324)),(to_sfixed_a(0.0001543516991659999)),(to_sfixed_a(1.8413658835925162e-05)),(to_sfixed_a(-0.00027713910094462335)),(to_sfixed_a(-4.657112731365487e-05)),(to_sfixed_a(-6.366134039126337e-05)),(to_sfixed_a(0.0002088224864564836)),(to_sfixed_a(-0.00021181323972996324)),(to_sfixed_a(5.017388320993632e-05)),(to_sfixed_a(0.00010078861669171602)),(to_sfixed_a(-0.00010923944500973448)),(to_sfixed_a(9.457598207518458e-05)),(to_sfixed_a(-0.00011075839574914426)),(to_sfixed_a(-9.125762153416872e-05)),(to_sfixed_a(-0.0001889562699943781)),(to_sfixed_a(0.00011841711966553703)),(to_sfixed_a(0.00017176297842524946)),(to_sfixed_a(6.527895311592147e-05)),(to_sfixed_a(1.663063812884502e-05)),(to_sfixed_a(-2.1813075363752432e-05)),(to_sfixed_a(-0.0003393535444047302)),(to_sfixed_a(9.649692219682038e-05)),(to_sfixed_a(0.00015609536785632372)),(to_sfixed_a(6.68663124088198e-05)),(to_sfixed_a(0.00011015294876415282)),(to_sfixed_a(0.00035080386442132294)),(to_sfixed_a(-8.841504313750193e-05)),(to_sfixed_a(-0.00011197580170119181)),(to_sfixed_a(6.589842814719304e-05)),(to_sfixed_a(0.00011928956519113854)),(to_sfixed_a(-8.37730840430595e-06)),(to_sfixed_a(-3.526087311911397e-05)),(to_sfixed_a(-0.0002713542489800602)),(to_sfixed_a(0.00017650096560828388)),(to_sfixed_a(-5.0056467443937436e-05)),(to_sfixed_a(-4.927627742290497e-05)),(to_sfixed_a(2.7038928237743676e-05)),(to_sfixed_a(0.00012057880667271093)),(to_sfixed_a(0.00020322861382737756)),(to_sfixed_a(7.179802923928946e-05)),(to_sfixed_a(-7.964765245560557e-05)),(to_sfixed_a(0.0001670651836320758)),(to_sfixed_a(0.0004008085234090686)),(to_sfixed_a(-0.00017720619507599622)),(to_sfixed_a(0.0002220917958766222)),(to_sfixed_a(-0.00010266016033710912)),(to_sfixed_a(-0.00030316252377815545)),(to_sfixed_a(0.00015634181909263134)),(to_sfixed_a(6.916494385222904e-06)),(to_sfixed_a(-0.00028837472200393677)),(to_sfixed_a(0.00015752417675685138)),(to_sfixed_a(-0.0001657687098486349)),(to_sfixed_a(-4.022021312266588e-05)),(to_sfixed_a(-0.00021018224651925266)),(to_sfixed_a(0.00021029167692176998)),(to_sfixed_a(3.2542091503273696e-05)),(to_sfixed_a(-6.269387813517824e-05)),(to_sfixed_a(-7.831077527953312e-05)),(to_sfixed_a(0.0001649375190027058)),(to_sfixed_a(0.0002684917417354882)),(to_sfixed_a(-9.279272489948198e-05)),(to_sfixed_a(6.524159834953025e-05)),(to_sfixed_a(-4.041708052682225e-06)),(to_sfixed_a(2.848364965757355e-05)),(to_sfixed_a(2.78526130159662e-07)),(to_sfixed_a(-0.0001628674945095554)),(to_sfixed_a(0.00011417608766350895)),(to_sfixed_a(0.020731793716549873)),(to_sfixed_a(0.00013067442341707647)),(to_sfixed_a(4.7408752834599e-06)),(to_sfixed_a(3.3257149425480748e-06)),(to_sfixed_a(-0.00014872632164042443)),(to_sfixed_a(-7.416649896185845e-05)),(to_sfixed_a(-6.777828093618155e-05)),(to_sfixed_a(0.0001661159039940685)),(to_sfixed_a(2.971970388898626e-05)),(to_sfixed_a(-5.659612361341715e-05)),(to_sfixed_a(2.022445187321864e-06)),(to_sfixed_a(-9.181410860037431e-05)),(to_sfixed_a(-9.58633390837349e-05)),(to_sfixed_a(-8.422565588261932e-05)),(to_sfixed_a(-5.276214506011456e-05)),(to_sfixed_a(-0.0001303970639128238)),(to_sfixed_a(-8.979684935184196e-05)),(to_sfixed_a(-0.00013921478239353746)),(to_sfixed_a(1.06934330688091e-05)),(to_sfixed_a(3.481965541141108e-05)),(to_sfixed_a(-0.0002319643390364945)),(to_sfixed_a(-0.00010119872604263946)),(to_sfixed_a(2.2172571334522218e-05)),(to_sfixed_a(0.02114614099264145)),(to_sfixed_a(-4.5644526835530996e-05)),(to_sfixed_a(0.02402200736105442)),(to_sfixed_a(0.16816526651382446)),(to_sfixed_a(-0.08665766566991806)),(to_sfixed_a(-0.25864025950431824)),(to_sfixed_a(0.02629758231341839)),(to_sfixed_a(-0.06450081616640091)),(to_sfixed_a(0.020615756511688232)),(to_sfixed_a(0.006823258940130472)),(to_sfixed_a(-0.0848432406783104)),(to_sfixed_a(0.17516814172267914)),(to_sfixed_a(0.0736784115433693)),(to_sfixed_a(0.14964225888252258)),(to_sfixed_a(-0.000106113038782496)),(to_sfixed_a(-2.4376671717618592e-05)),(to_sfixed_a(-4.281686051399447e-05)),(to_sfixed_a(5.0071452278643847e-05)),(to_sfixed_a(-2.1838670363649726e-05)),(to_sfixed_a(-3.216586264898069e-05)),(to_sfixed_a(-0.00015375774819403887)),(to_sfixed_a(-0.00013564353866968304)),(to_sfixed_a(1.3814572412229609e-05)),(to_sfixed_a(0.00011411993182264268)),(to_sfixed_a(1.6340776710421778e-05)),(to_sfixed_a(8.893773338058963e-05)),(to_sfixed_a(-0.0016889759572222829)),(to_sfixed_a(0.0654546394944191)),(to_sfixed_a(-0.02192692644894123)),(to_sfixed_a(0.033707451075315475)),(to_sfixed_a(0.1863986998796463)),(to_sfixed_a(-0.002993113361299038)),(to_sfixed_a(-0.10520419478416443)),(to_sfixed_a(-0.17218108475208282)),(to_sfixed_a(-0.046741362661123276)),(to_sfixed_a(-0.012073450721800327)),(to_sfixed_a(0.1589042991399765)),(to_sfixed_a(0.2239343822002411)),(to_sfixed_a(0.05719628185033798)),(to_sfixed_a(0.1579812467098236)),(to_sfixed_a(0.010103944689035416)),(to_sfixed_a(0.14838461577892303)),(to_sfixed_a(-0.03652704134583473)),(to_sfixed_a(-0.0003182607179041952)),(to_sfixed_a(-0.0008208940853364766)),(to_sfixed_a(-7.990470476215705e-05)),(to_sfixed_a(-3.264242332079448e-05)),(to_sfixed_a(-0.0001721284061204642)),(to_sfixed_a(-0.00033749337308108807)),(to_sfixed_a(0.00016832123219501227)),(to_sfixed_a(-0.0002294139558216557)),(to_sfixed_a(-0.00024661634233780205)),(to_sfixed_a(0.0034647518768906593)),(to_sfixed_a(0.10509857535362244)),(to_sfixed_a(0.0028025407809764147)),(to_sfixed_a(0.11999578028917313)),(to_sfixed_a(0.17238539457321167)),(to_sfixed_a(-0.021349869668483734)),(to_sfixed_a(0.10480624437332153)),(to_sfixed_a(0.17489291727542877)),(to_sfixed_a(0.08625710010528564)),(to_sfixed_a(0.11338923126459122)),(to_sfixed_a(0.2180739790201187)),(to_sfixed_a(0.14487044513225555)),(to_sfixed_a(0.4224502444267273)),(to_sfixed_a(0.45157429575920105)),(to_sfixed_a(0.19076862931251526)),(to_sfixed_a(0.35035058856010437)),(to_sfixed_a(0.08842478692531586)),(to_sfixed_a(0.08948833495378494)),(to_sfixed_a(-0.0003708317526616156)),(to_sfixed_a(0.1288789063692093)),(to_sfixed_a(-0.0013273287331685424)),(to_sfixed_a(-0.000514068640768528)),(to_sfixed_a(3.7733330827904865e-05)),(to_sfixed_a(0.0001370700483676046)),(to_sfixed_a(-0.00010832154657691717)),(to_sfixed_a(1.5758620065753348e-05)),(to_sfixed_a(8.201331365853548e-05)),(to_sfixed_a(-0.00014213850954547524)),(to_sfixed_a(0.0002627129724714905)),(to_sfixed_a(0.1003129705786705)),(to_sfixed_a(0.11535269021987915)),(to_sfixed_a(0.14293670654296875)),(to_sfixed_a(0.007121487986296415)),(to_sfixed_a(0.010845943354070187)),(to_sfixed_a(0.32034367322921753)),(to_sfixed_a(0.006528346799314022)),(to_sfixed_a(0.1489398032426834)),(to_sfixed_a(0.14516106247901917)),(to_sfixed_a(0.2577086091041565)),(to_sfixed_a(0.4914943277835846)),(to_sfixed_a(0.29626011848449707)),(to_sfixed_a(0.22447875142097473)),(to_sfixed_a(0.5142059326171875)),(to_sfixed_a(0.0788789838552475)),(to_sfixed_a(0.19540253281593323)),(to_sfixed_a(-0.07102052867412567)),(to_sfixed_a(-0.03992354869842529)),(to_sfixed_a(-0.06601934134960175)),(to_sfixed_a(-0.0033595524728298187)),(to_sfixed_a(-0.0031834004912525415)),(to_sfixed_a(-0.0030669751577079296)),(to_sfixed_a(-0.0001597972441231832)),(to_sfixed_a(0.00017218438733834773)),(to_sfixed_a(0.00016570673324167728)),(to_sfixed_a(9.608145046513528e-05)),(to_sfixed_a(-3.7188165151746944e-05)),(to_sfixed_a(-0.000118273361294996)),(to_sfixed_a(-0.029058918356895447)),(to_sfixed_a(-0.009145091287791729)),(to_sfixed_a(-0.07527601718902588)),(to_sfixed_a(-0.02600311115384102)),(to_sfixed_a(0.13149048388004303)),(to_sfixed_a(0.14198456704616547)),(to_sfixed_a(0.23024128377437592)),(to_sfixed_a(0.17256282269954681)),(to_sfixed_a(0.10675671696662903)),(to_sfixed_a(0.38832518458366394)),(to_sfixed_a(0.4266780912876129)),(to_sfixed_a(0.2766473889350891)),(to_sfixed_a(0.22703184187412262)),(to_sfixed_a(0.24523857235908508)),(to_sfixed_a(-0.08421419560909271)),(to_sfixed_a(-0.07405778765678406)),(to_sfixed_a(-0.005119544919580221)),(to_sfixed_a(-0.028585387393832207)),(to_sfixed_a(-0.05789804086089134)),(to_sfixed_a(-0.038974277675151825)),(to_sfixed_a(-0.003198661608621478)),(to_sfixed_a(-4.0503902710042894e-05)),(to_sfixed_a(0.0001498102064942941)),(to_sfixed_a(0.0001855759328464046)),(to_sfixed_a(0.00018641218775883317)),(to_sfixed_a(-5.5714117479510605e-05)),(to_sfixed_a(-0.00019315046665724367)),(to_sfixed_a(-0.007463808637112379)),(to_sfixed_a(-0.003391367383301258)),(to_sfixed_a(-0.115467868745327)),(to_sfixed_a(-0.08477974683046341)),(to_sfixed_a(-0.08393774926662445)),(to_sfixed_a(-0.08453406393527985)),(to_sfixed_a(-0.029673902317881584)),(to_sfixed_a(-0.031182214617729187)),(to_sfixed_a(-0.13987015187740326)),(to_sfixed_a(-0.2954123616218567)),(to_sfixed_a(-0.03706725314259529)),(to_sfixed_a(0.0034358520060777664)),(to_sfixed_a(-0.20534415543079376)),(to_sfixed_a(-0.09118463099002838)),(to_sfixed_a(-0.15483015775680542)),(to_sfixed_a(-0.08117490261793137)),(to_sfixed_a(-0.15660087764263153)),(to_sfixed_a(-0.06851989775896072)),(to_sfixed_a(-0.0981731116771698)),(to_sfixed_a(-0.14856542646884918)),(to_sfixed_a(-0.06542719900608063)),(to_sfixed_a(-0.015579692088067532)),(to_sfixed_a(-0.0001056996698025614)),(to_sfixed_a(-2.7843228963320144e-05)),(to_sfixed_a(0.00023498764494434)),(to_sfixed_a(-0.0002314852026756853)),(to_sfixed_a(0.00018363659910392016)),(to_sfixed_a(-2.868436240532901e-05)),(to_sfixed_a(-0.002129334257915616)),(to_sfixed_a(-0.09811974316835403)),(to_sfixed_a(-0.0587749108672142)),(to_sfixed_a(-0.17953379452228546)),(to_sfixed_a(-0.03398746997117996)),(to_sfixed_a(-0.13790634274482727)),(to_sfixed_a(-0.5683777332305908)),(to_sfixed_a(-0.3287181854248047)),(to_sfixed_a(-0.6515045166015625)),(to_sfixed_a(-0.9022272825241089)),(to_sfixed_a(-0.9436296820640564)),(to_sfixed_a(-0.484030157327652)),(to_sfixed_a(-0.6768970489501953)),(to_sfixed_a(-1.0100986957550049)),(to_sfixed_a(-0.710202693939209)),(to_sfixed_a(-0.7417339086532593)),(to_sfixed_a(-0.7909494638442993)),(to_sfixed_a(-0.7858597040176392)),(to_sfixed_a(-0.518357515335083)),(to_sfixed_a(-0.2943544387817383)),(to_sfixed_a(-0.2251480370759964)),(to_sfixed_a(-5.665911885444075e-05)),(to_sfixed_a(-2.227456570835784e-05)),(to_sfixed_a(0.00012857838009949774)),(to_sfixed_a(3.745685899048112e-05)),(to_sfixed_a(-0.00011971034837188199)),(to_sfixed_a(-4.591565448208712e-05)),(to_sfixed_a(-2.6405632524983957e-05)),(to_sfixed_a(-0.013342826627194881)),(to_sfixed_a(-0.09594004601240158)),(to_sfixed_a(-0.782444179058075)),(to_sfixed_a(-0.2686581015586853)),(to_sfixed_a(-0.32508087158203125)),(to_sfixed_a(-0.7216488718986511)),(to_sfixed_a(-0.77168208360672)),(to_sfixed_a(-0.7613273859024048)),(to_sfixed_a(-0.4246412217617035)),(to_sfixed_a(-0.638572096824646)),(to_sfixed_a(-0.318050742149353)),(to_sfixed_a(-0.34981271624565125)),(to_sfixed_a(-0.4111669957637787)),(to_sfixed_a(-0.07751524448394775)),(to_sfixed_a(-0.4956150949001312)),(to_sfixed_a(-0.6225377917289734)),(to_sfixed_a(-0.5328202247619629)),(to_sfixed_a(-0.49892768263816833)),(to_sfixed_a(-0.3124425411224365)),(to_sfixed_a(-0.35900411009788513)),(to_sfixed_a(-0.10415168851613998)),(to_sfixed_a(-0.05043879896402359)),(to_sfixed_a(-0.0002391927846474573)),(to_sfixed_a(0.00028746394673362374)),(to_sfixed_a(-0.00018970943347085267)),(to_sfixed_a(0.0002867663570214063)),(to_sfixed_a(-0.0002551196375861764)),(to_sfixed_a(-0.049563515931367874)),(to_sfixed_a(-0.14355270564556122)),(to_sfixed_a(-0.42047908902168274)),(to_sfixed_a(-0.34074100852012634)),(to_sfixed_a(-0.5554535984992981)),(to_sfixed_a(-0.24246279895305634)),(to_sfixed_a(-0.29196038842201233)),(to_sfixed_a(-0.33829814195632935)),(to_sfixed_a(-0.580596387386322)),(to_sfixed_a(-0.20466671884059906)),(to_sfixed_a(-0.23416684567928314)),(to_sfixed_a(0.028764938935637474)),(to_sfixed_a(-0.02906052954494953)),(to_sfixed_a(0.2005048394203186)),(to_sfixed_a(0.09754634648561478)),(to_sfixed_a(-0.06399887055158615)),(to_sfixed_a(-0.24399444460868835)),(to_sfixed_a(-0.24026831984519958)),(to_sfixed_a(-0.06754227727651596)),(to_sfixed_a(-0.12862013280391693)),(to_sfixed_a(-0.49871498346328735)),(to_sfixed_a(-0.14620617032051086)),(to_sfixed_a(1.7695541828288697e-05)),(to_sfixed_a(-6.523174670292065e-05)),(to_sfixed_a(-0.0003867769264616072)),(to_sfixed_a(1.3213361853559036e-05)),(to_sfixed_a(-2.4923243472585455e-05)),(to_sfixed_a(0.00011093638750026003)),(to_sfixed_a(0.0002517513348720968)),(to_sfixed_a(-0.23746994137763977)),(to_sfixed_a(-0.29226401448249817)),(to_sfixed_a(-0.2925817668437958)),(to_sfixed_a(-0.45931288599967957)),(to_sfixed_a(-0.5614559650421143)),(to_sfixed_a(-0.4252581000328064)),(to_sfixed_a(-0.06375610083341599)),(to_sfixed_a(0.10814139991998672)),(to_sfixed_a(0.6220471858978271)),(to_sfixed_a(0.7932753562927246)),(to_sfixed_a(0.19725272059440613)),(to_sfixed_a(-0.037684764713048935)),(to_sfixed_a(0.14244644343852997)),(to_sfixed_a(0.0896170437335968)),(to_sfixed_a(0.16358582675457)),(to_sfixed_a(-0.23067326843738556)),(to_sfixed_a(-0.005646985024213791)),(to_sfixed_a(-0.13222409784793854)),(to_sfixed_a(-0.2836230397224426)),(to_sfixed_a(-0.07025931030511856)),(to_sfixed_a(0.07344397157430649)),(to_sfixed_a(-2.9904886105214246e-05)),(to_sfixed_a(-0.0004996644565835595)),(to_sfixed_a(-4.859466935158707e-05)),(to_sfixed_a(-4.058025297126733e-05)),(to_sfixed_a(4.230684498907067e-05)),(to_sfixed_a(-0.000245893927058205)),(to_sfixed_a(0.000253221282036975)),(to_sfixed_a(-0.031243519857525826)),(to_sfixed_a(-0.4181487262248993)),(to_sfixed_a(-0.29952216148376465)),(to_sfixed_a(-0.043659888207912445)),(to_sfixed_a(-0.08718056976795197)),(to_sfixed_a(0.12403585761785507)),(to_sfixed_a(0.17413853108882904)),(to_sfixed_a(0.5091053247451782)),(to_sfixed_a(0.42101001739501953)),(to_sfixed_a(0.30718284845352173)),(to_sfixed_a(0.3000050485134125)),(to_sfixed_a(0.13307547569274902)),(to_sfixed_a(-0.004164527170360088)),(to_sfixed_a(0.176764115691185)),(to_sfixed_a(0.062286633998155594)),(to_sfixed_a(0.026717809960246086)),(to_sfixed_a(0.022173231467604637)),(to_sfixed_a(-0.05837210640311241)),(to_sfixed_a(-0.0448949821293354)),(to_sfixed_a(0.014732018113136292)),(to_sfixed_a(0.02546222321689129)),(to_sfixed_a(-0.0009883098537102342)),(to_sfixed_a(-0.001555315568111837)),(to_sfixed_a(0.00027396256336942315)),(to_sfixed_a(-3.797506360569969e-05)),(to_sfixed_a(0.00022310960048343986)),(to_sfixed_a(0.00018271422595717013)),(to_sfixed_a(0.00011565574095584452)),(to_sfixed_a(-0.0003585861704777926)),(to_sfixed_a(0.19203904271125793)),(to_sfixed_a(0.30101561546325684)),(to_sfixed_a(0.4674023687839508)),(to_sfixed_a(0.23841792345046997)),(to_sfixed_a(0.5084800124168396)),(to_sfixed_a(0.4727596044540405)),(to_sfixed_a(0.4995502531528473)),(to_sfixed_a(0.32994309067726135)),(to_sfixed_a(0.49020543694496155)),(to_sfixed_a(0.25515350699424744)),(to_sfixed_a(0.024880578741431236)),(to_sfixed_a(0.06697993725538254)),(to_sfixed_a(0.11091138422489166)),(to_sfixed_a(0.06563428044319153)),(to_sfixed_a(0.08052463829517365)),(to_sfixed_a(0.06390601396560669)),(to_sfixed_a(0.034753892570734024)),(to_sfixed_a(0.01970629394054413)),(to_sfixed_a(0.048370376229286194)),(to_sfixed_a(0.013839267194271088)),(to_sfixed_a(0.0004406693042255938)),(to_sfixed_a(0.00021143299818504602)),(to_sfixed_a(-5.012475958210416e-05)),(to_sfixed_a(-4.383442956168437e-06)),(to_sfixed_a(5.9544650866882876e-05)),(to_sfixed_a(-0.00012288587458897382)),(to_sfixed_a(-4.3630152504192665e-05)),(to_sfixed_a(-0.021045133471488953)),(to_sfixed_a(0.22924868762493134)),(to_sfixed_a(0.17977607250213623)),(to_sfixed_a(0.18231043219566345)),(to_sfixed_a(0.3419777750968933)),(to_sfixed_a(0.565719723701477)),(to_sfixed_a(0.33857792615890503)),(to_sfixed_a(0.08159187436103821)),(to_sfixed_a(0.09793422371149063)),(to_sfixed_a(0.23703406751155853)),(to_sfixed_a(0.15972639620304108)),(to_sfixed_a(0.10312002152204514)),(to_sfixed_a(0.15630947053432465)),(to_sfixed_a(0.0731920376420021)),(to_sfixed_a(0.0817660540342331)),(to_sfixed_a(-0.030182911083102226)),(to_sfixed_a(0.05704127997159958)),(to_sfixed_a(-0.016063572838902473)),(to_sfixed_a(-0.04313642904162407)),(to_sfixed_a(0.11428766697645187)),(to_sfixed_a(0.07284098863601685)),(to_sfixed_a(0.0007802959298714995)),(to_sfixed_a(-0.00022591307060793042)),(to_sfixed_a(-0.00026374933077022433)),(to_sfixed_a(1.8799368262989447e-05)),(to_sfixed_a(0.00015422466094605625)),(to_sfixed_a(-0.00042977751581929624)),(to_sfixed_a(-0.003562280675396323)),(to_sfixed_a(0.21484000980854034)),(to_sfixed_a(0.32530736923217773)),(to_sfixed_a(0.5706583857536316)),(to_sfixed_a(0.3986286520957947)),(to_sfixed_a(0.34113678336143494)),(to_sfixed_a(0.1153755784034729)),(to_sfixed_a(0.20200958847999573)),(to_sfixed_a(0.08971408009529114)),(to_sfixed_a(0.24849221110343933)),(to_sfixed_a(0.05793456360697746)),(to_sfixed_a(0.10672234743833542)),(to_sfixed_a(0.20609864592552185)),(to_sfixed_a(0.19386522471904755)),(to_sfixed_a(0.054870568215847015)),(to_sfixed_a(0.16223427653312683)),(to_sfixed_a(0.142709881067276)),(to_sfixed_a(0.11564107239246368)),(to_sfixed_a(0.2073180228471756)),(to_sfixed_a(-0.0021915524266660213)),(to_sfixed_a(-0.03498881310224533)),(to_sfixed_a(0.06406666338443756)),(to_sfixed_a(0.0026604016311466694)),(to_sfixed_a(6.796333309466718e-07)),(to_sfixed_a(-0.00026480239466764033)),(to_sfixed_a(-0.00016186067659873515)),(to_sfixed_a(6.948721420485526e-05)),(to_sfixed_a(-0.0024499697610735893)),(to_sfixed_a(-0.003228249726817012)),(to_sfixed_a(0.013325715437531471)),(to_sfixed_a(0.35161247849464417)),(to_sfixed_a(0.21444405615329742)),(to_sfixed_a(0.20929615199565887)),(to_sfixed_a(0.197675421833992)),(to_sfixed_a(0.3070380985736847)),(to_sfixed_a(0.30343446135520935)),(to_sfixed_a(0.32975614070892334)),(to_sfixed_a(0.2623361051082611)),(to_sfixed_a(0.0810299962759018)),(to_sfixed_a(0.10165682435035706)),(to_sfixed_a(0.009367025457322598)),(to_sfixed_a(0.18292075395584106)),(to_sfixed_a(0.13650791347026825)),(to_sfixed_a(-0.005404503084719181)),(to_sfixed_a(-0.19811700284481049)),(to_sfixed_a(0.0998600646853447)),(to_sfixed_a(0.05466221645474434)),(to_sfixed_a(0.04994521662592888)),(to_sfixed_a(-0.0011128144105896354)),(to_sfixed_a(0.00020822258375119418)),(to_sfixed_a(-9.250146831618622e-06)),(to_sfixed_a(0.00024524066247977316)),(to_sfixed_a(8.010287274373695e-05)),(to_sfixed_a(-9.121609036810696e-05)),(to_sfixed_a(-9.717144712340087e-05)),(to_sfixed_a(-0.0001651610800763592)),(to_sfixed_a(0.012622225098311901)),(to_sfixed_a(0.08427092432975769)),(to_sfixed_a(0.20324741303920746)),(to_sfixed_a(0.06614221632480621)),(to_sfixed_a(0.15580403804779053)),(to_sfixed_a(0.20720556378364563)),(to_sfixed_a(0.2660750448703766)),(to_sfixed_a(0.2967474162578583)),(to_sfixed_a(0.2991604506969452)),(to_sfixed_a(0.002396263414993882)),(to_sfixed_a(-0.1256694197654724)),(to_sfixed_a(0.0768035277724266)),(to_sfixed_a(0.15589693188667297)),(to_sfixed_a(0.16975171864032745)),(to_sfixed_a(-0.12307678163051605)),(to_sfixed_a(-0.023062001913785934)),(to_sfixed_a(0.12004802376031876)),(to_sfixed_a(0.015139041468501091)),(to_sfixed_a(-0.040748998522758484)),(to_sfixed_a(0.12604936957359314)),(to_sfixed_a(0.02590457908809185)),(to_sfixed_a(-0.0052773961797356606)),(to_sfixed_a(-0.00010595551430014893)),(to_sfixed_a(3.227484558010474e-05)),(to_sfixed_a(-9.889063221635297e-05)),(to_sfixed_a(3.945999560528435e-05)),(to_sfixed_a(-0.00015561094915028661)),(to_sfixed_a(-6.123002822278067e-05)),(to_sfixed_a(-0.04405658692121506)),(to_sfixed_a(0.0027754385955631733)),(to_sfixed_a(-0.06433537602424622)),(to_sfixed_a(0.04523308947682381)),(to_sfixed_a(-0.03835047781467438)),(to_sfixed_a(-0.09836599975824356)),(to_sfixed_a(0.09894601255655289)),(to_sfixed_a(0.33386310935020447)),(to_sfixed_a(0.04945991560816765)),(to_sfixed_a(0.002254074439406395)),(to_sfixed_a(0.09110281616449356)),(to_sfixed_a(0.17342475056648254)),(to_sfixed_a(0.2611145079135895)),(to_sfixed_a(0.0402083657681942)),(to_sfixed_a(0.004858565982431173)),(to_sfixed_a(0.0005954885855317116)),(to_sfixed_a(0.010732977651059628)),(to_sfixed_a(-0.10712483525276184)),(to_sfixed_a(0.07361508905887604)),(to_sfixed_a(0.04249975085258484)),(to_sfixed_a(0.06143728271126747)),(to_sfixed_a(1.8876873582485132e-05)),(to_sfixed_a(3.632170773926191e-05)),(to_sfixed_a(-7.838611054467037e-05)),(to_sfixed_a(-6.900208973092958e-05)),(to_sfixed_a(3.857529736706056e-05)),(to_sfixed_a(-0.00021142764308024198)),(to_sfixed_a(-0.00015139438619371504)),(to_sfixed_a(-0.00017142490833066404)),(to_sfixed_a(-0.0031051677651703358)),(to_sfixed_a(0.1865897923707962)),(to_sfixed_a(-0.12505526840686798)),(to_sfixed_a(0.061613090336322784)),(to_sfixed_a(0.02699410356581211)),(to_sfixed_a(0.01114222127944231)),(to_sfixed_a(0.19069449603557587)),(to_sfixed_a(-0.0689699798822403)),(to_sfixed_a(-0.030730310827493668)),(to_sfixed_a(-0.04347739368677139)),(to_sfixed_a(0.05641338601708412)),(to_sfixed_a(0.20540477335453033)),(to_sfixed_a(0.026152290403842926)),(to_sfixed_a(-0.019066983833909035)),(to_sfixed_a(0.014273206703364849)),(to_sfixed_a(-0.004342304076999426)),(to_sfixed_a(-0.0246873926371336)),(to_sfixed_a(0.24987201392650604)),(to_sfixed_a(-0.013778936117887497)),(to_sfixed_a(0.1460294872522354)),(to_sfixed_a(0.18413810431957245)),(to_sfixed_a(-0.00011050296598114073)),(to_sfixed_a(-9.554703865433112e-05)),(to_sfixed_a(9.438544111617375e-06)),(to_sfixed_a(-5.819587386213243e-05)),(to_sfixed_a(4.4785108912037686e-05)),(to_sfixed_a(8.279633766505867e-05)),(to_sfixed_a(5.998650522087701e-05)),(to_sfixed_a(-0.04678117111325264)),(to_sfixed_a(0.0019276695093140006)),(to_sfixed_a(0.0030909923370927572)),(to_sfixed_a(0.07719504833221436)),(to_sfixed_a(0.19746999442577362)),(to_sfixed_a(-0.02355898544192314)),(to_sfixed_a(-0.08759380877017975)),(to_sfixed_a(-0.1362997442483902)),(to_sfixed_a(0.14686085283756256)),(to_sfixed_a(0.11020242422819138)),(to_sfixed_a(-0.02444957196712494)),(to_sfixed_a(-0.1511434018611908)),(to_sfixed_a(0.05987479165196419)),(to_sfixed_a(0.1112048402428627)),(to_sfixed_a(-0.09439752995967865)),(to_sfixed_a(-0.02029591053724289)),(to_sfixed_a(-0.02927732653915882)),(to_sfixed_a(0.006718922406435013)),(to_sfixed_a(0.10028855502605438)),(to_sfixed_a(-0.00042835515341721475)),(to_sfixed_a(0.0028471776749938726)),(to_sfixed_a(-0.00020207598572596908)),(to_sfixed_a(-0.00010222529817838222)),(to_sfixed_a(6.200568896019831e-05)),(to_sfixed_a(-0.00017517991364002228)),(to_sfixed_a(-0.00022782571613788605)),(to_sfixed_a(-0.00037242809776216745)),(to_sfixed_a(0.00018629674741532654)),(to_sfixed_a(-0.00029048658325336874)),(to_sfixed_a(0.002324090339243412)),(to_sfixed_a(-0.03644729405641556)),(to_sfixed_a(0.03434479981660843)),(to_sfixed_a(-0.04252522438764572)),(to_sfixed_a(-0.08005873113870621)),(to_sfixed_a(-0.061878275126218796)),(to_sfixed_a(-0.11805269122123718)),(to_sfixed_a(-0.14424574375152588)),(to_sfixed_a(-0.12381958216428757)),(to_sfixed_a(-0.09210586547851562)),(to_sfixed_a(-0.12738199532032013)),(to_sfixed_a(0.01388560701161623)),(to_sfixed_a(-0.08494154363870621)),(to_sfixed_a(-0.15646892786026)),(to_sfixed_a(0.05834038928151131)),(to_sfixed_a(0.018519172444939613)),(to_sfixed_a(-0.0035039959475398064)),(to_sfixed_a(-0.01182587631046772)),(to_sfixed_a(-0.0044397879391908646)),(to_sfixed_a(3.0345534469233826e-05)),(to_sfixed_a(-4.372213879832998e-05)),(to_sfixed_a(-4.8951336793834344e-05)),(to_sfixed_a(0.00024495660909451544)),(to_sfixed_a(3.2222278605331667e-06)),(to_sfixed_a(0.0001817812299123034)),(to_sfixed_a(-1.6299685739795677e-05)),(to_sfixed_a(4.0056591387838125e-05)),(to_sfixed_a(-0.0002171992091462016)),(to_sfixed_a(0.03467772901058197)),(to_sfixed_a(-0.013830739073455334)),(to_sfixed_a(-0.09754141420125961)),(to_sfixed_a(-0.04208085685968399)),(to_sfixed_a(-0.07518705725669861)),(to_sfixed_a(-0.035423994064331055)),(to_sfixed_a(-0.1488436460494995)),(to_sfixed_a(-0.05921699479222298)),(to_sfixed_a(-0.012290765531361103)),(to_sfixed_a(-0.10907319188117981)),(to_sfixed_a(-0.08805801719427109)),(to_sfixed_a(-0.15510228276252747)),(to_sfixed_a(-0.273781418800354)),(to_sfixed_a(0.010954326950013638)),(to_sfixed_a(0.08152762055397034)),(to_sfixed_a(-0.03872513398528099)),(to_sfixed_a(0.04512681066989899)),(to_sfixed_a(-0.00913726631551981)),(to_sfixed_a(0.03631272166967392)),(to_sfixed_a(1.5185359188762959e-05)),(to_sfixed_a(-0.0002777451591100544)),(to_sfixed_a(-4.853971040574834e-05)),(to_sfixed_a(-7.838752208044752e-05)),(to_sfixed_a(-0.0001320158044109121)),(to_sfixed_a(-9.526123176328838e-05)),(to_sfixed_a(6.155212759040296e-05)),(to_sfixed_a(0.00039569599903188646)),(to_sfixed_a(-0.018475480377674103)),(to_sfixed_a(-0.005167090799659491)),(to_sfixed_a(-0.0774625837802887)),(to_sfixed_a(-0.15662360191345215)),(to_sfixed_a(-0.02474217861890793)),(to_sfixed_a(-0.058488018810749054)),(to_sfixed_a(-0.1347431093454361)),(to_sfixed_a(-0.11073268949985504)),(to_sfixed_a(-0.025152167305350304)),(to_sfixed_a(-0.12351754307746887)),(to_sfixed_a(0.023969030007719994)),(to_sfixed_a(-0.0710577443242073)),(to_sfixed_a(-0.12160123139619827)),(to_sfixed_a(-0.09309269487857819)),(to_sfixed_a(-0.049733810126781464)),(to_sfixed_a(0.002540945541113615)),(to_sfixed_a(0.007553454488515854)),(to_sfixed_a(0.04062014818191528)),(to_sfixed_a(0.020644180476665497)),(to_sfixed_a(-0.004541645757853985)),(to_sfixed_a(-7.145565905375406e-05)),(to_sfixed_a(-0.00013263133587315679)),(to_sfixed_a(4.879988409811631e-05)),(to_sfixed_a(7.007873500697315e-05)),(to_sfixed_a(-0.0001488867128500715)),(to_sfixed_a(4.6477467549266294e-05)),(to_sfixed_a(-0.00011222218017792329)),(to_sfixed_a(-1.5848099792492576e-05)),(to_sfixed_a(7.63185198593419e-06)),(to_sfixed_a(0.03373854234814644)),(to_sfixed_a(-0.04638248309493065)),(to_sfixed_a(-0.034742411226034164)),(to_sfixed_a(-0.07713870704174042)),(to_sfixed_a(-0.11945214122533798)),(to_sfixed_a(-0.13038285076618195)),(to_sfixed_a(-0.14050039649009705)),(to_sfixed_a(-0.14789558947086334)),(to_sfixed_a(-0.07467211037874222)),(to_sfixed_a(-0.10861971974372864)),(to_sfixed_a(-0.09988560527563095)),(to_sfixed_a(0.053839441388845444)),(to_sfixed_a(0.06811560690402985)),(to_sfixed_a(-0.004029766656458378)),(to_sfixed_a(-0.15045472979545593)),(to_sfixed_a(-0.13750296831130981)),(to_sfixed_a(-0.0005178157589398324)),(to_sfixed_a(-0.0020934317726641893)),(to_sfixed_a(-0.0019238459644839168)),(to_sfixed_a(5.3962907259119675e-05)),(to_sfixed_a(1.8472586816642433e-05)),(to_sfixed_a(-0.0002179389848606661)),(to_sfixed_a(-4.323423581809038e-06)),(to_sfixed_a(-0.0001522263919468969)),(to_sfixed_a(-1.9978326236014254e-05)),(to_sfixed_a(-0.0001606357836863026)),(to_sfixed_a(-3.901902891811915e-05)),(to_sfixed_a(-0.00025549117708578706)),(to_sfixed_a(-0.0006938977167010307)),(to_sfixed_a(-0.0005843286053277552)),(to_sfixed_a(0.0001195922086481005)),(to_sfixed_a(0.00027495500398799777)),(to_sfixed_a(-0.0003078771405853331)),(to_sfixed_a(-0.1571662276983261)),(to_sfixed_a(0.006679549813270569)),(to_sfixed_a(0.0024396213702857494)),(to_sfixed_a(-0.1254836618900299)),(to_sfixed_a(-0.03840235620737076)),(to_sfixed_a(-0.0038562119007110596)),(to_sfixed_a(0.007902667857706547)),(to_sfixed_a(-0.12734071910381317)),(to_sfixed_a(-0.17734937369823456)),(to_sfixed_a(-0.016485359519720078)),(to_sfixed_a(-0.008035533130168915)),(to_sfixed_a(1.0624953574733809e-05)),(to_sfixed_a(-9.468897769693285e-05)),(to_sfixed_a(-0.00013975132605992258)),(to_sfixed_a(-0.00012640542990993708)),(to_sfixed_a(4.216039087623358e-05)),(to_sfixed_a(0.0002908388269133866)),(to_sfixed_a(0.00013572048919741064)),(to_sfixed_a(0.00013676310481969267)),(to_sfixed_a(3.530913818394765e-05)),(to_sfixed_a(-0.00020636580302380025)),(to_sfixed_a(-0.000193793821381405)),(to_sfixed_a(-7.990095582499634e-06)),(to_sfixed_a(-0.0001664534502197057)),(to_sfixed_a(-0.00032449018908664584)),(to_sfixed_a(-0.00020002617384307086)),(to_sfixed_a(-0.00011235193233005702)),(to_sfixed_a(-3.889026993419975e-05)),(to_sfixed_a(-8.017985237529501e-06)),(to_sfixed_a(-0.00011497564264573157)),(to_sfixed_a(-0.00021515246771741658)),(to_sfixed_a(5.857953874510713e-05)),(to_sfixed_a(0.00014813833695370704)),(to_sfixed_a(-0.0001288533821934834)),(to_sfixed_a(-3.062051837332547e-05)),(to_sfixed_a(-0.00018591841217130423)),(to_sfixed_a(-8.599150169175118e-05)),(to_sfixed_a(-0.00043560811900533736)),(to_sfixed_a(0.000166442827321589)),(to_sfixed_a(0.0001672003127168864)),(to_sfixed_a(-0.00020812010916415602)),(to_sfixed_a(0.00018555000133346766)),(to_sfixed_a(0.00015918264398351312)),(to_sfixed_a(2.0333864085841924e-05)),(to_sfixed_a(-4.6335237129824236e-05)),(to_sfixed_a(5.8591878769220784e-05)));

    constant weight_n0_1 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(2.8026910513290204e-05)),(to_sfixed_a(0.00011689306847983971)),(to_sfixed_a(-7.835796714061871e-05)),(to_sfixed_a(0.00021529263176489621)),(to_sfixed_a(4.77654866699595e-05)),(to_sfixed_a(0.0003796041419263929)),(to_sfixed_a(6.72201786073856e-05)),(to_sfixed_a(-0.000275352067546919)),(to_sfixed_a(-0.0002417888172203675)),(to_sfixed_a(-0.00018258810450788587)),(to_sfixed_a(-0.00023059685190673918)),(to_sfixed_a(0.00017676022252999246)),(to_sfixed_a(8.310430712299421e-05)),(to_sfixed_a(-0.00015810086915735155)),(to_sfixed_a(-5.238113953964785e-05)),(to_sfixed_a(0.00014620364527218044)),(to_sfixed_a(0.00027088235947303474)),(to_sfixed_a(-2.2012409317540005e-06)),(to_sfixed_a(0.0002208653895650059)),(to_sfixed_a(0.0003293217741884291)),(to_sfixed_a(-0.0002059341495623812)),(to_sfixed_a(-3.963076596846804e-05)),(to_sfixed_a(-0.00019241744303144515)),(to_sfixed_a(-0.00012702356616500765)),(to_sfixed_a(0.00026569387409836054)),(to_sfixed_a(0.00024291501904372126)),(to_sfixed_a(-1.8699201973504387e-05)),(to_sfixed_a(0.00012232021254021674)),(to_sfixed_a(-0.0003026314952876419)),(to_sfixed_a(-0.0003763637214433402)),(to_sfixed_a(2.6509660528972745e-05)),(to_sfixed_a(-0.00010840978211490437)),(to_sfixed_a(-3.290191443738877e-06)),(to_sfixed_a(1.7431848391424865e-05)),(to_sfixed_a(6.404536543413997e-05)),(to_sfixed_a(0.00022294273367151618)),(to_sfixed_a(7.91292950452771e-06)),(to_sfixed_a(-2.44591137743555e-05)),(to_sfixed_a(0.00030697736656293273)),(to_sfixed_a(5.282364145386964e-05)),(to_sfixed_a(0.00017606947221793234)),(to_sfixed_a(9.004372986964881e-05)),(to_sfixed_a(-5.414868428488262e-05)),(to_sfixed_a(-6.061938256607391e-05)),(to_sfixed_a(-6.346141162794083e-05)),(to_sfixed_a(7.420904148602858e-05)),(to_sfixed_a(0.00010678958642529324)),(to_sfixed_a(5.1718365284614265e-05)),(to_sfixed_a(0.00015072687529027462)),(to_sfixed_a(1.483655159972841e-05)),(to_sfixed_a(8.733806316740811e-05)),(to_sfixed_a(-0.00028400865267030895)),(to_sfixed_a(-7.176964572863653e-06)),(to_sfixed_a(-0.00013840632163919508)),(to_sfixed_a(0.00010397801815997809)),(to_sfixed_a(-0.00012136343866586685)),(to_sfixed_a(0.0001699454733170569)),(to_sfixed_a(-0.00010661652777343988)),(to_sfixed_a(0.00038112830952741206)),(to_sfixed_a(2.898646698668017e-06)),(to_sfixed_a(-0.00014126382302492857)),(to_sfixed_a(0.00026109747705049813)),(to_sfixed_a(7.597352669108659e-05)),(to_sfixed_a(-6.362674321280792e-05)),(to_sfixed_a(-0.00011533348151715472)),(to_sfixed_a(-0.00014466764696408063)),(to_sfixed_a(0.0001244186278199777)),(to_sfixed_a(3.83363185392227e-05)),(to_sfixed_a(8.481028635287657e-05)),(to_sfixed_a(-0.0007431068224832416)),(to_sfixed_a(0.00017965921142604202)),(to_sfixed_a(-0.0002703071222640574)),(to_sfixed_a(6.287178985076025e-05)),(to_sfixed_a(6.244339601835236e-05)),(to_sfixed_a(7.257977267727256e-05)),(to_sfixed_a(-0.0001331331004621461)),(to_sfixed_a(0.0002701709163375199)),(to_sfixed_a(0.00011640129378065467)),(to_sfixed_a(-0.0002592082601040602)),(to_sfixed_a(-0.0004877984756603837)),(to_sfixed_a(-0.0001958230132004246)),(to_sfixed_a(5.927211532252841e-05)),(to_sfixed_a(-2.4464647140121087e-05)),(to_sfixed_a(6.535603461088613e-05)),(to_sfixed_a(-8.551415521651506e-05)),(to_sfixed_a(0.00015932254609651864)),(to_sfixed_a(-0.0002669181558303535)),(to_sfixed_a(0.0001588456507306546)),(to_sfixed_a(6.0430877056205645e-05)),(to_sfixed_a(3.639415808720514e-05)),(to_sfixed_a(3.609938721638173e-05)),(to_sfixed_a(6.549576937686652e-05)),(to_sfixed_a(-0.06361852586269379)),(to_sfixed_a(6.860539724584669e-05)),(to_sfixed_a(-0.07207644730806351)),(to_sfixed_a(0.1262901872396469)),(to_sfixed_a(-0.16117580235004425)),(to_sfixed_a(-0.12212809920310974)),(to_sfixed_a(-0.10771885514259338)),(to_sfixed_a(-0.058410048484802246)),(to_sfixed_a(0.010721931234002113)),(to_sfixed_a(0.023235013708472252)),(to_sfixed_a(-0.03738410398364067)),(to_sfixed_a(0.08526536822319031)),(to_sfixed_a(0.04780136048793793)),(to_sfixed_a(0.09702905267477036)),(to_sfixed_a(3.028110995728639e-06)),(to_sfixed_a(0.00017387466505169868)),(to_sfixed_a(-0.00013304405729286373)),(to_sfixed_a(-6.366286834236234e-05)),(to_sfixed_a(-0.00011968302715104073)),(to_sfixed_a(-0.00018209063273388892)),(to_sfixed_a(-3.860335345962085e-05)),(to_sfixed_a(1.130512828240171e-05)),(to_sfixed_a(0.00010474494774825871)),(to_sfixed_a(7.40577161195688e-05)),(to_sfixed_a(-3.0132503525237553e-05)),(to_sfixed_a(-5.215866258367896e-05)),(to_sfixed_a(-0.0005056363297626376)),(to_sfixed_a(0.050467535853385925)),(to_sfixed_a(0.06248586252331734)),(to_sfixed_a(-0.09455543756484985)),(to_sfixed_a(0.0298556350171566)),(to_sfixed_a(-0.07709259539842606)),(to_sfixed_a(-0.07499290257692337)),(to_sfixed_a(0.08807220309972763)),(to_sfixed_a(0.09479616582393646)),(to_sfixed_a(0.22756800055503845)),(to_sfixed_a(0.33931466937065125)),(to_sfixed_a(0.26518285274505615)),(to_sfixed_a(0.033111877739429474)),(to_sfixed_a(-0.005566807463765144)),(to_sfixed_a(-0.0006781172705814242)),(to_sfixed_a(0.12981344759464264)),(to_sfixed_a(0.09094754606485367)),(to_sfixed_a(-0.00026487221475690603)),(to_sfixed_a(0.0006302041583694518)),(to_sfixed_a(0.00022188492584973574)),(to_sfixed_a(-0.0001758369617164135)),(to_sfixed_a(-8.049087773542851e-05)),(to_sfixed_a(0.00023827256518416107)),(to_sfixed_a(0.00029221875593066216)),(to_sfixed_a(-7.508511316700606e-06)),(to_sfixed_a(2.4670842321938835e-05)),(to_sfixed_a(0.002899313811212778)),(to_sfixed_a(0.0820298045873642)),(to_sfixed_a(0.006982951425015926)),(to_sfixed_a(0.06441520154476166)),(to_sfixed_a(0.12201577425003052)),(to_sfixed_a(-0.006737720686942339)),(to_sfixed_a(0.08030728250741959)),(to_sfixed_a(0.236094668507576)),(to_sfixed_a(0.12738759815692902)),(to_sfixed_a(0.24604734778404236)),(to_sfixed_a(0.10271985083818436)),(to_sfixed_a(0.007558323442935944)),(to_sfixed_a(0.22524794936180115)),(to_sfixed_a(0.3071468770503998)),(to_sfixed_a(0.14144404232501984)),(to_sfixed_a(-0.029340147972106934)),(to_sfixed_a(0.050615303218364716)),(to_sfixed_a(0.08339126408100128)),(to_sfixed_a(0.003617824288085103)),(to_sfixed_a(0.11334837973117828)),(to_sfixed_a(-0.0009544803760945797)),(to_sfixed_a(-0.0001796358556021005)),(to_sfixed_a(-0.00022776360856369138)),(to_sfixed_a(-9.271353337680921e-05)),(to_sfixed_a(0.0001230130874319002)),(to_sfixed_a(-0.00032833864679560065)),(to_sfixed_a(1.7773616491467692e-05)),(to_sfixed_a(-0.00015893130330368876)),(to_sfixed_a(0.0008286083466373384)),(to_sfixed_a(0.07678481191396713)),(to_sfixed_a(0.051009878516197205)),(to_sfixed_a(0.03470972180366516)),(to_sfixed_a(0.0939006581902504)),(to_sfixed_a(0.24765826761722565)),(to_sfixed_a(0.4838480055332184)),(to_sfixed_a(0.21103209257125854)),(to_sfixed_a(0.36813223361968994)),(to_sfixed_a(0.2848922312259674)),(to_sfixed_a(0.3500087559223175)),(to_sfixed_a(0.4594041407108307)),(to_sfixed_a(0.1276887059211731)),(to_sfixed_a(0.277099609375)),(to_sfixed_a(0.5841360092163086)),(to_sfixed_a(0.25151699781417847)),(to_sfixed_a(0.28502339124679565)),(to_sfixed_a(0.12051480263471603)),(to_sfixed_a(0.02217959240078926)),(to_sfixed_a(-0.02245098352432251)),(to_sfixed_a(-0.004817829467356205)),(to_sfixed_a(-0.005100968759506941)),(to_sfixed_a(-0.002650028793141246)),(to_sfixed_a(-5.076059824205004e-05)),(to_sfixed_a(3.4053256968036294e-05)),(to_sfixed_a(-0.00012044158938806504)),(to_sfixed_a(-8.322882786160335e-05)),(to_sfixed_a(1.5091666682565119e-05)),(to_sfixed_a(-9.718937690195162e-06)),(to_sfixed_a(0.02355870045721531)),(to_sfixed_a(0.11973534524440765)),(to_sfixed_a(-0.02517259120941162)),(to_sfixed_a(0.1719667911529541)),(to_sfixed_a(0.10250457376241684)),(to_sfixed_a(0.31730011105537415)),(to_sfixed_a(0.0035293535329401493)),(to_sfixed_a(0.08314687013626099)),(to_sfixed_a(0.16380125284194946)),(to_sfixed_a(0.29394984245300293)),(to_sfixed_a(0.20514315366744995)),(to_sfixed_a(0.3405230641365051)),(to_sfixed_a(0.1345091164112091)),(to_sfixed_a(0.3622535169124603)),(to_sfixed_a(0.43287909030914307)),(to_sfixed_a(0.2713755667209625)),(to_sfixed_a(0.16872841119766235)),(to_sfixed_a(-0.01913141831755638)),(to_sfixed_a(0.17926737666130066)),(to_sfixed_a(-0.013554561883211136)),(to_sfixed_a(0.002055142307654023)),(to_sfixed_a(2.172904714825563e-05)),(to_sfixed_a(1.7133430446847342e-05)),(to_sfixed_a(5.761460852227174e-05)),(to_sfixed_a(0.0003459715226199478)),(to_sfixed_a(-9.039759606821463e-05)),(to_sfixed_a(-1.650562626309693e-05)),(to_sfixed_a(0.0610506534576416)),(to_sfixed_a(-0.01082637533545494)),(to_sfixed_a(0.016028642654418945)),(to_sfixed_a(0.13835135102272034)),(to_sfixed_a(0.04966849088668823)),(to_sfixed_a(-0.004673860035836697)),(to_sfixed_a(0.20344729721546173)),(to_sfixed_a(-0.0316188707947731)),(to_sfixed_a(0.0714062750339508)),(to_sfixed_a(-0.15679405629634857)),(to_sfixed_a(-0.12952712178230286)),(to_sfixed_a(0.020530184730887413)),(to_sfixed_a(-0.16688968241214752)),(to_sfixed_a(0.14329560101032257)),(to_sfixed_a(0.2508034408092499)),(to_sfixed_a(0.12980155646800995)),(to_sfixed_a(0.21180042624473572)),(to_sfixed_a(0.03246913105249405)),(to_sfixed_a(0.18720780313014984)),(to_sfixed_a(0.028604701161384583)),(to_sfixed_a(0.020743489265441895)),(to_sfixed_a(0.0037516586016863585)),(to_sfixed_a(0.0001995648053707555)),(to_sfixed_a(-8.696656550455373e-06)),(to_sfixed_a(3.3488009648863226e-05)),(to_sfixed_a(-8.754314330872148e-05)),(to_sfixed_a(-0.00016501828213222325)),(to_sfixed_a(-0.00012979144230484962)),(to_sfixed_a(-0.003933057188987732)),(to_sfixed_a(0.13091525435447693)),(to_sfixed_a(0.04764376953244209)),(to_sfixed_a(0.14933346211910248)),(to_sfixed_a(0.06481464207172394)),(to_sfixed_a(-0.05363186076283455)),(to_sfixed_a(-0.2108357846736908)),(to_sfixed_a(-0.06604219973087311)),(to_sfixed_a(-0.0013060095952823758)),(to_sfixed_a(-0.4513379633426666)),(to_sfixed_a(-0.4719831645488739)),(to_sfixed_a(-0.39383646845817566)),(to_sfixed_a(-0.539157509803772)),(to_sfixed_a(-0.810099720954895)),(to_sfixed_a(-0.4865310788154602)),(to_sfixed_a(-0.6402690410614014)),(to_sfixed_a(-0.4186071753501892)),(to_sfixed_a(-0.4383019208908081)),(to_sfixed_a(-0.37694448232650757)),(to_sfixed_a(-0.133114755153656)),(to_sfixed_a(-0.05440330505371094)),(to_sfixed_a(0.00010312928498024121)),(to_sfixed_a(-0.00019120216893497854)),(to_sfixed_a(0.0001228485634783283)),(to_sfixed_a(-2.1751056920038536e-05)),(to_sfixed_a(-0.00021029134222771972)),(to_sfixed_a(-4.687382897827774e-06)),(to_sfixed_a(6.770511390641332e-05)),(to_sfixed_a(-0.007502342574298382)),(to_sfixed_a(-0.007767036557197571)),(to_sfixed_a(-0.09277499467134476)),(to_sfixed_a(-0.15903374552726746)),(to_sfixed_a(-0.08137543499469757)),(to_sfixed_a(-0.24733705818653107)),(to_sfixed_a(-0.10377294570207596)),(to_sfixed_a(0.1265431046485901)),(to_sfixed_a(-0.183157280087471)),(to_sfixed_a(-0.05111822485923767)),(to_sfixed_a(-0.4364403486251831)),(to_sfixed_a(-0.47783246636390686)),(to_sfixed_a(-0.31564706563949585)),(to_sfixed_a(-0.03093445859849453)),(to_sfixed_a(-0.43343719840049744)),(to_sfixed_a(-0.5568534135818481)),(to_sfixed_a(-0.4158719778060913)),(to_sfixed_a(-0.20733849704265594)),(to_sfixed_a(-0.20126840472221375)),(to_sfixed_a(-0.012143697589635849)),(to_sfixed_a(-0.06948959082365036)),(to_sfixed_a(-0.03300303593277931)),(to_sfixed_a(9.093039989238605e-05)),(to_sfixed_a(2.0271396351745352e-05)),(to_sfixed_a(9.451396181248128e-05)),(to_sfixed_a(9.880889410851523e-05)),(to_sfixed_a(0.00017955248767975718)),(to_sfixed_a(-0.032276272773742676)),(to_sfixed_a(0.07833371311426163)),(to_sfixed_a(-0.09665881097316742)),(to_sfixed_a(-0.1420576572418213)),(to_sfixed_a(-0.06367572396993637)),(to_sfixed_a(0.08873985707759857)),(to_sfixed_a(0.16106373071670532)),(to_sfixed_a(0.18178507685661316)),(to_sfixed_a(0.43923690915107727)),(to_sfixed_a(0.42062991857528687)),(to_sfixed_a(-0.2073160707950592)),(to_sfixed_a(-0.41551119089126587)),(to_sfixed_a(-0.2596690356731415)),(to_sfixed_a(0.028678294271230698)),(to_sfixed_a(-0.007232842966914177)),(to_sfixed_a(-0.16606292128562927)),(to_sfixed_a(-0.22801466286182404)),(to_sfixed_a(-0.21410474181175232)),(to_sfixed_a(0.056685179471969604)),(to_sfixed_a(-0.05704149603843689)),(to_sfixed_a(-0.16324658691883087)),(to_sfixed_a(-0.11819890141487122)),(to_sfixed_a(-2.29928336921148e-05)),(to_sfixed_a(-0.00011730886035365984)),(to_sfixed_a(-9.76080700638704e-05)),(to_sfixed_a(0.0001902808144222945)),(to_sfixed_a(0.0002379633515374735)),(to_sfixed_a(-2.9682791137020104e-05)),(to_sfixed_a(-0.0002937235403805971)),(to_sfixed_a(0.11399678140878677)),(to_sfixed_a(0.15977010130882263)),(to_sfixed_a(0.018440881744027138)),(to_sfixed_a(0.29437512159347534)),(to_sfixed_a(0.2706339955329895)),(to_sfixed_a(0.3757200241088867)),(to_sfixed_a(0.42554202675819397)),(to_sfixed_a(0.32034972310066223)),(to_sfixed_a(-0.10635180026292801)),(to_sfixed_a(-1.000860333442688)),(to_sfixed_a(-0.6008201241493225)),(to_sfixed_a(-0.11862306296825409)),(to_sfixed_a(0.018231648951768875)),(to_sfixed_a(0.052389875054359436)),(to_sfixed_a(0.07628178596496582)),(to_sfixed_a(0.02600097842514515)),(to_sfixed_a(-0.21686479449272156)),(to_sfixed_a(-0.04192506521940231)),(to_sfixed_a(-0.11591257899999619)),(to_sfixed_a(0.1594526767730713)),(to_sfixed_a(-0.11596780270338058)),(to_sfixed_a(5.668173253070563e-05)),(to_sfixed_a(0.0001900708011817187)),(to_sfixed_a(3.5649256460601464e-05)),(to_sfixed_a(-1.9898388927686028e-05)),(to_sfixed_a(-1.5767949662404135e-05)),(to_sfixed_a(0.00026676655397750437)),(to_sfixed_a(-0.0004127770662307739)),(to_sfixed_a(0.02321324311196804)),(to_sfixed_a(-0.0016866248333826661)),(to_sfixed_a(0.33113500475883484)),(to_sfixed_a(0.2597621977329254)),(to_sfixed_a(0.3336586356163025)),(to_sfixed_a(0.2080952227115631)),(to_sfixed_a(0.07999636232852936)),(to_sfixed_a(-0.1564386487007141)),(to_sfixed_a(-0.4122641980648041)),(to_sfixed_a(-0.43461543321609497)),(to_sfixed_a(-0.3556008040904999)),(to_sfixed_a(-0.026410339400172234)),(to_sfixed_a(-0.01071267481893301)),(to_sfixed_a(-0.0017643653554841876)),(to_sfixed_a(-0.0146456528455019)),(to_sfixed_a(0.06759600341320038)),(to_sfixed_a(-0.09161705523729324)),(to_sfixed_a(0.13319160044193268)),(to_sfixed_a(-0.031752802431583405)),(to_sfixed_a(-0.2904398441314697)),(to_sfixed_a(-0.07993413507938385)),(to_sfixed_a(0.0007966634002514184)),(to_sfixed_a(-0.0008455410716123879)),(to_sfixed_a(1.876511305454187e-05)),(to_sfixed_a(0.0004196178924757987)),(to_sfixed_a(0.0001832255657063797)),(to_sfixed_a(-0.00027009204495698214)),(to_sfixed_a(0.0002587421622592956)),(to_sfixed_a(0.000734908040612936)),(to_sfixed_a(-0.23254770040512085)),(to_sfixed_a(-0.12900231778621674)),(to_sfixed_a(-0.12354456633329391)),(to_sfixed_a(0.08002981543540955)),(to_sfixed_a(-0.050598084926605225)),(to_sfixed_a(-0.27685460448265076)),(to_sfixed_a(-0.28867027163505554)),(to_sfixed_a(-0.5138734579086304)),(to_sfixed_a(-0.5518394112586975)),(to_sfixed_a(-0.1858844757080078)),(to_sfixed_a(-0.06592327356338501)),(to_sfixed_a(-0.12789438664913177)),(to_sfixed_a(0.025132769718766212)),(to_sfixed_a(-0.12052864581346512)),(to_sfixed_a(0.03476757928729057)),(to_sfixed_a(0.1386222392320633)),(to_sfixed_a(-0.05617844685912132)),(to_sfixed_a(-0.08323962986469269)),(to_sfixed_a(-0.10947932302951813)),(to_sfixed_a(-0.07580853998661041)),(to_sfixed_a(0.0006555430591106415)),(to_sfixed_a(-0.00037046981742605567)),(to_sfixed_a(8.10919955256395e-05)),(to_sfixed_a(-0.0003239293291699141)),(to_sfixed_a(8.923489804146811e-05)),(to_sfixed_a(-0.00010886693780776113)),(to_sfixed_a(4.5346987462835386e-05)),(to_sfixed_a(0.0006977407610975206)),(to_sfixed_a(-0.15281568467617035)),(to_sfixed_a(-0.22375638782978058)),(to_sfixed_a(-0.17278257012367249)),(to_sfixed_a(-0.42845526337623596)),(to_sfixed_a(-0.4640854001045227)),(to_sfixed_a(-0.3036110997200012)),(to_sfixed_a(-0.07617364078760147)),(to_sfixed_a(-0.6459639072418213)),(to_sfixed_a(-0.15584884583950043)),(to_sfixed_a(0.06428574025630951)),(to_sfixed_a(-0.033667005598545074)),(to_sfixed_a(-0.08052632957696915)),(to_sfixed_a(-0.20986899733543396)),(to_sfixed_a(-0.11983710527420044)),(to_sfixed_a(-0.19168798625469208)),(to_sfixed_a(0.01806975156068802)),(to_sfixed_a(-0.00012450020585674793)),(to_sfixed_a(-0.04183003306388855)),(to_sfixed_a(0.04232274740934372)),(to_sfixed_a(-0.15747040510177612)),(to_sfixed_a(0.0005398993962444365)),(to_sfixed_a(9.354955545859411e-05)),(to_sfixed_a(2.2261374397203326e-05)),(to_sfixed_a(-8.017701475182548e-05)),(to_sfixed_a(-0.0001699502463452518)),(to_sfixed_a(-0.0001221669081132859)),(to_sfixed_a(-0.002159229712560773)),(to_sfixed_a(-0.19812782108783722)),(to_sfixed_a(-0.4480918347835541)),(to_sfixed_a(-0.6613483428955078)),(to_sfixed_a(-0.581009566783905)),(to_sfixed_a(-0.5267136693000793)),(to_sfixed_a(-0.30225688219070435)),(to_sfixed_a(-0.44810354709625244)),(to_sfixed_a(-0.7196164131164551)),(to_sfixed_a(-0.2504248023033142)),(to_sfixed_a(0.044508811086416245)),(to_sfixed_a(0.1393503099679947)),(to_sfixed_a(-0.07189001888036728)),(to_sfixed_a(0.04663173109292984)),(to_sfixed_a(-0.12836997210979462)),(to_sfixed_a(-0.23244088888168335)),(to_sfixed_a(0.04037269204854965)),(to_sfixed_a(0.18392693996429443)),(to_sfixed_a(0.11272135376930237)),(to_sfixed_a(0.10293149948120117)),(to_sfixed_a(-0.08098559826612473)),(to_sfixed_a(-0.13517123460769653)),(to_sfixed_a(-0.013234675861895084)),(to_sfixed_a(-0.0001262612349819392)),(to_sfixed_a(0.00024274722090922296)),(to_sfixed_a(-2.0544584913295694e-05)),(to_sfixed_a(-2.0719391613965854e-05)),(to_sfixed_a(-0.00215563434176147)),(to_sfixed_a(-0.00194527895655483)),(to_sfixed_a(-0.05993359163403511)),(to_sfixed_a(-0.5237751603126526)),(to_sfixed_a(-0.25645625591278076)),(to_sfixed_a(-0.4120888113975525)),(to_sfixed_a(-0.5088644623756409)),(to_sfixed_a(-0.7517213225364685)),(to_sfixed_a(-0.5788984298706055)),(to_sfixed_a(-0.7244095802307129)),(to_sfixed_a(-0.6656739115715027)),(to_sfixed_a(-0.07347289472818375)),(to_sfixed_a(-0.03545298054814339)),(to_sfixed_a(-0.10990608483552933)),(to_sfixed_a(-0.09601181000471115)),(to_sfixed_a(-0.09125560522079468)),(to_sfixed_a(-0.22919398546218872)),(to_sfixed_a(0.2565149962902069)),(to_sfixed_a(0.08938101679086685)),(to_sfixed_a(0.03638884797692299)),(to_sfixed_a(0.16043893992900848)),(to_sfixed_a(-0.009102188050746918)),(to_sfixed_a(-1.0302101145498455e-05)),(to_sfixed_a(6.867766933282837e-05)),(to_sfixed_a(1.8436023310641758e-05)),(to_sfixed_a(4.262938455212861e-05)),(to_sfixed_a(2.3675616830587387e-05)),(to_sfixed_a(1.57069371198304e-05)),(to_sfixed_a(0.00038443284574896097)),(to_sfixed_a(-0.028439609333872795)),(to_sfixed_a(-0.17702417075634003)),(to_sfixed_a(-0.18953409790992737)),(to_sfixed_a(-0.04204221069812775)),(to_sfixed_a(-0.20586401224136353)),(to_sfixed_a(-0.3273661136627197)),(to_sfixed_a(-0.45884713530540466)),(to_sfixed_a(-0.7734923958778381)),(to_sfixed_a(-0.7309437394142151)),(to_sfixed_a(-0.5150865316390991)),(to_sfixed_a(-0.43175220489501953)),(to_sfixed_a(-0.4055514931678772)),(to_sfixed_a(0.003475509351119399)),(to_sfixed_a(-0.31474003195762634)),(to_sfixed_a(-0.09928193688392639)),(to_sfixed_a(0.16976475715637207)),(to_sfixed_a(0.10151174664497375)),(to_sfixed_a(0.0876607820391655)),(to_sfixed_a(0.2938157618045807)),(to_sfixed_a(0.05375074967741966)),(to_sfixed_a(-0.06873451918363571)),(to_sfixed_a(-0.011287215165793896)),(to_sfixed_a(0.00010612221376504749)),(to_sfixed_a(0.00030060269637033343)),(to_sfixed_a(2.8522459615487605e-05)),(to_sfixed_a(-7.77409368311055e-05)),(to_sfixed_a(8.260262984549627e-05)),(to_sfixed_a(3.626470515882829e-06)),(to_sfixed_a(0.08914974331855774)),(to_sfixed_a(0.0001037342517520301)),(to_sfixed_a(0.02924932911992073)),(to_sfixed_a(-0.05896342918276787)),(to_sfixed_a(0.01642242632806301)),(to_sfixed_a(-0.01596798561513424)),(to_sfixed_a(-0.09728001803159714)),(to_sfixed_a(-0.1807948648929596)),(to_sfixed_a(-0.15801341831684113)),(to_sfixed_a(0.05759567394852638)),(to_sfixed_a(-0.13427649438381195)),(to_sfixed_a(-0.2853466272354126)),(to_sfixed_a(-0.25214698910713196)),(to_sfixed_a(0.09719198197126389)),(to_sfixed_a(-0.06962606310844421)),(to_sfixed_a(0.0716254711151123)),(to_sfixed_a(0.08855385333299637)),(to_sfixed_a(0.19391320645809174)),(to_sfixed_a(0.1979150027036667)),(to_sfixed_a(0.2021053433418274)),(to_sfixed_a(0.06655176728963852)),(to_sfixed_a(-5.813956249767216e-06)),(to_sfixed_a(2.2953809093451127e-05)),(to_sfixed_a(-5.6618129747221246e-05)),(to_sfixed_a(-6.259892870730255e-06)),(to_sfixed_a(-2.970324203488417e-05)),(to_sfixed_a(-2.0466522983042523e-05)),(to_sfixed_a(-0.00025184356491081417)),(to_sfixed_a(2.4107859644573182e-05)),(to_sfixed_a(0.009199727326631546)),(to_sfixed_a(0.12377321720123291)),(to_sfixed_a(0.2548149824142456)),(to_sfixed_a(-0.10981564968824387)),(to_sfixed_a(-0.11924973875284195)),(to_sfixed_a(0.22951342165470123)),(to_sfixed_a(0.01673518493771553)),(to_sfixed_a(0.0755213275551796)),(to_sfixed_a(0.11319441348314285)),(to_sfixed_a(0.04479336738586426)),(to_sfixed_a(0.00435182498767972)),(to_sfixed_a(0.138851597905159)),(to_sfixed_a(0.07974381744861603)),(to_sfixed_a(0.11172237992286682)),(to_sfixed_a(0.17215567827224731)),(to_sfixed_a(0.19718578457832336)),(to_sfixed_a(0.2736396789550781)),(to_sfixed_a(0.18543580174446106)),(to_sfixed_a(0.09474550187587738)),(to_sfixed_a(0.009368030354380608)),(to_sfixed_a(-0.055667247623205185)),(to_sfixed_a(7.543966785306111e-05)),(to_sfixed_a(2.7144609703100286e-05)),(to_sfixed_a(-0.00017310146358795464)),(to_sfixed_a(-0.0003121832851320505)),(to_sfixed_a(-1.2830599189328495e-05)),(to_sfixed_a(-0.0001795871212380007)),(to_sfixed_a(7.063219527481124e-05)),(to_sfixed_a(0.007966653443872929)),(to_sfixed_a(-0.00013461419439408928)),(to_sfixed_a(0.07496341317892075)),(to_sfixed_a(-0.15035302937030792)),(to_sfixed_a(0.13481956720352173)),(to_sfixed_a(0.10090208053588867)),(to_sfixed_a(0.2863950729370117)),(to_sfixed_a(0.21036048233509064)),(to_sfixed_a(0.20808930695056915)),(to_sfixed_a(0.20014223456382751)),(to_sfixed_a(0.6231687664985657)),(to_sfixed_a(0.2527686655521393)),(to_sfixed_a(0.10916177928447723)),(to_sfixed_a(0.44955354928970337)),(to_sfixed_a(0.3046662509441376)),(to_sfixed_a(0.17162349820137024)),(to_sfixed_a(0.19825966656208038)),(to_sfixed_a(0.024780577048659325)),(to_sfixed_a(-0.008183087222278118)),(to_sfixed_a(-0.0011503173736855388)),(to_sfixed_a(0.010639741085469723)),(to_sfixed_a(-0.00012744682317133993)),(to_sfixed_a(0.00011702194024110213)),(to_sfixed_a(2.6003483071690425e-05)),(to_sfixed_a(4.7951427404768765e-05)),(to_sfixed_a(2.3158716430771165e-05)),(to_sfixed_a(-3.0310251531773247e-05)),(to_sfixed_a(-1.889622217277065e-05)),(to_sfixed_a(0.00018909707432612777)),(to_sfixed_a(0.028885290026664734)),(to_sfixed_a(-0.011383689939975739)),(to_sfixed_a(-0.005020097829401493)),(to_sfixed_a(0.10666989535093307)),(to_sfixed_a(-0.011287832632660866)),(to_sfixed_a(0.10193236917257309)),(to_sfixed_a(0.18331889808177948)),(to_sfixed_a(0.17235726118087769)),(to_sfixed_a(0.21106646955013275)),(to_sfixed_a(0.255526065826416)),(to_sfixed_a(0.18471920490264893)),(to_sfixed_a(0.3005519509315491)),(to_sfixed_a(0.1611267626285553)),(to_sfixed_a(0.5336921811103821)),(to_sfixed_a(0.3535763919353485)),(to_sfixed_a(-0.00873473659157753)),(to_sfixed_a(-0.031048541888594627)),(to_sfixed_a(-0.026737263426184654)),(to_sfixed_a(-0.0057756248861551285)),(to_sfixed_a(2.656649303389713e-05)),(to_sfixed_a(-1.8788439319905592e-06)),(to_sfixed_a(5.7445478887530044e-05)),(to_sfixed_a(4.2373059841338545e-05)),(to_sfixed_a(-7.102871313691139e-05)),(to_sfixed_a(0.00011870759772136807)),(to_sfixed_a(-2.1482193915289827e-05)),(to_sfixed_a(-5.112544386065565e-06)),(to_sfixed_a(0.00045476839295588434)),(to_sfixed_a(-0.02161298878490925)),(to_sfixed_a(-0.08644045144319534)),(to_sfixed_a(0.13033106923103333)),(to_sfixed_a(-0.1896180659532547)),(to_sfixed_a(0.021097207441926003)),(to_sfixed_a(0.17922717332839966)),(to_sfixed_a(0.35223641991615295)),(to_sfixed_a(0.12011507153511047)),(to_sfixed_a(0.11157641559839249)),(to_sfixed_a(0.18310566246509552)),(to_sfixed_a(0.23034271597862244)),(to_sfixed_a(0.3253977596759796)),(to_sfixed_a(0.4055330753326416)),(to_sfixed_a(0.23895718157291412)),(to_sfixed_a(0.04330919682979584)),(to_sfixed_a(0.12362223118543625)),(to_sfixed_a(-0.03736328333616257)),(to_sfixed_a(-0.01191723719239235)),(to_sfixed_a(-0.021005060523748398)),(to_sfixed_a(-0.00015735281340312213)),(to_sfixed_a(0.0001235272065969184)),(to_sfixed_a(8.38914347696118e-05)),(to_sfixed_a(9.663157106842846e-05)),(to_sfixed_a(1.8260918750456767e-06)),(to_sfixed_a(-0.00010815774294314906)),(to_sfixed_a(-0.0001483290980104357)),(to_sfixed_a(-1.8561002434580587e-05)),(to_sfixed_a(-0.006029751151800156)),(to_sfixed_a(-0.028321081772446632)),(to_sfixed_a(-0.02508191019296646)),(to_sfixed_a(0.23034480214118958)),(to_sfixed_a(0.29168587923049927)),(to_sfixed_a(0.14787410199642181)),(to_sfixed_a(0.02707662247121334)),(to_sfixed_a(0.1857692450284958)),(to_sfixed_a(0.3328527510166168)),(to_sfixed_a(0.2538491487503052)),(to_sfixed_a(0.19999614357948303)),(to_sfixed_a(0.11154606193304062)),(to_sfixed_a(0.30030977725982666)),(to_sfixed_a(0.17439693212509155)),(to_sfixed_a(0.08389919996261597)),(to_sfixed_a(0.04489239677786827)),(to_sfixed_a(0.005246683489531279)),(to_sfixed_a(-0.029396522790193558)),(to_sfixed_a(-0.01811262033879757)),(to_sfixed_a(-0.011996302753686905)),(to_sfixed_a(0.00018241227371618152)),(to_sfixed_a(1.164700461231405e-05)),(to_sfixed_a(6.037639832356945e-05)),(to_sfixed_a(-0.0002508853795006871)),(to_sfixed_a(9.305392450187355e-05)),(to_sfixed_a(-2.3494192191719776e-06)),(to_sfixed_a(3.0469391276710667e-05)),(to_sfixed_a(8.529268234269693e-05)),(to_sfixed_a(0.00019846041686832905)),(to_sfixed_a(-0.009621236473321915)),(to_sfixed_a(-0.015412342734634876)),(to_sfixed_a(0.012173130176961422)),(to_sfixed_a(0.1452757865190506)),(to_sfixed_a(0.04970735311508179)),(to_sfixed_a(0.16581737995147705)),(to_sfixed_a(-0.03705650568008423)),(to_sfixed_a(-0.04041766747832298)),(to_sfixed_a(0.016109030693769455)),(to_sfixed_a(0.05761362984776497)),(to_sfixed_a(0.1785314977169037)),(to_sfixed_a(0.004383646417409182)),(to_sfixed_a(0.11046615988016129)),(to_sfixed_a(-0.0028294799849390984)),(to_sfixed_a(-0.04008569195866585)),(to_sfixed_a(-0.03972348943352699)),(to_sfixed_a(-0.0009001002181321383)),(to_sfixed_a(-0.0037245501298457384)),(to_sfixed_a(-0.0038703589234501123)),(to_sfixed_a(-0.00010228257451672107)),(to_sfixed_a(8.944643195718527e-05)),(to_sfixed_a(8.734522998565808e-05)),(to_sfixed_a(-7.960800576256588e-05)),(to_sfixed_a(0.0001027667531161569)),(to_sfixed_a(9.2923546617385e-06)),(to_sfixed_a(0.00029011836159043014)),(to_sfixed_a(-7.368185470113531e-05)),(to_sfixed_a(-0.00015152647392824292)),(to_sfixed_a(-0.0008999009151011705)),(to_sfixed_a(-0.0009089261875487864)),(to_sfixed_a(-0.00011166262265760452)),(to_sfixed_a(-0.00015216761676128954)),(to_sfixed_a(0.0004235798551235348)),(to_sfixed_a(-0.049634821712970734)),(to_sfixed_a(-0.0012607596581801772)),(to_sfixed_a(-0.0027735892217606306)),(to_sfixed_a(-0.03318282961845398)),(to_sfixed_a(-0.010559783317148685)),(to_sfixed_a(4.1356088331667706e-05)),(to_sfixed_a(0.008374648168683052)),(to_sfixed_a(-0.03827548399567604)),(to_sfixed_a(-0.0535566620528698)),(to_sfixed_a(0.0005565852043218911)),(to_sfixed_a(0.0011358227347955108)),(to_sfixed_a(2.7171345209353603e-05)),(to_sfixed_a(-2.5299374101450667e-05)),(to_sfixed_a(-7.990535232238472e-05)),(to_sfixed_a(1.6984114381557447e-06)),(to_sfixed_a(-5.1848208386218175e-05)),(to_sfixed_a(9.672019950812683e-05)),(to_sfixed_a(-0.00026839543716050684)),(to_sfixed_a(-0.00023862232046667486)),(to_sfixed_a(-0.00021190183178987354)),(to_sfixed_a(0.0004985760897397995)),(to_sfixed_a(3.9228994864970446e-05)),(to_sfixed_a(1.5647106010874268e-07)),(to_sfixed_a(5.454788697534241e-05)),(to_sfixed_a(2.998302261403296e-05)),(to_sfixed_a(-0.0002606099587865174)),(to_sfixed_a(-5.116672764415853e-05)),(to_sfixed_a(0.0002094270457746461)),(to_sfixed_a(4.58380272903014e-05)),(to_sfixed_a(1.7410578948329203e-05)),(to_sfixed_a(-9.029382636072114e-05)),(to_sfixed_a(0.00010505507816560566)),(to_sfixed_a(-0.00040695126517675817)),(to_sfixed_a(0.0002714160946197808)),(to_sfixed_a(-0.0002544414019212127)),(to_sfixed_a(-0.00018399477994535118)),(to_sfixed_a(-2.4036153263296e-05)),(to_sfixed_a(-9.459985449211672e-05)),(to_sfixed_a(0.0001307574420934543)),(to_sfixed_a(4.7482702939305454e-05)),(to_sfixed_a(0.00023809749109204859)),(to_sfixed_a(2.8466511139413342e-05)),(to_sfixed_a(3.972628292103764e-06)),(to_sfixed_a(0.00020921436953358352)),(to_sfixed_a(9.12086688913405e-05)),(to_sfixed_a(-8.519346010871232e-05)));

    constant weight_n0_2 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-8.046497532632202e-05)),(to_sfixed_a(-0.00021497736452147365)),(to_sfixed_a(-7.800923776812851e-05)),(to_sfixed_a(-0.00034050093381665647)),(to_sfixed_a(-9.467040217714384e-05)),(to_sfixed_a(-0.00012576904555317014)),(to_sfixed_a(-4.1941399103961885e-05)),(to_sfixed_a(-0.000198495268705301)),(to_sfixed_a(-9.880152356345206e-05)),(to_sfixed_a(2.151266744476743e-05)),(to_sfixed_a(9.966000106942374e-06)),(to_sfixed_a(8.74432225828059e-05)),(to_sfixed_a(0.00027326084091328084)),(to_sfixed_a(1.6597075955360197e-05)),(to_sfixed_a(0.0002451194741297513)),(to_sfixed_a(1.3753705388808157e-05)),(to_sfixed_a(0.0002992683439515531)),(to_sfixed_a(-1.3271174793771934e-05)),(to_sfixed_a(1.5688727216911502e-05)),(to_sfixed_a(-0.00012186792446300387)),(to_sfixed_a(9.607452375348657e-05)),(to_sfixed_a(-8.294293365906924e-06)),(to_sfixed_a(-0.0001717723353067413)),(to_sfixed_a(-7.004081271588802e-05)),(to_sfixed_a(-0.00017270130047108978)),(to_sfixed_a(-0.00021547543292399496)),(to_sfixed_a(-0.00022217599325813353)),(to_sfixed_a(-6.959180609555915e-05)),(to_sfixed_a(-0.00015004960005171597)),(to_sfixed_a(-6.816672976128757e-05)),(to_sfixed_a(-2.2419179003918543e-05)),(to_sfixed_a(-0.00023070855240803212)),(to_sfixed_a(-3.7546433304669335e-05)),(to_sfixed_a(-0.00014923540584277362)),(to_sfixed_a(-0.00011305208317935467)),(to_sfixed_a(9.655670874053612e-05)),(to_sfixed_a(-6.0402544477256015e-05)),(to_sfixed_a(1.694825004960876e-05)),(to_sfixed_a(7.30056272004731e-05)),(to_sfixed_a(-1.996393984882161e-05)),(to_sfixed_a(-0.0001226376771228388)),(to_sfixed_a(0.00021990634559188038)),(to_sfixed_a(0.0002505687880329788)),(to_sfixed_a(0.00021125079365447164)),(to_sfixed_a(-3.330527397338301e-05)),(to_sfixed_a(3.287622530478984e-05)),(to_sfixed_a(-5.408283323049545e-05)),(to_sfixed_a(-2.629245318530593e-05)),(to_sfixed_a(7.622454722877592e-05)),(to_sfixed_a(6.552118429681286e-05)),(to_sfixed_a(1.83952615770977e-05)),(to_sfixed_a(-0.00016088184202089906)),(to_sfixed_a(-0.0001557412906549871)),(to_sfixed_a(-0.0002603639441076666)),(to_sfixed_a(6.61132944514975e-05)),(to_sfixed_a(3.4807835618266836e-05)),(to_sfixed_a(0.00020228014909662306)),(to_sfixed_a(5.392169623519294e-05)),(to_sfixed_a(-4.167861334281042e-05)),(to_sfixed_a(4.7956556954886764e-05)),(to_sfixed_a(-8.46033071866259e-05)),(to_sfixed_a(-0.0001766938657965511)),(to_sfixed_a(-3.502970139379613e-05)),(to_sfixed_a(0.00016178189252968878)),(to_sfixed_a(-5.382686867960729e-05)),(to_sfixed_a(-6.074002885725349e-05)),(to_sfixed_a(0.00012629076081793755)),(to_sfixed_a(2.435796159261372e-05)),(to_sfixed_a(-0.00013613338524010032)),(to_sfixed_a(-0.013901925645768642)),(to_sfixed_a(-4.230552076478489e-05)),(to_sfixed_a(6.718378426739946e-05)),(to_sfixed_a(2.7330186640028842e-05)),(to_sfixed_a(3.81971440219786e-05)),(to_sfixed_a(-3.588470281101763e-05)),(to_sfixed_a(0.00015569939569104463)),(to_sfixed_a(9.975124703487381e-05)),(to_sfixed_a(3.188827759004198e-05)),(to_sfixed_a(-6.339469837257639e-05)),(to_sfixed_a(0.00039511261275038123)),(to_sfixed_a(-1.053434971254319e-05)),(to_sfixed_a(0.00029609212651848793)),(to_sfixed_a(4.86536773678381e-05)),(to_sfixed_a(0.00019918310863431543)),(to_sfixed_a(-0.00020733449491672218)),(to_sfixed_a(0.0002410007145954296)),(to_sfixed_a(8.234195411205292e-05)),(to_sfixed_a(0.00015448257909156382)),(to_sfixed_a(0.00021931083756498992)),(to_sfixed_a(-2.571324102973449e-06)),(to_sfixed_a(0.00011838311183964834)),(to_sfixed_a(-0.0003543666680343449)),(to_sfixed_a(-0.03712580353021622)),(to_sfixed_a(-0.00013374697300605476)),(to_sfixed_a(-0.04202292859554291)),(to_sfixed_a(0.06483080238103867)),(to_sfixed_a(-0.010559549555182457)),(to_sfixed_a(-0.05946572870016098)),(to_sfixed_a(-0.06034732982516289)),(to_sfixed_a(0.006176332011818886)),(to_sfixed_a(-0.008178699761629105)),(to_sfixed_a(0.06311624497175217)),(to_sfixed_a(0.08187630772590637)),(to_sfixed_a(-0.07543785870075226)),(to_sfixed_a(-0.02619217522442341)),(to_sfixed_a(-0.05358433723449707)),(to_sfixed_a(5.26852672919631e-05)),(to_sfixed_a(-5.253153631201712e-06)),(to_sfixed_a(4.780920426128432e-05)),(to_sfixed_a(8.373360469704494e-05)),(to_sfixed_a(0.00015810722834430635)),(to_sfixed_a(0.00011613511014729738)),(to_sfixed_a(-0.00023160949058365077)),(to_sfixed_a(-5.660421606989985e-07)),(to_sfixed_a(1.2309151316003408e-05)),(to_sfixed_a(-3.1349183700513095e-05)),(to_sfixed_a(4.77614848932717e-05)),(to_sfixed_a(0.0001520778314443305)),(to_sfixed_a(4.114174589631148e-05)),(to_sfixed_a(0.033097922801971436)),(to_sfixed_a(0.04261365160346031)),(to_sfixed_a(-0.055285368114709854)),(to_sfixed_a(-0.15594437718391418)),(to_sfixed_a(0.11077339202165604)),(to_sfixed_a(-0.01772802136838436)),(to_sfixed_a(-0.17064614593982697)),(to_sfixed_a(0.030253687873482704)),(to_sfixed_a(-0.23340418934822083)),(to_sfixed_a(0.027274208143353462)),(to_sfixed_a(-0.18800504505634308)),(to_sfixed_a(-0.04667464643716812)),(to_sfixed_a(0.015226611867547035)),(to_sfixed_a(-0.014678815379738808)),(to_sfixed_a(-0.11159133911132812)),(to_sfixed_a(0.07231070101261139)),(to_sfixed_a(0.00011187101335963234)),(to_sfixed_a(0.0025297622196376324)),(to_sfixed_a(-0.0002649862435646355)),(to_sfixed_a(0.0001494980970164761)),(to_sfixed_a(-2.7254474844085053e-05)),(to_sfixed_a(-6.833514635218307e-05)),(to_sfixed_a(0.00014255658606998622)),(to_sfixed_a(-0.00016940044588409364)),(to_sfixed_a(2.5909550458891317e-05)),(to_sfixed_a(-0.0023092997726053)),(to_sfixed_a(0.030905690044164658)),(to_sfixed_a(-0.01643521524965763)),(to_sfixed_a(0.03400541469454765)),(to_sfixed_a(0.037405163049697876)),(to_sfixed_a(-0.03665921464562416)),(to_sfixed_a(-0.08572860807180405)),(to_sfixed_a(-0.07401634007692337)),(to_sfixed_a(0.0342421792447567)),(to_sfixed_a(0.2377559244632721)),(to_sfixed_a(0.04451458528637886)),(to_sfixed_a(0.06361914426088333)),(to_sfixed_a(-0.11630585789680481)),(to_sfixed_a(-0.19666670262813568)),(to_sfixed_a(-0.3075977861881256)),(to_sfixed_a(-0.43642354011535645)),(to_sfixed_a(0.042739301919937134)),(to_sfixed_a(-0.04871977120637894)),(to_sfixed_a(-0.0008894979837350547)),(to_sfixed_a(-0.02616673894226551)),(to_sfixed_a(0.002930411836132407)),(to_sfixed_a(0.00016453703574370593)),(to_sfixed_a(-4.172547778580338e-05)),(to_sfixed_a(-1.954985918928287e-06)),(to_sfixed_a(0.0001180809922516346)),(to_sfixed_a(-0.00018875881505664438)),(to_sfixed_a(-0.00012736588541883975)),(to_sfixed_a(-0.0002375811745878309)),(to_sfixed_a(0.00015834026271477342)),(to_sfixed_a(0.03381197527050972)),(to_sfixed_a(0.056657835841178894)),(to_sfixed_a(-0.09783504158258438)),(to_sfixed_a(-0.11964485049247742)),(to_sfixed_a(-0.08275943249464035)),(to_sfixed_a(-0.019037611782550812)),(to_sfixed_a(0.0663292407989502)),(to_sfixed_a(0.07175040245056152)),(to_sfixed_a(0.2025667130947113)),(to_sfixed_a(-0.06546350568532944)),(to_sfixed_a(-0.07795733213424683)),(to_sfixed_a(0.031704097986221313)),(to_sfixed_a(0.040597207844257355)),(to_sfixed_a(-0.19469930231571198)),(to_sfixed_a(-0.04377727955579758)),(to_sfixed_a(-0.13771909475326538)),(to_sfixed_a(-0.043989624828100204)),(to_sfixed_a(0.10480157285928726)),(to_sfixed_a(-0.031446199864149094)),(to_sfixed_a(0.004879345186054707)),(to_sfixed_a(0.006745800841599703)),(to_sfixed_a(0.0037883431650698185)),(to_sfixed_a(1.993447949644178e-05)),(to_sfixed_a(0.0003269196895416826)),(to_sfixed_a(-4.777437789016403e-05)),(to_sfixed_a(-0.00015534851991105825)),(to_sfixed_a(-0.00013779631990473717)),(to_sfixed_a(-0.0001030407875077799)),(to_sfixed_a(-0.04393536224961281)),(to_sfixed_a(0.21495819091796875)),(to_sfixed_a(0.04138920083642006)),(to_sfixed_a(-0.004495030269026756)),(to_sfixed_a(0.07532570511102676)),(to_sfixed_a(0.2809191942214966)),(to_sfixed_a(0.2525319755077362)),(to_sfixed_a(0.22708050906658173)),(to_sfixed_a(0.2351721227169037)),(to_sfixed_a(0.29321467876434326)),(to_sfixed_a(0.011112726293504238)),(to_sfixed_a(-0.04569646716117859)),(to_sfixed_a(-0.11200028657913208)),(to_sfixed_a(0.05242345109581947)),(to_sfixed_a(-0.09925518184900284)),(to_sfixed_a(0.03325355052947998)),(to_sfixed_a(0.13678669929504395)),(to_sfixed_a(0.07704155147075653)),(to_sfixed_a(0.24172794818878174)),(to_sfixed_a(-0.007461287081241608)),(to_sfixed_a(0.004747301805764437)),(to_sfixed_a(-0.000329188333125785)),(to_sfixed_a(2.8778180421795696e-05)),(to_sfixed_a(-0.00033925718162208796)),(to_sfixed_a(8.379239443456754e-05)),(to_sfixed_a(-0.000281765271211043)),(to_sfixed_a(7.52956184442155e-05)),(to_sfixed_a(0.03458494693040848)),(to_sfixed_a(-0.027823330834507942)),(to_sfixed_a(-0.05713890492916107)),(to_sfixed_a(0.04735632985830307)),(to_sfixed_a(-0.04746927320957184)),(to_sfixed_a(-0.04047684371471405)),(to_sfixed_a(0.20973296463489532)),(to_sfixed_a(-0.10083678364753723)),(to_sfixed_a(-0.040781084448099136)),(to_sfixed_a(0.021377356722950935)),(to_sfixed_a(0.23189713060855865)),(to_sfixed_a(0.2325848788022995)),(to_sfixed_a(0.18652120232582092)),(to_sfixed_a(0.16631188988685608)),(to_sfixed_a(0.2830381989479065)),(to_sfixed_a(0.03163385018706322)),(to_sfixed_a(0.23792065680027008)),(to_sfixed_a(0.06411122530698776)),(to_sfixed_a(0.07487621158361435)),(to_sfixed_a(0.14936280250549316)),(to_sfixed_a(0.12478097528219223)),(to_sfixed_a(-0.020670086145401)),(to_sfixed_a(-2.3126629457692616e-05)),(to_sfixed_a(-5.2696643251692876e-05)),(to_sfixed_a(0.00015985951176844537)),(to_sfixed_a(5.896803122595884e-05)),(to_sfixed_a(-2.750955354713369e-05)),(to_sfixed_a(2.1490042854566127e-05)),(to_sfixed_a(-6.0933591157663614e-05)),(to_sfixed_a(0.09548569470643997)),(to_sfixed_a(-0.005432402715086937)),(to_sfixed_a(0.04056327044963837)),(to_sfixed_a(-0.06314102560281754)),(to_sfixed_a(-0.09919778257608414)),(to_sfixed_a(-0.15032082796096802)),(to_sfixed_a(-0.24648135900497437)),(to_sfixed_a(-0.04296896606683731)),(to_sfixed_a(0.1606224924325943)),(to_sfixed_a(0.39095771312713623)),(to_sfixed_a(0.11053693294525146)),(to_sfixed_a(0.3789867162704468)),(to_sfixed_a(0.5841196179389954)),(to_sfixed_a(0.3954850435256958)),(to_sfixed_a(0.4626889228820801)),(to_sfixed_a(0.2674252390861511)),(to_sfixed_a(0.28185704350471497)),(to_sfixed_a(0.20767028629779816)),(to_sfixed_a(-0.02264704927802086)),(to_sfixed_a(0.06494763493537903)),(to_sfixed_a(-0.00012406756286509335)),(to_sfixed_a(9.675849287305027e-05)),(to_sfixed_a(-8.382752275792882e-05)),(to_sfixed_a(-0.00011441489186836407)),(to_sfixed_a(0.0001951876183738932)),(to_sfixed_a(-0.00018872212967835367)),(to_sfixed_a(-0.000111132234451361)),(to_sfixed_a(-0.0024721012450754642)),(to_sfixed_a(-0.08100222796201706)),(to_sfixed_a(-0.2883315682411194)),(to_sfixed_a(-0.1466139256954193)),(to_sfixed_a(-0.16924414038658142)),(to_sfixed_a(-0.2775673568248749)),(to_sfixed_a(-0.3293459713459015)),(to_sfixed_a(-0.38841524720191956)),(to_sfixed_a(-0.32050374150276184)),(to_sfixed_a(-0.004264062736183405)),(to_sfixed_a(-0.21746651828289032)),(to_sfixed_a(-0.17907555401325226)),(to_sfixed_a(0.015274935401976109)),(to_sfixed_a(-0.0668424442410469)),(to_sfixed_a(0.121919184923172)),(to_sfixed_a(0.23036399483680725)),(to_sfixed_a(0.2192114144563675)),(to_sfixed_a(0.1676129400730133)),(to_sfixed_a(0.03722633793950081)),(to_sfixed_a(0.10660218447446823)),(to_sfixed_a(0.008753941394388676)),(to_sfixed_a(0.031019551679491997)),(to_sfixed_a(7.85877782618627e-05)),(to_sfixed_a(4.6835135435685515e-05)),(to_sfixed_a(0.00015721269301138818)),(to_sfixed_a(-0.00026953144697472453)),(to_sfixed_a(-0.00010112202289747074)),(to_sfixed_a(0.027192698791623116)),(to_sfixed_a(-0.01659001223742962)),(to_sfixed_a(-0.19275610148906708)),(to_sfixed_a(-0.15221895277500153)),(to_sfixed_a(-0.2723161280155182)),(to_sfixed_a(-0.24958805739879608)),(to_sfixed_a(-0.14891625940799713)),(to_sfixed_a(-0.16902709007263184)),(to_sfixed_a(-0.04607589170336723)),(to_sfixed_a(-0.1990983784198761)),(to_sfixed_a(-0.1893664449453354)),(to_sfixed_a(-0.27921900153160095)),(to_sfixed_a(-0.39842742681503296)),(to_sfixed_a(-0.18280363082885742)),(to_sfixed_a(-0.1309550255537033)),(to_sfixed_a(-0.1157461404800415)),(to_sfixed_a(-0.23442144691944122)),(to_sfixed_a(-0.15195703506469727)),(to_sfixed_a(-0.08639512211084366)),(to_sfixed_a(-0.012178189121186733)),(to_sfixed_a(0.1751207560300827)),(to_sfixed_a(0.0539078563451767)),(to_sfixed_a(0.00013788664364255965)),(to_sfixed_a(0.00017814985767472535)),(to_sfixed_a(0.00021084527543280274)),(to_sfixed_a(0.0001413580175722018)),(to_sfixed_a(-0.00019976546172983944)),(to_sfixed_a(-0.0001841574558056891)),(to_sfixed_a(-1.986670667974977e-06)),(to_sfixed_a(-0.058800436556339264)),(to_sfixed_a(-0.034693293273448944)),(to_sfixed_a(-0.11884085088968277)),(to_sfixed_a(-0.2014032006263733)),(to_sfixed_a(-0.24271270632743835)),(to_sfixed_a(-0.016787396743893623)),(to_sfixed_a(0.15800654888153076)),(to_sfixed_a(0.023693235591053963)),(to_sfixed_a(0.26063627004623413)),(to_sfixed_a(0.07389640063047409)),(to_sfixed_a(-0.48365604877471924)),(to_sfixed_a(0.062062256038188934)),(to_sfixed_a(-0.33602288365364075)),(to_sfixed_a(-0.18108916282653809)),(to_sfixed_a(-0.11801356822252274)),(to_sfixed_a(-0.1866394579410553)),(to_sfixed_a(-0.19655410945415497)),(to_sfixed_a(-0.08423301577568054)),(to_sfixed_a(0.04571239650249481)),(to_sfixed_a(0.1237277090549469)),(to_sfixed_a(0.04933636635541916)),(to_sfixed_a(6.90786910126917e-05)),(to_sfixed_a(-0.0005909380852244794)),(to_sfixed_a(-0.00018172364798374474)),(to_sfixed_a(7.069685671012849e-05)),(to_sfixed_a(8.112679643090814e-05)),(to_sfixed_a(0.00041109442827291787)),(to_sfixed_a(-0.0003305696591269225)),(to_sfixed_a(-0.0032643405720591545)),(to_sfixed_a(-0.1053062304854393)),(to_sfixed_a(0.005343011114746332)),(to_sfixed_a(0.12474069744348526)),(to_sfixed_a(0.28573018312454224)),(to_sfixed_a(0.24998432397842407)),(to_sfixed_a(0.5403307676315308)),(to_sfixed_a(0.4954317808151245)),(to_sfixed_a(0.4076622426509857)),(to_sfixed_a(-0.5955532789230347)),(to_sfixed_a(-0.3282550275325775)),(to_sfixed_a(-0.1756996363401413)),(to_sfixed_a(-0.1378004401922226)),(to_sfixed_a(-0.04438969865441322)),(to_sfixed_a(-0.0016634096391499043)),(to_sfixed_a(-0.10675831884145737)),(to_sfixed_a(-0.05461210384964943)),(to_sfixed_a(0.09707241505384445)),(to_sfixed_a(-0.03127073869109154)),(to_sfixed_a(-0.03506944701075554)),(to_sfixed_a(-0.04916964843869209)),(to_sfixed_a(-0.0019361150916665792)),(to_sfixed_a(-0.0026076443027704954)),(to_sfixed_a(-0.00036698594340123236)),(to_sfixed_a(-9.736007632454857e-05)),(to_sfixed_a(4.092873859917745e-05)),(to_sfixed_a(-0.0005250826943665743)),(to_sfixed_a(9.256729390472174e-05)),(to_sfixed_a(-0.00021924928296357393)),(to_sfixed_a(0.23040498793125153)),(to_sfixed_a(0.3225906789302826)),(to_sfixed_a(0.4190056324005127)),(to_sfixed_a(0.4204423725605011)),(to_sfixed_a(0.562482476234436)),(to_sfixed_a(0.5719210505485535)),(to_sfixed_a(0.5826961994171143)),(to_sfixed_a(-0.06769419461488724)),(to_sfixed_a(-0.3103181719779968)),(to_sfixed_a(-0.16526155173778534)),(to_sfixed_a(0.06650129705667496)),(to_sfixed_a(0.062369588762521744)),(to_sfixed_a(0.02733718417584896)),(to_sfixed_a(0.02994246780872345)),(to_sfixed_a(0.03281114250421524)),(to_sfixed_a(0.01722577214241028)),(to_sfixed_a(-0.013224946334958076)),(to_sfixed_a(-0.04415766894817352)),(to_sfixed_a(-0.004257677588611841)),(to_sfixed_a(0.044752806425094604)),(to_sfixed_a(0.000503901916090399)),(to_sfixed_a(-0.00011381587682990357)),(to_sfixed_a(-5.6065571698127314e-05)),(to_sfixed_a(-0.00030445700394921005)),(to_sfixed_a(-0.0002947460161522031)),(to_sfixed_a(-6.281778769334778e-05)),(to_sfixed_a(8.773433364694938e-05)),(to_sfixed_a(0.0484701506793499)),(to_sfixed_a(0.37800872325897217)),(to_sfixed_a(0.32101765275001526)),(to_sfixed_a(0.6299644708633423)),(to_sfixed_a(0.9291806817054749)),(to_sfixed_a(1.0386760234832764)),(to_sfixed_a(0.6663742661476135)),(to_sfixed_a(0.0007215588702820241)),(to_sfixed_a(-0.327618807554245)),(to_sfixed_a(-0.3807973265647888)),(to_sfixed_a(-0.04639629274606705)),(to_sfixed_a(0.056364916265010834)),(to_sfixed_a(0.08513420820236206)),(to_sfixed_a(0.06269410252571106)),(to_sfixed_a(0.07793832570314407)),(to_sfixed_a(-0.07603270560503006)),(to_sfixed_a(-0.02268722839653492)),(to_sfixed_a(0.011316142044961452)),(to_sfixed_a(-0.03097177855670452)),(to_sfixed_a(0.03482230380177498)),(to_sfixed_a(0.001905175275169313)),(to_sfixed_a(0.0001255307870451361)),(to_sfixed_a(-4.900573185295798e-05)),(to_sfixed_a(0.00022155093029141426)),(to_sfixed_a(0.00023760604381095618)),(to_sfixed_a(0.00018918892601504922)),(to_sfixed_a(-0.0001670526253292337)),(to_sfixed_a(-0.0018200764898210764)),(to_sfixed_a(0.20260265469551086)),(to_sfixed_a(0.2041664868593216)),(to_sfixed_a(0.1646900624036789)),(to_sfixed_a(0.23022107779979706)),(to_sfixed_a(0.2692358195781708)),(to_sfixed_a(0.15761470794677734)),(to_sfixed_a(0.4294603765010834)),(to_sfixed_a(0.2442491203546524)),(to_sfixed_a(0.12715835869312286)),(to_sfixed_a(-0.260885089635849)),(to_sfixed_a(0.02979397401213646)),(to_sfixed_a(0.04429611191153526)),(to_sfixed_a(0.1401626169681549)),(to_sfixed_a(0.09262917935848236)),(to_sfixed_a(0.08194316923618317)),(to_sfixed_a(-0.06558866053819656)),(to_sfixed_a(-0.20541620254516602)),(to_sfixed_a(-0.09335830062627792)),(to_sfixed_a(-0.034963954240083694)),(to_sfixed_a(-0.08607024699449539)),(to_sfixed_a(-0.04137187451124191)),(to_sfixed_a(-0.009350634180009365)),(to_sfixed_a(-7.486460526706651e-05)),(to_sfixed_a(-0.00013390071399044245)),(to_sfixed_a(-7.736308180028573e-05)),(to_sfixed_a(2.5133011149591766e-05)),(to_sfixed_a(-0.0009249974391423166)),(to_sfixed_a(-0.001766917179338634)),(to_sfixed_a(-0.0070245093666017056)),(to_sfixed_a(0.09241864830255508)),(to_sfixed_a(-0.23230817914009094)),(to_sfixed_a(-0.07433094829320908)),(to_sfixed_a(-0.01894909143447876)),(to_sfixed_a(-0.3142315745353699)),(to_sfixed_a(-0.18847014009952545)),(to_sfixed_a(-0.4457690715789795)),(to_sfixed_a(-0.3911404311656952)),(to_sfixed_a(0.19959315657615662)),(to_sfixed_a(0.12443411350250244)),(to_sfixed_a(0.18592457473278046)),(to_sfixed_a(0.1941027045249939)),(to_sfixed_a(0.08940070867538452)),(to_sfixed_a(0.07256219536066055)),(to_sfixed_a(-0.25934872031211853)),(to_sfixed_a(0.06915844976902008)),(to_sfixed_a(-0.06839227676391602)),(to_sfixed_a(-0.0035718013532459736)),(to_sfixed_a(-0.020633768290281296)),(to_sfixed_a(0.00015886491746641695)),(to_sfixed_a(0.00016803173639345914)),(to_sfixed_a(0.00033704008092172444)),(to_sfixed_a(0.00022234077914617956)),(to_sfixed_a(0.0002423685509711504)),(to_sfixed_a(7.861519407015294e-05)),(to_sfixed_a(-0.00017766020027920604)),(to_sfixed_a(-0.019919883459806442)),(to_sfixed_a(-0.024144653230905533)),(to_sfixed_a(-0.3650911748409271)),(to_sfixed_a(-0.22970759868621826)),(to_sfixed_a(-0.33384859561920166)),(to_sfixed_a(-0.33790677785873413)),(to_sfixed_a(-0.28510168194770813)),(to_sfixed_a(-0.8431485295295715)),(to_sfixed_a(-0.8854100704193115)),(to_sfixed_a(-0.3472919464111328)),(to_sfixed_a(0.19373413920402527)),(to_sfixed_a(-0.08160882443189621)),(to_sfixed_a(0.006443879567086697)),(to_sfixed_a(0.10761118680238724)),(to_sfixed_a(0.1477985978126526)),(to_sfixed_a(0.03837200626730919)),(to_sfixed_a(-0.16545382142066956)),(to_sfixed_a(-0.119339719414711)),(to_sfixed_a(-0.19278641045093536)),(to_sfixed_a(-0.03764863684773445)),(to_sfixed_a(-0.04149581491947174)),(to_sfixed_a(-0.010692600160837173)),(to_sfixed_a(-0.00016982572560664266)),(to_sfixed_a(5.531066926778294e-05)),(to_sfixed_a(-5.5319596867775545e-05)),(to_sfixed_a(-0.00019888364477083087)),(to_sfixed_a(-7.789121445966884e-05)),(to_sfixed_a(1.9110364064545138e-06)),(to_sfixed_a(-0.1516575813293457)),(to_sfixed_a(-0.006032863166183233)),(to_sfixed_a(-0.2243906706571579)),(to_sfixed_a(-0.08093797415494919)),(to_sfixed_a(-0.4663037359714508)),(to_sfixed_a(-0.7248508930206299)),(to_sfixed_a(-0.8863752484321594)),(to_sfixed_a(-1.4572337865829468)),(to_sfixed_a(-1.137730360031128)),(to_sfixed_a(-0.2860887050628662)),(to_sfixed_a(-0.09264332056045532)),(to_sfixed_a(-0.17077238857746124)),(to_sfixed_a(0.023474276065826416)),(to_sfixed_a(0.06690755486488342)),(to_sfixed_a(-0.1074916273355484)),(to_sfixed_a(-0.1450517177581787)),(to_sfixed_a(-0.05052606388926506)),(to_sfixed_a(-0.03110494837164879)),(to_sfixed_a(-0.12183002382516861)),(to_sfixed_a(0.08059629052877426)),(to_sfixed_a(0.0022991937585175037)),(to_sfixed_a(-2.972048423544038e-05)),(to_sfixed_a(0.000147135928273201)),(to_sfixed_a(-1.4725319488206878e-05)),(to_sfixed_a(-1.995954880840145e-05)),(to_sfixed_a(-0.00025154746253974736)),(to_sfixed_a(-5.4544150771107525e-05)),(to_sfixed_a(-0.00016461446648463607)),(to_sfixed_a(0.00021302493405528367)),(to_sfixed_a(0.004434528294950724)),(to_sfixed_a(-0.06713977456092834)),(to_sfixed_a(0.018314452841877937)),(to_sfixed_a(-0.1638225018978119)),(to_sfixed_a(-0.38637179136276245)),(to_sfixed_a(-0.4070630669593811)),(to_sfixed_a(-0.15139715373516083)),(to_sfixed_a(-0.2987625300884247)),(to_sfixed_a(-0.24323756992816925)),(to_sfixed_a(0.09900982677936554)),(to_sfixed_a(-0.06776696443557739)),(to_sfixed_a(-0.08988314867019653)),(to_sfixed_a(-0.002392314374446869)),(to_sfixed_a(-0.06786487251520157)),(to_sfixed_a(0.11187281459569931)),(to_sfixed_a(-0.1903800666332245)),(to_sfixed_a(0.01735824905335903)),(to_sfixed_a(-0.14886565506458282)),(to_sfixed_a(0.028100036084651947)),(to_sfixed_a(0.0980968177318573)),(to_sfixed_a(0.05255606025457382)),(to_sfixed_a(-0.00025667191948741674)),(to_sfixed_a(0.00016693315410520881)),(to_sfixed_a(0.000226773860049434)),(to_sfixed_a(-0.0002832460158970207)),(to_sfixed_a(-0.0002512593928258866)),(to_sfixed_a(-2.364053443670855e-06)),(to_sfixed_a(8.018263906706125e-05)),(to_sfixed_a(-0.05757063254714012)),(to_sfixed_a(-0.0016995148034766316)),(to_sfixed_a(0.02244945988059044)),(to_sfixed_a(0.07496398687362671)),(to_sfixed_a(-0.23982706665992737)),(to_sfixed_a(-0.06793437153100967)),(to_sfixed_a(0.015533971600234509)),(to_sfixed_a(-0.012335703708231449)),(to_sfixed_a(-0.028682243078947067)),(to_sfixed_a(0.10628696531057358)),(to_sfixed_a(-0.0977889820933342)),(to_sfixed_a(0.07455267757177353)),(to_sfixed_a(-0.11840316653251648)),(to_sfixed_a(-0.09540949761867523)),(to_sfixed_a(0.07824186980724335)),(to_sfixed_a(-0.11120783537626266)),(to_sfixed_a(-0.10433313995599747)),(to_sfixed_a(-0.012709875591099262)),(to_sfixed_a(-0.0030977828428149223)),(to_sfixed_a(0.00021405558800324798)),(to_sfixed_a(0.006016483996063471)),(to_sfixed_a(9.463598689762875e-05)),(to_sfixed_a(0.00010261157876811922)),(to_sfixed_a(-7.006406667642295e-05)),(to_sfixed_a(0.0002101458521792665)),(to_sfixed_a(7.169522723415866e-05)),(to_sfixed_a(9.962506010197103e-05)),(to_sfixed_a(4.916903344565071e-05)),(to_sfixed_a(-0.00023495634377468377)),(to_sfixed_a(-0.06731029599905014)),(to_sfixed_a(-0.05929267406463623)),(to_sfixed_a(0.26889848709106445)),(to_sfixed_a(0.08742775768041611)),(to_sfixed_a(0.06097831949591637)),(to_sfixed_a(0.29942744970321655)),(to_sfixed_a(0.17048002779483795)),(to_sfixed_a(0.17461946606636047)),(to_sfixed_a(0.008656680583953857)),(to_sfixed_a(-0.0026094454806298018)),(to_sfixed_a(0.017354050651192665)),(to_sfixed_a(0.04584120586514473)),(to_sfixed_a(0.02488938346505165)),(to_sfixed_a(-0.19161321222782135)),(to_sfixed_a(0.03147251158952713)),(to_sfixed_a(-0.040665097534656525)),(to_sfixed_a(0.00982305034995079)),(to_sfixed_a(0.036931782960891724)),(to_sfixed_a(0.003814003197476268)),(to_sfixed_a(-2.5938975340977777e-06)),(to_sfixed_a(-7.979360088938847e-05)),(to_sfixed_a(7.249398913700134e-05)),(to_sfixed_a(0.00015894304669927806)),(to_sfixed_a(-0.0001375274732708931)),(to_sfixed_a(-3.51783492078539e-05)),(to_sfixed_a(0.0002271628036396578)),(to_sfixed_a(-0.00015005766181275249)),(to_sfixed_a(-0.0002216300490545109)),(to_sfixed_a(0.012102142907679081)),(to_sfixed_a(-0.022706257179379463)),(to_sfixed_a(0.07753495126962662)),(to_sfixed_a(0.038869716227054596)),(to_sfixed_a(0.0025414605624973774)),(to_sfixed_a(0.12585894763469696)),(to_sfixed_a(0.32070761919021606)),(to_sfixed_a(0.1121821403503418)),(to_sfixed_a(0.07074615359306335)),(to_sfixed_a(0.06059498339891434)),(to_sfixed_a(0.054268937557935715)),(to_sfixed_a(-0.07954640686511993)),(to_sfixed_a(-0.00650236289948225)),(to_sfixed_a(-0.18346145749092102)),(to_sfixed_a(-0.052729032933712006)),(to_sfixed_a(0.03610476851463318)),(to_sfixed_a(0.014195425435900688)),(to_sfixed_a(-0.0028494028374552727)),(to_sfixed_a(0.01951550878584385)),(to_sfixed_a(3.773831849684939e-05)),(to_sfixed_a(-4.324253950471757e-06)),(to_sfixed_a(6.086572102503851e-05)),(to_sfixed_a(0.00012094784324290231)),(to_sfixed_a(-2.3429196517099626e-05)),(to_sfixed_a(-0.00012264765973668545)),(to_sfixed_a(-0.00017427615239284933)),(to_sfixed_a(3.326096339151263e-05)),(to_sfixed_a(0.0077290041372179985)),(to_sfixed_a(-0.0050391932018101215)),(to_sfixed_a(0.0334060899913311)),(to_sfixed_a(0.3733423352241516)),(to_sfixed_a(0.3856814205646515)),(to_sfixed_a(0.2742951810359955)),(to_sfixed_a(0.1811385452747345)),(to_sfixed_a(0.05012256279587746)),(to_sfixed_a(0.09695800393819809)),(to_sfixed_a(0.024384373798966408)),(to_sfixed_a(0.12637114524841309)),(to_sfixed_a(-0.03763369843363762)),(to_sfixed_a(-0.15309745073318481)),(to_sfixed_a(-0.16887648403644562)),(to_sfixed_a(-0.05216968432068825)),(to_sfixed_a(0.006477156188338995)),(to_sfixed_a(-0.012431347742676735)),(to_sfixed_a(0.014160530641674995)),(to_sfixed_a(-0.003979541826993227)),(to_sfixed_a(-0.009529425762593746)),(to_sfixed_a(4.948767673340626e-05)),(to_sfixed_a(-0.000113427457108628)),(to_sfixed_a(7.70124916016357e-06)),(to_sfixed_a(-4.6311135520227253e-05)),(to_sfixed_a(0.00011210061347810552)),(to_sfixed_a(-0.00019227767188567668)),(to_sfixed_a(-0.00026339179021306336)),(to_sfixed_a(-0.000122235287562944)),(to_sfixed_a(-5.5100452300393954e-05)),(to_sfixed_a(0.02761063352227211)),(to_sfixed_a(0.019120773300528526)),(to_sfixed_a(0.008399982005357742)),(to_sfixed_a(0.06440547853708267)),(to_sfixed_a(0.04567387327551842)),(to_sfixed_a(0.1623685359954834)),(to_sfixed_a(-0.017623988911509514)),(to_sfixed_a(0.08512821048498154)),(to_sfixed_a(0.18154874444007874)),(to_sfixed_a(-0.003970075864344835)),(to_sfixed_a(-0.007344857789576054)),(to_sfixed_a(-0.09764513373374939)),(to_sfixed_a(-0.12581099569797516)),(to_sfixed_a(-0.00662554707378149)),(to_sfixed_a(-0.020727060735225677)),(to_sfixed_a(0.031363893300294876)),(to_sfixed_a(0.0004945399123243988)),(to_sfixed_a(0.0023943877313286066)),(to_sfixed_a(0.002347046509385109)),(to_sfixed_a(-0.00024174746067728847)),(to_sfixed_a(-9.584476356394589e-05)),(to_sfixed_a(-8.591649384470657e-05)),(to_sfixed_a(6.26443579676561e-05)),(to_sfixed_a(-0.00011283392086625099)),(to_sfixed_a(5.159827196621336e-05)),(to_sfixed_a(-2.1446170649142005e-05)),(to_sfixed_a(-0.0001398580352542922)),(to_sfixed_a(0.00014364701928570867)),(to_sfixed_a(-0.0012618079781532288)),(to_sfixed_a(-0.0010925240349024534)),(to_sfixed_a(0.00019187614088878036)),(to_sfixed_a(-8.03780130809173e-05)),(to_sfixed_a(0.00043829105561599135)),(to_sfixed_a(-0.027434056624770164)),(to_sfixed_a(-0.010929299518465996)),(to_sfixed_a(-0.00253581372089684)),(to_sfixed_a(-0.009148716926574707)),(to_sfixed_a(0.005851246416568756)),(to_sfixed_a(0.002665646141394973)),(to_sfixed_a(-0.00045704221702180803)),(to_sfixed_a(-0.015136979520320892)),(to_sfixed_a(-0.02110309526324272)),(to_sfixed_a(-0.0021100842859596014)),(to_sfixed_a(0.001147764502093196)),(to_sfixed_a(-0.00021157764422241598)),(to_sfixed_a(0.00014515366638079286)),(to_sfixed_a(-2.3911852622404695e-05)),(to_sfixed_a(4.949828507960774e-05)),(to_sfixed_a(5.3200270485831425e-05)),(to_sfixed_a(-1.2286249329918064e-05)),(to_sfixed_a(-0.0001999529340537265)),(to_sfixed_a(7.644020661246032e-05)),(to_sfixed_a(0.00018650785204954445)),(to_sfixed_a(-7.814873242750764e-05)),(to_sfixed_a(-4.9544411012902856e-05)),(to_sfixed_a(-7.978237408678979e-05)),(to_sfixed_a(6.762168050045148e-05)),(to_sfixed_a(0.0002771077852230519)),(to_sfixed_a(-0.00023781364143360406)),(to_sfixed_a(0.00020175687677692622)),(to_sfixed_a(5.51532612007577e-05)),(to_sfixed_a(-0.00019363328465260565)),(to_sfixed_a(2.1814401407027617e-05)),(to_sfixed_a(0.0001990980963455513)),(to_sfixed_a(-0.00022675780928693712)),(to_sfixed_a(0.00022376186097972095)),(to_sfixed_a(-8.020465611480176e-05)),(to_sfixed_a(8.151445217663422e-05)),(to_sfixed_a(4.962304956279695e-05)),(to_sfixed_a(3.898028353432892e-06)),(to_sfixed_a(4.2623378249118105e-05)),(to_sfixed_a(7.589693268528208e-05)),(to_sfixed_a(0.00030188242089934647)),(to_sfixed_a(-0.0001782383187673986)),(to_sfixed_a(0.0002671059046406299)),(to_sfixed_a(0.0002708226384129375)),(to_sfixed_a(-8.35738392197527e-05)),(to_sfixed_a(-0.00019242826965637505)),(to_sfixed_a(0.00017012552416417748)));

    constant weight_n0_3 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-0.00047038125921972096)),(to_sfixed_a(0.000456570356618613)),(to_sfixed_a(0.0002886892470996827)),(to_sfixed_a(-0.00010144486441276968)),(to_sfixed_a(-6.458765710704029e-05)),(to_sfixed_a(0.00010707275214372203)),(to_sfixed_a(-0.00015372117923106998)),(to_sfixed_a(-0.0003010535438079387)),(to_sfixed_a(-1.4452093637373764e-05)),(to_sfixed_a(-4.805752541869879e-05)),(to_sfixed_a(0.00012803431309293956)),(to_sfixed_a(-2.805524127325043e-05)),(to_sfixed_a(-9.764605783857405e-05)),(to_sfixed_a(-8.413878094870597e-05)),(to_sfixed_a(3.646447657956742e-05)),(to_sfixed_a(4.7459880079259165e-06)),(to_sfixed_a(-5.1317601901246235e-06)),(to_sfixed_a(9.5598996267654e-05)),(to_sfixed_a(-9.900581790134311e-05)),(to_sfixed_a(7.714274397585541e-05)),(to_sfixed_a(2.9812932552886195e-05)),(to_sfixed_a(0.00010994397598551586)),(to_sfixed_a(-1.3148601283319294e-05)),(to_sfixed_a(-0.00031155580654740334)),(to_sfixed_a(9.899849828798324e-06)),(to_sfixed_a(6.736734212609008e-05)),(to_sfixed_a(7.538869249401614e-05)),(to_sfixed_a(-0.00020769439288415015)),(to_sfixed_a(-2.005117858061567e-05)),(to_sfixed_a(0.00010865114018088207)),(to_sfixed_a(-7.329590152949095e-05)),(to_sfixed_a(0.0001919525529956445)),(to_sfixed_a(-8.083087595878169e-05)),(to_sfixed_a(9.512215910945088e-05)),(to_sfixed_a(2.5228206141036935e-05)),(to_sfixed_a(-0.00012830100604332983)),(to_sfixed_a(3.744774221559055e-05)),(to_sfixed_a(0.0002726102829910815)),(to_sfixed_a(7.237195677589625e-05)),(to_sfixed_a(0.00020860660879407078)),(to_sfixed_a(0.00021031302458141)),(to_sfixed_a(0.00020762898202519864)),(to_sfixed_a(0.0001757530408212915)),(to_sfixed_a(0.00011353824811521918)),(to_sfixed_a(0.0001365194475511089)),(to_sfixed_a(-0.00010273489897372201)),(to_sfixed_a(4.828813416679623e-06)),(to_sfixed_a(-0.00036840885877609253)),(to_sfixed_a(0.000534767925273627)),(to_sfixed_a(0.00022493276628665626)),(to_sfixed_a(-3.073348489124328e-05)),(to_sfixed_a(-0.00020949615282006562)),(to_sfixed_a(0.00018829536566045135)),(to_sfixed_a(-2.1957150238449685e-05)),(to_sfixed_a(-1.9988832718809135e-05)),(to_sfixed_a(-0.0002909466275013983)),(to_sfixed_a(-0.0003486363566480577)),(to_sfixed_a(0.00011382682714611292)),(to_sfixed_a(-0.00011453435581643134)),(to_sfixed_a(3.08569215121679e-05)),(to_sfixed_a(-3.572385321604088e-05)),(to_sfixed_a(4.434470974956639e-05)),(to_sfixed_a(-0.00016542307275813073)),(to_sfixed_a(0.000260679516941309)),(to_sfixed_a(-4.7791461838642135e-05)),(to_sfixed_a(-1.2075096492480952e-05)),(to_sfixed_a(-6.359891267493367e-05)),(to_sfixed_a(-1.848653846536763e-05)),(to_sfixed_a(-9.020455036079511e-05)),(to_sfixed_a(0.04475191608071327)),(to_sfixed_a(-3.987245145253837e-05)),(to_sfixed_a(1.0051922799902968e-05)),(to_sfixed_a(3.8818910979898646e-05)),(to_sfixed_a(-4.515548062045127e-05)),(to_sfixed_a(-0.0002601671149022877)),(to_sfixed_a(-0.00010633528290782124)),(to_sfixed_a(0.00012772483751177788)),(to_sfixed_a(9.227855480276048e-05)),(to_sfixed_a(4.1107836295850575e-05)),(to_sfixed_a(-0.00012180378689663485)),(to_sfixed_a(-4.603197885444388e-05)),(to_sfixed_a(7.456395542249084e-05)),(to_sfixed_a(2.8650491003645584e-05)),(to_sfixed_a(0.00010219793330179527)),(to_sfixed_a(-4.046282629133202e-05)),(to_sfixed_a(-2.99259463645285e-05)),(to_sfixed_a(-3.1155606848187745e-05)),(to_sfixed_a(0.0003503420448396355)),(to_sfixed_a(-2.5866945634334115e-06)),(to_sfixed_a(0.0001195675868075341)),(to_sfixed_a(-3.6643083149101585e-05)),(to_sfixed_a(-0.00023473285546060652)),(to_sfixed_a(0.06669211387634277)),(to_sfixed_a(7.409330282825977e-05)),(to_sfixed_a(0.07562926411628723)),(to_sfixed_a(-0.0544351190328598)),(to_sfixed_a(0.03143167495727539)),(to_sfixed_a(0.031501900404691696)),(to_sfixed_a(0.1130475252866745)),(to_sfixed_a(0.003349264618009329)),(to_sfixed_a(0.01438422966748476)),(to_sfixed_a(0.008946661837399006)),(to_sfixed_a(-0.21513858437538147)),(to_sfixed_a(0.12181991338729858)),(to_sfixed_a(0.018398547545075417)),(to_sfixed_a(0.03713665157556534)),(to_sfixed_a(8.1614576629363e-05)),(to_sfixed_a(9.160445188172162e-05)),(to_sfixed_a(0.00016118277562782168)),(to_sfixed_a(0.00015632351278327405)),(to_sfixed_a(-5.089083788334392e-05)),(to_sfixed_a(0.0001960258960025385)),(to_sfixed_a(-0.0002870687167160213)),(to_sfixed_a(8.507669008395169e-06)),(to_sfixed_a(-5.6933247833512723e-05)),(to_sfixed_a(-5.328109909896739e-05)),(to_sfixed_a(-0.00042537457193247974)),(to_sfixed_a(0.00017134888912551105)),(to_sfixed_a(-0.0003491994284559041)),(to_sfixed_a(-0.0016329552745446563)),(to_sfixed_a(0.05982019752264023)),(to_sfixed_a(0.09057814627885818)),(to_sfixed_a(-0.002355963923037052)),(to_sfixed_a(0.06979431957006454)),(to_sfixed_a(-0.0957731232047081)),(to_sfixed_a(-0.10555271059274673)),(to_sfixed_a(0.004874106030911207)),(to_sfixed_a(0.17840440571308136)),(to_sfixed_a(0.050197534263134)),(to_sfixed_a(0.05765928700566292)),(to_sfixed_a(-0.1035868301987648)),(to_sfixed_a(-0.09884300827980042)),(to_sfixed_a(-0.0022759244311600924)),(to_sfixed_a(0.04336882755160332)),(to_sfixed_a(0.029793981462717056)),(to_sfixed_a(-0.0005323665682226419)),(to_sfixed_a(0.001424369402229786)),(to_sfixed_a(0.00017072887567337602)),(to_sfixed_a(-0.0002497037930879742)),(to_sfixed_a(3.33863208652474e-05)),(to_sfixed_a(-0.0002077420795103535)),(to_sfixed_a(3.416087929508649e-05)),(to_sfixed_a(-8.730874833418056e-05)),(to_sfixed_a(0.00014109237235970795)),(to_sfixed_a(0.0018855552189052105)),(to_sfixed_a(0.013842187821865082)),(to_sfixed_a(0.015772150829434395)),(to_sfixed_a(0.12284009903669357)),(to_sfixed_a(-0.06437412649393082)),(to_sfixed_a(-0.035673465579748154)),(to_sfixed_a(0.014695750549435616)),(to_sfixed_a(-0.13270513713359833)),(to_sfixed_a(-0.09011121094226837)),(to_sfixed_a(0.1119374930858612)),(to_sfixed_a(0.019684243947267532)),(to_sfixed_a(0.14813776314258575)),(to_sfixed_a(-0.10968780517578125)),(to_sfixed_a(0.019374437630176544)),(to_sfixed_a(-0.17741765081882477)),(to_sfixed_a(-0.06674610823392868)),(to_sfixed_a(-0.05892971530556679)),(to_sfixed_a(-0.12970897555351257)),(to_sfixed_a(0.0007847927627153695)),(to_sfixed_a(0.057824622839689255)),(to_sfixed_a(0.0034320824779570103)),(to_sfixed_a(-7.649302278878167e-05)),(to_sfixed_a(-2.5046083464985713e-05)),(to_sfixed_a(4.9034447329177056e-06)),(to_sfixed_a(-2.3446576960850507e-05)),(to_sfixed_a(0.00013336013944353908)),(to_sfixed_a(-1.453360528103076e-05)),(to_sfixed_a(3.182346699759364e-05)),(to_sfixed_a(0.0002188866783399135)),(to_sfixed_a(0.010876033455133438)),(to_sfixed_a(0.01807115226984024)),(to_sfixed_a(-0.009453129023313522)),(to_sfixed_a(-0.06718812137842178)),(to_sfixed_a(-0.08161433041095734)),(to_sfixed_a(-0.3520870804786682)),(to_sfixed_a(-0.18941278755664825)),(to_sfixed_a(-0.2455061972141266)),(to_sfixed_a(-0.0649825781583786)),(to_sfixed_a(-0.12641099095344543)),(to_sfixed_a(-0.0717037171125412)),(to_sfixed_a(-0.0423603318631649)),(to_sfixed_a(-0.12971363961696625)),(to_sfixed_a(-0.0847514197230339)),(to_sfixed_a(-0.23994535207748413)),(to_sfixed_a(-0.2645759880542755)),(to_sfixed_a(-0.28336507081985474)),(to_sfixed_a(-0.0841335877776146)),(to_sfixed_a(-0.02044745348393917)),(to_sfixed_a(0.006032091565430164)),(to_sfixed_a(0.007404313888400793)),(to_sfixed_a(0.0028100418858230114)),(to_sfixed_a(0.00021755533816758543)),(to_sfixed_a(0.00010718061093939468)),(to_sfixed_a(-7.394022395601496e-05)),(to_sfixed_a(-0.00016064097872003913)),(to_sfixed_a(-1.9968359993072227e-05)),(to_sfixed_a(-0.0001855394075391814)),(to_sfixed_a(-0.026794586330652237)),(to_sfixed_a(0.058309100568294525)),(to_sfixed_a(0.028908690437674522)),(to_sfixed_a(-0.09364311397075653)),(to_sfixed_a(-0.12036523967981339)),(to_sfixed_a(-0.476841002702713)),(to_sfixed_a(-0.24959522485733032)),(to_sfixed_a(-0.26326024532318115)),(to_sfixed_a(-0.4696711599826813)),(to_sfixed_a(-0.14766128361225128)),(to_sfixed_a(-0.24518005549907684)),(to_sfixed_a(0.07365927845239639)),(to_sfixed_a(-0.12206661701202393)),(to_sfixed_a(-0.24565017223358154)),(to_sfixed_a(-0.6684373021125793)),(to_sfixed_a(-0.43355438113212585)),(to_sfixed_a(-0.3644111454486847)),(to_sfixed_a(-0.09465258568525314)),(to_sfixed_a(-0.3372337818145752)),(to_sfixed_a(0.022931409999728203)),(to_sfixed_a(-0.004108642227947712)),(to_sfixed_a(4.6460227167699486e-05)),(to_sfixed_a(3.742316403076984e-05)),(to_sfixed_a(-0.0001810725370887667)),(to_sfixed_a(-3.303991979919374e-05)),(to_sfixed_a(-1.5022785191831645e-05)),(to_sfixed_a(7.907221151981503e-05)),(to_sfixed_a(0.049196891486644745)),(to_sfixed_a(-0.0033694826997816563)),(to_sfixed_a(0.008712566457688808)),(to_sfixed_a(-0.22725805640220642)),(to_sfixed_a(-0.1294662058353424)),(to_sfixed_a(-0.2129485160112381)),(to_sfixed_a(-0.1374877691268921)),(to_sfixed_a(-0.23048008978366852)),(to_sfixed_a(-0.19227582216262817)),(to_sfixed_a(-0.287274569272995)),(to_sfixed_a(-0.05061723664402962)),(to_sfixed_a(-0.30627578496932983)),(to_sfixed_a(-0.3508332669734955)),(to_sfixed_a(-0.5539825558662415)),(to_sfixed_a(-0.714851438999176)),(to_sfixed_a(-0.44618961215019226)),(to_sfixed_a(-0.3216479420661926)),(to_sfixed_a(-0.07394609600305557)),(to_sfixed_a(-0.44528234004974365)),(to_sfixed_a(-0.19933359324932098)),(to_sfixed_a(-0.09793626517057419)),(to_sfixed_a(-0.018296170979738235)),(to_sfixed_a(-4.67460222353111e-06)),(to_sfixed_a(-1.2720194717985578e-05)),(to_sfixed_a(0.00020049541490152478)),(to_sfixed_a(5.280677942209877e-05)),(to_sfixed_a(1.369138317386387e-05)),(to_sfixed_a(-0.0002364930260227993)),(to_sfixed_a(0.0003404368762858212)),(to_sfixed_a(0.06470324844121933)),(to_sfixed_a(-0.06661653518676758)),(to_sfixed_a(-0.03480851277709007)),(to_sfixed_a(-0.07622507959604263)),(to_sfixed_a(-0.04271840304136276)),(to_sfixed_a(-0.16384774446487427)),(to_sfixed_a(-0.05112534761428833)),(to_sfixed_a(-0.028840893879532814)),(to_sfixed_a(-0.021884111687541008)),(to_sfixed_a(-0.0060133980587124825)),(to_sfixed_a(-0.12894919514656067)),(to_sfixed_a(-0.585265040397644)),(to_sfixed_a(-0.5414776802062988)),(to_sfixed_a(-0.4998356103897095)),(to_sfixed_a(-0.591149091720581)),(to_sfixed_a(-0.3555888235569)),(to_sfixed_a(-0.2659251391887665)),(to_sfixed_a(-0.23378242552280426)),(to_sfixed_a(-0.016974681988358498)),(to_sfixed_a(-0.10351002961397171)),(to_sfixed_a(1.712291305011604e-05)),(to_sfixed_a(6.0599588323384523e-05)),(to_sfixed_a(5.558563498198055e-05)),(to_sfixed_a(-0.00011850317969219759)),(to_sfixed_a(0.0002005762653425336)),(to_sfixed_a(-0.00015349537716247141)),(to_sfixed_a(0.0003711808822117746)),(to_sfixed_a(-0.004345930181443691)),(to_sfixed_a(-0.006671068724244833)),(to_sfixed_a(0.09322851896286011)),(to_sfixed_a(-0.00219640857540071)),(to_sfixed_a(-0.038335170596838)),(to_sfixed_a(0.050477899610996246)),(to_sfixed_a(-0.09104088693857193)),(to_sfixed_a(0.35483652353286743)),(to_sfixed_a(0.09934277832508087)),(to_sfixed_a(0.7114606499671936)),(to_sfixed_a(0.7984837889671326)),(to_sfixed_a(0.29117605090141296)),(to_sfixed_a(-0.03259938210248947)),(to_sfixed_a(-0.028997281566262245)),(to_sfixed_a(-0.2313365936279297)),(to_sfixed_a(-0.1482093781232834)),(to_sfixed_a(-0.04651299864053726)),(to_sfixed_a(-0.08850077539682388)),(to_sfixed_a(0.17211832106113434)),(to_sfixed_a(-0.15085430443286896)),(to_sfixed_a(-0.014002185314893723)),(to_sfixed_a(-0.014449363574385643)),(to_sfixed_a(-8.76274352776818e-05)),(to_sfixed_a(-0.0001818762393668294)),(to_sfixed_a(0.00035376628511585295)),(to_sfixed_a(2.082045830320567e-05)),(to_sfixed_a(-1.5978315786924213e-05)),(to_sfixed_a(0.008145100437104702)),(to_sfixed_a(0.17028430104255676)),(to_sfixed_a(0.2191743701696396)),(to_sfixed_a(0.036928314715623856)),(to_sfixed_a(0.22605153918266296)),(to_sfixed_a(0.1782340556383133)),(to_sfixed_a(0.2942701280117035)),(to_sfixed_a(0.35646435618400574)),(to_sfixed_a(0.5627197027206421)),(to_sfixed_a(0.7857637405395508)),(to_sfixed_a(0.6899304389953613)),(to_sfixed_a(0.3890565037727356)),(to_sfixed_a(0.16848969459533691)),(to_sfixed_a(0.1313125044107437)),(to_sfixed_a(0.20929813385009766)),(to_sfixed_a(0.21315135061740875)),(to_sfixed_a(0.2800613045692444)),(to_sfixed_a(0.31983163952827454)),(to_sfixed_a(0.10919013619422913)),(to_sfixed_a(0.07560615241527557)),(to_sfixed_a(-0.1531175673007965)),(to_sfixed_a(-0.03848070278763771)),(to_sfixed_a(2.346702558497782e-06)),(to_sfixed_a(3.455347177805379e-05)),(to_sfixed_a(8.036835060920566e-05)),(to_sfixed_a(3.3766409615054727e-05)),(to_sfixed_a(6.274801125982776e-05)),(to_sfixed_a(-1.5552150216535665e-05)),(to_sfixed_a(-3.984935028711334e-05)),(to_sfixed_a(0.09933222085237503)),(to_sfixed_a(0.12648409605026245)),(to_sfixed_a(0.15683752298355103)),(to_sfixed_a(0.3518942892551422)),(to_sfixed_a(0.5132710337638855)),(to_sfixed_a(0.5539117455482483)),(to_sfixed_a(0.3854782283306122)),(to_sfixed_a(0.6330752968788147)),(to_sfixed_a(0.23103827238082886)),(to_sfixed_a(0.14341439306735992)),(to_sfixed_a(0.15769974887371063)),(to_sfixed_a(0.17428624629974365)),(to_sfixed_a(0.13109393417835236)),(to_sfixed_a(0.1807524710893631)),(to_sfixed_a(0.15916316211223602)),(to_sfixed_a(0.5476757884025574)),(to_sfixed_a(0.47648337483406067)),(to_sfixed_a(0.15563321113586426)),(to_sfixed_a(0.05299399420619011)),(to_sfixed_a(-0.21756485104560852)),(to_sfixed_a(0.02816510945558548)),(to_sfixed_a(0.00015074289694894105)),(to_sfixed_a(0.0004924439126625657)),(to_sfixed_a(-5.788338967249729e-05)),(to_sfixed_a(0.00022875801369082183)),(to_sfixed_a(-3.712287434609607e-05)),(to_sfixed_a(5.292299101711251e-05)),(to_sfixed_a(-5.9343179600546136e-05)),(to_sfixed_a(-0.023116547614336014)),(to_sfixed_a(0.3609989881515503)),(to_sfixed_a(0.236455500125885)),(to_sfixed_a(0.36350786685943604)),(to_sfixed_a(0.24764253199100494)),(to_sfixed_a(0.22712787985801697)),(to_sfixed_a(0.2628035247325897)),(to_sfixed_a(0.38540711998939514)),(to_sfixed_a(0.13871249556541443)),(to_sfixed_a(-0.11616013944149017)),(to_sfixed_a(-0.0591459684073925)),(to_sfixed_a(-0.01578269526362419)),(to_sfixed_a(0.2396164834499359)),(to_sfixed_a(0.10479182004928589)),(to_sfixed_a(0.18093328177928925)),(to_sfixed_a(0.2265351563692093)),(to_sfixed_a(0.3160912096500397)),(to_sfixed_a(0.04362925514578819)),(to_sfixed_a(-0.06448567658662796)),(to_sfixed_a(0.18676608800888062)),(to_sfixed_a(0.08812405169010162)),(to_sfixed_a(0.002805558033287525)),(to_sfixed_a(0.0042111254297196865)),(to_sfixed_a(8.135782991303131e-05)),(to_sfixed_a(0.0002022746339207515)),(to_sfixed_a(-0.0001998182269744575)),(to_sfixed_a(-0.00031751260394230485)),(to_sfixed_a(8.676861762069166e-05)),(to_sfixed_a(0.0016215642681345344)),(to_sfixed_a(0.20407922565937042)),(to_sfixed_a(0.16564218699932098)),(to_sfixed_a(-0.13439905643463135)),(to_sfixed_a(0.1270667314529419)),(to_sfixed_a(-0.11102218925952911)),(to_sfixed_a(0.2801143229007721)),(to_sfixed_a(-0.15339647233486176)),(to_sfixed_a(0.052739713340997696)),(to_sfixed_a(-0.08853216469287872)),(to_sfixed_a(-0.09292677789926529)),(to_sfixed_a(0.09866614639759064)),(to_sfixed_a(0.05804640054702759)),(to_sfixed_a(0.1792934387922287)),(to_sfixed_a(0.3328661024570465)),(to_sfixed_a(0.11521166563034058)),(to_sfixed_a(-0.021175451576709747)),(to_sfixed_a(0.15104955434799194)),(to_sfixed_a(0.12757404148578644)),(to_sfixed_a(0.13531889021396637)),(to_sfixed_a(0.040009185671806335)),(to_sfixed_a(-0.0002527447941247374)),(to_sfixed_a(1.837455783970654e-05)),(to_sfixed_a(8.264637290267274e-05)),(to_sfixed_a(9.160336048807949e-05)),(to_sfixed_a(-9.216742000717204e-06)),(to_sfixed_a(0.0004075336910318583)),(to_sfixed_a(0.0001526240521343425)),(to_sfixed_a(-0.0025308970361948013)),(to_sfixed_a(-0.03704330697655678)),(to_sfixed_a(-0.04215754568576813)),(to_sfixed_a(-0.08693671226501465)),(to_sfixed_a(0.1324441283941269)),(to_sfixed_a(-0.0376151017844677)),(to_sfixed_a(-0.03460836783051491)),(to_sfixed_a(0.1330481618642807)),(to_sfixed_a(0.1294083595275879)),(to_sfixed_a(0.16248847544193268)),(to_sfixed_a(0.15969403088092804)),(to_sfixed_a(0.16325883567333221)),(to_sfixed_a(0.18519198894500732)),(to_sfixed_a(0.31722983717918396)),(to_sfixed_a(0.10922367125749588)),(to_sfixed_a(0.15685443580150604)),(to_sfixed_a(0.1790885329246521)),(to_sfixed_a(0.06932659447193146)),(to_sfixed_a(-0.014193644747138023)),(to_sfixed_a(0.060209836810827255)),(to_sfixed_a(0.174446702003479)),(to_sfixed_a(0.00014014384942129254)),(to_sfixed_a(0.00010056450992124155)),(to_sfixed_a(0.0002563262823969126)),(to_sfixed_a(8.312018326250836e-05)),(to_sfixed_a(-0.00030413427157327533)),(to_sfixed_a(0.0003789174370467663)),(to_sfixed_a(-0.0006285619456321001)),(to_sfixed_a(0.011988927610218525)),(to_sfixed_a(-0.05380101501941681)),(to_sfixed_a(-0.35113248229026794)),(to_sfixed_a(-0.08878809958696365)),(to_sfixed_a(-0.09170141816139221)),(to_sfixed_a(-0.08807067573070526)),(to_sfixed_a(0.0452721081674099)),(to_sfixed_a(-0.08470042794942856)),(to_sfixed_a(-0.10932207852602005)),(to_sfixed_a(-0.09991197288036346)),(to_sfixed_a(0.16069553792476654)),(to_sfixed_a(0.3149528503417969)),(to_sfixed_a(0.29899147152900696)),(to_sfixed_a(0.31690627336502075)),(to_sfixed_a(0.14728602766990662)),(to_sfixed_a(-0.25800755620002747)),(to_sfixed_a(-0.0456952229142189)),(to_sfixed_a(0.11401760578155518)),(to_sfixed_a(-0.0324486643075943)),(to_sfixed_a(0.12424518167972565)),(to_sfixed_a(0.15701143443584442)),(to_sfixed_a(-0.008314905688166618)),(to_sfixed_a(-0.0002325113455299288)),(to_sfixed_a(-1.4282039956015069e-05)),(to_sfixed_a(0.0001124443078879267)),(to_sfixed_a(0.0001275520189665258)),(to_sfixed_a(-0.0001240330602740869)),(to_sfixed_a(-0.0006150074186734855)),(to_sfixed_a(0.024193933233618736)),(to_sfixed_a(-0.05278350040316582)),(to_sfixed_a(-0.22455395758152008)),(to_sfixed_a(-0.06275849789381027)),(to_sfixed_a(-0.059536412358284)),(to_sfixed_a(-0.20298567414283752)),(to_sfixed_a(-0.5248786807060242)),(to_sfixed_a(-0.5909352898597717)),(to_sfixed_a(-0.43630295991897583)),(to_sfixed_a(0.15237802267074585)),(to_sfixed_a(0.04626370221376419)),(to_sfixed_a(0.4806484282016754)),(to_sfixed_a(0.31044164299964905)),(to_sfixed_a(0.24695435166358948)),(to_sfixed_a(0.31064334511756897)),(to_sfixed_a(-0.04236193001270294)),(to_sfixed_a(-0.07019932568073273)),(to_sfixed_a(0.03246535733342171)),(to_sfixed_a(-0.05419417843222618)),(to_sfixed_a(-0.024977173656225204)),(to_sfixed_a(0.00021399669640231878)),(to_sfixed_a(-0.00030576749122701585)),(to_sfixed_a(-4.6689267037436366e-05)),(to_sfixed_a(-0.00030042926664464176)),(to_sfixed_a(0.0003390912024769932)),(to_sfixed_a(-0.00016295195382554084)),(to_sfixed_a(-3.8690508517902344e-05)),(to_sfixed_a(-0.017163172364234924)),(to_sfixed_a(0.13796789944171906)),(to_sfixed_a(-0.020485535264015198)),(to_sfixed_a(0.04183721914887428)),(to_sfixed_a(-0.26660799980163574)),(to_sfixed_a(-0.25004157423973083)),(to_sfixed_a(-0.375862181186676)),(to_sfixed_a(-0.41347917914390564)),(to_sfixed_a(-0.4264949858188629)),(to_sfixed_a(-0.49167853593826294)),(to_sfixed_a(0.12717781960964203)),(to_sfixed_a(0.475713849067688)),(to_sfixed_a(0.4493933320045471)),(to_sfixed_a(0.49235132336616516)),(to_sfixed_a(0.11437491327524185)),(to_sfixed_a(-0.01864646188914776)),(to_sfixed_a(-0.26966577768325806)),(to_sfixed_a(-0.040433987975120544)),(to_sfixed_a(-0.08425456285476685)),(to_sfixed_a(-0.005965373944491148)),(to_sfixed_a(0.05044352263212204)),(to_sfixed_a(-0.005353562068194151)),(to_sfixed_a(-8.852559403749183e-05)),(to_sfixed_a(0.00018377906235400587)),(to_sfixed_a(9.330758621217683e-05)),(to_sfixed_a(-0.00011253597040195018)),(to_sfixed_a(0.0001434840087313205)),(to_sfixed_a(-0.0003020661824848503)),(to_sfixed_a(0.009008606895804405)),(to_sfixed_a(-0.001257814816199243)),(to_sfixed_a(0.13818393647670746)),(to_sfixed_a(0.011682912707328796)),(to_sfixed_a(-0.09034302830696106)),(to_sfixed_a(-0.2728208899497986)),(to_sfixed_a(-0.20216451585292816)),(to_sfixed_a(-0.3294016718864441)),(to_sfixed_a(-0.34613415598869324)),(to_sfixed_a(-0.16418051719665527)),(to_sfixed_a(0.031027978286147118)),(to_sfixed_a(0.5203559994697571)),(to_sfixed_a(0.7409859895706177)),(to_sfixed_a(0.1518891155719757)),(to_sfixed_a(-0.036476749926805496)),(to_sfixed_a(-0.11012599617242813)),(to_sfixed_a(0.01779812015593052)),(to_sfixed_a(0.025519652292132378)),(to_sfixed_a(-0.06585822254419327)),(to_sfixed_a(-0.04605657979846001)),(to_sfixed_a(-0.011348078958690166)),(to_sfixed_a(-9.350349864689633e-05)),(to_sfixed_a(3.0293034797068685e-05)),(to_sfixed_a(0.0001493444142397493)),(to_sfixed_a(0.00031425507040694356)),(to_sfixed_a(4.17650408053305e-05)),(to_sfixed_a(9.689133003121242e-05)),(to_sfixed_a(-0.00015507084026467055)),(to_sfixed_a(-2.515415872039739e-05)),(to_sfixed_a(-0.009141919203102589)),(to_sfixed_a(0.045919269323349)),(to_sfixed_a(-0.31217458844184875)),(to_sfixed_a(-0.1856674700975418)),(to_sfixed_a(-0.06742294132709503)),(to_sfixed_a(-0.11849883943796158)),(to_sfixed_a(-0.15925854444503784)),(to_sfixed_a(0.001744202570989728)),(to_sfixed_a(-0.19559772312641144)),(to_sfixed_a(0.11033407598733902)),(to_sfixed_a(0.31240925192832947)),(to_sfixed_a(0.1293725073337555)),(to_sfixed_a(0.05789627879858017)),(to_sfixed_a(-0.0520051047205925)),(to_sfixed_a(-0.08068881183862686)),(to_sfixed_a(-0.011976132169365883)),(to_sfixed_a(0.006426139734685421)),(to_sfixed_a(0.1160479187965393)),(to_sfixed_a(0.08789781481027603)),(to_sfixed_a(-0.0811217799782753)),(to_sfixed_a(-0.18352645635604858)),(to_sfixed_a(0.00013092630251776427)),(to_sfixed_a(-9.323786071036011e-05)),(to_sfixed_a(-5.999305722070858e-05)),(to_sfixed_a(9.329211752628908e-05)),(to_sfixed_a(-0.00022871453256811947)),(to_sfixed_a(-0.00021819073299411684)),(to_sfixed_a(-8.593225356889889e-05)),(to_sfixed_a(-0.02109639160335064)),(to_sfixed_a(0.0006613050354644656)),(to_sfixed_a(0.08946914970874786)),(to_sfixed_a(-0.1422547698020935)),(to_sfixed_a(-0.15697650611400604)),(to_sfixed_a(-0.27899619936943054)),(to_sfixed_a(0.043643999844789505)),(to_sfixed_a(-0.03725932538509369)),(to_sfixed_a(0.040101561695337296)),(to_sfixed_a(-0.0819699615240097)),(to_sfixed_a(-0.2921290099620819)),(to_sfixed_a(-0.25715169310569763)),(to_sfixed_a(-0.08786174654960632)),(to_sfixed_a(-0.08726818114519119)),(to_sfixed_a(-0.0016560147050768137)),(to_sfixed_a(-0.1499534696340561)),(to_sfixed_a(-0.09504082053899765)),(to_sfixed_a(-0.02013908326625824)),(to_sfixed_a(-0.04128492996096611)),(to_sfixed_a(0.0007494311430491507)),(to_sfixed_a(0.0015138507587835193)),(to_sfixed_a(-0.00015084799088072032)),(to_sfixed_a(-0.00011101687414338812)),(to_sfixed_a(0.00022571189037989825)),(to_sfixed_a(1.602858719707001e-05)),(to_sfixed_a(-0.00025328612537123263)),(to_sfixed_a(-5.581010555033572e-05)),(to_sfixed_a(-0.00018558920419309288)),(to_sfixed_a(0.00011481817637104541)),(to_sfixed_a(-0.06006071716547012)),(to_sfixed_a(0.03451960161328316)),(to_sfixed_a(-0.11582870781421661)),(to_sfixed_a(-0.023005085065960884)),(to_sfixed_a(0.042033035308122635)),(to_sfixed_a(-0.13312271237373352)),(to_sfixed_a(0.08083092421293259)),(to_sfixed_a(-0.10255441069602966)),(to_sfixed_a(-0.16321395337581635)),(to_sfixed_a(-0.25981757044792175)),(to_sfixed_a(-0.1837257742881775)),(to_sfixed_a(-0.3958896994590759)),(to_sfixed_a(-0.2785471975803375)),(to_sfixed_a(-0.4238939583301544)),(to_sfixed_a(0.012718180194497108)),(to_sfixed_a(0.03561316058039665)),(to_sfixed_a(0.015504356473684311)),(to_sfixed_a(0.007950404658913612)),(to_sfixed_a(0.010154915042221546)),(to_sfixed_a(-6.721255340380594e-05)),(to_sfixed_a(8.039462409215048e-05)),(to_sfixed_a(0.00019922512001357973)),(to_sfixed_a(-0.00011699606693582609)),(to_sfixed_a(3.884183388436213e-05)),(to_sfixed_a(-9.968189988285303e-05)),(to_sfixed_a(0.00026350290863774717)),(to_sfixed_a(-0.00011456644278950989)),(to_sfixed_a(0.00030105505720712245)),(to_sfixed_a(-0.06019197404384613)),(to_sfixed_a(-0.05147837474942207)),(to_sfixed_a(-0.06339258700609207)),(to_sfixed_a(-0.16842813789844513)),(to_sfixed_a(0.0110018914565444)),(to_sfixed_a(0.04773196205496788)),(to_sfixed_a(-0.1294011026620865)),(to_sfixed_a(-0.11954689025878906)),(to_sfixed_a(-0.19854463636875153)),(to_sfixed_a(-0.17683693766593933)),(to_sfixed_a(-0.22597834467887878)),(to_sfixed_a(-0.3242974877357483)),(to_sfixed_a(-0.27542126178741455)),(to_sfixed_a(-0.22918067872524261)),(to_sfixed_a(0.1485200971364975)),(to_sfixed_a(-0.1119157075881958)),(to_sfixed_a(-0.004390973597764969)),(to_sfixed_a(0.005222694482654333)),(to_sfixed_a(-0.010764642618596554)),(to_sfixed_a(-9.400754061061889e-05)),(to_sfixed_a(0.00019888645329046994)),(to_sfixed_a(-3.8889753341209143e-05)),(to_sfixed_a(0.00023548118770122528)),(to_sfixed_a(0.00013355014380067587)),(to_sfixed_a(-0.0001856147573562339)),(to_sfixed_a(3.898708746419288e-05)),(to_sfixed_a(4.528364661382511e-05)),(to_sfixed_a(-0.0087739871814847)),(to_sfixed_a(-0.040925510227680206)),(to_sfixed_a(-0.03784802183508873)),(to_sfixed_a(-0.016519585624337196)),(to_sfixed_a(-0.01573696918785572)),(to_sfixed_a(-0.10006456822156906)),(to_sfixed_a(-0.12638331949710846)),(to_sfixed_a(0.029651738703250885)),(to_sfixed_a(-0.40473228693008423)),(to_sfixed_a(-0.41839542984962463)),(to_sfixed_a(-0.13956618309020996)),(to_sfixed_a(-0.1194157674908638)),(to_sfixed_a(-0.4322773814201355)),(to_sfixed_a(-0.06300903111696243)),(to_sfixed_a(0.07154732942581177)),(to_sfixed_a(-0.06231777369976044)),(to_sfixed_a(0.011319879442453384)),(to_sfixed_a(-0.020864155143499374)),(to_sfixed_a(-0.01153524313122034)),(to_sfixed_a(-0.011321269907057285)),(to_sfixed_a(0.00021754432236775756)),(to_sfixed_a(-7.35582725610584e-05)),(to_sfixed_a(-0.000188371108379215)),(to_sfixed_a(-0.00011511091724969447)),(to_sfixed_a(0.0001341936003882438)),(to_sfixed_a(-3.3572247048141435e-05)),(to_sfixed_a(-9.604050137568265e-05)),(to_sfixed_a(-6.212234438862652e-05)),(to_sfixed_a(-4.825551877729595e-05)),(to_sfixed_a(0.008818652480840683)),(to_sfixed_a(-0.022652091458439827)),(to_sfixed_a(-0.016707731410861015)),(to_sfixed_a(-0.1794336587190628)),(to_sfixed_a(-0.23008780181407928)),(to_sfixed_a(0.054832957684993744)),(to_sfixed_a(-0.027205608785152435)),(to_sfixed_a(-0.11889538913965225)),(to_sfixed_a(0.027108626440167427)),(to_sfixed_a(0.010467614978551865)),(to_sfixed_a(-0.09877119958400726)),(to_sfixed_a(-0.2366970032453537)),(to_sfixed_a(0.0029587061144411564)),(to_sfixed_a(-0.0022696317173540592)),(to_sfixed_a(-0.15320894122123718)),(to_sfixed_a(-0.02338729240000248)),(to_sfixed_a(0.0001505899999756366)),(to_sfixed_a(-0.0017683913465589285)),(to_sfixed_a(-0.002007395261898637)),(to_sfixed_a(-2.0718385712825693e-05)),(to_sfixed_a(0.00013950178981758654)),(to_sfixed_a(3.2167397876037285e-05)),(to_sfixed_a(-2.4820717953843996e-05)),(to_sfixed_a(-0.00019515701569616795)),(to_sfixed_a(-8.870320743881166e-05)),(to_sfixed_a(0.00020155051606707275)),(to_sfixed_a(-0.00010271209612255916)),(to_sfixed_a(6.891693192301318e-05)),(to_sfixed_a(0.002111306181177497)),(to_sfixed_a(0.0022422648034989834)),(to_sfixed_a(-3.943747287848964e-05)),(to_sfixed_a(-0.0002686037332750857)),(to_sfixed_a(-0.0002528050390537828)),(to_sfixed_a(-0.06244007498025894)),(to_sfixed_a(0.0011108259204775095)),(to_sfixed_a(0.00026344083016738296)),(to_sfixed_a(-0.04045188054442406)),(to_sfixed_a(0.024952035397291183)),(to_sfixed_a(0.0022766750771552324)),(to_sfixed_a(-0.03808616101741791)),(to_sfixed_a(-0.049814071506261826)),(to_sfixed_a(-0.07029025256633759)),(to_sfixed_a(-0.004401484504342079)),(to_sfixed_a(-0.0033759961370378733)),(to_sfixed_a(5.9304216847522184e-05)),(to_sfixed_a(-0.0002965606690850109)),(to_sfixed_a(-1.2059574146405794e-05)),(to_sfixed_a(6.309857326414203e-06)),(to_sfixed_a(-0.0002967215550597757)),(to_sfixed_a(-0.00033310847356915474)),(to_sfixed_a(-0.00013737642439082265)),(to_sfixed_a(-1.0172200745728333e-05)),(to_sfixed_a(0.0002105957828462124)),(to_sfixed_a(-4.932330557494424e-05)),(to_sfixed_a(-0.00018165321671403944)),(to_sfixed_a(7.918354094726965e-05)),(to_sfixed_a(-0.00021070399088785052)),(to_sfixed_a(-6.898937135701999e-05)),(to_sfixed_a(2.9677710699616e-05)),(to_sfixed_a(-8.090554183581844e-05)),(to_sfixed_a(0.00015589497343171388)),(to_sfixed_a(0.00014743955398444086)),(to_sfixed_a(-3.916327841579914e-05)),(to_sfixed_a(0.00010380456660641357)),(to_sfixed_a(-0.0001161669788416475)),(to_sfixed_a(0.0004258671251591295)),(to_sfixed_a(-9.850660717347637e-05)),(to_sfixed_a(0.00011431801249273121)),(to_sfixed_a(0.00024421015405096114)),(to_sfixed_a(4.2831878090510145e-05)),(to_sfixed_a(-9.272168972529471e-05)),(to_sfixed_a(0.0002792907180264592)),(to_sfixed_a(-0.00011097916285507381)),(to_sfixed_a(9.460924047743902e-05)),(to_sfixed_a(0.00011091191845480353)),(to_sfixed_a(-3.382677050467464e-06)),(to_sfixed_a(0.0003192428848706186)),(to_sfixed_a(0.00025444512721151114)),(to_sfixed_a(-8.653772965772077e-05)));

    constant weight_n0_4 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(8.787620026851073e-05)),(to_sfixed_a(-0.00017054950876627117)),(to_sfixed_a(5.306629100232385e-05)),(to_sfixed_a(-5.1087874453514814e-05)),(to_sfixed_a(1.6343272363883443e-05)),(to_sfixed_a(-0.00024505952023901045)),(to_sfixed_a(0.0001605019497219473)),(to_sfixed_a(2.926665729319211e-05)),(to_sfixed_a(7.814656419213861e-05)),(to_sfixed_a(-0.00015648544649593532)),(to_sfixed_a(6.725953426212072e-06)),(to_sfixed_a(-7.639380783075467e-05)),(to_sfixed_a(0.0001865629747044295)),(to_sfixed_a(5.286953819449991e-05)),(to_sfixed_a(-1.533579961687792e-05)),(to_sfixed_a(4.4427953980630264e-05)),(to_sfixed_a(-0.00023168780899140984)),(to_sfixed_a(-4.70418126496952e-05)),(to_sfixed_a(-9.638974006520584e-05)),(to_sfixed_a(-6.006733747199178e-05)),(to_sfixed_a(8.07135584182106e-05)),(to_sfixed_a(0.00010778414434753358)),(to_sfixed_a(-5.3843821660848334e-05)),(to_sfixed_a(-4.333728793426417e-05)),(to_sfixed_a(0.00022118468768894672)),(to_sfixed_a(-6.526745710289106e-05)),(to_sfixed_a(-2.578536805231124e-05)),(to_sfixed_a(-0.0001238560362253338)),(to_sfixed_a(6.663325621047989e-05)),(to_sfixed_a(-0.00015408528270199895)),(to_sfixed_a(0.00017049061716534197)),(to_sfixed_a(-0.00039915184606797993)),(to_sfixed_a(2.6975634682457894e-05)),(to_sfixed_a(0.00034483266063034534)),(to_sfixed_a(0.00020509428577497602)),(to_sfixed_a(-6.553481216542423e-05)),(to_sfixed_a(-7.397344597848132e-05)),(to_sfixed_a(-0.00013827814836986363)),(to_sfixed_a(-2.0120880435570143e-05)),(to_sfixed_a(1.3681547898158897e-05)),(to_sfixed_a(-0.00012212173896841705)),(to_sfixed_a(-6.889408541610464e-05)),(to_sfixed_a(-5.173031604499556e-05)),(to_sfixed_a(9.600264456821606e-05)),(to_sfixed_a(0.00015969092783052474)),(to_sfixed_a(-0.00020631169900298119)),(to_sfixed_a(-7.414721039822325e-05)),(to_sfixed_a(4.7077621275093406e-05)),(to_sfixed_a(0.0002394648763583973)),(to_sfixed_a(7.790126255713403e-05)),(to_sfixed_a(8.155377145158127e-05)),(to_sfixed_a(-0.0001889566919999197)),(to_sfixed_a(0.00023916742065921426)),(to_sfixed_a(-0.0001892975706141442)),(to_sfixed_a(-5.737765968660824e-05)),(to_sfixed_a(6.866428157081828e-05)),(to_sfixed_a(9.12912146304734e-05)),(to_sfixed_a(5.016239811084233e-05)),(to_sfixed_a(7.769263902446255e-05)),(to_sfixed_a(-0.00017811887664720416)),(to_sfixed_a(1.2706384040939156e-05)),(to_sfixed_a(-4.2637700971681625e-05)),(to_sfixed_a(-0.00017512412159703672)),(to_sfixed_a(-0.0003358552057761699)),(to_sfixed_a(0.00015260826330631971)),(to_sfixed_a(5.83978726353962e-05)),(to_sfixed_a(-0.00010012755228672177)),(to_sfixed_a(0.0003330692707095295)),(to_sfixed_a(-8.738015458220616e-05)),(to_sfixed_a(-0.0030559345614165068)),(to_sfixed_a(-4.379355232231319e-05)),(to_sfixed_a(-0.0002320361672900617)),(to_sfixed_a(-7.401392213068902e-05)),(to_sfixed_a(-3.9138718420872465e-05)),(to_sfixed_a(9.183982183458284e-05)),(to_sfixed_a(0.00017557704995851964)),(to_sfixed_a(-5.0024231313727796e-05)),(to_sfixed_a(1.125848211813718e-05)),(to_sfixed_a(1.078887544281315e-05)),(to_sfixed_a(0.00024559267330914736)),(to_sfixed_a(-0.00021952978568151593)),(to_sfixed_a(-6.008012860547751e-05)),(to_sfixed_a(0.00015815113147255033)),(to_sfixed_a(-3.019632822542917e-05)),(to_sfixed_a(6.383329309755936e-05)),(to_sfixed_a(0.00010029589611804113)),(to_sfixed_a(0.00030610451358370483)),(to_sfixed_a(3.488975562504493e-05)),(to_sfixed_a(5.8071502280654386e-05)),(to_sfixed_a(0.00012886531476397067)),(to_sfixed_a(8.69951782078715e-06)),(to_sfixed_a(0.00015125762729439884)),(to_sfixed_a(0.01530761830508709)),(to_sfixed_a(0.00012302870163694024)),(to_sfixed_a(0.01739456318318844)),(to_sfixed_a(-0.052260879427194595)),(to_sfixed_a(0.038495901972055435)),(to_sfixed_a(-0.0015186553355306387)),(to_sfixed_a(0.025550518184900284)),(to_sfixed_a(0.0439247228205204)),(to_sfixed_a(0.013084886595606804)),(to_sfixed_a(0.012962357141077518)),(to_sfixed_a(-0.036978334188461304)),(to_sfixed_a(-0.008096719160676003)),(to_sfixed_a(-0.000985989230684936)),(to_sfixed_a(-0.0020333644933998585)),(to_sfixed_a(-0.0003051296225748956)),(to_sfixed_a(-1.9195944332750514e-05)),(to_sfixed_a(-0.00013066134124528617)),(to_sfixed_a(5.487454836838879e-05)),(to_sfixed_a(2.3926555513753556e-05)),(to_sfixed_a(-3.072273830184713e-05)),(to_sfixed_a(0.00017483922420069575)),(to_sfixed_a(1.9111317669739947e-05)),(to_sfixed_a(0.00012347781739663333)),(to_sfixed_a(5.421613604994491e-05)),(to_sfixed_a(6.512026448035613e-05)),(to_sfixed_a(-0.0001505302352597937)),(to_sfixed_a(0.0009411094943061471)),(to_sfixed_a(-0.03877285122871399)),(to_sfixed_a(-0.03464126214385033)),(to_sfixed_a(0.028827453032135963)),(to_sfixed_a(0.041681043803691864)),(to_sfixed_a(-0.00826707761734724)),(to_sfixed_a(0.08515701442956924)),(to_sfixed_a(-0.027736255899071693)),(to_sfixed_a(-0.1002606526017189)),(to_sfixed_a(-0.050233665853738785)),(to_sfixed_a(-0.19903236627578735)),(to_sfixed_a(-0.026201320812106133)),(to_sfixed_a(-0.02708347514271736)),(to_sfixed_a(-0.024700473994016647)),(to_sfixed_a(-0.0008886433206498623)),(to_sfixed_a(-0.013579891063272953)),(to_sfixed_a(0.11883045732975006)),(to_sfixed_a(0.0006189111154526472)),(to_sfixed_a(-0.0015441245632246137)),(to_sfixed_a(-0.0001284575992031023)),(to_sfixed_a(-8.306924428325146e-05)),(to_sfixed_a(-5.036377478973009e-05)),(to_sfixed_a(-1.8424991139909253e-05)),(to_sfixed_a(3.266832572990097e-05)),(to_sfixed_a(7.124871626729146e-05)),(to_sfixed_a(-4.805091884918511e-05)),(to_sfixed_a(-0.0002442077675368637)),(to_sfixed_a(-0.05655904486775398)),(to_sfixed_a(0.0022357236593961716)),(to_sfixed_a(-0.003367482451722026)),(to_sfixed_a(-0.007235497701913118)),(to_sfixed_a(0.011345403268933296)),(to_sfixed_a(0.015434247441589832)),(to_sfixed_a(-0.0473177507519722)),(to_sfixed_a(0.060696568340063095)),(to_sfixed_a(0.00477168383076787)),(to_sfixed_a(-0.016307901591062546)),(to_sfixed_a(0.05899424105882645)),(to_sfixed_a(0.10242073982954025)),(to_sfixed_a(-0.00656833965331316)),(to_sfixed_a(0.09887068718671799)),(to_sfixed_a(0.25658100843429565)),(to_sfixed_a(-0.1763029545545578)),(to_sfixed_a(-0.0022247808519750834)),(to_sfixed_a(-0.0011928811436519027)),(to_sfixed_a(0.02398993819952011)),(to_sfixed_a(-0.001838325522840023)),(to_sfixed_a(-0.00016664747090544552)),(to_sfixed_a(-0.00025870130048133433)),(to_sfixed_a(0.00016963158850558102)),(to_sfixed_a(0.00020284643687773496)),(to_sfixed_a(-2.387950189586263e-05)),(to_sfixed_a(0.0002204533520853147)),(to_sfixed_a(0.00021139481395948678)),(to_sfixed_a(-3.480273517197929e-05)),(to_sfixed_a(-0.05440009385347366)),(to_sfixed_a(-0.0774373933672905)),(to_sfixed_a(-0.14072692394256592)),(to_sfixed_a(0.028892850503325462)),(to_sfixed_a(0.15775711834430695)),(to_sfixed_a(0.15421618521213531)),(to_sfixed_a(0.04205198958516121)),(to_sfixed_a(-0.09612391144037247)),(to_sfixed_a(0.13488012552261353)),(to_sfixed_a(0.12325671315193176)),(to_sfixed_a(0.03726740553975105)),(to_sfixed_a(-0.03808722645044327)),(to_sfixed_a(0.0772676169872284)),(to_sfixed_a(-0.039477575570344925)),(to_sfixed_a(-0.06990876793861389)),(to_sfixed_a(-0.0812973901629448)),(to_sfixed_a(0.03765900805592537)),(to_sfixed_a(0.03501644730567932)),(to_sfixed_a(0.07095120847225189)),(to_sfixed_a(0.002173582324758172)),(to_sfixed_a(0.003534207120537758)),(to_sfixed_a(0.0026899485383182764)),(to_sfixed_a(-0.00029067305149510503)),(to_sfixed_a(6.84548940625973e-05)),(to_sfixed_a(8.551392966182902e-05)),(to_sfixed_a(-0.00022038949828129262)),(to_sfixed_a(0.00011950332554988563)),(to_sfixed_a(-0.00010405087959952652)),(to_sfixed_a(0.007279667071998119)),(to_sfixed_a(-0.19681155681610107)),(to_sfixed_a(-0.040355779230594635)),(to_sfixed_a(0.20263159275054932)),(to_sfixed_a(-0.06664068251848221)),(to_sfixed_a(0.0687689259648323)),(to_sfixed_a(0.05991298332810402)),(to_sfixed_a(-0.07795164734125137)),(to_sfixed_a(0.13415074348449707)),(to_sfixed_a(-0.02453635446727276)),(to_sfixed_a(0.06508401036262512)),(to_sfixed_a(0.19579510390758514)),(to_sfixed_a(-0.05980316177010536)),(to_sfixed_a(-0.09261955320835114)),(to_sfixed_a(0.11000511050224304)),(to_sfixed_a(-0.01660323143005371)),(to_sfixed_a(-0.11315418779850006)),(to_sfixed_a(-0.04187105968594551)),(to_sfixed_a(-0.1317170113325119)),(to_sfixed_a(0.014492218382656574)),(to_sfixed_a(-0.004547080025076866)),(to_sfixed_a(-0.0001423338399035856)),(to_sfixed_a(6.21810759184882e-05)),(to_sfixed_a(-5.994784805807285e-05)),(to_sfixed_a(6.026200935593806e-05)),(to_sfixed_a(-0.0001174578137579374)),(to_sfixed_a(-4.4710068323183805e-06)),(to_sfixed_a(-0.03708851337432861)),(to_sfixed_a(-0.02707359567284584)),(to_sfixed_a(-0.011078638024628162)),(to_sfixed_a(-0.0008552400395274162)),(to_sfixed_a(0.03438305854797363)),(to_sfixed_a(0.09786690771579742)),(to_sfixed_a(-0.0586048848927021)),(to_sfixed_a(-0.05296164005994797)),(to_sfixed_a(0.02842932753264904)),(to_sfixed_a(0.16212771832942963)),(to_sfixed_a(0.0330694206058979)),(to_sfixed_a(0.014056835323572159)),(to_sfixed_a(-0.02325424738228321)),(to_sfixed_a(-0.03112785518169403)),(to_sfixed_a(-0.25131410360336304)),(to_sfixed_a(-0.058589816093444824)),(to_sfixed_a(-0.24529361724853516)),(to_sfixed_a(-0.08814627677202225)),(to_sfixed_a(-0.027782144024968147)),(to_sfixed_a(-0.135166198015213)),(to_sfixed_a(-0.10218683630228043)),(to_sfixed_a(0.005430268589407206)),(to_sfixed_a(0.00010640854452503845)),(to_sfixed_a(8.630665251985192e-05)),(to_sfixed_a(-8.73929457156919e-05)),(to_sfixed_a(8.649959636386484e-05)),(to_sfixed_a(0.0002142989105777815)),(to_sfixed_a(-0.00027523087919689715)),(to_sfixed_a(-0.002630175556987524)),(to_sfixed_a(-0.13740967214107513)),(to_sfixed_a(-0.011720886453986168)),(to_sfixed_a(0.03902135789394379)),(to_sfixed_a(0.08730890601873398)),(to_sfixed_a(0.05163514241576195)),(to_sfixed_a(0.33610203862190247)),(to_sfixed_a(0.12029118090867996)),(to_sfixed_a(0.05906405299901962)),(to_sfixed_a(0.008559919893741608)),(to_sfixed_a(-0.08327639102935791)),(to_sfixed_a(-0.10150658339262009)),(to_sfixed_a(-0.12361779063940048)),(to_sfixed_a(-0.10439526289701462)),(to_sfixed_a(-0.10258867591619492)),(to_sfixed_a(-0.17651259899139404)),(to_sfixed_a(-0.061791062355041504)),(to_sfixed_a(0.008265256881713867)),(to_sfixed_a(0.055819492787122726)),(to_sfixed_a(0.07558337599039078)),(to_sfixed_a(0.014041541144251823)),(to_sfixed_a(1.6212050468311645e-05)),(to_sfixed_a(3.9915015804581344e-05)),(to_sfixed_a(-7.238405669340864e-05)),(to_sfixed_a(-0.0002609950315672904)),(to_sfixed_a(5.485540532390587e-05)),(to_sfixed_a(-8.006291318451986e-05)),(to_sfixed_a(-6.122421473264694e-05)),(to_sfixed_a(-0.003420049324631691)),(to_sfixed_a(0.024706825613975525)),(to_sfixed_a(0.14981158077716827)),(to_sfixed_a(0.1272558867931366)),(to_sfixed_a(0.11345984041690826)),(to_sfixed_a(0.1570689082145691)),(to_sfixed_a(0.17536453902721405)),(to_sfixed_a(-0.08707393705844879)),(to_sfixed_a(0.10728418081998825)),(to_sfixed_a(-0.3943382799625397)),(to_sfixed_a(0.10410575568675995)),(to_sfixed_a(0.10397767275571823)),(to_sfixed_a(-0.03369555622339249)),(to_sfixed_a(-0.019189029932022095)),(to_sfixed_a(0.0073820059187710285)),(to_sfixed_a(-0.12757356464862823)),(to_sfixed_a(-0.03195947781205177)),(to_sfixed_a(-0.023398293182253838)),(to_sfixed_a(-0.017512256279587746)),(to_sfixed_a(-0.1321568787097931)),(to_sfixed_a(-0.04992067813873291)),(to_sfixed_a(-0.013630918227136135)),(to_sfixed_a(-1.9531646103132516e-05)),(to_sfixed_a(-0.00017658236902207136)),(to_sfixed_a(-0.0001942522794706747)),(to_sfixed_a(-0.00011272619303781539)),(to_sfixed_a(-3.1554754968965426e-05)),(to_sfixed_a(-0.025524262338876724)),(to_sfixed_a(-0.05825059488415718)),(to_sfixed_a(0.1507936418056488)),(to_sfixed_a(0.06828440725803375)),(to_sfixed_a(0.144905224442482)),(to_sfixed_a(0.1670515388250351)),(to_sfixed_a(-0.07190432399511337)),(to_sfixed_a(0.016506023705005646)),(to_sfixed_a(-0.28556063771247864)),(to_sfixed_a(-0.25110334157943726)),(to_sfixed_a(-0.09325777739286423)),(to_sfixed_a(0.29593005776405334)),(to_sfixed_a(0.16375212371349335)),(to_sfixed_a(0.06947116553783417)),(to_sfixed_a(0.139716237783432)),(to_sfixed_a(0.3026503026485443)),(to_sfixed_a(0.07837969064712524)),(to_sfixed_a(0.08261554688215256)),(to_sfixed_a(0.018416576087474823)),(to_sfixed_a(0.08348531275987625)),(to_sfixed_a(-0.12040030211210251)),(to_sfixed_a(-0.1328846514225006)),(to_sfixed_a(0.00016397054423578084)),(to_sfixed_a(-0.00020049001614097506)),(to_sfixed_a(-1.4047141121409368e-05)),(to_sfixed_a(0.00017692643450573087)),(to_sfixed_a(-0.0001371804828522727)),(to_sfixed_a(-8.235479617724195e-05)),(to_sfixed_a(0.00024499985738657415)),(to_sfixed_a(0.08801811933517456)),(to_sfixed_a(-0.13267774879932404)),(to_sfixed_a(0.023026159033179283)),(to_sfixed_a(0.08585222065448761)),(to_sfixed_a(-0.1248839795589447)),(to_sfixed_a(-0.179705411195755)),(to_sfixed_a(-0.3451401889324188)),(to_sfixed_a(-0.48460525274276733)),(to_sfixed_a(-0.10328494012355804)),(to_sfixed_a(0.3362245261669159)),(to_sfixed_a(0.40577295422554016)),(to_sfixed_a(0.16959671676158905)),(to_sfixed_a(0.39597660303115845)),(to_sfixed_a(0.19720865786075592)),(to_sfixed_a(0.05307799205183983)),(to_sfixed_a(0.20923376083374023)),(to_sfixed_a(-0.15232935547828674)),(to_sfixed_a(0.10891222208738327)),(to_sfixed_a(0.1428280919790268)),(to_sfixed_a(0.18652580678462982)),(to_sfixed_a(-0.013934366405010223)),(to_sfixed_a(2.3534914362244308e-05)),(to_sfixed_a(0.0001888537226477638)),(to_sfixed_a(-5.6979361033882014e-06)),(to_sfixed_a(4.517783236224204e-05)),(to_sfixed_a(-0.00015147592057473958)),(to_sfixed_a(-0.0005281860940158367)),(to_sfixed_a(0.00040188271668739617)),(to_sfixed_a(-0.04811546206474304)),(to_sfixed_a(-0.08020062744617462)),(to_sfixed_a(-0.3807150423526764)),(to_sfixed_a(-0.15898190438747406)),(to_sfixed_a(-0.2967652678489685)),(to_sfixed_a(-0.0003530653193593025)),(to_sfixed_a(-0.20092599093914032)),(to_sfixed_a(-0.050545889884233475)),(to_sfixed_a(0.08394407480955124)),(to_sfixed_a(0.7017003297805786)),(to_sfixed_a(0.6984500288963318)),(to_sfixed_a(0.3139721155166626)),(to_sfixed_a(0.08659657835960388)),(to_sfixed_a(0.13425883650779724)),(to_sfixed_a(0.011562059633433819)),(to_sfixed_a(0.08789759874343872)),(to_sfixed_a(0.11300652474164963)),(to_sfixed_a(-0.015270703472197056)),(to_sfixed_a(0.018162697553634644)),(to_sfixed_a(0.08521861582994461)),(to_sfixed_a(0.018592489883303642)),(to_sfixed_a(-0.001974242739379406)),(to_sfixed_a(-0.0014610814396291971)),(to_sfixed_a(-0.00013687221508007497)),(to_sfixed_a(9.851808135863394e-05)),(to_sfixed_a(0.0001770943053998053)),(to_sfixed_a(0.00047789435484446585)),(to_sfixed_a(1.573509507579729e-05)),(to_sfixed_a(0.002792647108435631)),(to_sfixed_a(-0.2881230413913727)),(to_sfixed_a(-0.012018912471830845)),(to_sfixed_a(-0.2443704754114151)),(to_sfixed_a(0.06305251270532608)),(to_sfixed_a(-0.31366679072380066)),(to_sfixed_a(-0.11395639181137085)),(to_sfixed_a(-0.07742960751056671)),(to_sfixed_a(0.6339347958564758)),(to_sfixed_a(0.8740556240081787)),(to_sfixed_a(0.5783506631851196)),(to_sfixed_a(0.1786992847919464)),(to_sfixed_a(0.1763010025024414)),(to_sfixed_a(0.011392548680305481)),(to_sfixed_a(-0.02583269774913788)),(to_sfixed_a(-0.2218881994485855)),(to_sfixed_a(-0.10101714730262756)),(to_sfixed_a(0.0230987761169672)),(to_sfixed_a(0.003595740767195821)),(to_sfixed_a(-0.17363010346889496)),(to_sfixed_a(-0.0477563701570034)),(to_sfixed_a(0.0003261837409809232)),(to_sfixed_a(-0.00026134151266887784)),(to_sfixed_a(-5.234383206698112e-05)),(to_sfixed_a(-5.419543958851136e-05)),(to_sfixed_a(-3.1356299587059766e-05)),(to_sfixed_a(-0.0003146465460304171)),(to_sfixed_a(-1.4635253137385007e-05)),(to_sfixed_a(-0.0663464292883873)),(to_sfixed_a(0.11716368794441223)),(to_sfixed_a(0.02592514082789421)),(to_sfixed_a(-0.007994428277015686)),(to_sfixed_a(0.11468308418989182)),(to_sfixed_a(0.24508598446846008)),(to_sfixed_a(0.36160096526145935)),(to_sfixed_a(0.41815879940986633)),(to_sfixed_a(0.7680930495262146)),(to_sfixed_a(1.099413275718689)),(to_sfixed_a(0.30665698647499084)),(to_sfixed_a(0.07539442181587219)),(to_sfixed_a(0.022368818521499634)),(to_sfixed_a(-0.09621212631464005)),(to_sfixed_a(-0.22238974273204803)),(to_sfixed_a(-0.07422903180122375)),(to_sfixed_a(-0.16413404047489166)),(to_sfixed_a(-0.011669122613966465)),(to_sfixed_a(-0.07698168605566025)),(to_sfixed_a(-0.1321507841348648)),(to_sfixed_a(-0.08559054136276245)),(to_sfixed_a(-3.5360259062144905e-05)),(to_sfixed_a(-0.00018960569286718965)),(to_sfixed_a(5.083410724182613e-05)),(to_sfixed_a(-3.318617382319644e-05)),(to_sfixed_a(0.0001284214959014207)),(to_sfixed_a(0.0002250920661026612)),(to_sfixed_a(0.0022421949543058872)),(to_sfixed_a(-0.08191442489624023)),(to_sfixed_a(-0.4929720461368561)),(to_sfixed_a(-0.8551101684570312)),(to_sfixed_a(-0.7730817794799805)),(to_sfixed_a(-0.5114004611968994)),(to_sfixed_a(-0.05886045843362808)),(to_sfixed_a(0.4791634678840637)),(to_sfixed_a(0.858680009841919)),(to_sfixed_a(0.9318419098854065)),(to_sfixed_a(0.8701635003089905)),(to_sfixed_a(0.06955938786268234)),(to_sfixed_a(0.018238091841340065)),(to_sfixed_a(-0.020690850913524628)),(to_sfixed_a(-0.1570218801498413)),(to_sfixed_a(-0.1962096244096756)),(to_sfixed_a(-0.21940593421459198)),(to_sfixed_a(-0.14668554067611694)),(to_sfixed_a(-0.10471811145544052)),(to_sfixed_a(-0.023071544244885445)),(to_sfixed_a(0.08551717549562454)),(to_sfixed_a(-0.012539416551589966)),(to_sfixed_a(0.025698835030198097)),(to_sfixed_a(-1.266224353457801e-05)),(to_sfixed_a(3.993534846813418e-05)),(to_sfixed_a(7.270458445418626e-05)),(to_sfixed_a(0.00022157053172122687)),(to_sfixed_a(0.001363943563774228)),(to_sfixed_a(0.002338459948077798)),(to_sfixed_a(-0.09504784643650055)),(to_sfixed_a(-0.4974280595779419)),(to_sfixed_a(-0.46288391947746277)),(to_sfixed_a(-0.46332257986068726)),(to_sfixed_a(-0.7034745216369629)),(to_sfixed_a(-0.5525832176208496)),(to_sfixed_a(-0.31866174936294556)),(to_sfixed_a(0.1948811411857605)),(to_sfixed_a(0.6929913759231567)),(to_sfixed_a(0.08670610934495926)),(to_sfixed_a(0.1176997646689415)),(to_sfixed_a(-0.129945307970047)),(to_sfixed_a(-0.26000550389289856)),(to_sfixed_a(-0.2542911767959595)),(to_sfixed_a(-0.1824500560760498)),(to_sfixed_a(-0.13637107610702515)),(to_sfixed_a(-0.005219238344579935)),(to_sfixed_a(0.014620005153119564)),(to_sfixed_a(-0.20157048106193542)),(to_sfixed_a(0.01599884405732155)),(to_sfixed_a(2.4993087208713405e-05)),(to_sfixed_a(0.00024605970247648656)),(to_sfixed_a(2.7717131160898134e-05)),(to_sfixed_a(3.7139041523914784e-05)),(to_sfixed_a(0.00023168823099695146)),(to_sfixed_a(6.555200525326654e-05)),(to_sfixed_a(0.0002765218960121274)),(to_sfixed_a(-0.007238788530230522)),(to_sfixed_a(-0.0828440934419632)),(to_sfixed_a(-0.23670382797718048)),(to_sfixed_a(-0.341502845287323)),(to_sfixed_a(-0.5041407942771912)),(to_sfixed_a(-0.7192566394805908)),(to_sfixed_a(-0.42975449562072754)),(to_sfixed_a(-0.44492942094802856)),(to_sfixed_a(-0.012487259693443775)),(to_sfixed_a(-0.3519546091556549)),(to_sfixed_a(-0.21682897210121155)),(to_sfixed_a(-0.27314335107803345)),(to_sfixed_a(-0.19386659562587738)),(to_sfixed_a(-0.10941048711538315)),(to_sfixed_a(-0.2532217502593994)),(to_sfixed_a(-0.21519528329372406)),(to_sfixed_a(-0.07684449106454849)),(to_sfixed_a(-0.060518402606248856)),(to_sfixed_a(0.054151374846696854)),(to_sfixed_a(-0.056372977793216705)),(to_sfixed_a(0.04380811005830765)),(to_sfixed_a(0.04076313227415085)),(to_sfixed_a(-1.931504266394768e-05)),(to_sfixed_a(0.00015851360512897372)),(to_sfixed_a(-5.5164797231554985e-05)),(to_sfixed_a(-4.844474824494682e-05)),(to_sfixed_a(-0.0002402470272500068)),(to_sfixed_a(-3.3865471777971834e-06)),(to_sfixed_a(-0.0806097462773323)),(to_sfixed_a(0.0067386687733232975)),(to_sfixed_a(-0.026609258726239204)),(to_sfixed_a(-0.11406739801168442)),(to_sfixed_a(-0.27274563908576965)),(to_sfixed_a(-0.5033494830131531)),(to_sfixed_a(-0.3867948055267334)),(to_sfixed_a(-0.50958251953125)),(to_sfixed_a(-0.2761036157608032)),(to_sfixed_a(-0.45051899552345276)),(to_sfixed_a(-0.3384341299533844)),(to_sfixed_a(-0.4835829734802246)),(to_sfixed_a(-0.23414190113544464)),(to_sfixed_a(0.0010956694604828954)),(to_sfixed_a(-0.12130679190158844)),(to_sfixed_a(-0.05901676416397095)),(to_sfixed_a(0.030435768887400627)),(to_sfixed_a(-0.12398918718099594)),(to_sfixed_a(0.10628359019756317)),(to_sfixed_a(-0.06491631269454956)),(to_sfixed_a(0.08117055892944336)),(to_sfixed_a(-1.1860302038257942e-05)),(to_sfixed_a(7.950594590511173e-05)),(to_sfixed_a(-0.00011696250294335186)),(to_sfixed_a(-0.0002827302960213274)),(to_sfixed_a(-8.173652895493433e-05)),(to_sfixed_a(0.00014762200589757413)),(to_sfixed_a(-0.0001609580940566957)),(to_sfixed_a(-1.4970541997172404e-05)),(to_sfixed_a(-0.025208568200469017)),(to_sfixed_a(-0.01669572852551937)),(to_sfixed_a(0.005627643316984177)),(to_sfixed_a(-0.026982471346855164)),(to_sfixed_a(0.1530425250530243)),(to_sfixed_a(0.056081973016262054)),(to_sfixed_a(-0.050770096480846405)),(to_sfixed_a(0.1436711847782135)),(to_sfixed_a(-0.2060716152191162)),(to_sfixed_a(0.04029807075858116)),(to_sfixed_a(-0.13411982357501984)),(to_sfixed_a(-0.04169582203030586)),(to_sfixed_a(-0.05428003519773483)),(to_sfixed_a(-0.1492260843515396)),(to_sfixed_a(0.25457361340522766)),(to_sfixed_a(0.12357297539710999)),(to_sfixed_a(0.1683197170495987)),(to_sfixed_a(0.07221904397010803)),(to_sfixed_a(0.010315821506083012)),(to_sfixed_a(-0.023033279925584793)),(to_sfixed_a(-0.04314405471086502)),(to_sfixed_a(5.306177627062425e-05)),(to_sfixed_a(0.00014437880599871278)),(to_sfixed_a(-2.901791231124662e-05)),(to_sfixed_a(-9.507335562375374e-06)),(to_sfixed_a(-0.00010987371933879331)),(to_sfixed_a(5.683866766048595e-05)),(to_sfixed_a(5.396932829171419e-05)),(to_sfixed_a(0.009485830552875996)),(to_sfixed_a(0.0013109594583511353)),(to_sfixed_a(0.21567003428936005)),(to_sfixed_a(0.2271811068058014)),(to_sfixed_a(0.27613791823387146)),(to_sfixed_a(0.05897637456655502)),(to_sfixed_a(0.1636492908000946)),(to_sfixed_a(-0.17657937109470367)),(to_sfixed_a(0.06898273527622223)),(to_sfixed_a(0.05393499135971069)),(to_sfixed_a(0.15671131014823914)),(to_sfixed_a(-0.1385146677494049)),(to_sfixed_a(-0.07297348231077194)),(to_sfixed_a(-0.19835643470287323)),(to_sfixed_a(-0.1220538467168808)),(to_sfixed_a(-0.009430167265236378)),(to_sfixed_a(0.0006692706956528127)),(to_sfixed_a(-0.015927158296108246)),(to_sfixed_a(0.034946952015161514)),(to_sfixed_a(3.3814620110206306e-05)),(to_sfixed_a(-0.04351118206977844)),(to_sfixed_a(-9.497849532635882e-05)),(to_sfixed_a(0.0001726293412502855)),(to_sfixed_a(-0.00018578552408143878)),(to_sfixed_a(2.6305880965082906e-05)),(to_sfixed_a(-8.628270006738603e-05)),(to_sfixed_a(-0.00026184055604971945)),(to_sfixed_a(1.4823305718891788e-05)),(to_sfixed_a(0.00010256865061819553)),(to_sfixed_a(0.08671201765537262)),(to_sfixed_a(0.02674955315887928)),(to_sfixed_a(0.19483745098114014)),(to_sfixed_a(-0.13987068831920624)),(to_sfixed_a(0.015204837545752525)),(to_sfixed_a(0.05914444103837013)),(to_sfixed_a(0.2946401834487915)),(to_sfixed_a(0.159925639629364)),(to_sfixed_a(-0.05182661861181259)),(to_sfixed_a(0.09300442039966583)),(to_sfixed_a(-0.06840449571609497)),(to_sfixed_a(-0.08113081753253937)),(to_sfixed_a(-0.06412898749113083)),(to_sfixed_a(0.15717048943042755)),(to_sfixed_a(-0.11043644696474075)),(to_sfixed_a(-0.059043969959020615)),(to_sfixed_a(0.0015612904680892825)),(to_sfixed_a(-0.05266325920820236)),(to_sfixed_a(-0.0037293711211532354)),(to_sfixed_a(2.78753195743775e-05)),(to_sfixed_a(0.0001804641360649839)),(to_sfixed_a(-1.5290919463950559e-06)),(to_sfixed_a(5.6096541811712086e-05)),(to_sfixed_a(4.4825388613389805e-05)),(to_sfixed_a(-3.925415512640029e-05)),(to_sfixed_a(0.0001089619254344143)),(to_sfixed_a(0.00013140295050106943)),(to_sfixed_a(-0.00020654873515013605)),(to_sfixed_a(0.029850687831640244)),(to_sfixed_a(0.07493841648101807)),(to_sfixed_a(0.16081275045871735)),(to_sfixed_a(0.2676430344581604)),(to_sfixed_a(0.017016591504216194)),(to_sfixed_a(0.20095811784267426)),(to_sfixed_a(0.20036587119102478)),(to_sfixed_a(0.17078550159931183)),(to_sfixed_a(0.07811007648706436)),(to_sfixed_a(0.061929743736982346)),(to_sfixed_a(-0.08676473796367645)),(to_sfixed_a(0.10752596706151962)),(to_sfixed_a(-0.04140423238277435)),(to_sfixed_a(0.2001209408044815)),(to_sfixed_a(0.026122933253645897)),(to_sfixed_a(0.01083647646009922)),(to_sfixed_a(-0.02093498408794403)),(to_sfixed_a(0.0003679529472719878)),(to_sfixed_a(-0.017314204946160316)),(to_sfixed_a(0.0001523983955848962)),(to_sfixed_a(-7.085997640388086e-05)),(to_sfixed_a(-8.590820652898401e-05)),(to_sfixed_a(2.2460148102254607e-05)),(to_sfixed_a(0.0002581265289336443)),(to_sfixed_a(-0.00011953144712606445)),(to_sfixed_a(6.874031532788649e-05)),(to_sfixed_a(-8.279242319986224e-05)),(to_sfixed_a(0.0029292346443980932)),(to_sfixed_a(0.03842722997069359)),(to_sfixed_a(0.013373153284192085)),(to_sfixed_a(0.44316431879997253)),(to_sfixed_a(0.15931063890457153)),(to_sfixed_a(0.1456969678401947)),(to_sfixed_a(0.16689366102218628)),(to_sfixed_a(0.26876100897789)),(to_sfixed_a(0.17598359286785126)),(to_sfixed_a(0.06049279123544693)),(to_sfixed_a(0.1969141811132431)),(to_sfixed_a(-0.011284515261650085)),(to_sfixed_a(-0.17889058589935303)),(to_sfixed_a(-0.19769248366355896)),(to_sfixed_a(-0.08152379095554352)),(to_sfixed_a(-0.04755260795354843)),(to_sfixed_a(0.004151606000959873)),(to_sfixed_a(0.0005208759102970362)),(to_sfixed_a(0.00693786283954978)),(to_sfixed_a(0.015639502555131912)),(to_sfixed_a(0.00010281798313371837)),(to_sfixed_a(0.00039131080848164856)),(to_sfixed_a(0.00020977313397452235)),(to_sfixed_a(-0.00019348481146153063)),(to_sfixed_a(-1.6612517356406897e-05)),(to_sfixed_a(5.9711335779866204e-05)),(to_sfixed_a(0.00017740437760949135)),(to_sfixed_a(-0.0002414429181953892)),(to_sfixed_a(2.1022671717219055e-05)),(to_sfixed_a(-0.03143544867634773)),(to_sfixed_a(0.0073585971258580685)),(to_sfixed_a(0.005700818728655577)),(to_sfixed_a(0.04392817243933678)),(to_sfixed_a(0.038702115416526794)),(to_sfixed_a(0.2967463433742523)),(to_sfixed_a(0.0675833597779274)),(to_sfixed_a(0.15129464864730835)),(to_sfixed_a(0.09071912616491318)),(to_sfixed_a(0.05269646272063255)),(to_sfixed_a(-0.02879047580063343)),(to_sfixed_a(0.014229784719645977)),(to_sfixed_a(-0.04686935618519783)),(to_sfixed_a(0.004279920365661383)),(to_sfixed_a(-0.002462460659444332)),(to_sfixed_a(0.017702946439385414)),(to_sfixed_a(-0.0002223859919467941)),(to_sfixed_a(0.0011417618952691555)),(to_sfixed_a(0.0018813071073964238)),(to_sfixed_a(-4.8819591029314324e-05)),(to_sfixed_a(-4.262573929736391e-05)),(to_sfixed_a(5.1761333452304825e-05)),(to_sfixed_a(-3.1045427022036165e-05)),(to_sfixed_a(5.306800403559464e-07)),(to_sfixed_a(9.748661796038505e-06)),(to_sfixed_a(-6.235428736545146e-05)),(to_sfixed_a(-6.400190613931045e-05)),(to_sfixed_a(0.0001802421174943447)),(to_sfixed_a(0.0006016689003445208)),(to_sfixed_a(0.0008700813050381839)),(to_sfixed_a(-6.913980178069323e-05)),(to_sfixed_a(5.912251435802318e-05)),(to_sfixed_a(-0.00045990385115146637)),(to_sfixed_a(0.011611344292759895)),(to_sfixed_a(0.01082556787878275)),(to_sfixed_a(0.0034256211947649717)),(to_sfixed_a(0.006350786425173283)),(to_sfixed_a(-0.0317838080227375)),(to_sfixed_a(-0.016840185970067978)),(to_sfixed_a(0.0022131777368485928)),(to_sfixed_a(0.004172558430582285)),(to_sfixed_a(0.006357417441904545)),(to_sfixed_a(-0.0026588912587612867)),(to_sfixed_a(-0.001680342829786241)),(to_sfixed_a(3.0724315820407355e-06)),(to_sfixed_a(-6.21935396338813e-05)),(to_sfixed_a(-0.00029881118098273873)),(to_sfixed_a(9.345349099021405e-05)),(to_sfixed_a(0.00041911975131370127)),(to_sfixed_a(8.388271766079924e-08)),(to_sfixed_a(-3.7346901081036776e-05)),(to_sfixed_a(-0.00018816019291989505)),(to_sfixed_a(1.4796527466387488e-05)),(to_sfixed_a(2.8733389626722783e-05)),(to_sfixed_a(-0.0001387201191391796)),(to_sfixed_a(-0.00013165167183615267)),(to_sfixed_a(4.592942786985077e-05)),(to_sfixed_a(-0.0004272855294402689)),(to_sfixed_a(-0.0001726381160551682)),(to_sfixed_a(-0.0002727170358411968)),(to_sfixed_a(-0.0002978566335514188)),(to_sfixed_a(4.866273229708895e-05)),(to_sfixed_a(5.8874931710306555e-05)),(to_sfixed_a(-0.00011460899986559525)),(to_sfixed_a(-2.9449503927025944e-05)),(to_sfixed_a(0.00020045759447384626)),(to_sfixed_a(0.00020525498257484287)),(to_sfixed_a(0.00011804773384938017)),(to_sfixed_a(-0.00017761685012374073)),(to_sfixed_a(-3.523439590935595e-05)),(to_sfixed_a(-4.241497299517505e-05)),(to_sfixed_a(5.550554487854242e-05)),(to_sfixed_a(-7.125730189727619e-05)),(to_sfixed_a(-0.0001115965933422558)),(to_sfixed_a(0.0001856360031524673)),(to_sfixed_a(1.454877474316163e-05)),(to_sfixed_a(-9.650673746364191e-05)),(to_sfixed_a(0.0003728304582182318)),(to_sfixed_a(0.00012913935643155128)));

    constant weight_n0_5 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-3.7188088754191995e-05)),(to_sfixed_a(0.00011999334674328566)),(to_sfixed_a(-0.00027145270723849535)),(to_sfixed_a(-1.327226073044585e-05)),(to_sfixed_a(-0.000290295371087268)),(to_sfixed_a(0.00014644261682406068)),(to_sfixed_a(0.00030866972520016134)),(to_sfixed_a(8.72340242494829e-05)),(to_sfixed_a(-8.373514720005915e-05)),(to_sfixed_a(-0.0001380344183417037)),(to_sfixed_a(0.00018439417181070894)),(to_sfixed_a(9.36814922170015e-06)),(to_sfixed_a(-0.0002955399395432323)),(to_sfixed_a(-0.0003171995631419122)),(to_sfixed_a(-3.9468719478463754e-05)),(to_sfixed_a(-0.00014349090633913875)),(to_sfixed_a(0.00010798087168950588)),(to_sfixed_a(-0.00011273650306975469)),(to_sfixed_a(0.0001690464123385027)),(to_sfixed_a(-0.0002501932031009346)),(to_sfixed_a(7.17645525583066e-05)),(to_sfixed_a(0.00036440257099457085)),(to_sfixed_a(-5.3310450311983004e-05)),(to_sfixed_a(-2.026220272455248e-06)),(to_sfixed_a(-0.00031021019094623625)),(to_sfixed_a(0.00010703325824579224)),(to_sfixed_a(0.0001867789978859946)),(to_sfixed_a(-5.203639011597261e-05)),(to_sfixed_a(-6.132336420705542e-05)),(to_sfixed_a(-0.00016452120325993747)),(to_sfixed_a(-0.00014206650666892529)),(to_sfixed_a(0.00027501076692715287)),(to_sfixed_a(8.86806592461653e-05)),(to_sfixed_a(0.00023443518148269504)),(to_sfixed_a(0.00013629432942252606)),(to_sfixed_a(0.0002823840477503836)),(to_sfixed_a(-2.869901800295338e-05)),(to_sfixed_a(8.05448871687986e-05)),(to_sfixed_a(-0.00019893705029971898)),(to_sfixed_a(0.00034174160100519657)),(to_sfixed_a(-0.00019159297517035156)),(to_sfixed_a(-1.193377647723537e-05)),(to_sfixed_a(0.00012703986431006342)),(to_sfixed_a(0.00020908254373352975)),(to_sfixed_a(0.0003853580274153501)),(to_sfixed_a(1.7004809706122614e-05)),(to_sfixed_a(0.0002653926203493029)),(to_sfixed_a(-4.840076144319028e-05)),(to_sfixed_a(-0.00016365245392080396)),(to_sfixed_a(-0.00024037595721893013)),(to_sfixed_a(5.553944720304571e-05)),(to_sfixed_a(-4.561927562463097e-05)),(to_sfixed_a(9.518268052488565e-05)),(to_sfixed_a(5.653141488437541e-05)),(to_sfixed_a(-0.00015377564704976976)),(to_sfixed_a(-0.00031114197918213904)),(to_sfixed_a(-0.00020932703046128154)),(to_sfixed_a(1.0545427358010784e-05)),(to_sfixed_a(0.00011467421427369118)),(to_sfixed_a(-1.1118547263322398e-05)),(to_sfixed_a(-4.510654980549589e-05)),(to_sfixed_a(0.00010003977513406426)),(to_sfixed_a(0.00010351373930461705)),(to_sfixed_a(-0.00011682027979986742)),(to_sfixed_a(-0.00011464174167485908)),(to_sfixed_a(-8.808085840428248e-05)),(to_sfixed_a(7.404005737043917e-05)),(to_sfixed_a(7.258963887579739e-05)),(to_sfixed_a(8.665659697726369e-05)),(to_sfixed_a(-0.0031410115770995617)),(to_sfixed_a(-0.00017235710402019322)),(to_sfixed_a(-0.00011667313810903579)),(to_sfixed_a(4.282635927665979e-05)),(to_sfixed_a(0.0001109372969949618)),(to_sfixed_a(-0.00015013226948212832)),(to_sfixed_a(3.105675568804145e-05)),(to_sfixed_a(0.0001427763345418498)),(to_sfixed_a(6.044406472938135e-05)),(to_sfixed_a(-5.739813786931336e-05)),(to_sfixed_a(0.00016421113105025142)),(to_sfixed_a(-0.0001457293110433966)),(to_sfixed_a(-0.0002058929967461154)),(to_sfixed_a(-0.000222287853830494)),(to_sfixed_a(0.00013699931150767952)),(to_sfixed_a(-2.2236226868699305e-05)),(to_sfixed_a(-0.00032409370760433376)),(to_sfixed_a(-0.00012587924720719457)),(to_sfixed_a(-9.917958959704265e-05)),(to_sfixed_a(6.295085040619597e-05)),(to_sfixed_a(5.587925625150092e-05)),(to_sfixed_a(3.4214146580779925e-05)),(to_sfixed_a(-0.00018148777598980814)),(to_sfixed_a(0.006907588802278042)),(to_sfixed_a(-0.00011147913028253242)),(to_sfixed_a(0.007789220195263624)),(to_sfixed_a(0.16116482019424438)),(to_sfixed_a(0.03712513670325279)),(to_sfixed_a(0.010274265892803669)),(to_sfixed_a(0.03774411976337433)),(to_sfixed_a(0.028034484013915062)),(to_sfixed_a(-0.002628721296787262)),(to_sfixed_a(0.29004761576652527)),(to_sfixed_a(0.03272704780101776)),(to_sfixed_a(-0.08132384717464447)),(to_sfixed_a(-0.040871504694223404)),(to_sfixed_a(-0.08281077444553375)),(to_sfixed_a(-6.228881102288142e-05)),(to_sfixed_a(3.6527737847791286e-06)),(to_sfixed_a(0.00018716974591370672)),(to_sfixed_a(-2.3490827516070567e-05)),(to_sfixed_a(-9.245728142559528e-05)),(to_sfixed_a(0.00013312780356500298)),(to_sfixed_a(-9.518479055259377e-05)),(to_sfixed_a(-2.7287993361824192e-05)),(to_sfixed_a(3.5559069146984257e-06)),(to_sfixed_a(0.00028675489011220634)),(to_sfixed_a(-5.096746463095769e-05)),(to_sfixed_a(-8.322126814164221e-05)),(to_sfixed_a(0.00021048150665592402)),(to_sfixed_a(0.0817185491323471)),(to_sfixed_a(-0.01126138400286436)),(to_sfixed_a(0.013307121582329273)),(to_sfixed_a(-0.5988447070121765)),(to_sfixed_a(0.2082771211862564)),(to_sfixed_a(0.02318062260746956)),(to_sfixed_a(0.3021210730075836)),(to_sfixed_a(0.29588234424591064)),(to_sfixed_a(0.2995806336402893)),(to_sfixed_a(0.15812626481056213)),(to_sfixed_a(-0.33729761838912964)),(to_sfixed_a(-0.2568790316581726)),(to_sfixed_a(-0.054900918155908585)),(to_sfixed_a(0.012100842781364918)),(to_sfixed_a(-0.2996458411216736)),(to_sfixed_a(0.013808735646307468)),(to_sfixed_a(0.00015889581118244678)),(to_sfixed_a(-0.0012697090860456228)),(to_sfixed_a(3.3078715205192566e-05)),(to_sfixed_a(-9.994328866014257e-05)),(to_sfixed_a(-2.6941930627799593e-05)),(to_sfixed_a(-8.944082946982235e-05)),(to_sfixed_a(0.00012525836064014584)),(to_sfixed_a(0.0001004336736514233)),(to_sfixed_a(-0.00024536080309189856)),(to_sfixed_a(-0.0017802607035264373)),(to_sfixed_a(0.11910706758499146)),(to_sfixed_a(-2.397886191829457e-07)),(to_sfixed_a(0.13800089061260223)),(to_sfixed_a(0.15229538083076477)),(to_sfixed_a(-0.19284044206142426)),(to_sfixed_a(-0.23307475447654724)),(to_sfixed_a(0.14301356673240662)),(to_sfixed_a(0.36907291412353516)),(to_sfixed_a(0.39476606249809265)),(to_sfixed_a(0.21152247488498688)),(to_sfixed_a(0.44103628396987915)),(to_sfixed_a(0.09835170954465866)),(to_sfixed_a(-0.17218372225761414)),(to_sfixed_a(-0.2445690780878067)),(to_sfixed_a(0.1104075089097023)),(to_sfixed_a(0.025327453389763832)),(to_sfixed_a(0.02830309420824051)),(to_sfixed_a(-0.00045774245518259704)),(to_sfixed_a(-0.052202705293893814)),(to_sfixed_a(-0.0018646372482180595)),(to_sfixed_a(-0.00034637239878065884)),(to_sfixed_a(4.089579306310043e-05)),(to_sfixed_a(-0.00013374752597883344)),(to_sfixed_a(0.00010764309263322502)),(to_sfixed_a(7.70422411733307e-05)),(to_sfixed_a(0.00015572491975035518)),(to_sfixed_a(-9.592405695002526e-05)),(to_sfixed_a(-0.0006044666515663266)),(to_sfixed_a(0.11637944728136063)),(to_sfixed_a(0.0564689002931118)),(to_sfixed_a(-0.2872686982154846)),(to_sfixed_a(-0.5537518262863159)),(to_sfixed_a(-0.46845221519470215)),(to_sfixed_a(-0.028392262756824493)),(to_sfixed_a(0.03858570754528046)),(to_sfixed_a(0.29772770404815674)),(to_sfixed_a(0.4164024889469147)),(to_sfixed_a(0.4448007643222809)),(to_sfixed_a(0.2832200825214386)),(to_sfixed_a(-0.16454598307609558)),(to_sfixed_a(-0.19174017012119293)),(to_sfixed_a(-0.312639981508255)),(to_sfixed_a(-0.13699765503406525)),(to_sfixed_a(-0.27575576305389404)),(to_sfixed_a(0.033260881900787354)),(to_sfixed_a(0.3035152554512024)),(to_sfixed_a(0.33105480670928955)),(to_sfixed_a(0.00013775276602245867)),(to_sfixed_a(8.560645073885098e-05)),(to_sfixed_a(0.0005348548293113708)),(to_sfixed_a(3.673411129057058e-06)),(to_sfixed_a(0.00019716167298611253)),(to_sfixed_a(0.0001475809986004606)),(to_sfixed_a(-0.00014764844672754407)),(to_sfixed_a(-0.00019262525893282145)),(to_sfixed_a(-0.00022571250156033784)),(to_sfixed_a(-0.012606301344931126)),(to_sfixed_a(-0.013916922733187675)),(to_sfixed_a(-0.045500498265028)),(to_sfixed_a(-0.4186767637729645)),(to_sfixed_a(-0.022625651210546494)),(to_sfixed_a(-0.17282602190971375)),(to_sfixed_a(0.31978726387023926)),(to_sfixed_a(0.26724934577941895)),(to_sfixed_a(0.7020347714424133)),(to_sfixed_a(0.5072035789489746)),(to_sfixed_a(-0.049383606761693954)),(to_sfixed_a(-0.16264621913433075)),(to_sfixed_a(-0.24455192685127258)),(to_sfixed_a(0.026792369782924652)),(to_sfixed_a(-0.07405406981706619)),(to_sfixed_a(-0.16698682308197021)),(to_sfixed_a(0.054979875683784485)),(to_sfixed_a(0.012522786855697632)),(to_sfixed_a(0.15194964408874512)),(to_sfixed_a(0.04954303428530693)),(to_sfixed_a(0.001311011495999992)),(to_sfixed_a(-3.9469330658903345e-05)),(to_sfixed_a(9.228581802744884e-06)),(to_sfixed_a(-4.423040445544757e-05)),(to_sfixed_a(-0.0002127340849256143)),(to_sfixed_a(2.384052459092345e-05)),(to_sfixed_a(-1.8995282516698353e-05)),(to_sfixed_a(-0.028383951634168625)),(to_sfixed_a(-0.1613880842924118)),(to_sfixed_a(-0.10846884548664093)),(to_sfixed_a(-0.1873386651277542)),(to_sfixed_a(-0.5271762609481812)),(to_sfixed_a(-0.3254018723964691)),(to_sfixed_a(-0.1967001110315323)),(to_sfixed_a(-0.0374416820704937)),(to_sfixed_a(0.015377922914922237)),(to_sfixed_a(0.4184104800224304)),(to_sfixed_a(0.34765225648880005)),(to_sfixed_a(-0.05586320534348488)),(to_sfixed_a(-0.2924375534057617)),(to_sfixed_a(-0.24926410615444183)),(to_sfixed_a(-0.19623620808124542)),(to_sfixed_a(-0.1533878892660141)),(to_sfixed_a(-0.10737854242324829)),(to_sfixed_a(0.1965663582086563)),(to_sfixed_a(0.0028193993493914604)),(to_sfixed_a(-0.056390926241874695)),(to_sfixed_a(0.038096919655799866)),(to_sfixed_a(0.025724926963448524)),(to_sfixed_a(2.151534999939031e-06)),(to_sfixed_a(0.00032367228413932025)),(to_sfixed_a(8.491174230584875e-05)),(to_sfixed_a(-1.35143664010684e-05)),(to_sfixed_a(2.8490783734014258e-05)),(to_sfixed_a(0.0005260472535155714)),(to_sfixed_a(0.0004516408662311733)),(to_sfixed_a(0.004869373980909586)),(to_sfixed_a(0.04530596733093262)),(to_sfixed_a(-0.135306254029274)),(to_sfixed_a(-0.24131062626838684)),(to_sfixed_a(-0.34315401315689087)),(to_sfixed_a(-0.5664849877357483)),(to_sfixed_a(-0.38531726598739624)),(to_sfixed_a(-0.3386123478412628)),(to_sfixed_a(0.09533660113811493)),(to_sfixed_a(0.4599137604236603)),(to_sfixed_a(0.0879586786031723)),(to_sfixed_a(-0.032901741564273834)),(to_sfixed_a(0.3012137711048126)),(to_sfixed_a(0.3274075984954834)),(to_sfixed_a(0.3358830511569977)),(to_sfixed_a(0.3173236846923828)),(to_sfixed_a(0.32844609022140503)),(to_sfixed_a(0.171473428606987)),(to_sfixed_a(0.2468927800655365)),(to_sfixed_a(0.13880325853824615)),(to_sfixed_a(4.354469638201408e-05)),(to_sfixed_a(7.129992445698008e-05)),(to_sfixed_a(-5.823604624310974e-06)),(to_sfixed_a(0.00029615004314109683)),(to_sfixed_a(7.459214248228818e-05)),(to_sfixed_a(-0.00017313534044660628)),(to_sfixed_a(0.0002741178614087403)),(to_sfixed_a(0.0036392132751643658)),(to_sfixed_a(-0.06143615022301674)),(to_sfixed_a(-0.277217298746109)),(to_sfixed_a(-0.342950701713562)),(to_sfixed_a(-0.4656330645084381)),(to_sfixed_a(-0.8907003998756409)),(to_sfixed_a(-0.8033604025840759)),(to_sfixed_a(-0.7809858918190002)),(to_sfixed_a(-0.32106268405914307)),(to_sfixed_a(0.20942150056362152)),(to_sfixed_a(0.39309176802635193)),(to_sfixed_a(0.010353874415159225)),(to_sfixed_a(-0.22452332079410553)),(to_sfixed_a(-0.1496959924697876)),(to_sfixed_a(0.3457874655723572)),(to_sfixed_a(0.4806446433067322)),(to_sfixed_a(0.37790554761886597)),(to_sfixed_a(0.3158530592918396)),(to_sfixed_a(0.34449371695518494)),(to_sfixed_a(0.15316538512706757)),(to_sfixed_a(0.07423713803291321)),(to_sfixed_a(0.012573955580592155)),(to_sfixed_a(-8.379917562706396e-05)),(to_sfixed_a(4.3214178731432185e-05)),(to_sfixed_a(-0.00011155472748214379)),(to_sfixed_a(-1.4731349438079633e-05)),(to_sfixed_a(0.00014214350085239857)),(to_sfixed_a(0.02817424200475216)),(to_sfixed_a(-0.08156860619783401)),(to_sfixed_a(-0.22895756363868713)),(to_sfixed_a(-0.3570556640625)),(to_sfixed_a(-0.3321892023086548)),(to_sfixed_a(-0.30957603454589844)),(to_sfixed_a(-0.2946203351020813)),(to_sfixed_a(0.022268330678343773)),(to_sfixed_a(0.12044715136289597)),(to_sfixed_a(0.26170653104782104)),(to_sfixed_a(0.09511690586805344)),(to_sfixed_a(0.17312508821487427)),(to_sfixed_a(-0.04053167626261711)),(to_sfixed_a(-0.04968196526169777)),(to_sfixed_a(-0.0488334521651268)),(to_sfixed_a(0.22592386603355408)),(to_sfixed_a(0.24440321326255798)),(to_sfixed_a(0.0906311497092247)),(to_sfixed_a(0.011219422332942486)),(to_sfixed_a(0.11949530988931656)),(to_sfixed_a(0.2980339825153351)),(to_sfixed_a(0.17231881618499756)),(to_sfixed_a(-2.3012456949800253e-05)),(to_sfixed_a(0.00014761851343791932)),(to_sfixed_a(0.00021518937137443572)),(to_sfixed_a(5.6773031246848404e-05)),(to_sfixed_a(9.484906331636012e-05)),(to_sfixed_a(7.173137419158593e-05)),(to_sfixed_a(7.258597906911746e-05)),(to_sfixed_a(0.041923705488443375)),(to_sfixed_a(-0.07641243934631348)),(to_sfixed_a(-0.15285241603851318)),(to_sfixed_a(0.08476956188678741)),(to_sfixed_a(0.13825492560863495)),(to_sfixed_a(0.07041645795106888)),(to_sfixed_a(0.3557383120059967)),(to_sfixed_a(0.3407164514064789)),(to_sfixed_a(0.7196459174156189)),(to_sfixed_a(0.5156542062759399)),(to_sfixed_a(0.26099249720573425)),(to_sfixed_a(0.05676611140370369)),(to_sfixed_a(0.007071299012750387)),(to_sfixed_a(-0.21691718697547913)),(to_sfixed_a(-0.13803833723068237)),(to_sfixed_a(0.17416605353355408)),(to_sfixed_a(-0.00410766527056694)),(to_sfixed_a(0.0637449398636818)),(to_sfixed_a(0.10472021251916885)),(to_sfixed_a(-0.05294756218791008)),(to_sfixed_a(-0.016746867448091507)),(to_sfixed_a(0.00010691594798117876)),(to_sfixed_a(-0.0001049134079948999)),(to_sfixed_a(7.501566869905218e-05)),(to_sfixed_a(-7.208478200482205e-05)),(to_sfixed_a(0.00020379443594720215)),(to_sfixed_a(8.662130130687729e-05)),(to_sfixed_a(0.00015840416017454118)),(to_sfixed_a(-0.00949887651950121)),(to_sfixed_a(-0.12314584851264954)),(to_sfixed_a(0.008110626600682735)),(to_sfixed_a(0.2875392735004425)),(to_sfixed_a(0.021064141765236855)),(to_sfixed_a(0.21081222593784332)),(to_sfixed_a(0.28566092252731323)),(to_sfixed_a(0.3492269515991211)),(to_sfixed_a(0.289195716381073)),(to_sfixed_a(0.41440144181251526)),(to_sfixed_a(0.17119145393371582)),(to_sfixed_a(-0.10953123867511749)),(to_sfixed_a(0.001420157845132053)),(to_sfixed_a(-0.1810631901025772)),(to_sfixed_a(-0.03253709524869919)),(to_sfixed_a(-0.08958691358566284)),(to_sfixed_a(0.03499028831720352)),(to_sfixed_a(0.000391782057704404)),(to_sfixed_a(-0.06036143749952316)),(to_sfixed_a(-0.16716432571411133)),(to_sfixed_a(0.006383569911122322)),(to_sfixed_a(-0.0029483328107744455)),(to_sfixed_a(-0.0014680592576041818)),(to_sfixed_a(-0.0001674196100793779)),(to_sfixed_a(-0.00014304605429060757)),(to_sfixed_a(-0.00018335445201955736)),(to_sfixed_a(0.0002437657822156325)),(to_sfixed_a(-6.130198016762733e-05)),(to_sfixed_a(0.0025576187763363123)),(to_sfixed_a(-0.03377417474985123)),(to_sfixed_a(0.0662437379360199)),(to_sfixed_a(0.04872327670454979)),(to_sfixed_a(0.15747615694999695)),(to_sfixed_a(0.20010758936405182)),(to_sfixed_a(-0.025788625702261925)),(to_sfixed_a(-0.13572609424591064)),(to_sfixed_a(0.08412634581327438)),(to_sfixed_a(0.3264017105102539)),(to_sfixed_a(0.07457727938890457)),(to_sfixed_a(-0.04261104762554169)),(to_sfixed_a(-0.03791337087750435)),(to_sfixed_a(-0.11099500209093094)),(to_sfixed_a(-0.254379004240036)),(to_sfixed_a(-0.27733272314071655)),(to_sfixed_a(-0.1370367556810379)),(to_sfixed_a(0.04488052427768707)),(to_sfixed_a(0.013692094013094902)),(to_sfixed_a(-0.06386180222034454)),(to_sfixed_a(-0.08228959143161774)),(to_sfixed_a(0.0001156088401330635)),(to_sfixed_a(-6.79361037327908e-05)),(to_sfixed_a(-0.00023362782667391002)),(to_sfixed_a(-0.00018458654813002795)),(to_sfixed_a(-0.000212126033147797)),(to_sfixed_a(-2.8447660952224396e-05)),(to_sfixed_a(-0.00027071262593381107)),(to_sfixed_a(-0.01382340770214796)),(to_sfixed_a(-0.034897733479738235)),(to_sfixed_a(-0.18377673625946045)),(to_sfixed_a(-0.39208507537841797)),(to_sfixed_a(-0.4290488660335541)),(to_sfixed_a(-0.42067548632621765)),(to_sfixed_a(-0.39280831813812256)),(to_sfixed_a(-0.0283208005130291)),(to_sfixed_a(0.1566978394985199)),(to_sfixed_a(0.18677304685115814)),(to_sfixed_a(0.0035469799768179655)),(to_sfixed_a(-0.05691495165228844)),(to_sfixed_a(-0.021019725129008293)),(to_sfixed_a(-0.3377007842063904)),(to_sfixed_a(-0.20932894945144653)),(to_sfixed_a(-0.2767668068408966)),(to_sfixed_a(-0.3352068066596985)),(to_sfixed_a(-0.07878590375185013)),(to_sfixed_a(-0.13719329237937927)),(to_sfixed_a(0.08163312822580338)),(to_sfixed_a(0.01956363581120968)),(to_sfixed_a(0.00047552440082654357)),(to_sfixed_a(-1.08168069345993e-06)),(to_sfixed_a(0.00013290120114106685)),(to_sfixed_a(-7.19031595508568e-05)),(to_sfixed_a(-0.00017604295862838626)),(to_sfixed_a(-0.0005080262199044228)),(to_sfixed_a(-0.004301921464502811)),(to_sfixed_a(0.018253007903695107)),(to_sfixed_a(-0.03297989070415497)),(to_sfixed_a(-0.3032784163951874)),(to_sfixed_a(-0.25269490480422974)),(to_sfixed_a(-0.3114909827709198)),(to_sfixed_a(-0.3832527697086334)),(to_sfixed_a(-0.33403775095939636)),(to_sfixed_a(-0.3764675259590149)),(to_sfixed_a(-0.12299548834562302)),(to_sfixed_a(-0.2239801287651062)),(to_sfixed_a(-0.020399386063218117)),(to_sfixed_a(-0.09887152165174484)),(to_sfixed_a(0.006390768103301525)),(to_sfixed_a(-0.1362125724554062)),(to_sfixed_a(-0.04713362455368042)),(to_sfixed_a(-0.16562685370445251)),(to_sfixed_a(-0.31346943974494934)),(to_sfixed_a(-0.17833948135375977)),(to_sfixed_a(-0.07821281254291534)),(to_sfixed_a(0.031121963635087013)),(to_sfixed_a(-0.0003775997320190072)),(to_sfixed_a(-0.008348776958882809)),(to_sfixed_a(9.795738878892735e-05)),(to_sfixed_a(-3.9779428334441036e-05)),(to_sfixed_a(-3.0165621865307912e-05)),(to_sfixed_a(-7.313026435440406e-05)),(to_sfixed_a(-0.003091531340032816)),(to_sfixed_a(-0.004368796478956938)),(to_sfixed_a(0.05834272876381874)),(to_sfixed_a(-0.052444275468587875)),(to_sfixed_a(-0.16461093723773956)),(to_sfixed_a(-0.41981497406959534)),(to_sfixed_a(-0.39168524742126465)),(to_sfixed_a(-0.2556931674480438)),(to_sfixed_a(-0.2817992866039276)),(to_sfixed_a(-0.21951040625572205)),(to_sfixed_a(-0.1038510650396347)),(to_sfixed_a(-0.25185999274253845)),(to_sfixed_a(-0.20057746767997742)),(to_sfixed_a(-0.012861013412475586)),(to_sfixed_a(-0.1972108632326126)),(to_sfixed_a(-0.17939479649066925)),(to_sfixed_a(-0.07499968260526657)),(to_sfixed_a(0.015916112810373306)),(to_sfixed_a(-0.08702737092971802)),(to_sfixed_a(-0.05821675434708595)),(to_sfixed_a(-0.12621362507343292)),(to_sfixed_a(0.01223091408610344)),(to_sfixed_a(8.829708531266078e-05)),(to_sfixed_a(-0.00020546004816424102)),(to_sfixed_a(-0.00015690909640397877)),(to_sfixed_a(7.705471944063902e-05)),(to_sfixed_a(0.00010852582636289299)),(to_sfixed_a(9.842812687566038e-06)),(to_sfixed_a(-0.00010756112169474363)),(to_sfixed_a(-0.024992570281028748)),(to_sfixed_a(-0.010601385496556759)),(to_sfixed_a(-0.12541373074054718)),(to_sfixed_a(0.13420720398426056)),(to_sfixed_a(0.08924365043640137)),(to_sfixed_a(0.0030241275671869516)),(to_sfixed_a(-0.07521340250968933)),(to_sfixed_a(-0.023056041449308395)),(to_sfixed_a(0.18028096854686737)),(to_sfixed_a(0.046131595969200134)),(to_sfixed_a(0.026459142565727234)),(to_sfixed_a(-0.14334595203399658)),(to_sfixed_a(-0.15103782713413239)),(to_sfixed_a(-0.052779775112867355)),(to_sfixed_a(0.05114230513572693)),(to_sfixed_a(-0.03598886728286743)),(to_sfixed_a(-0.13955625891685486)),(to_sfixed_a(-0.08840282261371613)),(to_sfixed_a(-0.31444859504699707)),(to_sfixed_a(0.08054269850254059)),(to_sfixed_a(0.022464998066425323)),(to_sfixed_a(-0.02157719060778618)),(to_sfixed_a(-0.0001182173436973244)),(to_sfixed_a(0.0002224157942691818)),(to_sfixed_a(0.00013499327178578824)),(to_sfixed_a(0.0001653452345635742)),(to_sfixed_a(2.6975876608048566e-05)),(to_sfixed_a(0.00029764900682494044)),(to_sfixed_a(0.11883673816919327)),(to_sfixed_a(0.0014637401327490807)),(to_sfixed_a(0.14859138429164886)),(to_sfixed_a(0.004100314807146788)),(to_sfixed_a(0.1419575959444046)),(to_sfixed_a(0.3499457836151123)),(to_sfixed_a(0.47355496883392334)),(to_sfixed_a(0.5554585456848145)),(to_sfixed_a(0.500778317451477)),(to_sfixed_a(0.11115308105945587)),(to_sfixed_a(-0.02454819157719612)),(to_sfixed_a(-0.21018587052822113)),(to_sfixed_a(-0.10345666855573654)),(to_sfixed_a(0.06029509752988815)),(to_sfixed_a(0.07290593534708023)),(to_sfixed_a(-0.05496659874916077)),(to_sfixed_a(-0.040491633117198944)),(to_sfixed_a(-0.11584043502807617)),(to_sfixed_a(-0.22380158305168152)),(to_sfixed_a(0.009037981741130352)),(to_sfixed_a(0.14280813932418823)),(to_sfixed_a(-0.00021264680253807455)),(to_sfixed_a(0.00021808876772411168)),(to_sfixed_a(5.038256131228991e-05)),(to_sfixed_a(6.328007293632254e-05)),(to_sfixed_a(-0.00010033968283096328)),(to_sfixed_a(-0.00017161430150736123)),(to_sfixed_a(0.00012098121078452095)),(to_sfixed_a(-0.0001327422505710274)),(to_sfixed_a(0.005759736057370901)),(to_sfixed_a(-0.09818597882986069)),(to_sfixed_a(0.19218452274799347)),(to_sfixed_a(-0.03855369985103607)),(to_sfixed_a(0.16681616008281708)),(to_sfixed_a(0.25852710008621216)),(to_sfixed_a(0.20725196599960327)),(to_sfixed_a(0.4221634268760681)),(to_sfixed_a(0.6437061429023743)),(to_sfixed_a(0.07019469141960144)),(to_sfixed_a(0.09786750376224518)),(to_sfixed_a(-0.2150007039308548)),(to_sfixed_a(-0.01034192182123661)),(to_sfixed_a(0.04421096667647362)),(to_sfixed_a(-0.03338940441608429)),(to_sfixed_a(-0.12260360270738602)),(to_sfixed_a(-0.1544676125049591)),(to_sfixed_a(-0.09450546652078629)),(to_sfixed_a(0.059115100651979446)),(to_sfixed_a(0.015761632472276688)),(to_sfixed_a(-0.0443238839507103)),(to_sfixed_a(0.00017971242778003216)),(to_sfixed_a(0.00011729358811862767)),(to_sfixed_a(7.783316686982289e-05)),(to_sfixed_a(0.00010151378228329122)),(to_sfixed_a(0.00018537003779783845)),(to_sfixed_a(0.00019654854258988053)),(to_sfixed_a(-7.655958324903622e-05)),(to_sfixed_a(-0.0403573177754879)),(to_sfixed_a(0.0006527399527840316)),(to_sfixed_a(0.11424650251865387)),(to_sfixed_a(0.03732510283589363)),(to_sfixed_a(0.28842201828956604)),(to_sfixed_a(0.17073263227939606)),(to_sfixed_a(0.03694659471511841)),(to_sfixed_a(0.2407216578722)),(to_sfixed_a(0.1214291900396347)),(to_sfixed_a(0.2224152386188507)),(to_sfixed_a(0.21740323305130005)),(to_sfixed_a(0.169432133436203)),(to_sfixed_a(-0.01720050349831581)),(to_sfixed_a(-0.11280380189418793)),(to_sfixed_a(-0.167866051197052)),(to_sfixed_a(-0.12481288611888885)),(to_sfixed_a(0.05252351611852646)),(to_sfixed_a(0.036602746695280075)),(to_sfixed_a(0.10201902687549591)),(to_sfixed_a(0.0006508406950160861)),(to_sfixed_a(0.0033166727516800165)),(to_sfixed_a(-0.0001271173096029088)),(to_sfixed_a(-0.0001428963296348229)),(to_sfixed_a(-6.442003359552473e-05)),(to_sfixed_a(9.117544686887413e-05)),(to_sfixed_a(0.00011348298721713945)),(to_sfixed_a(4.191010884824209e-05)),(to_sfixed_a(0.0002676969161257148)),(to_sfixed_a(0.0003170620184391737)),(to_sfixed_a(0.05765247344970703)),(to_sfixed_a(0.026974590495228767)),(to_sfixed_a(-0.08262206614017487)),(to_sfixed_a(0.041770514100790024)),(to_sfixed_a(0.029049767181277275)),(to_sfixed_a(0.11276302486658096)),(to_sfixed_a(0.011141642928123474)),(to_sfixed_a(0.1415920853614807)),(to_sfixed_a(0.14220720529556274)),(to_sfixed_a(0.02640020288527012)),(to_sfixed_a(-0.08321323245763779)),(to_sfixed_a(0.0004144422127865255)),(to_sfixed_a(-0.09216775000095367)),(to_sfixed_a(-0.1573190689086914)),(to_sfixed_a(-0.05823371186852455)),(to_sfixed_a(0.02661173604428768)),(to_sfixed_a(0.01623767614364624)),(to_sfixed_a(0.014208945445716381)),(to_sfixed_a(-0.0009426442557014525)),(to_sfixed_a(8.617995626991615e-05)),(to_sfixed_a(-2.4320117518072948e-05)),(to_sfixed_a(-3.2293512049363926e-05)),(to_sfixed_a(2.9516479116864502e-05)),(to_sfixed_a(-4.421867924975231e-05)),(to_sfixed_a(0.00010430523252580315)),(to_sfixed_a(0.00011339634511386976)),(to_sfixed_a(0.0001923446252476424)),(to_sfixed_a(0.0003223238745704293)),(to_sfixed_a(-0.020347684621810913)),(to_sfixed_a(0.04256894439458847)),(to_sfixed_a(-0.03311355412006378)),(to_sfixed_a(0.270630806684494)),(to_sfixed_a(0.11499390006065369)),(to_sfixed_a(0.09887140244245529)),(to_sfixed_a(0.18346068263053894)),(to_sfixed_a(0.21349062025547028)),(to_sfixed_a(0.12792138755321503)),(to_sfixed_a(0.021981768310070038)),(to_sfixed_a(0.028670087456703186)),(to_sfixed_a(-0.1654846966266632)),(to_sfixed_a(0.13195009529590607)),(to_sfixed_a(-0.011870761401951313)),(to_sfixed_a(-0.05857829749584198)),(to_sfixed_a(-0.010058330371975899)),(to_sfixed_a(-0.0026149435434490442)),(to_sfixed_a(0.0018717956263571978)),(to_sfixed_a(-0.0028636003844439983)),(to_sfixed_a(4.971984162693843e-05)),(to_sfixed_a(0.0002141716395271942)),(to_sfixed_a(-9.090201638173312e-05)),(to_sfixed_a(-9.833845251705498e-05)),(to_sfixed_a(2.966773899970576e-05)),(to_sfixed_a(-0.00011593438102863729)),(to_sfixed_a(-0.0001467390829930082)),(to_sfixed_a(-6.200699863256887e-05)),(to_sfixed_a(-0.010717455297708511)),(to_sfixed_a(0.0009901040466502309)),(to_sfixed_a(-0.044525764882564545)),(to_sfixed_a(-0.11448167264461517)),(to_sfixed_a(0.09331724047660828)),(to_sfixed_a(0.003933391533792019)),(to_sfixed_a(-0.15737248957157135)),(to_sfixed_a(0.18518966436386108)),(to_sfixed_a(-0.01735365204513073)),(to_sfixed_a(-0.0581195168197155)),(to_sfixed_a(0.037312328815460205)),(to_sfixed_a(-0.02068439871072769)),(to_sfixed_a(-0.20038630068302155)),(to_sfixed_a(-0.19508406519889832)),(to_sfixed_a(-0.020229022949934006)),(to_sfixed_a(-0.015347808599472046)),(to_sfixed_a(-0.0006531209801323712)),(to_sfixed_a(0.03336165100336075)),(to_sfixed_a(0.001606243778951466)),(to_sfixed_a(0.006993868388235569)),(to_sfixed_a(5.293890353641473e-05)),(to_sfixed_a(-0.00014274970453698188)),(to_sfixed_a(-4.142847501498181e-06)),(to_sfixed_a(-6.575903535122052e-05)),(to_sfixed_a(4.439146141521633e-05)),(to_sfixed_a(3.3690583222778514e-05)),(to_sfixed_a(-0.0002748899278230965)),(to_sfixed_a(2.472215965099167e-05)),(to_sfixed_a(-0.0001334729604423046)),(to_sfixed_a(-0.032012030482292175)),(to_sfixed_a(-0.026657385751605034)),(to_sfixed_a(-0.11749137192964554)),(to_sfixed_a(-0.08695296198129654)),(to_sfixed_a(0.029635637998580933)),(to_sfixed_a(0.020827200263738632)),(to_sfixed_a(-0.019696572795510292)),(to_sfixed_a(-0.08824504911899567)),(to_sfixed_a(-0.13633807003498077)),(to_sfixed_a(-0.06322069466114044)),(to_sfixed_a(0.019946828484535217)),(to_sfixed_a(-0.1374737024307251)),(to_sfixed_a(-0.027765441685914993)),(to_sfixed_a(0.008717759512364864)),(to_sfixed_a(-0.010994741693139076)),(to_sfixed_a(0.18472379446029663)),(to_sfixed_a(0.0007211664924398065)),(to_sfixed_a(0.002532368991523981)),(to_sfixed_a(0.0032362458296120167)),(to_sfixed_a(-8.584505849285051e-05)),(to_sfixed_a(3.1944222428137437e-05)),(to_sfixed_a(2.6128678655368276e-05)),(to_sfixed_a(1.4163410014589317e-05)),(to_sfixed_a(5.5129770771600306e-05)),(to_sfixed_a(-0.0001864587829913944)),(to_sfixed_a(-4.076805635122582e-05)),(to_sfixed_a(0.00018479360733181238)),(to_sfixed_a(-5.647914076689631e-05)),(to_sfixed_a(0.0008601979352533817)),(to_sfixed_a(0.0007414942374452949)),(to_sfixed_a(0.00013712537474930286)),(to_sfixed_a(7.890420420153532e-06)),(to_sfixed_a(0.0005760134081356227)),(to_sfixed_a(-0.04998370260000229)),(to_sfixed_a(0.008272337727248669)),(to_sfixed_a(0.0006302589317783713)),(to_sfixed_a(-0.05321749299764633)),(to_sfixed_a(-0.08778636157512665)),(to_sfixed_a(-0.015724467113614082)),(to_sfixed_a(-0.0058187199756503105)),(to_sfixed_a(-0.04444893077015877)),(to_sfixed_a(-0.05465426295995712)),(to_sfixed_a(0.005368019919842482)),(to_sfixed_a(0.002926150569692254)),(to_sfixed_a(7.706048199906945e-05)),(to_sfixed_a(1.615869769011624e-05)),(to_sfixed_a(-7.42625561542809e-05)),(to_sfixed_a(7.277143140527187e-06)),(to_sfixed_a(-2.501397284504492e-05)),(to_sfixed_a(5.073900683782995e-05)),(to_sfixed_a(-0.0003033427055925131)),(to_sfixed_a(0.00013931706780567765)),(to_sfixed_a(2.0669062905653846e-06)),(to_sfixed_a(5.816919292556122e-05)),(to_sfixed_a(-6.882168577249104e-07)),(to_sfixed_a(0.00012424511078279465)),(to_sfixed_a(0.00023461320961359888)),(to_sfixed_a(4.6883833419997245e-05)),(to_sfixed_a(0.00014508231834042817)),(to_sfixed_a(-6.691214366583154e-05)),(to_sfixed_a(-0.00039422494592145085)),(to_sfixed_a(-0.00010085824033012614)),(to_sfixed_a(4.576351784635335e-05)),(to_sfixed_a(0.00019451466505415738)),(to_sfixed_a(0.0001656607782933861)),(to_sfixed_a(-4.5895907533122227e-05)),(to_sfixed_a(-8.351868018507957e-05)),(to_sfixed_a(0.00013263979053590447)),(to_sfixed_a(-2.181807576562278e-05)),(to_sfixed_a(2.735757880145684e-05)),(to_sfixed_a(0.0003217394696548581)),(to_sfixed_a(0.00015724643890280277)),(to_sfixed_a(3.0877972676535137e-06)),(to_sfixed_a(-0.00010828946687979624)),(to_sfixed_a(4.5048062020214275e-05)),(to_sfixed_a(4.063676533405669e-05)),(to_sfixed_a(8.510494080837816e-05)),(to_sfixed_a(6.31449802313e-05)),(to_sfixed_a(-0.00013282512372825295)));

    constant weight_n0_6 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(3.0395709472941235e-05)),(to_sfixed_a(-8.95069824764505e-05)),(to_sfixed_a(0.000274300662567839)),(to_sfixed_a(0.00025640931562520564)),(to_sfixed_a(-0.000217588254599832)),(to_sfixed_a(0.00017481284157838672)),(to_sfixed_a(0.0001607134036021307)),(to_sfixed_a(-0.00018224109953735024)),(to_sfixed_a(8.135809184750542e-05)),(to_sfixed_a(-0.0002142704470315948)),(to_sfixed_a(-0.00011403766256989911)),(to_sfixed_a(0.00021327940339688212)),(to_sfixed_a(-9.027728083310649e-05)),(to_sfixed_a(6.546192889800295e-05)),(to_sfixed_a(-1.3197481166571379e-05)),(to_sfixed_a(0.00011255548452027142)),(to_sfixed_a(-0.0003237272903788835)),(to_sfixed_a(0.0003945560602005571)),(to_sfixed_a(0.00025398738216608763)),(to_sfixed_a(-0.0001403731876052916)),(to_sfixed_a(-3.847212792607024e-05)),(to_sfixed_a(0.0002200876479037106)),(to_sfixed_a(1.8851153072318994e-05)),(to_sfixed_a(3.369141631992534e-05)),(to_sfixed_a(2.3402570150210522e-05)),(to_sfixed_a(9.911793767969357e-07)),(to_sfixed_a(-0.0001016769529087469)),(to_sfixed_a(3.389867197256535e-05)),(to_sfixed_a(9.6303949248977e-05)),(to_sfixed_a(5.005598359275609e-05)),(to_sfixed_a(-0.00013752171071246266)),(to_sfixed_a(8.074272045632824e-05)),(to_sfixed_a(-0.00015439536946360022)),(to_sfixed_a(3.2238134735962376e-05)),(to_sfixed_a(0.00015661980432923883)),(to_sfixed_a(0.00020457922073546797)),(to_sfixed_a(1.3348966604098678e-05)),(to_sfixed_a(-1.4906309843354393e-05)),(to_sfixed_a(-4.192988490103744e-05)),(to_sfixed_a(-5.976479224045761e-05)),(to_sfixed_a(0.000103439437225461)),(to_sfixed_a(0.00033955968683585525)),(to_sfixed_a(-0.00011298764729872346)),(to_sfixed_a(0.00011104049190180376)),(to_sfixed_a(-1.443286510038888e-05)),(to_sfixed_a(0.00027643784414976835)),(to_sfixed_a(-0.00036402783007360995)),(to_sfixed_a(9.838202822720632e-05)),(to_sfixed_a(1.0960293366224505e-05)),(to_sfixed_a(4.4823095777246635e-06)),(to_sfixed_a(1.1837608326459303e-05)),(to_sfixed_a(7.271313370438293e-05)),(to_sfixed_a(0.0002182535972679034)),(to_sfixed_a(0.00032597320387139916)),(to_sfixed_a(-0.00012850819621235132)),(to_sfixed_a(-0.0002923424472101033)),(to_sfixed_a(0.00016220870020333678)),(to_sfixed_a(0.00015039087156765163)),(to_sfixed_a(6.144172220956534e-05)),(to_sfixed_a(0.00018525772611610591)),(to_sfixed_a(-0.0001605181023478508)),(to_sfixed_a(-3.4249122109031305e-05)),(to_sfixed_a(-8.90519550011959e-06)),(to_sfixed_a(-0.0001980162487598136)),(to_sfixed_a(-0.0001520555088063702)),(to_sfixed_a(-3.125102739431895e-05)),(to_sfixed_a(4.1795366996666417e-05)),(to_sfixed_a(6.0465365095296875e-05)),(to_sfixed_a(-6.24826570856385e-05)),(to_sfixed_a(0.006525924429297447)),(to_sfixed_a(-5.1521848945412785e-05)),(to_sfixed_a(-0.00022564164828509092)),(to_sfixed_a(-1.4240753444028087e-05)),(to_sfixed_a(-8.18444459582679e-05)),(to_sfixed_a(0.0001428911928087473)),(to_sfixed_a(0.0002563309681136161)),(to_sfixed_a(-4.018304753117263e-05)),(to_sfixed_a(-0.00021972488320898265)),(to_sfixed_a(-0.00026624943711794913)),(to_sfixed_a(-0.00031468659290112555)),(to_sfixed_a(0.0001323064643656835)),(to_sfixed_a(-9.301696991315112e-05)),(to_sfixed_a(-4.949167123413645e-05)),(to_sfixed_a(0.0002551699581090361)),(to_sfixed_a(-2.4168120944523253e-05)),(to_sfixed_a(0.00014379076310433447)),(to_sfixed_a(-0.00011066931620007381)),(to_sfixed_a(-8.44118621898815e-05)),(to_sfixed_a(0.00017795244639273733)),(to_sfixed_a(-8.437132055405527e-05)),(to_sfixed_a(1.8487751731299795e-05)),(to_sfixed_a(0.00018786959117278457)),(to_sfixed_a(0.01966591365635395)),(to_sfixed_a(1.8401365196041297e-06)),(to_sfixed_a(0.022080928087234497)),(to_sfixed_a(-0.07979941368103027)),(to_sfixed_a(0.05783900246024132)),(to_sfixed_a(-0.09577881544828415)),(to_sfixed_a(0.053074903786182404)),(to_sfixed_a(0.013761552050709724)),(to_sfixed_a(0.0065650129690766335)),(to_sfixed_a(-0.07014849036931992)),(to_sfixed_a(0.04154995083808899)),(to_sfixed_a(0.01540424395352602)),(to_sfixed_a(0.0019373540999367833)),(to_sfixed_a(0.003808088367804885)),(to_sfixed_a(1.297518792853225e-05)),(to_sfixed_a(0.0002411807217868045)),(to_sfixed_a(5.686611984856427e-06)),(to_sfixed_a(-0.0002480590483173728)),(to_sfixed_a(7.984180410858244e-05)),(to_sfixed_a(-0.00010879419278353453)),(to_sfixed_a(-8.761295248405077e-06)),(to_sfixed_a(-0.0001488486013840884)),(to_sfixed_a(-6.303624832071364e-05)),(to_sfixed_a(0.00014467042637988925)),(to_sfixed_a(-0.00020083793788217008)),(to_sfixed_a(3.0062290534260683e-05)),(to_sfixed_a(-0.00013311323709785938)),(to_sfixed_a(-0.045551642775535583)),(to_sfixed_a(0.08937850594520569)),(to_sfixed_a(0.022059326991438866)),(to_sfixed_a(-0.10845924913883209)),(to_sfixed_a(-0.03081672079861164)),(to_sfixed_a(-0.016226675361394882)),(to_sfixed_a(-0.06854758411645889)),(to_sfixed_a(-0.19377289712429047)),(to_sfixed_a(-0.07738149911165237)),(to_sfixed_a(-0.23249483108520508)),(to_sfixed_a(-0.18486294150352478)),(to_sfixed_a(-0.06369452178478241)),(to_sfixed_a(0.08444149047136307)),(to_sfixed_a(0.006569272838532925)),(to_sfixed_a(0.024347377941012383)),(to_sfixed_a(0.046863097697496414)),(to_sfixed_a(-0.0007911635329946876)),(to_sfixed_a(0.0008670171373523772)),(to_sfixed_a(1.5179771253315266e-05)),(to_sfixed_a(0.00017785267846193165)),(to_sfixed_a(0.0001802062470233068)),(to_sfixed_a(0.00011551205534487963)),(to_sfixed_a(-0.00010531464067753404)),(to_sfixed_a(9.177320862363558e-06)),(to_sfixed_a(-8.345975948031992e-05)),(to_sfixed_a(0.00016412511467933655)),(to_sfixed_a(-0.07521022111177444)),(to_sfixed_a(-0.008883114904165268)),(to_sfixed_a(-0.12290763109922409)),(to_sfixed_a(-0.06492313742637634)),(to_sfixed_a(0.0042696078307926655)),(to_sfixed_a(0.06381848454475403)),(to_sfixed_a(0.06471405923366547)),(to_sfixed_a(-0.18196791410446167)),(to_sfixed_a(-0.30427253246307373)),(to_sfixed_a(-0.12174597382545471)),(to_sfixed_a(-0.1464894413948059)),(to_sfixed_a(-0.07217787206172943)),(to_sfixed_a(-0.2952911853790283)),(to_sfixed_a(0.049318667501211166)),(to_sfixed_a(-0.13024906814098358)),(to_sfixed_a(0.1272583156824112)),(to_sfixed_a(0.04632310941815376)),(to_sfixed_a(0.0022314111702144146)),(to_sfixed_a(0.03746296837925911)),(to_sfixed_a(0.0013586065033450723)),(to_sfixed_a(-0.0003334882785566151)),(to_sfixed_a(-1.2998280908504967e-05)),(to_sfixed_a(-0.00015047818305902183)),(to_sfixed_a(0.00011571971845114604)),(to_sfixed_a(0.00032021975493989885)),(to_sfixed_a(0.00015474979591090232)),(to_sfixed_a(0.00016298021364491433)),(to_sfixed_a(0.00018138455925509334)),(to_sfixed_a(-0.07148797065019608)),(to_sfixed_a(-0.02378256618976593)),(to_sfixed_a(-0.12957637012004852)),(to_sfixed_a(-0.11172798275947571)),(to_sfixed_a(-0.2807255685329437)),(to_sfixed_a(-0.08213426917791367)),(to_sfixed_a(-0.004383102059364319)),(to_sfixed_a(0.0102931447327137)),(to_sfixed_a(0.0013681304408237338)),(to_sfixed_a(-0.12799832224845886)),(to_sfixed_a(-0.14002859592437744)),(to_sfixed_a(-0.18175584077835083)),(to_sfixed_a(-0.054825592786073685)),(to_sfixed_a(-0.11091817915439606)),(to_sfixed_a(-0.02016325481235981)),(to_sfixed_a(0.03274756669998169)),(to_sfixed_a(-0.07682155817747116)),(to_sfixed_a(0.06629350036382675)),(to_sfixed_a(-0.005873859394341707)),(to_sfixed_a(0.0009139921749010682)),(to_sfixed_a(0.0006640341016463935)),(to_sfixed_a(-0.0005587747436948121)),(to_sfixed_a(8.62807864905335e-05)),(to_sfixed_a(-0.0001604203716851771)),(to_sfixed_a(0.00014978795661590993)),(to_sfixed_a(2.20471356442431e-05)),(to_sfixed_a(5.5181015341077e-05)),(to_sfixed_a(-0.00011348248517606407)),(to_sfixed_a(0.026981797069311142)),(to_sfixed_a(0.07792846113443375)),(to_sfixed_a(0.03587159141898155)),(to_sfixed_a(-0.23161229491233826)),(to_sfixed_a(0.0801997184753418)),(to_sfixed_a(0.507469117641449)),(to_sfixed_a(0.12196832150220871)),(to_sfixed_a(0.2311597615480423)),(to_sfixed_a(0.09453552216291428)),(to_sfixed_a(-0.03274872899055481)),(to_sfixed_a(-0.06967086344957352)),(to_sfixed_a(-0.1370249092578888)),(to_sfixed_a(-0.0301347728818655)),(to_sfixed_a(-0.13097131252288818)),(to_sfixed_a(-0.10589928925037384)),(to_sfixed_a(0.07338853180408478)),(to_sfixed_a(0.035269297659397125)),(to_sfixed_a(0.12149418145418167)),(to_sfixed_a(0.018473105505108833)),(to_sfixed_a(0.03844580426812172)),(to_sfixed_a(-0.00013689820480067283)),(to_sfixed_a(0.00014070590259507298)),(to_sfixed_a(-5.436842911876738e-05)),(to_sfixed_a(-5.668488665833138e-05)),(to_sfixed_a(3.614449951783172e-06)),(to_sfixed_a(-0.00017194289830513299)),(to_sfixed_a(-0.00015253754099830985)),(to_sfixed_a(0.09001140296459198)),(to_sfixed_a(0.028936129063367844)),(to_sfixed_a(0.12063068896532059)),(to_sfixed_a(0.03708454966545105)),(to_sfixed_a(-0.13240256905555725)),(to_sfixed_a(0.21527297794818878)),(to_sfixed_a(0.23124472796916962)),(to_sfixed_a(0.36271533370018005)),(to_sfixed_a(0.20165352523326874)),(to_sfixed_a(0.01694202981889248)),(to_sfixed_a(0.002640628023073077)),(to_sfixed_a(0.016660116612911224)),(to_sfixed_a(-0.21732443571090698)),(to_sfixed_a(0.0016476697055622935)),(to_sfixed_a(0.10147187113761902)),(to_sfixed_a(0.06857497245073318)),(to_sfixed_a(0.004760755226016045)),(to_sfixed_a(-0.16608084738254547)),(to_sfixed_a(0.041348423808813095)),(to_sfixed_a(-0.02027813531458378)),(to_sfixed_a(0.027461780235171318)),(to_sfixed_a(-0.047302115708589554)),(to_sfixed_a(-5.41487243026495e-05)),(to_sfixed_a(-0.0003466065682005137)),(to_sfixed_a(3.326519072288647e-05)),(to_sfixed_a(8.758810145081952e-05)),(to_sfixed_a(0.00025749055203050375)),(to_sfixed_a(-0.00012499258446041495)),(to_sfixed_a(0.0014644768089056015)),(to_sfixed_a(0.11251004040241241)),(to_sfixed_a(-0.004056022502481937)),(to_sfixed_a(0.011063742451369762)),(to_sfixed_a(-0.0031783210579305887)),(to_sfixed_a(0.14200998842716217)),(to_sfixed_a(0.14751949906349182)),(to_sfixed_a(0.2877964675426483)),(to_sfixed_a(0.4234919548034668)),(to_sfixed_a(0.2265208512544632)),(to_sfixed_a(0.17335167527198792)),(to_sfixed_a(-0.2092256397008896)),(to_sfixed_a(-0.23566177487373352)),(to_sfixed_a(-0.03264590725302696)),(to_sfixed_a(0.019915509968996048)),(to_sfixed_a(0.09419945627450943)),(to_sfixed_a(-0.06066533550620079)),(to_sfixed_a(-0.12356717884540558)),(to_sfixed_a(0.07244791090488434)),(to_sfixed_a(-0.07110845297574997)),(to_sfixed_a(-0.06741169095039368)),(to_sfixed_a(-5.375825276132673e-05)),(to_sfixed_a(0.0005011419416405261)),(to_sfixed_a(-4.110762893105857e-05)),(to_sfixed_a(0.00014617727720178664)),(to_sfixed_a(-2.7367283109924756e-05)),(to_sfixed_a(-6.969608512008563e-05)),(to_sfixed_a(-9.041729936143383e-05)),(to_sfixed_a(0.004089794587343931)),(to_sfixed_a(0.026947999373078346)),(to_sfixed_a(0.1694774627685547)),(to_sfixed_a(0.18789178133010864)),(to_sfixed_a(0.05075865238904953)),(to_sfixed_a(-0.048517219722270966)),(to_sfixed_a(0.21699677407741547)),(to_sfixed_a(0.1581266075372696)),(to_sfixed_a(0.19950968027114868)),(to_sfixed_a(-0.09076827019453049)),(to_sfixed_a(-0.6430677175521851)),(to_sfixed_a(-0.15137958526611328)),(to_sfixed_a(-0.08285657316446304)),(to_sfixed_a(-0.06134886294603348)),(to_sfixed_a(0.03348277509212494)),(to_sfixed_a(0.09444904327392578)),(to_sfixed_a(0.07399318367242813)),(to_sfixed_a(0.042622216045856476)),(to_sfixed_a(-0.005606100894510746)),(to_sfixed_a(-0.08606112748384476)),(to_sfixed_a(0.08950693905353546)),(to_sfixed_a(0.0022538178600370884)),(to_sfixed_a(-8.149092536768876e-06)),(to_sfixed_a(-0.00021676642063539475)),(to_sfixed_a(-0.00029337088926695287)),(to_sfixed_a(-6.0804035456385463e-05)),(to_sfixed_a(8.658194565214217e-05)),(to_sfixed_a(-0.009045582264661789)),(to_sfixed_a(0.08213196694850922)),(to_sfixed_a(-0.06863187998533249)),(to_sfixed_a(0.13094183802604675)),(to_sfixed_a(-0.01809871941804886)),(to_sfixed_a(-0.0701829344034195)),(to_sfixed_a(-0.23677337169647217)),(to_sfixed_a(-0.4401986598968506)),(to_sfixed_a(-0.6336374878883362)),(to_sfixed_a(-0.7770739793777466)),(to_sfixed_a(-0.4217340052127838)),(to_sfixed_a(-0.2513499855995178)),(to_sfixed_a(-0.03104257397353649)),(to_sfixed_a(-0.1508507877588272)),(to_sfixed_a(0.16969837248325348)),(to_sfixed_a(0.16475586593151093)),(to_sfixed_a(-0.01729607582092285)),(to_sfixed_a(0.15738508105278015)),(to_sfixed_a(-0.10250884294509888)),(to_sfixed_a(0.038112886250019073)),(to_sfixed_a(-0.21685731410980225)),(to_sfixed_a(0.0927174836397171)),(to_sfixed_a(3.814190858975053e-05)),(to_sfixed_a(-4.6546654630219564e-05)),(to_sfixed_a(-1.9515759049681947e-05)),(to_sfixed_a(-6.0512134950840846e-05)),(to_sfixed_a(0.00024615516304038465)),(to_sfixed_a(9.86452869256027e-05)),(to_sfixed_a(0.00013731361832469702)),(to_sfixed_a(-0.15225209295749664)),(to_sfixed_a(-0.39670467376708984)),(to_sfixed_a(-0.19490092992782593)),(to_sfixed_a(-0.30749568343162537)),(to_sfixed_a(-0.6825044751167297)),(to_sfixed_a(-0.9241513609886169)),(to_sfixed_a(-0.6510217785835266)),(to_sfixed_a(-0.378390371799469)),(to_sfixed_a(-0.16507922112941742)),(to_sfixed_a(-0.16259784996509552)),(to_sfixed_a(0.0927780494093895)),(to_sfixed_a(0.3486827313899994)),(to_sfixed_a(0.05981110408902168)),(to_sfixed_a(0.2226448357105255)),(to_sfixed_a(0.09818382561206818)),(to_sfixed_a(-0.18215814232826233)),(to_sfixed_a(0.07659375667572021)),(to_sfixed_a(-0.046918611973524094)),(to_sfixed_a(-0.0022842136677354574)),(to_sfixed_a(-0.20519542694091797)),(to_sfixed_a(-0.02111894264817238)),(to_sfixed_a(9.810725168790668e-05)),(to_sfixed_a(-0.00012009042256977409)),(to_sfixed_a(0.00019403325859457254)),(to_sfixed_a(2.6868436179938726e-05)),(to_sfixed_a(3.483239925117232e-05)),(to_sfixed_a(0.00019020619220100343)),(to_sfixed_a(0.00035361506161279976)),(to_sfixed_a(-0.05971458554267883)),(to_sfixed_a(-0.3373408019542694)),(to_sfixed_a(-0.6490280628204346)),(to_sfixed_a(-0.5964956879615784)),(to_sfixed_a(-0.5448429584503174)),(to_sfixed_a(-0.32859131693840027)),(to_sfixed_a(-0.03199498727917671)),(to_sfixed_a(0.004333360120654106)),(to_sfixed_a(0.2796191871166229)),(to_sfixed_a(0.0791744738817215)),(to_sfixed_a(0.01955498196184635)),(to_sfixed_a(0.020897267386317253)),(to_sfixed_a(0.16484121978282928)),(to_sfixed_a(0.0837986096739769)),(to_sfixed_a(0.08157862722873688)),(to_sfixed_a(0.2067469358444214)),(to_sfixed_a(-0.14757494628429413)),(to_sfixed_a(0.039940692484378815)),(to_sfixed_a(0.027006186544895172)),(to_sfixed_a(-0.12437504529953003)),(to_sfixed_a(0.025480415672063828)),(to_sfixed_a(0.0011911385226994753)),(to_sfixed_a(0.0002483983989804983)),(to_sfixed_a(0.00025339657440781593)),(to_sfixed_a(-0.000172352374647744)),(to_sfixed_a(-0.00019416998839005828)),(to_sfixed_a(-7.586884748889133e-05)),(to_sfixed_a(-5.4657783039147034e-05)),(to_sfixed_a(0.0011479295790195465)),(to_sfixed_a(-0.8248506784439087)),(to_sfixed_a(-0.31364312767982483)),(to_sfixed_a(0.02133130468428135)),(to_sfixed_a(0.021990787237882614)),(to_sfixed_a(0.061766479164361954)),(to_sfixed_a(0.0962604507803917)),(to_sfixed_a(0.4927321970462799)),(to_sfixed_a(0.12778715789318085)),(to_sfixed_a(0.14251069724559784)),(to_sfixed_a(0.07929942011833191)),(to_sfixed_a(0.1843484342098236)),(to_sfixed_a(0.112239308655262)),(to_sfixed_a(0.16782639920711517)),(to_sfixed_a(0.27094724774360657)),(to_sfixed_a(0.2066914141178131)),(to_sfixed_a(0.09478896856307983)),(to_sfixed_a(0.02033940516412258)),(to_sfixed_a(-0.01775440201163292)),(to_sfixed_a(0.011157194152474403)),(to_sfixed_a(0.06116848438978195)),(to_sfixed_a(-0.00018619332695379853)),(to_sfixed_a(7.851214468246326e-05)),(to_sfixed_a(3.181712963851169e-05)),(to_sfixed_a(-5.817205965286121e-05)),(to_sfixed_a(-0.0001345552154816687)),(to_sfixed_a(-4.5832352043362334e-05)),(to_sfixed_a(-0.00013315636897459626)),(to_sfixed_a(-0.027740437537431717)),(to_sfixed_a(-0.19264841079711914)),(to_sfixed_a(-0.1701764464378357)),(to_sfixed_a(-0.3479699194431305)),(to_sfixed_a(-0.4836372137069702)),(to_sfixed_a(-0.3144383132457733)),(to_sfixed_a(0.05113893747329712)),(to_sfixed_a(-0.12476257234811783)),(to_sfixed_a(-0.044502563774585724)),(to_sfixed_a(0.0977495014667511)),(to_sfixed_a(0.14856624603271484)),(to_sfixed_a(0.10541199892759323)),(to_sfixed_a(0.19363142549991608)),(to_sfixed_a(0.2893243432044983)),(to_sfixed_a(0.29966050386428833)),(to_sfixed_a(0.25188055634498596)),(to_sfixed_a(0.08056971430778503)),(to_sfixed_a(0.034700021147727966)),(to_sfixed_a(-0.050402138382196426)),(to_sfixed_a(-0.11914409697055817)),(to_sfixed_a(0.05494266748428345)),(to_sfixed_a(-0.0003206364926882088)),(to_sfixed_a(0.0003725358110386878)),(to_sfixed_a(-8.194560359697789e-05)),(to_sfixed_a(-6.620187923545018e-05)),(to_sfixed_a(0.00040137808537110686)),(to_sfixed_a(-9.131272236118093e-05)),(to_sfixed_a(0.002061376115307212)),(to_sfixed_a(-0.03611105680465698)),(to_sfixed_a(-0.008734025992453098)),(to_sfixed_a(-0.16915208101272583)),(to_sfixed_a(-0.42190271615982056)),(to_sfixed_a(-0.35259583592414856)),(to_sfixed_a(-0.19781585037708282)),(to_sfixed_a(-0.251567542552948)),(to_sfixed_a(-0.7062748670578003)),(to_sfixed_a(-0.2821027934551239)),(to_sfixed_a(-0.2514653503894806)),(to_sfixed_a(0.10620984435081482)),(to_sfixed_a(0.07100661844015121)),(to_sfixed_a(0.280193030834198)),(to_sfixed_a(0.23043422400951385)),(to_sfixed_a(0.39539191126823425)),(to_sfixed_a(0.23164649307727814)),(to_sfixed_a(0.18388722836971283)),(to_sfixed_a(0.044738609343767166)),(to_sfixed_a(-0.09750577807426453)),(to_sfixed_a(0.01882159523665905)),(to_sfixed_a(0.05612851306796074)),(to_sfixed_a(0.019235895946621895)),(to_sfixed_a(-0.00010848198871826753)),(to_sfixed_a(0.00016377314750570804)),(to_sfixed_a(1.2777002666553017e-05)),(to_sfixed_a(0.00019055882876273245)),(to_sfixed_a(0.0015048040077090263)),(to_sfixed_a(0.0019359933212399483)),(to_sfixed_a(0.13296106457710266)),(to_sfixed_a(-0.11843894422054291)),(to_sfixed_a(-0.13869939744472504)),(to_sfixed_a(-0.2771451771259308)),(to_sfixed_a(-0.2357965111732483)),(to_sfixed_a(-0.4172861874103546)),(to_sfixed_a(-0.49053511023521423)),(to_sfixed_a(-0.7793645858764648)),(to_sfixed_a(-0.7620854377746582)),(to_sfixed_a(-0.2686692774295807)),(to_sfixed_a(-0.0372784398496151)),(to_sfixed_a(0.293748140335083)),(to_sfixed_a(0.34280478954315186)),(to_sfixed_a(0.17640377581119537)),(to_sfixed_a(0.2122942954301834)),(to_sfixed_a(-0.025505904108285904)),(to_sfixed_a(0.0544389933347702)),(to_sfixed_a(-0.06928449124097824)),(to_sfixed_a(-0.1754426807165146)),(to_sfixed_a(-0.026833996176719666)),(to_sfixed_a(2.0298572053434327e-05)),(to_sfixed_a(0.00011342045036144555)),(to_sfixed_a(4.689088382292539e-05)),(to_sfixed_a(2.445317295496352e-05)),(to_sfixed_a(4.018512845505029e-05)),(to_sfixed_a(-7.351356180151924e-05)),(to_sfixed_a(-0.0004884491208940744)),(to_sfixed_a(-0.022908220067620277)),(to_sfixed_a(0.021939139813184738)),(to_sfixed_a(0.23980402946472168)),(to_sfixed_a(0.3109489679336548)),(to_sfixed_a(0.24931256473064423)),(to_sfixed_a(0.13463720679283142)),(to_sfixed_a(-0.4517902433872223)),(to_sfixed_a(-0.6639541983604431)),(to_sfixed_a(-0.510284423828125)),(to_sfixed_a(-0.36520111560821533)),(to_sfixed_a(-0.04059463366866112)),(to_sfixed_a(0.14787700772285461)),(to_sfixed_a(0.32416850328445435)),(to_sfixed_a(0.29606106877326965)),(to_sfixed_a(0.23177620768547058)),(to_sfixed_a(0.034267544746398926)),(to_sfixed_a(-0.06660417467355728)),(to_sfixed_a(-0.17361357808113098)),(to_sfixed_a(-0.2318829894065857)),(to_sfixed_a(-0.11862213909626007)),(to_sfixed_a(-0.005637396592646837)),(to_sfixed_a(0.030243005603551865)),(to_sfixed_a(9.55586729105562e-05)),(to_sfixed_a(2.38904631260084e-05)),(to_sfixed_a(-0.00016841063916217536)),(to_sfixed_a(-0.00036919835838489234)),(to_sfixed_a(-4.752446329803206e-05)),(to_sfixed_a(0.0002173713583033532)),(to_sfixed_a(0.1444992572069168)),(to_sfixed_a(-0.0008884271373972297)),(to_sfixed_a(0.06377433985471725)),(to_sfixed_a(0.08036402612924576)),(to_sfixed_a(0.4066859483718872)),(to_sfixed_a(0.239628866314888)),(to_sfixed_a(0.2912803590297699)),(to_sfixed_a(0.1283291131258011)),(to_sfixed_a(0.12957291305065155)),(to_sfixed_a(-0.10351034253835678)),(to_sfixed_a(0.05507507547736168)),(to_sfixed_a(0.18656671047210693)),(to_sfixed_a(0.35196810960769653)),(to_sfixed_a(0.03396570309996605)),(to_sfixed_a(-0.009477372281253338)),(to_sfixed_a(-0.07775068283081055)),(to_sfixed_a(-0.05375419929623604)),(to_sfixed_a(-0.2554636299610138)),(to_sfixed_a(-0.20066945254802704)),(to_sfixed_a(0.01646040566265583)),(to_sfixed_a(-0.06461597234010696)),(to_sfixed_a(-9.25465501495637e-05)),(to_sfixed_a(1.3106372534821276e-05)),(to_sfixed_a(0.00025975616881623864)),(to_sfixed_a(0.00032358523458242416)),(to_sfixed_a(-7.55710425437428e-05)),(to_sfixed_a(-0.0001427673560101539)),(to_sfixed_a(-6.94321101946116e-07)),(to_sfixed_a(0.0001473509328207001)),(to_sfixed_a(-0.0005935126100666821)),(to_sfixed_a(-0.000994959264062345)),(to_sfixed_a(-0.1186266839504242)),(to_sfixed_a(-0.0671471655368805)),(to_sfixed_a(-0.10905057936906815)),(to_sfixed_a(0.12530827522277832)),(to_sfixed_a(0.047750648111104965)),(to_sfixed_a(0.13810928165912628)),(to_sfixed_a(0.11320837587118149)),(to_sfixed_a(0.06817682832479477)),(to_sfixed_a(0.1391735076904297)),(to_sfixed_a(0.23330187797546387)),(to_sfixed_a(-0.003944766242057085)),(to_sfixed_a(0.045249562710523605)),(to_sfixed_a(-0.2805020809173584)),(to_sfixed_a(-0.29749828577041626)),(to_sfixed_a(-0.3246769309043884)),(to_sfixed_a(-0.09118032455444336)),(to_sfixed_a(0.014646715484559536)),(to_sfixed_a(0.13705530762672424)),(to_sfixed_a(0.13505317270755768)),(to_sfixed_a(7.828141679055989e-05)),(to_sfixed_a(0.00012204711674712598)),(to_sfixed_a(-0.00029724958585575223)),(to_sfixed_a(-0.000123709934996441)),(to_sfixed_a(-0.0001586561556905508)),(to_sfixed_a(-0.00019589340081438422)),(to_sfixed_a(-0.00013831017713528126)),(to_sfixed_a(0.042121220380067825)),(to_sfixed_a(0.0003454398538451642)),(to_sfixed_a(0.08994308859109879)),(to_sfixed_a(-0.3127180337905884)),(to_sfixed_a(-0.06735486537218094)),(to_sfixed_a(-0.19447484612464905)),(to_sfixed_a(0.1072099506855011)),(to_sfixed_a(0.217965766787529)),(to_sfixed_a(-0.021092401817440987)),(to_sfixed_a(0.27881306409835815)),(to_sfixed_a(-0.10811129212379456)),(to_sfixed_a(-0.1412239372730255)),(to_sfixed_a(-0.03563293069601059)),(to_sfixed_a(0.011940118856728077)),(to_sfixed_a(-0.02003517746925354)),(to_sfixed_a(-0.21479961276054382)),(to_sfixed_a(-0.3627113699913025)),(to_sfixed_a(-0.09929929673671722)),(to_sfixed_a(-0.10934460163116455)),(to_sfixed_a(-1.591359068697784e-05)),(to_sfixed_a(-0.012275397777557373)),(to_sfixed_a(-5.730247721658088e-05)),(to_sfixed_a(-0.0001355269196210429)),(to_sfixed_a(0.00023796249297447503)),(to_sfixed_a(0.00019554361642803997)),(to_sfixed_a(-0.00013234541984274983)),(to_sfixed_a(1.9738405171665363e-05)),(to_sfixed_a(0.00015372376947198063)),(to_sfixed_a(-1.4795693459745962e-05)),(to_sfixed_a(-0.033596549183130264)),(to_sfixed_a(-0.0418565459549427)),(to_sfixed_a(-0.2926080822944641)),(to_sfixed_a(0.049096763134002686)),(to_sfixed_a(-0.06924083083868027)),(to_sfixed_a(-0.09097307920455933)),(to_sfixed_a(0.09020373970270157)),(to_sfixed_a(0.03798767179250717)),(to_sfixed_a(-0.06267620623111725)),(to_sfixed_a(-0.11024990677833557)),(to_sfixed_a(-0.002295867772772908)),(to_sfixed_a(-0.1147545799612999)),(to_sfixed_a(-0.1285981982946396)),(to_sfixed_a(-0.5356552004814148)),(to_sfixed_a(0.05914422497153282)),(to_sfixed_a(-0.10628443211317062)),(to_sfixed_a(-0.02208823151886463)),(to_sfixed_a(-0.018808655440807343)),(to_sfixed_a(-0.005724884103983641)),(to_sfixed_a(5.014162525185384e-05)),(to_sfixed_a(-6.0133588704047725e-05)),(to_sfixed_a(0.000264825823251158)),(to_sfixed_a(-0.00010533159365877509)),(to_sfixed_a(1.991387762245722e-05)),(to_sfixed_a(3.0187646189006045e-05)),(to_sfixed_a(0.00012462720042094588)),(to_sfixed_a(0.00018924663891084492)),(to_sfixed_a(-6.364323053276166e-05)),(to_sfixed_a(0.0817948430776596)),(to_sfixed_a(-0.016788864508271217)),(to_sfixed_a(-0.08855997025966644)),(to_sfixed_a(-0.07884731888771057)),(to_sfixed_a(-0.03780105337500572)),(to_sfixed_a(0.06020171195268631)),(to_sfixed_a(0.007516284007579088)),(to_sfixed_a(0.0014070235192775726)),(to_sfixed_a(-0.04614710435271263)),(to_sfixed_a(-0.11439199000597)),(to_sfixed_a(-0.09054621309041977)),(to_sfixed_a(-0.32369309663772583)),(to_sfixed_a(-0.29719123244285583)),(to_sfixed_a(-0.12115299701690674)),(to_sfixed_a(0.022245444357395172)),(to_sfixed_a(-0.03967327997088432)),(to_sfixed_a(-0.06372194737195969)),(to_sfixed_a(-0.003512375522404909)),(to_sfixed_a(-0.040654052048921585)),(to_sfixed_a(0.00010282263247063383)),(to_sfixed_a(1.8726046619121917e-05)),(to_sfixed_a(8.806256664684042e-05)),(to_sfixed_a(2.4201559426728636e-05)),(to_sfixed_a(0.00019416975555941463)),(to_sfixed_a(-0.00021119344455655664)),(to_sfixed_a(7.969700163812377e-06)),(to_sfixed_a(4.309593350626528e-05)),(to_sfixed_a(0.007899126969277859)),(to_sfixed_a(-0.013161910697817802)),(to_sfixed_a(0.03303218632936478)),(to_sfixed_a(-0.08334527909755707)),(to_sfixed_a(-0.12688840925693512)),(to_sfixed_a(-0.1734331101179123)),(to_sfixed_a(-0.3579603433609009)),(to_sfixed_a(-0.0952097699046135)),(to_sfixed_a(-0.11134207993745804)),(to_sfixed_a(-0.14350098371505737)),(to_sfixed_a(-0.30657094717025757)),(to_sfixed_a(-0.0969928652048111)),(to_sfixed_a(0.015619689598679543)),(to_sfixed_a(-0.12264657765626907)),(to_sfixed_a(-0.1601054072380066)),(to_sfixed_a(-0.07203991711139679)),(to_sfixed_a(-0.007173285819590092)),(to_sfixed_a(-0.03190970420837402)),(to_sfixed_a(-0.020289301872253418)),(to_sfixed_a(0.0060400934889912605)),(to_sfixed_a(0.0001949887373484671)),(to_sfixed_a(0.0002465302241034806)),(to_sfixed_a(0.00013124373799655586)),(to_sfixed_a(3.4598524507600814e-05)),(to_sfixed_a(0.00022337598784361035)),(to_sfixed_a(-1.2435517646736116e-06)),(to_sfixed_a(0.00024855579249560833)),(to_sfixed_a(-5.201229214435443e-05)),(to_sfixed_a(-5.3238010877976194e-05)),(to_sfixed_a(0.031340718269348145)),(to_sfixed_a(0.01990327425301075)),(to_sfixed_a(0.00046244022087194026)),(to_sfixed_a(0.0070635308511555195)),(to_sfixed_a(-0.06328606605529785)),(to_sfixed_a(0.1075875535607338)),(to_sfixed_a(0.04568988084793091)),(to_sfixed_a(-0.0075518605299293995)),(to_sfixed_a(0.014319737441837788)),(to_sfixed_a(-0.06475569307804108)),(to_sfixed_a(-0.02535792626440525)),(to_sfixed_a(0.2575763761997223)),(to_sfixed_a(0.015194736421108246)),(to_sfixed_a(-0.0018810373730957508)),(to_sfixed_a(0.04901614412665367)),(to_sfixed_a(0.027325022965669632)),(to_sfixed_a(-1.2173334653198253e-05)),(to_sfixed_a(0.0026124166324734688)),(to_sfixed_a(0.003013793844729662)),(to_sfixed_a(1.694200182100758e-05)),(to_sfixed_a(0.00018536459538154304)),(to_sfixed_a(-0.0002362500672461465)),(to_sfixed_a(6.24457243247889e-05)),(to_sfixed_a(0.00018864076992031187)),(to_sfixed_a(0.0002618557773530483)),(to_sfixed_a(-3.09342794935219e-05)),(to_sfixed_a(0.0001246091560460627)),(to_sfixed_a(6.856859727122355e-06)),(to_sfixed_a(-3.206944165867753e-05)),(to_sfixed_a(-0.00034255048376508057)),(to_sfixed_a(4.1365972720086575e-05)),(to_sfixed_a(-0.0004091597511433065)),(to_sfixed_a(-0.00036736318725161254)),(to_sfixed_a(0.0633343979716301)),(to_sfixed_a(-0.0002665386418811977)),(to_sfixed_a(-0.0030532937962561846)),(to_sfixed_a(0.046884484589099884)),(to_sfixed_a(0.05316336825489998)),(to_sfixed_a(0.008448158390820026)),(to_sfixed_a(0.01513570174574852)),(to_sfixed_a(0.04973280057311058)),(to_sfixed_a(0.06822039186954498)),(to_sfixed_a(0.003710707649588585)),(to_sfixed_a(0.001971346791833639)),(to_sfixed_a(-6.197894254000857e-05)),(to_sfixed_a(4.639910184778273e-05)),(to_sfixed_a(-5.828493522130884e-05)),(to_sfixed_a(0.0002310072595719248)),(to_sfixed_a(-5.808407149743289e-05)),(to_sfixed_a(5.2478586439974606e-05)),(to_sfixed_a(3.9037931856000796e-05)),(to_sfixed_a(0.00016063575458247215)),(to_sfixed_a(-0.00027966973721049726)),(to_sfixed_a(0.00011473378981463611)),(to_sfixed_a(-0.00010913109144894406)),(to_sfixed_a(2.6245414119330235e-05)),(to_sfixed_a(2.484536889824085e-05)),(to_sfixed_a(-0.0002554908278398216)),(to_sfixed_a(0.0002938829711638391)),(to_sfixed_a(-0.00017505098367109895)),(to_sfixed_a(-0.0001192488634842448)),(to_sfixed_a(-0.00026925260317511857)),(to_sfixed_a(0.0002356726472498849)),(to_sfixed_a(7.052694127196446e-05)),(to_sfixed_a(-0.00014940736582502723)),(to_sfixed_a(-0.00010758429561974481)),(to_sfixed_a(4.997547875973396e-05)),(to_sfixed_a(0.0001393870625179261)),(to_sfixed_a(-2.3765538571751676e-05)),(to_sfixed_a(8.407342102145776e-05)),(to_sfixed_a(-0.000170427534612827)),(to_sfixed_a(0.00023145614250097424)),(to_sfixed_a(8.589561184635386e-05)),(to_sfixed_a(0.00012726565182674676)),(to_sfixed_a(0.00013395925634540617)),(to_sfixed_a(-9.46805375861004e-05)),(to_sfixed_a(-2.2269228793447837e-05)),(to_sfixed_a(-0.00027143029728904366)),(to_sfixed_a(3.944928175769746e-05)));

    constant weight_n0_7 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(9.989850696001668e-06)),(to_sfixed_a(8.636365964775905e-05)),(to_sfixed_a(6.988312816247344e-05)),(to_sfixed_a(5.9813606640091166e-05)),(to_sfixed_a(-2.0550178305711597e-05)),(to_sfixed_a(-7.963008101796731e-05)),(to_sfixed_a(-6.663558451691642e-05)),(to_sfixed_a(0.00015662526129744947)),(to_sfixed_a(0.00020838248019572347)),(to_sfixed_a(9.581031918060035e-05)),(to_sfixed_a(-0.00024597058654762805)),(to_sfixed_a(-3.9851845940575004e-05)),(to_sfixed_a(0.00014876284694764763)),(to_sfixed_a(0.0003693017642945051)),(to_sfixed_a(0.00019285180314909667)),(to_sfixed_a(0.0002274524886161089)),(to_sfixed_a(-0.00027175850118510425)),(to_sfixed_a(0.00021467896294780076)),(to_sfixed_a(-0.0001493167510489002)),(to_sfixed_a(-3.120343171758577e-05)),(to_sfixed_a(-7.422240742016584e-05)),(to_sfixed_a(-0.00012967389193363488)),(to_sfixed_a(0.00019845170027110726)),(to_sfixed_a(-0.00037517197779379785)),(to_sfixed_a(0.0001953742903424427)),(to_sfixed_a(0.00016528739070054144)),(to_sfixed_a(8.414646435994655e-05)),(to_sfixed_a(-0.00020893869805149734)),(to_sfixed_a(2.2327076294459403e-05)),(to_sfixed_a(0.0002869957825168967)),(to_sfixed_a(0.00029255871777422726)),(to_sfixed_a(-5.990233694319613e-05)),(to_sfixed_a(-0.00015771272592246532)),(to_sfixed_a(-0.00011141527647851035)),(to_sfixed_a(0.0001856002927524969)),(to_sfixed_a(-0.00018748770526144654)),(to_sfixed_a(0.00012594496365636587)),(to_sfixed_a(-0.00019483872165437788)),(to_sfixed_a(0.0002284893998876214)),(to_sfixed_a(-0.00021221015776973218)),(to_sfixed_a(-7.748949428787455e-05)),(to_sfixed_a(-0.00010901391215156764)),(to_sfixed_a(-4.9642083467915654e-05)),(to_sfixed_a(1.5532261841144646e-06)),(to_sfixed_a(-1.5035378737593419e-06)),(to_sfixed_a(-0.0002769177663139999)),(to_sfixed_a(-7.722172449575737e-05)),(to_sfixed_a(0.00013856746954843402)),(to_sfixed_a(-9.598812903277576e-05)),(to_sfixed_a(-8.13467413536273e-05)),(to_sfixed_a(0.00017060484969988465)),(to_sfixed_a(0.00017863832181319594)),(to_sfixed_a(0.0001171723852166906)),(to_sfixed_a(-1.629727012186777e-05)),(to_sfixed_a(5.669312668032944e-05)),(to_sfixed_a(-0.0001401591143803671)),(to_sfixed_a(0.00015240484208334237)),(to_sfixed_a(-5.607316779787652e-05)),(to_sfixed_a(5.787869667983614e-05)),(to_sfixed_a(-7.523712702095509e-05)),(to_sfixed_a(-1.5256246115313843e-05)),(to_sfixed_a(-0.00024305173428729177)),(to_sfixed_a(5.060206967755221e-05)),(to_sfixed_a(-0.00019663436978589743)),(to_sfixed_a(9.104825585382059e-05)),(to_sfixed_a(-4.2684470827225596e-05)),(to_sfixed_a(-0.00019393773982301354)),(to_sfixed_a(-2.7732778562494786e-06)),(to_sfixed_a(-3.6670851841336116e-05)),(to_sfixed_a(-0.04710233956575394)),(to_sfixed_a(4.7368044761242345e-05)),(to_sfixed_a(4.318701758165844e-05)),(to_sfixed_a(-1.9459048417047597e-05)),(to_sfixed_a(9.398034308105707e-05)),(to_sfixed_a(0.0001821917830966413)),(to_sfixed_a(0.00010223377466900274)),(to_sfixed_a(5.4706353694200516e-05)),(to_sfixed_a(0.0002665107022039592)),(to_sfixed_a(0.00010447706881677732)),(to_sfixed_a(-0.0001625983277335763)),(to_sfixed_a(-4.5770942961098626e-05)),(to_sfixed_a(5.833229806739837e-05)),(to_sfixed_a(0.0001938327623065561)),(to_sfixed_a(-3.283767000539228e-05)),(to_sfixed_a(5.730747216148302e-05)),(to_sfixed_a(-0.00020338327158242464)),(to_sfixed_a(0.00013412104453891516)),(to_sfixed_a(-4.0669670852366835e-05)),(to_sfixed_a(-0.00010789353837026283)),(to_sfixed_a(-6.421911621146137e-06)),(to_sfixed_a(-0.00022808446374256164)),(to_sfixed_a(-0.00013650204346049577)),(to_sfixed_a(-0.03659605607390404)),(to_sfixed_a(9.448199853068218e-05)),(to_sfixed_a(-0.04118715599179268)),(to_sfixed_a(0.041003093123435974)),(to_sfixed_a(-0.10226769745349884)),(to_sfixed_a(0.056810710579156876)),(to_sfixed_a(-0.13206060230731964)),(to_sfixed_a(0.023096904158592224)),(to_sfixed_a(-0.003994896076619625)),(to_sfixed_a(-0.1091671958565712)),(to_sfixed_a(0.20783820748329163)),(to_sfixed_a(-0.07952279597520828)),(to_sfixed_a(0.0074414946138858795)),(to_sfixed_a(0.015359196811914444)),(to_sfixed_a(-4.037962935399264e-05)),(to_sfixed_a(-0.0002433123008813709)),(to_sfixed_a(-0.00016343273455277085)),(to_sfixed_a(-0.00010464361548656598)),(to_sfixed_a(-0.00012106842041248456)),(to_sfixed_a(9.459778812015429e-05)),(to_sfixed_a(-0.00028183363610878587)),(to_sfixed_a(0.0002255822764709592)),(to_sfixed_a(-0.00011334034206811339)),(to_sfixed_a(-4.541236557997763e-05)),(to_sfixed_a(0.00013080492499284446)),(to_sfixed_a(6.316799408523366e-05)),(to_sfixed_a(0.0011137938126921654)),(to_sfixed_a(0.018727727234363556)),(to_sfixed_a(-0.0166368056088686)),(to_sfixed_a(-0.05473916232585907)),(to_sfixed_a(-0.011184928007423878)),(to_sfixed_a(-0.10559305548667908)),(to_sfixed_a(0.0018097517313435674)),(to_sfixed_a(-0.21065488457679749)),(to_sfixed_a(0.20333251357078552)),(to_sfixed_a(0.18931923806667328)),(to_sfixed_a(0.1776919662952423)),(to_sfixed_a(0.08936650305986404)),(to_sfixed_a(0.16515301167964935)),(to_sfixed_a(-0.04255625233054161)),(to_sfixed_a(-0.023313170298933983)),(to_sfixed_a(0.09310978651046753)),(to_sfixed_a(0.007615505717694759)),(to_sfixed_a(0.00012974190758541226)),(to_sfixed_a(-0.0003469669900368899)),(to_sfixed_a(7.58001406211406e-05)),(to_sfixed_a(3.934365668101236e-05)),(to_sfixed_a(-0.0001441097992938012)),(to_sfixed_a(-6.803293217672035e-05)),(to_sfixed_a(-0.0001368314551655203)),(to_sfixed_a(-0.0002200684102717787)),(to_sfixed_a(0.00032139665563590825)),(to_sfixed_a(-5.1476392400218174e-05)),(to_sfixed_a(0.017805466428399086)),(to_sfixed_a(-0.0067808423191308975)),(to_sfixed_a(-0.014003215357661247)),(to_sfixed_a(-0.008894327096641064)),(to_sfixed_a(0.03971179574728012)),(to_sfixed_a(-0.007561307866126299)),(to_sfixed_a(-0.12319128215312958)),(to_sfixed_a(-0.0849074050784111)),(to_sfixed_a(-0.09949160367250443)),(to_sfixed_a(0.036941055208444595)),(to_sfixed_a(-0.1822584867477417)),(to_sfixed_a(-0.15007685124874115)),(to_sfixed_a(0.09136602282524109)),(to_sfixed_a(0.15783679485321045)),(to_sfixed_a(-0.015116598457098007)),(to_sfixed_a(-0.023318028077483177)),(to_sfixed_a(-0.04921712353825569)),(to_sfixed_a(-0.00045301084173843265)),(to_sfixed_a(0.033697862178087234)),(to_sfixed_a(0.0005398727371357381)),(to_sfixed_a(0.0010005063377320766)),(to_sfixed_a(7.826725777704269e-05)),(to_sfixed_a(8.716033335076645e-05)),(to_sfixed_a(8.159858407452703e-05)),(to_sfixed_a(7.964677206473425e-05)),(to_sfixed_a(5.834956027683802e-05)),(to_sfixed_a(-3.061724783037789e-05)),(to_sfixed_a(-1.0463287253514864e-05)),(to_sfixed_a(0.015112304128706455)),(to_sfixed_a(0.0008646539645269513)),(to_sfixed_a(0.13611142337322235)),(to_sfixed_a(0.2282264083623886)),(to_sfixed_a(0.05256270617246628)),(to_sfixed_a(-0.035184405744075775)),(to_sfixed_a(-0.08293650299310684)),(to_sfixed_a(-0.11758724600076675)),(to_sfixed_a(-0.17611850798130035)),(to_sfixed_a(-0.30736732482910156)),(to_sfixed_a(0.03767375275492668)),(to_sfixed_a(0.25506019592285156)),(to_sfixed_a(0.10295780748128891)),(to_sfixed_a(0.20420551300048828)),(to_sfixed_a(0.10254564136266708)),(to_sfixed_a(0.08595051616430283)),(to_sfixed_a(0.046103786677122116)),(to_sfixed_a(-0.1517799347639084)),(to_sfixed_a(-0.22674110531806946)),(to_sfixed_a(-0.0041154976934194565)),(to_sfixed_a(-0.0053142583929002285)),(to_sfixed_a(-0.003539640922099352)),(to_sfixed_a(-2.1441232092911378e-05)),(to_sfixed_a(-6.665155524387956e-06)),(to_sfixed_a(-0.00023306756338570267)),(to_sfixed_a(-0.00014434430340770632)),(to_sfixed_a(6.210459105204791e-05)),(to_sfixed_a(-1.3955273061583284e-05)),(to_sfixed_a(-0.011960635893046856)),(to_sfixed_a(-0.18135088682174683)),(to_sfixed_a(0.011081679724156857)),(to_sfixed_a(0.013846267946064472)),(to_sfixed_a(0.06068409979343414)),(to_sfixed_a(-0.5846296548843384)),(to_sfixed_a(-0.3320189416408539)),(to_sfixed_a(-0.26070648431777954)),(to_sfixed_a(-0.31915706396102905)),(to_sfixed_a(-0.17576570808887482)),(to_sfixed_a(0.07982759177684784)),(to_sfixed_a(0.14387483894824982)),(to_sfixed_a(0.4339224100112915)),(to_sfixed_a(0.4458525478839874)),(to_sfixed_a(0.6282455921173096)),(to_sfixed_a(0.5433234572410583)),(to_sfixed_a(0.02644924819469452)),(to_sfixed_a(-0.11550413072109222)),(to_sfixed_a(0.27003055810928345)),(to_sfixed_a(-0.14839376509189606)),(to_sfixed_a(0.0031083920039236546)),(to_sfixed_a(-8.037497173063457e-05)),(to_sfixed_a(-5.6390581448795274e-05)),(to_sfixed_a(0.00021020670828875154)),(to_sfixed_a(-8.114675438264385e-06)),(to_sfixed_a(-0.0002832794561982155)),(to_sfixed_a(-7.622322300449014e-05)),(to_sfixed_a(0.016489610075950623)),(to_sfixed_a(0.052407097071409225)),(to_sfixed_a(-0.0174026470631361)),(to_sfixed_a(-0.17993591725826263)),(to_sfixed_a(-0.15961511433124542)),(to_sfixed_a(-0.06977177411317825)),(to_sfixed_a(-0.12005021423101425)),(to_sfixed_a(-0.03942515701055527)),(to_sfixed_a(-0.15040679275989532)),(to_sfixed_a(-0.18975110352039337)),(to_sfixed_a(-0.3821408450603485)),(to_sfixed_a(0.33218592405319214)),(to_sfixed_a(0.6144606471061707)),(to_sfixed_a(0.6969485878944397)),(to_sfixed_a(0.753994345664978)),(to_sfixed_a(0.2634252905845642)),(to_sfixed_a(0.32720810174942017)),(to_sfixed_a(0.13728943467140198)),(to_sfixed_a(0.05019476264715195)),(to_sfixed_a(0.2073381543159485)),(to_sfixed_a(0.10371678322553635)),(to_sfixed_a(0.02348993718624115)),(to_sfixed_a(-0.00022588649881072342)),(to_sfixed_a(7.275116513483226e-05)),(to_sfixed_a(-0.00010304696479579434)),(to_sfixed_a(-6.0411424783524126e-05)),(to_sfixed_a(-4.083953535882756e-05)),(to_sfixed_a(0.00013613661576528102)),(to_sfixed_a(-0.0017529733013361692)),(to_sfixed_a(-0.036009274423122406)),(to_sfixed_a(-0.07080525159835815)),(to_sfixed_a(-0.06163753196597099)),(to_sfixed_a(-0.04749852791428566)),(to_sfixed_a(-0.022788990288972855)),(to_sfixed_a(-0.3586407005786896)),(to_sfixed_a(-0.08646883815526962)),(to_sfixed_a(-0.3226136565208435)),(to_sfixed_a(-0.3868980407714844)),(to_sfixed_a(-0.2735556960105896)),(to_sfixed_a(0.08857160061597824)),(to_sfixed_a(0.43058186769485474)),(to_sfixed_a(0.5635559558868408)),(to_sfixed_a(0.27304607629776)),(to_sfixed_a(0.11060771346092224)),(to_sfixed_a(0.23223379254341125)),(to_sfixed_a(0.077410988509655)),(to_sfixed_a(-0.03804505988955498)),(to_sfixed_a(-0.18842893838882446)),(to_sfixed_a(0.16328087449073792)),(to_sfixed_a(0.0001301816082559526)),(to_sfixed_a(-2.518824112485163e-05)),(to_sfixed_a(3.407138865441084e-05)),(to_sfixed_a(-0.00016435857105534524)),(to_sfixed_a(-0.00023613194935023785)),(to_sfixed_a(-7.127502613002434e-05)),(to_sfixed_a(-0.0002547767071519047)),(to_sfixed_a(-0.005462760105729103)),(to_sfixed_a(-0.0018928417703136802)),(to_sfixed_a(0.007477376610040665)),(to_sfixed_a(-0.07710921764373779)),(to_sfixed_a(-0.06323876976966858)),(to_sfixed_a(-0.14517125487327576)),(to_sfixed_a(0.054759431630373)),(to_sfixed_a(0.2137620896100998)),(to_sfixed_a(-0.016889503225684166)),(to_sfixed_a(0.06069266051054001)),(to_sfixed_a(0.05501345172524452)),(to_sfixed_a(-0.18967831134796143)),(to_sfixed_a(0.33538374304771423)),(to_sfixed_a(0.133027583360672)),(to_sfixed_a(-0.26764389872550964)),(to_sfixed_a(-0.3070669174194336)),(to_sfixed_a(-0.35006991028785706)),(to_sfixed_a(-0.378428190946579)),(to_sfixed_a(-0.1779116988182068)),(to_sfixed_a(-0.07599500566720963)),(to_sfixed_a(0.1267681121826172)),(to_sfixed_a(0.03725823014974594)),(to_sfixed_a(2.667253829713445e-05)),(to_sfixed_a(8.961780258687213e-05)),(to_sfixed_a(0.00037821015575900674)),(to_sfixed_a(0.00013832544209435582)),(to_sfixed_a(3.723072950378992e-05)),(to_sfixed_a(-0.02301104925572872)),(to_sfixed_a(0.037927255034446716)),(to_sfixed_a(0.06494104117155075)),(to_sfixed_a(-0.07925281673669815)),(to_sfixed_a(0.09073343127965927)),(to_sfixed_a(0.15835337340831757)),(to_sfixed_a(0.00836233887821436)),(to_sfixed_a(0.16112059354782104)),(to_sfixed_a(0.3280060589313507)),(to_sfixed_a(0.3359488248825073)),(to_sfixed_a(0.2490128129720688)),(to_sfixed_a(0.24955567717552185)),(to_sfixed_a(0.36291852593421936)),(to_sfixed_a(0.15719924867153168)),(to_sfixed_a(-0.288984090089798)),(to_sfixed_a(-0.34330251812934875)),(to_sfixed_a(-0.7253929972648621)),(to_sfixed_a(-0.7384796142578125)),(to_sfixed_a(-0.16852545738220215)),(to_sfixed_a(-0.27451854944229126)),(to_sfixed_a(-0.036166001111269)),(to_sfixed_a(0.05450662225484848)),(to_sfixed_a(0.00011544494918780401)),(to_sfixed_a(0.0002503185532987118)),(to_sfixed_a(-0.00010865743388421834)),(to_sfixed_a(0.00035075965570285916)),(to_sfixed_a(-0.0001994837512029335)),(to_sfixed_a(-0.00031757421675138175)),(to_sfixed_a(3.5562530683819205e-05)),(to_sfixed_a(0.02022121287882328)),(to_sfixed_a(-0.02449127472937107)),(to_sfixed_a(-0.012911995872855186)),(to_sfixed_a(0.12641116976737976)),(to_sfixed_a(0.2078903764486313)),(to_sfixed_a(0.1637527346611023)),(to_sfixed_a(0.2262912541627884)),(to_sfixed_a(0.30587267875671387)),(to_sfixed_a(0.06544665992259979)),(to_sfixed_a(0.20878590643405914)),(to_sfixed_a(0.3156565725803375)),(to_sfixed_a(0.480609267950058)),(to_sfixed_a(-0.0037865566555410624)),(to_sfixed_a(-0.2876240611076355)),(to_sfixed_a(-0.04038863256573677)),(to_sfixed_a(-0.7460634112358093)),(to_sfixed_a(-0.7427223324775696)),(to_sfixed_a(-0.3431084156036377)),(to_sfixed_a(-0.270659476518631)),(to_sfixed_a(-0.24543559551239014)),(to_sfixed_a(-0.03404773026704788)),(to_sfixed_a(-8.891889592632651e-06)),(to_sfixed_a(0.0005426777061074972)),(to_sfixed_a(9.751960169523954e-05)),(to_sfixed_a(-2.693876376724802e-05)),(to_sfixed_a(1.8244727471028455e-05)),(to_sfixed_a(1.989251177292317e-05)),(to_sfixed_a(-1.4512858797388617e-05)),(to_sfixed_a(-0.05370179936289787)),(to_sfixed_a(-0.02074463479220867)),(to_sfixed_a(-0.05142960324883461)),(to_sfixed_a(0.1090671643614769)),(to_sfixed_a(-0.07938345521688461)),(to_sfixed_a(0.03138292208313942)),(to_sfixed_a(0.09029722958803177)),(to_sfixed_a(0.18823176622390747)),(to_sfixed_a(0.08371800929307938)),(to_sfixed_a(0.04998881369829178)),(to_sfixed_a(0.5268518328666687)),(to_sfixed_a(0.1931643784046173)),(to_sfixed_a(0.36224162578582764)),(to_sfixed_a(-0.0416206531226635)),(to_sfixed_a(-0.06574772298336029)),(to_sfixed_a(-0.6296451091766357)),(to_sfixed_a(-0.09819938242435455)),(to_sfixed_a(-0.1745855063199997)),(to_sfixed_a(-0.12940625846385956)),(to_sfixed_a(-0.4643233120441437)),(to_sfixed_a(-0.046469464898109436)),(to_sfixed_a(-0.0011996770044788718)),(to_sfixed_a(-0.0010207847226411104)),(to_sfixed_a(-9.481099550612271e-05)),(to_sfixed_a(-4.820668436877895e-06)),(to_sfixed_a(8.453202462987974e-05)),(to_sfixed_a(0.00014279705646913499)),(to_sfixed_a(5.954031439614482e-05)),(to_sfixed_a(0.00012847040488850325)),(to_sfixed_a(-0.012260419316589832)),(to_sfixed_a(0.023635154590010643)),(to_sfixed_a(-0.1548001766204834)),(to_sfixed_a(0.06918363273143768)),(to_sfixed_a(-0.2191488891839981)),(to_sfixed_a(0.06587602198123932)),(to_sfixed_a(-0.06824245303869247)),(to_sfixed_a(0.11527277529239655)),(to_sfixed_a(0.12917280197143555)),(to_sfixed_a(0.28171613812446594)),(to_sfixed_a(0.218711256980896)),(to_sfixed_a(0.02392471581697464)),(to_sfixed_a(0.045307956635951996)),(to_sfixed_a(0.05586106330156326)),(to_sfixed_a(-0.2360992580652237)),(to_sfixed_a(-0.2909332513809204)),(to_sfixed_a(-0.21399465203285217)),(to_sfixed_a(-0.11793205887079239)),(to_sfixed_a(0.10441475361585617)),(to_sfixed_a(-0.0021528240758925676)),(to_sfixed_a(0.00045753279118798673)),(to_sfixed_a(0.000433504581451416)),(to_sfixed_a(-1.9550063370843418e-05)),(to_sfixed_a(-1.3668541214428842e-05)),(to_sfixed_a(-0.0001657638931646943)),(to_sfixed_a(0.00021714599279221147)),(to_sfixed_a(-0.00010078057675855234)),(to_sfixed_a(-0.06804337352514267)),(to_sfixed_a(-0.11550246924161911)),(to_sfixed_a(-0.15320667624473572)),(to_sfixed_a(-0.22379440069198608)),(to_sfixed_a(-0.3221435844898224)),(to_sfixed_a(-0.29117950797080994)),(to_sfixed_a(-0.19204263389110565)),(to_sfixed_a(-0.04805522412061691)),(to_sfixed_a(0.17502813041210175)),(to_sfixed_a(0.2407078742980957)),(to_sfixed_a(-0.037592608481645584)),(to_sfixed_a(0.1982152760028839)),(to_sfixed_a(0.1395387500524521)),(to_sfixed_a(0.1971089243888855)),(to_sfixed_a(0.0706084743142128)),(to_sfixed_a(-0.19277946650981903)),(to_sfixed_a(-0.17810994386672974)),(to_sfixed_a(-0.06268763542175293)),(to_sfixed_a(0.014036192558705807)),(to_sfixed_a(0.03179760277271271)),(to_sfixed_a(0.12812426686286926)),(to_sfixed_a(0.0007169125601649284)),(to_sfixed_a(5.357964982977137e-05)),(to_sfixed_a(-0.00012285365664865822)),(to_sfixed_a(0.00014444009866565466)),(to_sfixed_a(-4.888178955297917e-05)),(to_sfixed_a(0.0004004263610113412)),(to_sfixed_a(-0.0012610489502549171)),(to_sfixed_a(-0.06713616847991943)),(to_sfixed_a(-0.11528833210468292)),(to_sfixed_a(-0.27303147315979004)),(to_sfixed_a(-0.08495793491601944)),(to_sfixed_a(-0.24350379407405853)),(to_sfixed_a(-0.17078973352909088)),(to_sfixed_a(-0.0871969684958458)),(to_sfixed_a(-0.23288215696811676)),(to_sfixed_a(0.1000923365354538)),(to_sfixed_a(0.11369099467992783)),(to_sfixed_a(-0.009934375062584877)),(to_sfixed_a(0.20165406167507172)),(to_sfixed_a(0.20972391963005066)),(to_sfixed_a(0.17125995457172394)),(to_sfixed_a(-0.20264990627765656)),(to_sfixed_a(-0.2081654816865921)),(to_sfixed_a(-0.3270747661590576)),(to_sfixed_a(-0.3157344162464142)),(to_sfixed_a(-0.2575269639492035)),(to_sfixed_a(-0.21157510578632355)),(to_sfixed_a(0.00043812417425215244)),(to_sfixed_a(0.0003938322770409286)),(to_sfixed_a(-0.00022330551291815937)),(to_sfixed_a(0.0002719048352446407)),(to_sfixed_a(7.322433521039784e-05)),(to_sfixed_a(0.00018485740292817354)),(to_sfixed_a(-0.0004200237162876874)),(to_sfixed_a(-0.001161509775556624)),(to_sfixed_a(0.07134570926427841)),(to_sfixed_a(-0.045052431523799896)),(to_sfixed_a(-0.09645023941993713)),(to_sfixed_a(-0.13226447999477386)),(to_sfixed_a(-0.10821402817964554)),(to_sfixed_a(-0.06771770119667053)),(to_sfixed_a(-0.06071940064430237)),(to_sfixed_a(-0.1056700125336647)),(to_sfixed_a(-0.011107636615633965)),(to_sfixed_a(-0.23883502185344696)),(to_sfixed_a(-0.1956343948841095)),(to_sfixed_a(0.18213266134262085)),(to_sfixed_a(0.444266676902771)),(to_sfixed_a(-0.09865197539329529)),(to_sfixed_a(0.07040101289749146)),(to_sfixed_a(-0.0635942742228508)),(to_sfixed_a(0.18935778737068176)),(to_sfixed_a(-0.14509131014347076)),(to_sfixed_a(-0.06798356771469116)),(to_sfixed_a(0.00037357458495534956)),(to_sfixed_a(7.910021668067202e-05)),(to_sfixed_a(-6.521523027913645e-05)),(to_sfixed_a(3.9861824916442856e-05)),(to_sfixed_a(-0.00019364804029464722)),(to_sfixed_a(-0.00016032769053708762)),(to_sfixed_a(0.00015105555939953774)),(to_sfixed_a(-0.00045154025428928435)),(to_sfixed_a(0.008219867013394833)),(to_sfixed_a(0.1254035383462906)),(to_sfixed_a(-0.0026947648730129004)),(to_sfixed_a(0.09686443954706192)),(to_sfixed_a(0.0035705009941011667)),(to_sfixed_a(-0.11864917725324631)),(to_sfixed_a(-0.1273868978023529)),(to_sfixed_a(-0.07837755233049393)),(to_sfixed_a(0.11250346153974533)),(to_sfixed_a(-0.12508215010166168)),(to_sfixed_a(-0.05731174349784851)),(to_sfixed_a(0.07789064198732376)),(to_sfixed_a(0.12423841655254364)),(to_sfixed_a(0.17686788737773895)),(to_sfixed_a(-0.06150643527507782)),(to_sfixed_a(-0.12278342992067337)),(to_sfixed_a(-0.3745637834072113)),(to_sfixed_a(-0.1722583770751953)),(to_sfixed_a(-0.5033408999443054)),(to_sfixed_a(-0.06269601732492447)),(to_sfixed_a(-0.06708145141601562)),(to_sfixed_a(-0.005824373569339514)),(to_sfixed_a(-5.171444354346022e-05)),(to_sfixed_a(2.656702599779237e-05)),(to_sfixed_a(0.000178164045792073)),(to_sfixed_a(-0.0003347157617099583)),(to_sfixed_a(9.14238189579919e-05)),(to_sfixed_a(-1.4549264051311184e-05)),(to_sfixed_a(0.07673340290784836)),(to_sfixed_a(-0.0015036464901641011)),(to_sfixed_a(-0.16289718449115753)),(to_sfixed_a(0.0019509118283167481)),(to_sfixed_a(0.010706599801778793)),(to_sfixed_a(0.05222669616341591)),(to_sfixed_a(0.08773652464151382)),(to_sfixed_a(-0.046502236276865005)),(to_sfixed_a(-0.13808013498783112)),(to_sfixed_a(0.31899455189704895)),(to_sfixed_a(0.026815271005034447)),(to_sfixed_a(0.032920755445957184)),(to_sfixed_a(0.24765434861183167)),(to_sfixed_a(-0.014459755271673203)),(to_sfixed_a(-0.09530985355377197)),(to_sfixed_a(-0.1947789192199707)),(to_sfixed_a(-0.05553567036986351)),(to_sfixed_a(-0.10946419090032578)),(to_sfixed_a(-0.14182016253471375)),(to_sfixed_a(-0.17191585898399353)),(to_sfixed_a(-0.06321059912443161)),(to_sfixed_a(-8.566153701394796e-05)),(to_sfixed_a(2.1214253138168715e-05)),(to_sfixed_a(-0.00018223478400614113)),(to_sfixed_a(5.385353142628446e-05)),(to_sfixed_a(0.00028266868321225047)),(to_sfixed_a(5.6682124522922095e-06)),(to_sfixed_a(0.0002837134525179863)),(to_sfixed_a(-3.1465293432120234e-05)),(to_sfixed_a(0.006497920490801334)),(to_sfixed_a(0.007905940525233746)),(to_sfixed_a(0.10090084373950958)),(to_sfixed_a(-0.058926478028297424)),(to_sfixed_a(-0.048143479973077774)),(to_sfixed_a(-0.30792340636253357)),(to_sfixed_a(-0.07721257954835892)),(to_sfixed_a(-0.03299502283334732)),(to_sfixed_a(-0.11830353736877441)),(to_sfixed_a(-0.10906516760587692)),(to_sfixed_a(-0.1535053700208664)),(to_sfixed_a(-0.13003884255886078)),(to_sfixed_a(-0.1116548553109169)),(to_sfixed_a(-0.11774399131536484)),(to_sfixed_a(-0.4280914068222046)),(to_sfixed_a(-0.3865424394607544)),(to_sfixed_a(-0.4123353064060211)),(to_sfixed_a(-0.14851988852024078)),(to_sfixed_a(-0.03831741586327553)),(to_sfixed_a(-0.0930105447769165)),(to_sfixed_a(-0.07479733228683472)),(to_sfixed_a(-0.00012425325985532254)),(to_sfixed_a(4.043221633764915e-05)),(to_sfixed_a(2.5818200811045244e-05)),(to_sfixed_a(4.4109747250331566e-06)),(to_sfixed_a(3.06756301142741e-05)),(to_sfixed_a(-0.0001157484803115949)),(to_sfixed_a(2.3822401544748573e-06)),(to_sfixed_a(-0.022456839680671692)),(to_sfixed_a(-3.116795778623782e-05)),(to_sfixed_a(0.05228105187416077)),(to_sfixed_a(-0.04248904064297676)),(to_sfixed_a(0.0530475452542305)),(to_sfixed_a(-0.05738500505685806)),(to_sfixed_a(-0.04334885999560356)),(to_sfixed_a(-0.04363498091697693)),(to_sfixed_a(-0.131078839302063)),(to_sfixed_a(-0.03542352095246315)),(to_sfixed_a(-0.22769534587860107)),(to_sfixed_a(-0.09437961876392365)),(to_sfixed_a(-0.09940970689058304)),(to_sfixed_a(-0.25190848112106323)),(to_sfixed_a(-0.2855066657066345)),(to_sfixed_a(-0.2792110741138458)),(to_sfixed_a(-0.39567798376083374)),(to_sfixed_a(-0.0784459188580513)),(to_sfixed_a(-0.06058753654360771)),(to_sfixed_a(-7.192184421001002e-05)),(to_sfixed_a(-0.02404506504535675)),(to_sfixed_a(3.386203752597794e-05)),(to_sfixed_a(0.00025438351440243423)),(to_sfixed_a(-0.00020744539506267756)),(to_sfixed_a(-6.74906259519048e-05)),(to_sfixed_a(-2.953280636575073e-05)),(to_sfixed_a(0.0001267585321329534)),(to_sfixed_a(0.00013178130029700696)),(to_sfixed_a(7.793854456394911e-05)),(to_sfixed_a(-0.08406517654657364)),(to_sfixed_a(-0.027334172278642654)),(to_sfixed_a(0.0763900876045227)),(to_sfixed_a(0.06894358992576599)),(to_sfixed_a(-0.10066196322441101)),(to_sfixed_a(0.021947836503386497)),(to_sfixed_a(0.027107803151011467)),(to_sfixed_a(0.02169088087975979)),(to_sfixed_a(-0.08697565644979477)),(to_sfixed_a(-0.07342362403869629)),(to_sfixed_a(0.07876835018396378)),(to_sfixed_a(-0.06802720576524734)),(to_sfixed_a(-0.00315558142028749)),(to_sfixed_a(-0.4709527790546417)),(to_sfixed_a(-0.14915108680725098)),(to_sfixed_a(-0.042580895125865936)),(to_sfixed_a(-0.023520562797784805)),(to_sfixed_a(-0.03856196627020836)),(to_sfixed_a(-0.0011651146924123168)),(to_sfixed_a(3.205938992323354e-05)),(to_sfixed_a(1.2178494216641411e-05)),(to_sfixed_a(6.147510430309922e-05)),(to_sfixed_a(9.332823537988588e-05)),(to_sfixed_a(0.0001618341339053586)),(to_sfixed_a(-0.00019153555331286043)),(to_sfixed_a(-1.2857452020398341e-05)),(to_sfixed_a(0.00016769669309724122)),(to_sfixed_a(-0.00022266083396971226)),(to_sfixed_a(-0.011488557793200016)),(to_sfixed_a(0.10011261701583862)),(to_sfixed_a(-0.16493305563926697)),(to_sfixed_a(0.09074985980987549)),(to_sfixed_a(0.03586301952600479)),(to_sfixed_a(0.010635718703269958)),(to_sfixed_a(-0.047080039978027344)),(to_sfixed_a(-0.1314888745546341)),(to_sfixed_a(0.05424228310585022)),(to_sfixed_a(0.038520462810993195)),(to_sfixed_a(-0.0027468150947242975)),(to_sfixed_a(-0.29269134998321533)),(to_sfixed_a(-0.016299663111567497)),(to_sfixed_a(-0.13411159813404083)),(to_sfixed_a(-0.18638890981674194)),(to_sfixed_a(-0.0024033666122704744)),(to_sfixed_a(-0.02419973909854889)),(to_sfixed_a(-0.0026549750473350286)),(to_sfixed_a(-0.00877541396766901)),(to_sfixed_a(-4.6644574467791244e-05)),(to_sfixed_a(-5.7464603742118925e-05)),(to_sfixed_a(0.00015636705211363733)),(to_sfixed_a(0.00024633045541122556)),(to_sfixed_a(-2.276031591463834e-05)),(to_sfixed_a(-0.00012163039355073124)),(to_sfixed_a(-0.00011028915469069034)),(to_sfixed_a(9.574587602401152e-05)),(to_sfixed_a(-0.001151047763414681)),(to_sfixed_a(0.031601179391145706)),(to_sfixed_a(-0.004257158376276493)),(to_sfixed_a(-0.08434806764125824)),(to_sfixed_a(0.07570000737905502)),(to_sfixed_a(-0.06414542347192764)),(to_sfixed_a(-0.07661404460668564)),(to_sfixed_a(-0.15995290875434875)),(to_sfixed_a(0.04813404381275177)),(to_sfixed_a(0.025156661868095398)),(to_sfixed_a(-0.07880523800849915)),(to_sfixed_a(-0.10504601150751114)),(to_sfixed_a(-0.337491899728775)),(to_sfixed_a(-0.22513920068740845)),(to_sfixed_a(-0.10096415132284164)),(to_sfixed_a(-0.11284760385751724)),(to_sfixed_a(-0.009320194832980633)),(to_sfixed_a(-0.05159607157111168)),(to_sfixed_a(-0.007123782765120268)),(to_sfixed_a(0.002407516585662961)),(to_sfixed_a(0.0002308950643055141)),(to_sfixed_a(-0.0001180005565402098)),(to_sfixed_a(2.6016999981948175e-05)),(to_sfixed_a(8.85589251993224e-05)),(to_sfixed_a(7.189423922682181e-05)),(to_sfixed_a(-1.6114356185426004e-05)),(to_sfixed_a(-9.336380753666162e-05)),(to_sfixed_a(0.00012577345478348434)),(to_sfixed_a(-5.226022403803654e-05)),(to_sfixed_a(-0.012630220502614975)),(to_sfixed_a(-0.0035497762728482485)),(to_sfixed_a(0.02335815317928791)),(to_sfixed_a(-0.14552725851535797)),(to_sfixed_a(0.07352352887392044)),(to_sfixed_a(-0.017762428149580956)),(to_sfixed_a(-0.08391468971967697)),(to_sfixed_a(0.262164831161499)),(to_sfixed_a(-0.09919174015522003)),(to_sfixed_a(0.005554261151701212)),(to_sfixed_a(-0.09175453335046768)),(to_sfixed_a(-0.10866854339838028)),(to_sfixed_a(-0.08810370415449142)),(to_sfixed_a(-0.020008176565170288)),(to_sfixed_a(-0.0658775269985199)),(to_sfixed_a(-0.1332894265651703)),(to_sfixed_a(0.00043521783663891256)),(to_sfixed_a(-0.0008026102441363037)),(to_sfixed_a(-0.0006387089379131794)),(to_sfixed_a(-6.359385224641301e-06)),(to_sfixed_a(7.234516669996083e-05)),(to_sfixed_a(-8.230052480939776e-05)),(to_sfixed_a(0.00014695213758386672)),(to_sfixed_a(0.0002278978208778426)),(to_sfixed_a(-3.677606946439482e-05)),(to_sfixed_a(-0.0001900314528029412)),(to_sfixed_a(-9.13301992113702e-05)),(to_sfixed_a(8.053793862927705e-05)),(to_sfixed_a(-0.003653760300949216)),(to_sfixed_a(-0.003577382303774357)),(to_sfixed_a(0.0001749862713040784)),(to_sfixed_a(5.8916397392749786e-05)),(to_sfixed_a(-0.00020408810814842582)),(to_sfixed_a(-0.056399278342723846)),(to_sfixed_a(0.006911148317158222)),(to_sfixed_a(0.0008487740997225046)),(to_sfixed_a(-0.04605657234787941)),(to_sfixed_a(0.03530697897076607)),(to_sfixed_a(0.017112214118242264)),(to_sfixed_a(0.01223767176270485)),(to_sfixed_a(-0.04791608452796936)),(to_sfixed_a(-0.06695671379566193)),(to_sfixed_a(-0.002476373454555869)),(to_sfixed_a(-0.0012200456112623215)),(to_sfixed_a(-2.8399259463185444e-05)),(to_sfixed_a(0.00021620946063194424)),(to_sfixed_a(-5.492142736329697e-05)),(to_sfixed_a(0.0003375927626620978)),(to_sfixed_a(2.735570660661324e-06)),(to_sfixed_a(9.437272819923237e-05)),(to_sfixed_a(8.990825881483033e-05)),(to_sfixed_a(9.889450302580371e-05)),(to_sfixed_a(-0.00035305265919305384)),(to_sfixed_a(0.0003071081591770053)),(to_sfixed_a(5.3247789765009657e-05)),(to_sfixed_a(-3.068975274800323e-05)),(to_sfixed_a(0.00024292949819937348)),(to_sfixed_a(0.0002980482531711459)),(to_sfixed_a(-3.277371433796361e-05)),(to_sfixed_a(-2.725774720602203e-06)),(to_sfixed_a(1.9270788470748812e-05)),(to_sfixed_a(-0.00014452725008595735)),(to_sfixed_a(-0.0002331523282919079)),(to_sfixed_a(0.00011292680574115366)),(to_sfixed_a(-0.00013615888019558042)),(to_sfixed_a(6.901488086441532e-05)),(to_sfixed_a(5.9477479226188734e-05)),(to_sfixed_a(8.013081242097542e-05)),(to_sfixed_a(-0.00015570315008517355)),(to_sfixed_a(0.0002133841480826959)),(to_sfixed_a(-9.975777356885374e-05)),(to_sfixed_a(-3.7396275729406625e-05)),(to_sfixed_a(5.279316610540263e-06)),(to_sfixed_a(-7.453048601746559e-05)),(to_sfixed_a(-1.2240712749189697e-05)),(to_sfixed_a(1.2631498975679278e-05)),(to_sfixed_a(-2.622408646857366e-05)),(to_sfixed_a(-2.4338696675840765e-05)),(to_sfixed_a(-0.00016315981338266283)));

    constant weight_n0_8 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-8.027817239053547e-05)),(to_sfixed_a(-0.0001779182639438659)),(to_sfixed_a(5.740418782806955e-05)),(to_sfixed_a(-0.00025814620312303305)),(to_sfixed_a(-9.186509851133451e-05)),(to_sfixed_a(2.6639503630576655e-05)),(to_sfixed_a(-0.0001845584629336372)),(to_sfixed_a(-4.824778807233088e-05)),(to_sfixed_a(-0.00023897642677184194)),(to_sfixed_a(-0.00018504809122532606)),(to_sfixed_a(9.216705802828074e-05)),(to_sfixed_a(1.6507547115907073e-05)),(to_sfixed_a(0.00010208826279267669)),(to_sfixed_a(0.00016998180944938213)),(to_sfixed_a(-0.00019617821089923382)),(to_sfixed_a(-0.00048267285455949605)),(to_sfixed_a(2.5840496164164506e-05)),(to_sfixed_a(0.00020182691514492035)),(to_sfixed_a(-0.0002562941226642579)),(to_sfixed_a(0.0004087837296538055)),(to_sfixed_a(-4.7197198000503704e-05)),(to_sfixed_a(-0.00014404227840714157)),(to_sfixed_a(0.00024696276523172855)),(to_sfixed_a(1.226612221216783e-05)),(to_sfixed_a(6.771805055905133e-05)),(to_sfixed_a(-4.399612225824967e-05)),(to_sfixed_a(-2.176636189687997e-05)),(to_sfixed_a(8.427107241004705e-05)),(to_sfixed_a(0.00021097825083415955)),(to_sfixed_a(2.6043875550385565e-05)),(to_sfixed_a(-0.0001189934991998598)),(to_sfixed_a(-0.0002811859012581408)),(to_sfixed_a(0.00016162566316779703)),(to_sfixed_a(3.946093420381658e-05)),(to_sfixed_a(9.497901373833884e-06)),(to_sfixed_a(5.397526911110617e-05)),(to_sfixed_a(-3.799913974944502e-05)),(to_sfixed_a(0.0001257135154446587)),(to_sfixed_a(-9.464655886404216e-05)),(to_sfixed_a(4.4093849282944575e-05)),(to_sfixed_a(-9.405700984643772e-05)),(to_sfixed_a(2.3551599952043034e-05)),(to_sfixed_a(0.00010372180986450985)),(to_sfixed_a(-0.00016167579451575875)),(to_sfixed_a(-0.0002044605789706111)),(to_sfixed_a(-6.314524944173172e-05)),(to_sfixed_a(-0.00036887041642330587)),(to_sfixed_a(0.00012909685028716922)),(to_sfixed_a(-0.00013658481475431472)),(to_sfixed_a(-0.00013997517817188054)),(to_sfixed_a(0.00027171007241122425)),(to_sfixed_a(4.9372676585335284e-05)),(to_sfixed_a(0.0003522112383507192)),(to_sfixed_a(0.0001524869294371456)),(to_sfixed_a(0.00010658948303898796)),(to_sfixed_a(-5.3170097089605406e-05)),(to_sfixed_a(7.492223085137084e-05)),(to_sfixed_a(-4.486854959395714e-05)),(to_sfixed_a(-7.909085979918018e-05)),(to_sfixed_a(-0.00010061285138363019)),(to_sfixed_a(0.00012849748600274324)),(to_sfixed_a(0.0001566547289257869)),(to_sfixed_a(3.6630935937864706e-05)),(to_sfixed_a(-4.7846915549598634e-06)),(to_sfixed_a(0.00010781432501971722)),(to_sfixed_a(-0.0003331504121888429)),(to_sfixed_a(-0.0001195521472254768)),(to_sfixed_a(-0.00019619782688096166)),(to_sfixed_a(4.3569885747274384e-05)),(to_sfixed_a(0.011020860634744167)),(to_sfixed_a(3.076966822845861e-05)),(to_sfixed_a(0.000162653173902072)),(to_sfixed_a(5.355858593247831e-05)),(to_sfixed_a(-3.372194623807445e-05)),(to_sfixed_a(5.5694526963634416e-05)),(to_sfixed_a(-1.9777546640398214e-06)),(to_sfixed_a(0.00020608775957953185)),(to_sfixed_a(-4.59186703665182e-05)),(to_sfixed_a(1.4373334124684334e-05)),(to_sfixed_a(5.575160321313888e-05)),(to_sfixed_a(3.587512401281856e-05)),(to_sfixed_a(2.9665543479495682e-05)),(to_sfixed_a(-5.877104194951244e-05)),(to_sfixed_a(-0.00019848087686114013)),(to_sfixed_a(-0.0002135978575097397)),(to_sfixed_a(6.153613503556699e-05)),(to_sfixed_a(-0.0001702152512734756)),(to_sfixed_a(0.00026331402477808297)),(to_sfixed_a(8.78728533280082e-05)),(to_sfixed_a(0.00028003082843497396)),(to_sfixed_a(0.0001556509087095037)),(to_sfixed_a(2.405181476206053e-05)),(to_sfixed_a(-0.08078541606664658)),(to_sfixed_a(-0.00016070243145804852)),(to_sfixed_a(-0.09161288291215897)),(to_sfixed_a(-0.17467063665390015)),(to_sfixed_a(-0.18177583813667297)),(to_sfixed_a(-0.06182728335261345)),(to_sfixed_a(-0.1119978204369545)),(to_sfixed_a(0.28234177827835083)),(to_sfixed_a(0.009207000024616718)),(to_sfixed_a(0.28833022713661194)),(to_sfixed_a(-0.08212126046419144)),(to_sfixed_a(0.11142493039369583)),(to_sfixed_a(0.049404338002204895)),(to_sfixed_a(0.10024593025445938)),(to_sfixed_a(-0.00011789436393883079)),(to_sfixed_a(-0.00010733901581261307)),(to_sfixed_a(-9.842697909334674e-05)),(to_sfixed_a(0.00010008479875978082)),(to_sfixed_a(-0.00021051095973234624)),(to_sfixed_a(0.00012853452062699944)),(to_sfixed_a(0.0002455800131428987)),(to_sfixed_a(1.7961961930268444e-05)),(to_sfixed_a(0.0002695558359846473)),(to_sfixed_a(0.00012826766760554165)),(to_sfixed_a(-0.00022364968026522547)),(to_sfixed_a(-2.0172825315967202e-05)),(to_sfixed_a(-0.0006271810852922499)),(to_sfixed_a(-0.09615956246852875)),(to_sfixed_a(-0.017966289073228836)),(to_sfixed_a(-0.11767257750034332)),(to_sfixed_a(-0.7011717557907104)),(to_sfixed_a(-0.09309080243110657)),(to_sfixed_a(-0.19433963298797607)),(to_sfixed_a(0.11252090334892273)),(to_sfixed_a(0.1564398556947708)),(to_sfixed_a(0.15618158876895905)),(to_sfixed_a(0.2134656012058258)),(to_sfixed_a(-0.16935224831104279)),(to_sfixed_a(-0.2538347840309143)),(to_sfixed_a(-0.021581510081887245)),(to_sfixed_a(-0.0031187995336949825)),(to_sfixed_a(-0.17778758704662323)),(to_sfixed_a(-0.006902165245264769)),(to_sfixed_a(-0.00021243821538519114)),(to_sfixed_a(-0.0011646868661046028)),(to_sfixed_a(0.0002409973822068423)),(to_sfixed_a(0.0001248340413440019)),(to_sfixed_a(-4.1428203985560685e-05)),(to_sfixed_a(0.00027174269780516624)),(to_sfixed_a(3.1713407224742696e-05)),(to_sfixed_a(0.0003357250243425369)),(to_sfixed_a(-0.00010746165935415775)),(to_sfixed_a(-4.2041832784889266e-05)),(to_sfixed_a(-0.1517234593629837)),(to_sfixed_a(-0.011248617433011532)),(to_sfixed_a(-0.028102710843086243)),(to_sfixed_a(-0.17534901201725006)),(to_sfixed_a(-0.1997665911912918)),(to_sfixed_a(-0.1149665117263794)),(to_sfixed_a(-0.20275941491127014)),(to_sfixed_a(-0.22584104537963867)),(to_sfixed_a(-0.0620703399181366)),(to_sfixed_a(0.19334882497787476)),(to_sfixed_a(0.2323833703994751)),(to_sfixed_a(-0.05149143934249878)),(to_sfixed_a(-0.4161478579044342)),(to_sfixed_a(-0.1731647104024887)),(to_sfixed_a(-0.002387840999290347)),(to_sfixed_a(-0.05736016482114792)),(to_sfixed_a(-0.04405727609992027)),(to_sfixed_a(-0.0007115720654837787)),(to_sfixed_a(0.048811424523591995)),(to_sfixed_a(-0.00031317578395828605)),(to_sfixed_a(-0.0004189342726022005)),(to_sfixed_a(-3.381946589797735e-05)),(to_sfixed_a(0.00026083545526489615)),(to_sfixed_a(0.00014005131379235536)),(to_sfixed_a(-0.00017895929340738803)),(to_sfixed_a(7.588130756630562e-06)),(to_sfixed_a(-7.86831442383118e-05)),(to_sfixed_a(8.81154410308227e-05)),(to_sfixed_a(-0.14387045800685883)),(to_sfixed_a(-0.12975527346134186)),(to_sfixed_a(-0.556299090385437)),(to_sfixed_a(-0.48441460728645325)),(to_sfixed_a(-0.7182724475860596)),(to_sfixed_a(0.045874737203121185)),(to_sfixed_a(-0.07186654955148697)),(to_sfixed_a(0.1632237434387207)),(to_sfixed_a(0.1572737693786621)),(to_sfixed_a(0.44198834896087646)),(to_sfixed_a(0.4876742959022522)),(to_sfixed_a(-0.22163107991218567)),(to_sfixed_a(0.02060130052268505)),(to_sfixed_a(0.29920247197151184)),(to_sfixed_a(0.05382338911294937)),(to_sfixed_a(-0.1409807652235031)),(to_sfixed_a(0.019876761361956596)),(to_sfixed_a(0.14768141508102417)),(to_sfixed_a(0.19828002154827118)),(to_sfixed_a(-0.0026223058812320232)),(to_sfixed_a(-0.003024761565029621)),(to_sfixed_a(-0.0023569397162646055)),(to_sfixed_a(0.00022078704205341637)),(to_sfixed_a(-2.2274178263614886e-05)),(to_sfixed_a(0.00016296170360874385)),(to_sfixed_a(8.430145680904388e-05)),(to_sfixed_a(3.457403363427147e-05)),(to_sfixed_a(3.746154470718466e-05)),(to_sfixed_a(0.02955366112291813)),(to_sfixed_a(-0.16036242246627808)),(to_sfixed_a(-0.09708157926797867)),(to_sfixed_a(-0.3421209156513214)),(to_sfixed_a(-0.2801368534564972)),(to_sfixed_a(0.08756493031978607)),(to_sfixed_a(-0.1990489661693573)),(to_sfixed_a(-0.06811004132032394)),(to_sfixed_a(0.7129780054092407)),(to_sfixed_a(0.4165950119495392)),(to_sfixed_a(0.31673502922058105)),(to_sfixed_a(0.04154481366276741)),(to_sfixed_a(-0.08922003209590912)),(to_sfixed_a(0.03524917736649513)),(to_sfixed_a(0.06333241611719131)),(to_sfixed_a(-0.1026851236820221)),(to_sfixed_a(0.07407710701227188)),(to_sfixed_a(0.06054156646132469)),(to_sfixed_a(0.5685696601867676)),(to_sfixed_a(0.04864312335848808)),(to_sfixed_a(0.00794818252325058)),(to_sfixed_a(8.673813863424584e-05)),(to_sfixed_a(-3.70552770618815e-05)),(to_sfixed_a(0.00011697788431774825)),(to_sfixed_a(-3.9224243664648384e-05)),(to_sfixed_a(0.0003286535502411425)),(to_sfixed_a(8.794433961156756e-05)),(to_sfixed_a(-0.041264086961746216)),(to_sfixed_a(-0.15671060979366302)),(to_sfixed_a(0.07520901411771774)),(to_sfixed_a(-0.11069347709417343)),(to_sfixed_a(-0.21786683797836304)),(to_sfixed_a(-0.24283422529697418)),(to_sfixed_a(-0.35243159532546997)),(to_sfixed_a(0.16225220263004303)),(to_sfixed_a(0.2669175863265991)),(to_sfixed_a(0.4781559407711029)),(to_sfixed_a(0.5245923399925232)),(to_sfixed_a(0.2934834063053131)),(to_sfixed_a(-0.07727329432964325)),(to_sfixed_a(0.07692364603281021)),(to_sfixed_a(0.03254340589046478)),(to_sfixed_a(-0.01359505020081997)),(to_sfixed_a(0.14410124719142914)),(to_sfixed_a(0.13891243934631348)),(to_sfixed_a(0.2851096987724304)),(to_sfixed_a(0.16256839036941528)),(to_sfixed_a(0.14331622421741486)),(to_sfixed_a(0.004907465539872646)),(to_sfixed_a(-0.00014459695375990123)),(to_sfixed_a(6.011580626363866e-05)),(to_sfixed_a(-0.00032415249734185636)),(to_sfixed_a(8.403517858823761e-05)),(to_sfixed_a(4.78928122902289e-05)),(to_sfixed_a(-6.961406324990094e-05)),(to_sfixed_a(0.002237249631434679)),(to_sfixed_a(0.015567705035209656)),(to_sfixed_a(-0.0024424628354609013)),(to_sfixed_a(-0.13583189249038696)),(to_sfixed_a(-0.10283530503511429)),(to_sfixed_a(-0.08587870746850967)),(to_sfixed_a(0.05081258341670036)),(to_sfixed_a(0.23851323127746582)),(to_sfixed_a(0.4842953681945801)),(to_sfixed_a(0.76866614818573)),(to_sfixed_a(0.4823560416698456)),(to_sfixed_a(-0.030311839655041695)),(to_sfixed_a(-0.5008273124694824)),(to_sfixed_a(-0.5381326079368591)),(to_sfixed_a(-0.42552855610847473)),(to_sfixed_a(-0.6226681470870972)),(to_sfixed_a(-0.3197179436683655)),(to_sfixed_a(-0.30572161078453064)),(to_sfixed_a(-0.28368425369262695)),(to_sfixed_a(-0.10885647684335709)),(to_sfixed_a(0.12236594408750534)),(to_sfixed_a(-2.9668135539395735e-05)),(to_sfixed_a(-0.00027452618815004826)),(to_sfixed_a(-9.540147584630176e-05)),(to_sfixed_a(0.00024935483816079795)),(to_sfixed_a(1.29570025819703e-05)),(to_sfixed_a(7.446909876307473e-05)),(to_sfixed_a(0.00011774688755394891)),(to_sfixed_a(0.013044779188930988)),(to_sfixed_a(0.08437395840883255)),(to_sfixed_a(0.25982794165611267)),(to_sfixed_a(0.3009050190448761)),(to_sfixed_a(0.22840452194213867)),(to_sfixed_a(0.10736849904060364)),(to_sfixed_a(0.22447188198566437)),(to_sfixed_a(0.12869253754615784)),(to_sfixed_a(0.4112175703048706)),(to_sfixed_a(0.6899430751800537)),(to_sfixed_a(0.3793645203113556)),(to_sfixed_a(0.05639728158712387)),(to_sfixed_a(-0.3695269525051117)),(to_sfixed_a(-0.4614432752132416)),(to_sfixed_a(-0.5522042512893677)),(to_sfixed_a(-0.4737744629383087)),(to_sfixed_a(-0.3010529577732086)),(to_sfixed_a(-0.12292661517858505)),(to_sfixed_a(0.002818579552695155)),(to_sfixed_a(0.026453200727701187)),(to_sfixed_a(0.07985007017850876)),(to_sfixed_a(0.006362683139741421)),(to_sfixed_a(-7.464875670848414e-05)),(to_sfixed_a(-4.711801739176735e-05)),(to_sfixed_a(-0.00011325920786475763)),(to_sfixed_a(8.995865937322378e-05)),(to_sfixed_a(3.62815881089773e-05)),(to_sfixed_a(-0.04035695642232895)),(to_sfixed_a(0.023896558210253716)),(to_sfixed_a(0.3059476912021637)),(to_sfixed_a(0.3121967911720276)),(to_sfixed_a(0.36185145378112793)),(to_sfixed_a(-0.08879035711288452)),(to_sfixed_a(0.015307598747313023)),(to_sfixed_a(0.020576495677232742)),(to_sfixed_a(0.21530646085739136)),(to_sfixed_a(0.15436390042304993)),(to_sfixed_a(0.22765441238880157)),(to_sfixed_a(0.075535848736763)),(to_sfixed_a(-0.17826586961746216)),(to_sfixed_a(-0.09556742757558823)),(to_sfixed_a(-0.3273387849330902)),(to_sfixed_a(-0.5068155527114868)),(to_sfixed_a(-0.36059147119522095)),(to_sfixed_a(-0.2924594283103943)),(to_sfixed_a(-0.11332210898399353)),(to_sfixed_a(0.0463075116276741)),(to_sfixed_a(-0.19829832017421722)),(to_sfixed_a(0.005659584421664476)),(to_sfixed_a(-4.199136310489848e-05)),(to_sfixed_a(1.633891588426195e-05)),(to_sfixed_a(0.0001919768692459911)),(to_sfixed_a(4.260774949216284e-05)),(to_sfixed_a(0.00011939335672650486)),(to_sfixed_a(0.0002288015530211851)),(to_sfixed_a(-0.00018184476357419044)),(to_sfixed_a(0.13552691042423248)),(to_sfixed_a(-0.045893337577581406)),(to_sfixed_a(0.14886093139648438)),(to_sfixed_a(0.021573368459939957)),(to_sfixed_a(-0.00926445797085762)),(to_sfixed_a(-0.11625827103853226)),(to_sfixed_a(-0.16001783311367035)),(to_sfixed_a(-0.14510378241539001)),(to_sfixed_a(-0.2676658034324646)),(to_sfixed_a(0.03806082904338837)),(to_sfixed_a(-0.0012495683040469885)),(to_sfixed_a(0.11646775901317596)),(to_sfixed_a(0.06568120419979095)),(to_sfixed_a(-0.09350109100341797)),(to_sfixed_a(0.011775967665016651)),(to_sfixed_a(-0.12358946353197098)),(to_sfixed_a(-0.2982068359851837)),(to_sfixed_a(-0.1540437787771225)),(to_sfixed_a(-0.16024206578731537)),(to_sfixed_a(0.12140175700187683)),(to_sfixed_a(0.11625214666128159)),(to_sfixed_a(7.90160265751183e-05)),(to_sfixed_a(0.00015732081374153495)),(to_sfixed_a(-3.371978164068423e-05)),(to_sfixed_a(0.00010481235949555412)),(to_sfixed_a(-4.6877743443474174e-05)),(to_sfixed_a(4.275551327737048e-05)),(to_sfixed_a(0.00031153627787716687)),(to_sfixed_a(-0.027184659615159035)),(to_sfixed_a(0.15268179774284363)),(to_sfixed_a(-0.11761797219514847)),(to_sfixed_a(-0.30198872089385986)),(to_sfixed_a(-0.21292829513549805)),(to_sfixed_a(-0.34781408309936523)),(to_sfixed_a(-0.21041446924209595)),(to_sfixed_a(-0.04454375430941582)),(to_sfixed_a(0.15455219149589539)),(to_sfixed_a(-0.16284964978694916)),(to_sfixed_a(0.02305419184267521)),(to_sfixed_a(0.06729012727737427)),(to_sfixed_a(0.05948716029524803)),(to_sfixed_a(0.07601951062679291)),(to_sfixed_a(0.02502073347568512)),(to_sfixed_a(0.03701478987932205)),(to_sfixed_a(0.20156456530094147)),(to_sfixed_a(-0.03558020666241646)),(to_sfixed_a(-0.05588063225150108)),(to_sfixed_a(-0.19943904876708984)),(to_sfixed_a(-0.10163155198097229)),(to_sfixed_a(0.0005640725721605122)),(to_sfixed_a(0.0018905358156189322)),(to_sfixed_a(-0.00026352255372330546)),(to_sfixed_a(2.974546623590868e-05)),(to_sfixed_a(0.0002692940179258585)),(to_sfixed_a(3.189139533787966e-05)),(to_sfixed_a(-0.00021047583140898496)),(to_sfixed_a(-0.0009155725711025298)),(to_sfixed_a(-0.14569368958473206)),(to_sfixed_a(-0.15581609308719635)),(to_sfixed_a(-0.37259119749069214)),(to_sfixed_a(-0.2764037549495697)),(to_sfixed_a(-0.3186235725879669)),(to_sfixed_a(0.0367971770465374)),(to_sfixed_a(-0.05951705202460289)),(to_sfixed_a(-0.01092727854847908)),(to_sfixed_a(-0.24742738902568817)),(to_sfixed_a(-0.06558740139007568)),(to_sfixed_a(-0.003217325545847416)),(to_sfixed_a(0.053841035813093185)),(to_sfixed_a(0.002392788417637348)),(to_sfixed_a(0.11535030603408813)),(to_sfixed_a(-0.03340040147304535)),(to_sfixed_a(-0.002634804928675294)),(to_sfixed_a(-0.004447621293365955)),(to_sfixed_a(-0.12185931950807571)),(to_sfixed_a(-0.05371568724513054)),(to_sfixed_a(-0.04951867088675499)),(to_sfixed_a(-0.0001165943467640318)),(to_sfixed_a(0.0003563273057807237)),(to_sfixed_a(-0.00022465281654149294)),(to_sfixed_a(0.00014331942657008767)),(to_sfixed_a(-0.0005632569082081318)),(to_sfixed_a(-3.928426303900778e-05)),(to_sfixed_a(0.0002565465110819787)),(to_sfixed_a(-0.040273137390613556)),(to_sfixed_a(-0.11071103066205978)),(to_sfixed_a(0.09592203795909882)),(to_sfixed_a(0.12930911779403687)),(to_sfixed_a(0.2021220624446869)),(to_sfixed_a(0.16709047555923462)),(to_sfixed_a(0.236394464969635)),(to_sfixed_a(-0.10748069733381271)),(to_sfixed_a(0.019447142258286476)),(to_sfixed_a(-0.09571422636508942)),(to_sfixed_a(0.06682126969099045)),(to_sfixed_a(0.0863458663225174)),(to_sfixed_a(0.009240134619176388)),(to_sfixed_a(0.05834579840302467)),(to_sfixed_a(-0.028581062331795692)),(to_sfixed_a(0.03520772606134415)),(to_sfixed_a(-0.15142671763896942)),(to_sfixed_a(-0.07015594094991684)),(to_sfixed_a(-0.029134739190340042)),(to_sfixed_a(-0.19702684879302979)),(to_sfixed_a(-0.04448448494076729)),(to_sfixed_a(-0.0005737764877267182)),(to_sfixed_a(-0.0002234861603938043)),(to_sfixed_a(-0.0003496047283988446)),(to_sfixed_a(0.00010953433957183734)),(to_sfixed_a(-4.8240872274618596e-05)),(to_sfixed_a(0.0002268858952447772)),(to_sfixed_a(0.004698226228356361)),(to_sfixed_a(0.07585379481315613)),(to_sfixed_a(0.14959150552749634)),(to_sfixed_a(0.07225265353918076)),(to_sfixed_a(0.3143567144870758)),(to_sfixed_a(0.24709834158420563)),(to_sfixed_a(0.32133394479751587)),(to_sfixed_a(0.23610781133174896)),(to_sfixed_a(0.038994304835796356)),(to_sfixed_a(0.14143253862857819)),(to_sfixed_a(0.04270223155617714)),(to_sfixed_a(0.01667257584631443)),(to_sfixed_a(0.045291777700185776)),(to_sfixed_a(-0.060839466750621796)),(to_sfixed_a(-0.1461976170539856)),(to_sfixed_a(-0.010714891366660595)),(to_sfixed_a(-0.16326439380645752)),(to_sfixed_a(-0.19518034160137177)),(to_sfixed_a(-0.08035564422607422)),(to_sfixed_a(-0.06185542047023773)),(to_sfixed_a(-0.13863752782344818)),(to_sfixed_a(-0.09958904981613159)),(to_sfixed_a(-0.004123803693801165)),(to_sfixed_a(-1.7857870261650532e-05)),(to_sfixed_a(9.519092418486252e-05)),(to_sfixed_a(5.427095675258897e-05)),(to_sfixed_a(0.00017348004621453583)),(to_sfixed_a(0.002985199447721243)),(to_sfixed_a(0.004755242727696896)),(to_sfixed_a(0.10239151120185852)),(to_sfixed_a(0.2315390557050705)),(to_sfixed_a(0.15036430954933167)),(to_sfixed_a(0.19012276828289032)),(to_sfixed_a(0.28702861070632935)),(to_sfixed_a(0.22712348401546478)),(to_sfixed_a(0.26321539282798767)),(to_sfixed_a(0.2253301739692688)),(to_sfixed_a(0.14943070709705353)),(to_sfixed_a(0.23359835147857666)),(to_sfixed_a(-0.012846832163631916)),(to_sfixed_a(0.0970199853181839)),(to_sfixed_a(-0.16728636622428894)),(to_sfixed_a(-0.09643810242414474)),(to_sfixed_a(-0.16287937760353088)),(to_sfixed_a(-0.25423818826675415)),(to_sfixed_a(0.11846332252025604)),(to_sfixed_a(-0.08140550553798676)),(to_sfixed_a(-0.15437497198581696)),(to_sfixed_a(0.010326811112463474)),(to_sfixed_a(-5.0579801609274e-05)),(to_sfixed_a(-8.048825111472979e-05)),(to_sfixed_a(-0.0001597562659299001)),(to_sfixed_a(-6.306709838099778e-05)),(to_sfixed_a(0.00020263523038011044)),(to_sfixed_a(-9.639812196837738e-05)),(to_sfixed_a(-0.00015006888133939356)),(to_sfixed_a(-0.0030187941156327724)),(to_sfixed_a(-0.0426642969250679)),(to_sfixed_a(0.2538605332374573)),(to_sfixed_a(0.0940888375043869)),(to_sfixed_a(0.1584448218345642)),(to_sfixed_a(0.02178931050002575)),(to_sfixed_a(0.20554450154304504)),(to_sfixed_a(0.04982622712850571)),(to_sfixed_a(0.04041607305407524)),(to_sfixed_a(0.061211250722408295)),(to_sfixed_a(0.0770256295800209)),(to_sfixed_a(-0.028099901974201202)),(to_sfixed_a(0.13047830760478973)),(to_sfixed_a(-0.03811338543891907)),(to_sfixed_a(-0.20216800272464752)),(to_sfixed_a(-0.10954176634550095)),(to_sfixed_a(-0.19945548474788666)),(to_sfixed_a(-0.0016539905918762088)),(to_sfixed_a(-0.2442111223936081)),(to_sfixed_a(-0.11811548471450806)),(to_sfixed_a(-0.09139206260442734)),(to_sfixed_a(-0.0052703064866364)),(to_sfixed_a(4.229539990774356e-05)),(to_sfixed_a(6.494222361652646e-06)),(to_sfixed_a(-8.871745376382023e-05)),(to_sfixed_a(9.234805474989116e-06)),(to_sfixed_a(4.199198428977979e-06)),(to_sfixed_a(1.3521933396987151e-05)),(to_sfixed_a(-0.057482264935970306)),(to_sfixed_a(0.0024564487393945456)),(to_sfixed_a(-0.1271660327911377)),(to_sfixed_a(0.02500057779252529)),(to_sfixed_a(0.06727729737758636)),(to_sfixed_a(0.10315429419279099)),(to_sfixed_a(-0.00967432837933302)),(to_sfixed_a(-0.14684626460075378)),(to_sfixed_a(-0.35393214225769043)),(to_sfixed_a(0.02372077852487564)),(to_sfixed_a(-0.113378144800663)),(to_sfixed_a(0.03391969949007034)),(to_sfixed_a(0.04643351957201958)),(to_sfixed_a(-0.06949333101511002)),(to_sfixed_a(-0.16337022185325623)),(to_sfixed_a(-0.12947224080562592)),(to_sfixed_a(-0.06279558688402176)),(to_sfixed_a(-0.061449430882930756)),(to_sfixed_a(-0.03742947056889534)),(to_sfixed_a(-0.0668795257806778)),(to_sfixed_a(0.045685525983572006)),(to_sfixed_a(-0.0001381884649163112)),(to_sfixed_a(-0.00018256356997881085)),(to_sfixed_a(0.00016304271412082016)),(to_sfixed_a(3.069380181841552e-05)),(to_sfixed_a(-0.0002074139192700386)),(to_sfixed_a(4.555857231025584e-05)),(to_sfixed_a(-0.00010505444515729323)),(to_sfixed_a(-0.00010109585855389014)),(to_sfixed_a(0.015489491634070873)),(to_sfixed_a(0.12183120101690292)),(to_sfixed_a(0.10964648425579071)),(to_sfixed_a(0.07481341809034348)),(to_sfixed_a(0.07392612844705582)),(to_sfixed_a(-0.06958829611539841)),(to_sfixed_a(-0.021879572421312332)),(to_sfixed_a(-0.2538294494152069)),(to_sfixed_a(0.02977737970650196)),(to_sfixed_a(-0.000529878365341574)),(to_sfixed_a(-0.014969836920499802)),(to_sfixed_a(0.00503853615373373)),(to_sfixed_a(0.05125783383846283)),(to_sfixed_a(-0.06008857488632202)),(to_sfixed_a(-0.061911869794130325)),(to_sfixed_a(-0.20730042457580566)),(to_sfixed_a(-0.15691089630126953)),(to_sfixed_a(-0.026667539030313492)),(to_sfixed_a(-0.011850769631564617)),(to_sfixed_a(-0.08611395210027695)),(to_sfixed_a(-0.08550362288951874)),(to_sfixed_a(-0.000158897673827596)),(to_sfixed_a(7.33094202587381e-05)),(to_sfixed_a(-1.8190528862760402e-05)),(to_sfixed_a(-9.823583241086453e-05)),(to_sfixed_a(-5.681643960997462e-05)),(to_sfixed_a(0.00025100994389504194)),(to_sfixed_a(-2.1177040252950974e-05)),(to_sfixed_a(0.053290434181690216)),(to_sfixed_a(0.0008318062173202634)),(to_sfixed_a(-0.060596100986003876)),(to_sfixed_a(0.06228536367416382)),(to_sfixed_a(0.0023856009356677532)),(to_sfixed_a(0.14174631237983704)),(to_sfixed_a(0.029624460265040398)),(to_sfixed_a(0.10758674889802933)),(to_sfixed_a(0.013456042855978012)),(to_sfixed_a(0.0433175154030323)),(to_sfixed_a(0.12478252500295639)),(to_sfixed_a(0.04704807698726654)),(to_sfixed_a(-0.008375264704227448)),(to_sfixed_a(0.087699756026268)),(to_sfixed_a(-0.10170037299394608)),(to_sfixed_a(-0.0665561631321907)),(to_sfixed_a(-0.0856349840760231)),(to_sfixed_a(-0.010252485983073711)),(to_sfixed_a(0.14618924260139465)),(to_sfixed_a(0.000805896648671478)),(to_sfixed_a(-0.0042138416320085526)),(to_sfixed_a(1.5232901205308735e-05)),(to_sfixed_a(-1.620156763237901e-05)),(to_sfixed_a(-5.612206587102264e-05)),(to_sfixed_a(0.0003437938285060227)),(to_sfixed_a(-0.0002118271659128368)),(to_sfixed_a(1.4453060430241749e-05)),(to_sfixed_a(0.0001293635432375595)),(to_sfixed_a(0.000379089149646461)),(to_sfixed_a(-0.03481822833418846)),(to_sfixed_a(0.06324080377817154)),(to_sfixed_a(0.2710548937320709)),(to_sfixed_a(0.065520741045475)),(to_sfixed_a(-0.060365814715623856)),(to_sfixed_a(0.07234593480825424)),(to_sfixed_a(0.002992567140609026)),(to_sfixed_a(0.059311751276254654)),(to_sfixed_a(0.046737123280763626)),(to_sfixed_a(0.0289025716483593)),(to_sfixed_a(-0.05940721929073334)),(to_sfixed_a(0.09493078291416168)),(to_sfixed_a(-0.051221128553152084)),(to_sfixed_a(-0.12114138156175613)),(to_sfixed_a(0.07168672978878021)),(to_sfixed_a(0.04611385613679886)),(to_sfixed_a(-0.010156574659049511)),(to_sfixed_a(-0.018577808514237404)),(to_sfixed_a(-0.0017082494450733066)),(to_sfixed_a(0.00041056584450416267)),(to_sfixed_a(9.734800551086664e-05)),(to_sfixed_a(0.00020440870139282197)),(to_sfixed_a(7.787944923620671e-05)),(to_sfixed_a(-0.0001174578137579374)),(to_sfixed_a(-1.266894832951948e-05)),(to_sfixed_a(0.0001445391826564446)),(to_sfixed_a(1.4940547771402635e-05)),(to_sfixed_a(0.0005648066871799529)),(to_sfixed_a(0.003788106609135866)),(to_sfixed_a(-0.006981207989156246)),(to_sfixed_a(-0.13855257630348206)),(to_sfixed_a(0.005440525710582733)),(to_sfixed_a(0.09004515409469604)),(to_sfixed_a(-0.004522812087088823)),(to_sfixed_a(0.21670225262641907)),(to_sfixed_a(0.1554996818304062)),(to_sfixed_a(0.11489054560661316)),(to_sfixed_a(0.19023139774799347)),(to_sfixed_a(0.21182164549827576)),(to_sfixed_a(-0.10320553183555603)),(to_sfixed_a(0.2549281418323517)),(to_sfixed_a(0.02867971919476986)),(to_sfixed_a(-0.003656096290796995)),(to_sfixed_a(0.11629167199134827)),(to_sfixed_a(0.11945617944002151)),(to_sfixed_a(0.009482979774475098)),(to_sfixed_a(0.08716142922639847)),(to_sfixed_a(-0.00013678795949090272)),(to_sfixed_a(-0.00013785585178993642)),(to_sfixed_a(-7.213825301732868e-05)),(to_sfixed_a(9.697264613350853e-05)),(to_sfixed_a(-5.646575300488621e-05)),(to_sfixed_a(8.319252083310857e-05)),(to_sfixed_a(-2.325079003639985e-05)),(to_sfixed_a(0.00014321778144221753)),(to_sfixed_a(-0.018854163587093353)),(to_sfixed_a(-0.00896712951362133)),(to_sfixed_a(-0.07912164181470871)),(to_sfixed_a(-0.0022232651244848967)),(to_sfixed_a(-0.09749948233366013)),(to_sfixed_a(0.09541607648134232)),(to_sfixed_a(-0.09476964175701141)),(to_sfixed_a(0.06639360636472702)),(to_sfixed_a(0.21705414354801178)),(to_sfixed_a(0.19019092619419098)),(to_sfixed_a(-0.14306072890758514)),(to_sfixed_a(-0.0871240571141243)),(to_sfixed_a(-0.17280052602291107)),(to_sfixed_a(-0.056078143417835236)),(to_sfixed_a(-0.02279525250196457)),(to_sfixed_a(0.09797167032957077)),(to_sfixed_a(-0.0041624088771641254)),(to_sfixed_a(0.09272401034832001)),(to_sfixed_a(0.06811824440956116)),(to_sfixed_a(0.025739433243870735)),(to_sfixed_a(-5.716251507692505e-06)),(to_sfixed_a(-0.0004169595777057111)),(to_sfixed_a(-0.0003707119030877948)),(to_sfixed_a(-0.0003377805114723742)),(to_sfixed_a(0.00024829150061123073)),(to_sfixed_a(2.1199766706558876e-05)),(to_sfixed_a(-2.830201992765069e-05)),(to_sfixed_a(0.00016572648019064218)),(to_sfixed_a(-0.00012666317343246192)),(to_sfixed_a(-0.01558313425630331)),(to_sfixed_a(-0.04761633649468422)),(to_sfixed_a(-0.12347226589918137)),(to_sfixed_a(-0.01605394296348095)),(to_sfixed_a(0.06539206951856613)),(to_sfixed_a(-0.03423783928155899)),(to_sfixed_a(0.1309618204832077)),(to_sfixed_a(0.08485568314790726)),(to_sfixed_a(0.04658433422446251)),(to_sfixed_a(0.05882592126727104)),(to_sfixed_a(0.0033865340519696474)),(to_sfixed_a(0.15037359297275543)),(to_sfixed_a(0.0845896452665329)),(to_sfixed_a(0.02357003651559353)),(to_sfixed_a(0.1850147843360901)),(to_sfixed_a(0.3425489068031311)),(to_sfixed_a(0.0011587276821956038)),(to_sfixed_a(0.007617767434567213)),(to_sfixed_a(0.008761908859014511)),(to_sfixed_a(8.410366717725992e-06)),(to_sfixed_a(-0.00014018680667504668)),(to_sfixed_a(8.208499639295042e-05)),(to_sfixed_a(0.0001767755748005584)),(to_sfixed_a(0.000467666337499395)),(to_sfixed_a(-0.00043778461986221373)),(to_sfixed_a(0.00014023251424077898)),(to_sfixed_a(4.20839660364436e-06)),(to_sfixed_a(-0.0001223614817718044)),(to_sfixed_a(-0.0022083919029682875)),(to_sfixed_a(-0.0023850887082517147)),(to_sfixed_a(-0.0002003631816478446)),(to_sfixed_a(0.00026368076214566827)),(to_sfixed_a(0.0001884228113340214)),(to_sfixed_a(0.11912243813276291)),(to_sfixed_a(-0.002161689568310976)),(to_sfixed_a(-0.00015445776807609946)),(to_sfixed_a(0.08741314709186554)),(to_sfixed_a(0.0007930469000712037)),(to_sfixed_a(-0.00456821545958519)),(to_sfixed_a(0.05431560426950455)),(to_sfixed_a(0.09510636329650879)),(to_sfixed_a(0.13544996082782745)),(to_sfixed_a(0.0140537079423666)),(to_sfixed_a(0.006125984247773886)),(to_sfixed_a(-3.511572867864743e-05)),(to_sfixed_a(-0.000213828549021855)),(to_sfixed_a(8.768396219238639e-05)),(to_sfixed_a(-0.00013636561925522983)),(to_sfixed_a(-0.0002747252583503723)),(to_sfixed_a(-3.6587043723557144e-05)),(to_sfixed_a(-0.00015296867059078068)),(to_sfixed_a(-0.00015683681704103947)),(to_sfixed_a(5.030681859352626e-05)),(to_sfixed_a(2.444674464641139e-05)),(to_sfixed_a(-0.00024439216940663755)),(to_sfixed_a(1.7297563317697495e-05)),(to_sfixed_a(0.0002132506633643061)),(to_sfixed_a(-0.00020707417570520192)),(to_sfixed_a(5.391117520048283e-05)),(to_sfixed_a(7.106327393557876e-05)),(to_sfixed_a(8.422850805800408e-05)),(to_sfixed_a(0.00023877638159319758)),(to_sfixed_a(-0.00016648462042212486)),(to_sfixed_a(0.0001660399866523221)),(to_sfixed_a(-0.00019109982531517744)),(to_sfixed_a(1.704659553070087e-05)),(to_sfixed_a(-2.0835492250625975e-05)),(to_sfixed_a(6.01816936978139e-05)),(to_sfixed_a(-0.00013794911501463503)),(to_sfixed_a(7.430370897054672e-05)),(to_sfixed_a(-0.00016928237164393067)),(to_sfixed_a(3.31060764438007e-05)),(to_sfixed_a(0.00023217200941871852)),(to_sfixed_a(-0.00029575263033621013)),(to_sfixed_a(-6.348107854137197e-05)),(to_sfixed_a(-8.15338862594217e-05)),(to_sfixed_a(7.34271498004091e-06)),(to_sfixed_a(-7.191274926299229e-05)),(to_sfixed_a(-4.2393953663122375e-06)));

    constant weight_n0_9 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(2.0984269212931395e-05)),(to_sfixed_a(1.4450354683503974e-05)),(to_sfixed_a(-0.00011874364281538874)),(to_sfixed_a(-0.00010843716881936416)),(to_sfixed_a(-0.00017418591596651822)),(to_sfixed_a(2.7874164516106248e-05)),(to_sfixed_a(-5.119626621308271e-06)),(to_sfixed_a(0.00013752795348409563)),(to_sfixed_a(-0.00011551416537258774)),(to_sfixed_a(0.00012296324712224305)),(to_sfixed_a(-5.880647677258821e-06)),(to_sfixed_a(-7.352302054641768e-05)),(to_sfixed_a(0.00014514864597003907)),(to_sfixed_a(-0.00018547331274021417)),(to_sfixed_a(0.00021044156164862216)),(to_sfixed_a(0.00012719916412606835)),(to_sfixed_a(0.00023778261675033718)),(to_sfixed_a(-8.311334386235103e-05)),(to_sfixed_a(-6.035900514689274e-05)),(to_sfixed_a(-0.00010982232925016433)),(to_sfixed_a(0.00022390371304936707)),(to_sfixed_a(-0.000430155050707981)),(to_sfixed_a(0.00017130687774624676)),(to_sfixed_a(0.0001248455373570323)),(to_sfixed_a(-0.00026373527362011373)),(to_sfixed_a(-7.540236401837319e-05)),(to_sfixed_a(-9.352347115054727e-05)),(to_sfixed_a(-0.00026651768712326884)),(to_sfixed_a(0.00019470010010991246)),(to_sfixed_a(0.00010700813436415046)),(to_sfixed_a(0.00010046739771496505)),(to_sfixed_a(0.00012148469249950722)),(to_sfixed_a(8.779398922342807e-05)),(to_sfixed_a(-0.0001231069618370384)),(to_sfixed_a(0.00011515461665112525)),(to_sfixed_a(0.00020865126862190664)),(to_sfixed_a(7.036617898847908e-05)),(to_sfixed_a(0.00011818778148153797)),(to_sfixed_a(8.522471034666523e-05)),(to_sfixed_a(-5.89160435993108e-06)),(to_sfixed_a(4.4085256377002224e-05)),(to_sfixed_a(0.00015205328236334026)),(to_sfixed_a(0.00029637670377269387)),(to_sfixed_a(-7.082163210725412e-05)),(to_sfixed_a(0.00024358952941838652)),(to_sfixed_a(5.4290492698783055e-05)),(to_sfixed_a(-9.271472663385794e-06)),(to_sfixed_a(2.1876796381548047e-05)),(to_sfixed_a(-6.91647655912675e-05)),(to_sfixed_a(4.472670116228983e-05)),(to_sfixed_a(-1.1331709174555726e-05)),(to_sfixed_a(0.00011861546954605728)),(to_sfixed_a(2.1009727788623422e-05)),(to_sfixed_a(9.539982420392334e-05)),(to_sfixed_a(-0.000127259103464894)),(to_sfixed_a(-0.00012367728049866855)),(to_sfixed_a(-0.00031561136711388826)),(to_sfixed_a(0.0001334719854639843)),(to_sfixed_a(-0.0001664679730311036)),(to_sfixed_a(-1.9465747755020857e-05)),(to_sfixed_a(7.63673015171662e-05)),(to_sfixed_a(0.00014440531958825886)),(to_sfixed_a(-0.00026126729790121317)),(to_sfixed_a(6.00382627453655e-05)),(to_sfixed_a(-7.423589067911962e-06)),(to_sfixed_a(-9.486687486059964e-05)),(to_sfixed_a(5.817870260216296e-05)),(to_sfixed_a(0.00020815845346078277)),(to_sfixed_a(1.1249320778006222e-05)),(to_sfixed_a(0.0013031598646193743)),(to_sfixed_a(-0.00013160076923668385)),(to_sfixed_a(-1.4674506928713527e-05)),(to_sfixed_a(-6.868323544040322e-05)),(to_sfixed_a(-0.00017264786583837122)),(to_sfixed_a(-3.2904001272981986e-05)),(to_sfixed_a(-6.385637789207976e-06)),(to_sfixed_a(-0.00018364543211646378)),(to_sfixed_a(-7.018325413810089e-05)),(to_sfixed_a(0.00012218303163535893)),(to_sfixed_a(-8.544189768144861e-05)),(to_sfixed_a(-0.00016006742953322828)),(to_sfixed_a(-1.9592938770074397e-05)),(to_sfixed_a(-4.816171349375509e-05)),(to_sfixed_a(-3.5760811442742124e-05)),(to_sfixed_a(-0.0001357859291601926)),(to_sfixed_a(-2.8174263206892647e-06)),(to_sfixed_a(-0.00011727963283192366)),(to_sfixed_a(-0.00029104796703904867)),(to_sfixed_a(0.0001980755478143692)),(to_sfixed_a(9.266090637538582e-05)),(to_sfixed_a(-8.363906090380624e-05)),(to_sfixed_a(0.0002642099279910326)),(to_sfixed_a(-0.018702000379562378)),(to_sfixed_a(-1.7540909539093263e-05)),(to_sfixed_a(-0.02109602652490139)),(to_sfixed_a(-0.01988104172050953)),(to_sfixed_a(0.0029106508009135723)),(to_sfixed_a(0.05991661176085472)),(to_sfixed_a(0.005812405608594418)),(to_sfixed_a(-0.061825934797525406)),(to_sfixed_a(0.02856607362627983)),(to_sfixed_a(-0.07536963373422623)),(to_sfixed_a(0.3225984573364258)),(to_sfixed_a(-0.05069710314273834)),(to_sfixed_a(-0.03094135783612728)),(to_sfixed_a(-0.062476761639118195)),(to_sfixed_a(3.36375851475168e-05)),(to_sfixed_a(-5.4546075261896476e-05)),(to_sfixed_a(-8.659232116769999e-05)),(to_sfixed_a(-3.675838161143474e-05)),(to_sfixed_a(0.00011876533972099423)),(to_sfixed_a(0.00015111347602214664)),(to_sfixed_a(-6.255455809878185e-05)),(to_sfixed_a(-0.00011350140266586095)),(to_sfixed_a(-0.00019848020747303963)),(to_sfixed_a(0.00010420253238407895)),(to_sfixed_a(-7.294574606930837e-05)),(to_sfixed_a(0.00019042800704482943)),(to_sfixed_a(0.0003911272797267884)),(to_sfixed_a(-0.011408815160393715)),(to_sfixed_a(-0.014564640820026398)),(to_sfixed_a(-0.02955162711441517)),(to_sfixed_a(-0.631264865398407)),(to_sfixed_a(-0.17742152512073517)),(to_sfixed_a(0.16370248794555664)),(to_sfixed_a(0.3179040253162384)),(to_sfixed_a(0.3204334080219269)),(to_sfixed_a(0.005373596679419279)),(to_sfixed_a(0.1774224191904068)),(to_sfixed_a(-0.032730650156736374)),(to_sfixed_a(0.05738150328397751)),(to_sfixed_a(-0.03958498686552048)),(to_sfixed_a(0.009546798653900623)),(to_sfixed_a(0.09731633961200714)),(to_sfixed_a(-0.02146962471306324)),(to_sfixed_a(4.030067793792114e-05)),(to_sfixed_a(-0.0008172827656380832)),(to_sfixed_a(0.0002065750741166994)),(to_sfixed_a(-0.000157345668412745)),(to_sfixed_a(0.0002840676752384752)),(to_sfixed_a(6.613949517486617e-05)),(to_sfixed_a(1.1753514627343975e-05)),(to_sfixed_a(-0.00010286768520018086)),(to_sfixed_a(-0.00010537898924667388)),(to_sfixed_a(0.0013359898002818227)),(to_sfixed_a(-0.020725497975945473)),(to_sfixed_a(-0.004109921399503946)),(to_sfixed_a(-0.2022199034690857)),(to_sfixed_a(0.001972166821360588)),(to_sfixed_a(-0.039628297090530396)),(to_sfixed_a(0.040633611381053925)),(to_sfixed_a(-0.08476667106151581)),(to_sfixed_a(0.3133244812488556)),(to_sfixed_a(0.10671508312225342)),(to_sfixed_a(-0.0024058306589722633)),(to_sfixed_a(-0.1810886263847351)),(to_sfixed_a(0.254666268825531)),(to_sfixed_a(0.006910430733114481)),(to_sfixed_a(0.4862278997898102)),(to_sfixed_a(0.12040764093399048)),(to_sfixed_a(0.31083640456199646)),(to_sfixed_a(0.22086875140666962)),(to_sfixed_a(-0.0001595369540154934)),(to_sfixed_a(-0.06561823934316635)),(to_sfixed_a(-0.00035320065217092633)),(to_sfixed_a(-2.181562922487501e-05)),(to_sfixed_a(-0.00017285504145547748)),(to_sfixed_a(-0.00013487219985108823)),(to_sfixed_a(3.2133171771420166e-05)),(to_sfixed_a(9.683562893769704e-06)),(to_sfixed_a(-0.00017102411948144436)),(to_sfixed_a(-9.980829054256901e-05)),(to_sfixed_a(2.4983653474919265e-06)),(to_sfixed_a(-0.018656127154827118)),(to_sfixed_a(-0.0020954704377800226)),(to_sfixed_a(-0.03841428831219673)),(to_sfixed_a(-0.17428447306156158)),(to_sfixed_a(-0.2877950370311737)),(to_sfixed_a(0.16472406685352325)),(to_sfixed_a(-0.03433908149600029)),(to_sfixed_a(0.09395178407430649)),(to_sfixed_a(-0.06427812576293945)),(to_sfixed_a(0.029936932027339935)),(to_sfixed_a(0.12502051889896393)),(to_sfixed_a(-0.15587542951107025)),(to_sfixed_a(0.0010675224475562572)),(to_sfixed_a(0.24697494506835938)),(to_sfixed_a(0.37759438157081604)),(to_sfixed_a(0.5107161402702332)),(to_sfixed_a(-0.012105444446206093)),(to_sfixed_a(0.20453768968582153)),(to_sfixed_a(0.16211800277233124)),(to_sfixed_a(0.0033039364498108625)),(to_sfixed_a(0.004768497310578823)),(to_sfixed_a(0.002471987856552005)),(to_sfixed_a(-0.0001312729000346735)),(to_sfixed_a(-0.00022549797722604126)),(to_sfixed_a(1.9273851648904383e-05)),(to_sfixed_a(-9.530072929919697e-06)),(to_sfixed_a(4.585004717228003e-06)),(to_sfixed_a(0.00013821732136420906)),(to_sfixed_a(0.002267307136207819)),(to_sfixed_a(0.013799455016851425)),(to_sfixed_a(0.004145369399338961)),(to_sfixed_a(-0.042501673102378845)),(to_sfixed_a(0.01656114123761654)),(to_sfixed_a(0.00669997651129961)),(to_sfixed_a(0.09634711593389511)),(to_sfixed_a(0.2417265623807907)),(to_sfixed_a(-0.2180083692073822)),(to_sfixed_a(-0.4259404242038727)),(to_sfixed_a(-0.33683523535728455)),(to_sfixed_a(-0.22216321527957916)),(to_sfixed_a(0.013819589279592037)),(to_sfixed_a(0.4069550037384033)),(to_sfixed_a(0.4606263041496277)),(to_sfixed_a(0.28964900970458984)),(to_sfixed_a(0.278142511844635)),(to_sfixed_a(0.06763570010662079)),(to_sfixed_a(0.1365336924791336)),(to_sfixed_a(0.0654519647359848)),(to_sfixed_a(0.002077357843518257)),(to_sfixed_a(-0.00017355747695546597)),(to_sfixed_a(-0.00013899691111873835)),(to_sfixed_a(1.4195946278050542e-05)),(to_sfixed_a(3.491920142550953e-05)),(to_sfixed_a(0.00022187376453075558)),(to_sfixed_a(3.477687869235524e-06)),(to_sfixed_a(-0.003414195030927658)),(to_sfixed_a(0.0423286147415638)),(to_sfixed_a(-0.003106127493083477)),(to_sfixed_a(-0.04369984567165375)),(to_sfixed_a(-0.6213170289993286)),(to_sfixed_a(-0.051106758415699005)),(to_sfixed_a(-0.029287410899996758)),(to_sfixed_a(-0.196283757686615)),(to_sfixed_a(0.14211662113666534)),(to_sfixed_a(-0.21992605924606323)),(to_sfixed_a(-0.6460056900978088)),(to_sfixed_a(-0.6827647686004639)),(to_sfixed_a(-0.5365216732025146)),(to_sfixed_a(-0.2372266948223114)),(to_sfixed_a(0.43960586190223694)),(to_sfixed_a(0.37675273418426514)),(to_sfixed_a(-0.17606692016124725)),(to_sfixed_a(0.22737610340118408)),(to_sfixed_a(0.08226215839385986)),(to_sfixed_a(-0.026382438838481903)),(to_sfixed_a(0.031115982681512833)),(to_sfixed_a(-0.013257330283522606)),(to_sfixed_a(4.391116453916766e-05)),(to_sfixed_a(0.00012443296145647764)),(to_sfixed_a(4.6112891141092405e-05)),(to_sfixed_a(0.00013203101116232574)),(to_sfixed_a(-0.0001753647084115073)),(to_sfixed_a(0.00016491132555529475)),(to_sfixed_a(-0.003829676192253828)),(to_sfixed_a(-0.050400957465171814)),(to_sfixed_a(-0.05937657877802849)),(to_sfixed_a(-0.19433185458183289)),(to_sfixed_a(-0.18555988371372223)),(to_sfixed_a(-0.0034415211994200945)),(to_sfixed_a(-0.057579156011343)),(to_sfixed_a(0.39031872153282166)),(to_sfixed_a(0.3618676960468292)),(to_sfixed_a(-0.09392976015806198)),(to_sfixed_a(-0.47232088446617126)),(to_sfixed_a(-0.7437951564788818)),(to_sfixed_a(-0.5834929943084717)),(to_sfixed_a(-0.37823519110679626)),(to_sfixed_a(0.16353212296962738)),(to_sfixed_a(0.45227766036987305)),(to_sfixed_a(0.5510830879211426)),(to_sfixed_a(-0.05377049744129181)),(to_sfixed_a(0.0015218165935948491)),(to_sfixed_a(0.13531583547592163)),(to_sfixed_a(-0.0024724549148231745)),(to_sfixed_a(-0.00016866762598510832)),(to_sfixed_a(-6.907482747919858e-05)),(to_sfixed_a(-3.176855170750059e-05)),(to_sfixed_a(-6.261494854697958e-05)),(to_sfixed_a(-0.0001622113777557388)),(to_sfixed_a(-0.00022211510804481804)),(to_sfixed_a(-0.00024189293617382646)),(to_sfixed_a(-0.001496839802712202)),(to_sfixed_a(0.009257839992642403)),(to_sfixed_a(0.04148666560649872)),(to_sfixed_a(-0.011289683170616627)),(to_sfixed_a(0.08498148620128632)),(to_sfixed_a(-0.22850291430950165)),(to_sfixed_a(0.18747468292713165)),(to_sfixed_a(0.2952699363231659)),(to_sfixed_a(0.17280876636505127)),(to_sfixed_a(0.06312423199415207)),(to_sfixed_a(-0.46002912521362305)),(to_sfixed_a(-0.5041407346725464)),(to_sfixed_a(-0.3323698043823242)),(to_sfixed_a(0.012131883762776852)),(to_sfixed_a(0.14102210104465485)),(to_sfixed_a(0.37914860248565674)),(to_sfixed_a(0.33102837204933167)),(to_sfixed_a(0.09345311671495438)),(to_sfixed_a(0.07576829940080643)),(to_sfixed_a(-0.03632107377052307)),(to_sfixed_a(-0.009735851548612118)),(to_sfixed_a(-0.040622565895318985)),(to_sfixed_a(-0.00021344788547139615)),(to_sfixed_a(0.00012257517664693296)),(to_sfixed_a(0.0002534123486839235)),(to_sfixed_a(-5.614766996586695e-05)),(to_sfixed_a(0.00021317928622011095)),(to_sfixed_a(-0.0037288509774953127)),(to_sfixed_a(-0.01446612924337387)),(to_sfixed_a(0.0005287356907501817)),(to_sfixed_a(0.02094174176454544)),(to_sfixed_a(0.054096415638923645)),(to_sfixed_a(-0.03861235827207565)),(to_sfixed_a(-0.03308403491973877)),(to_sfixed_a(0.11495181173086166)),(to_sfixed_a(0.18543463945388794)),(to_sfixed_a(0.19752176105976105)),(to_sfixed_a(-0.13490194082260132)),(to_sfixed_a(-0.3595799505710602)),(to_sfixed_a(-0.43932515382766724)),(to_sfixed_a(-0.21890750527381897)),(to_sfixed_a(0.3427281081676483)),(to_sfixed_a(0.6671648025512695)),(to_sfixed_a(0.3735533058643341)),(to_sfixed_a(0.40875837206840515)),(to_sfixed_a(0.3305959701538086)),(to_sfixed_a(0.07106751203536987)),(to_sfixed_a(0.004491683095693588)),(to_sfixed_a(0.07634502649307251)),(to_sfixed_a(0.00010018133616540581)),(to_sfixed_a(1.676039391895756e-05)),(to_sfixed_a(0.0002769230050034821)),(to_sfixed_a(-7.91212878539227e-05)),(to_sfixed_a(-0.00020923494594171643)),(to_sfixed_a(-6.0164624301251024e-05)),(to_sfixed_a(-0.0001634021318750456)),(to_sfixed_a(0.05665719509124756)),(to_sfixed_a(0.04971706494688988)),(to_sfixed_a(0.016946133226156235)),(to_sfixed_a(0.12172510474920273)),(to_sfixed_a(0.1793559491634369)),(to_sfixed_a(0.12433163821697235)),(to_sfixed_a(0.30782899260520935)),(to_sfixed_a(0.2350776642560959)),(to_sfixed_a(-0.04054134339094162)),(to_sfixed_a(-0.03698946535587311)),(to_sfixed_a(-0.1824275106191635)),(to_sfixed_a(-0.20833539962768555)),(to_sfixed_a(0.19689282774925232)),(to_sfixed_a(0.2568875551223755)),(to_sfixed_a(0.06425287574529648)),(to_sfixed_a(0.39954033493995667)),(to_sfixed_a(0.37924957275390625)),(to_sfixed_a(0.06291631609201431)),(to_sfixed_a(0.007976638153195381)),(to_sfixed_a(0.10115905851125717)),(to_sfixed_a(0.03167270869016647)),(to_sfixed_a(7.461529094143771e-06)),(to_sfixed_a(-0.0002779635542538017)),(to_sfixed_a(0.00018788882880471647)),(to_sfixed_a(-0.00011946378799621016)),(to_sfixed_a(0.0003127158561255783)),(to_sfixed_a(-5.15900319442153e-05)),(to_sfixed_a(-0.0001858925970736891)),(to_sfixed_a(-0.011776714585721493)),(to_sfixed_a(0.09778256714344025)),(to_sfixed_a(0.02881789021193981)),(to_sfixed_a(0.03979605436325073)),(to_sfixed_a(-0.009028258733451366)),(to_sfixed_a(-0.0885571613907814)),(to_sfixed_a(0.04352394491434097)),(to_sfixed_a(0.10436410456895828)),(to_sfixed_a(0.08658342808485031)),(to_sfixed_a(-0.14595872163772583)),(to_sfixed_a(-0.011142627336084843)),(to_sfixed_a(0.11622395366430283)),(to_sfixed_a(-0.14575035870075226)),(to_sfixed_a(0.16881337761878967)),(to_sfixed_a(-0.005745599512010813)),(to_sfixed_a(0.02941901609301567)),(to_sfixed_a(-0.32737624645233154)),(to_sfixed_a(0.11445077508687973)),(to_sfixed_a(-0.07719989120960236)),(to_sfixed_a(-0.05024467036128044)),(to_sfixed_a(-0.021829264238476753)),(to_sfixed_a(0.002045055152848363)),(to_sfixed_a(0.0004855548031628132)),(to_sfixed_a(-0.00014539618859998882)),(to_sfixed_a(-0.0003515417920425534)),(to_sfixed_a(6.777081580366939e-06)),(to_sfixed_a(-0.00020043364202138036)),(to_sfixed_a(-0.00021649232076015323)),(to_sfixed_a(-0.0009310093591921031)),(to_sfixed_a(0.21719591319561005)),(to_sfixed_a(0.04877357557415962)),(to_sfixed_a(-0.15103358030319214)),(to_sfixed_a(-0.24143126606941223)),(to_sfixed_a(-0.11936268955469131)),(to_sfixed_a(-0.09162009507417679)),(to_sfixed_a(-0.16786924004554749)),(to_sfixed_a(-0.03343626484274864)),(to_sfixed_a(0.10930871963500977)),(to_sfixed_a(0.10641175508499146)),(to_sfixed_a(0.15213137865066528)),(to_sfixed_a(0.04973196983337402)),(to_sfixed_a(0.08986075222492218)),(to_sfixed_a(0.0390046201646328)),(to_sfixed_a(-0.0697411298751831)),(to_sfixed_a(0.023041866719722748)),(to_sfixed_a(-0.38850709795951843)),(to_sfixed_a(-0.14053769409656525)),(to_sfixed_a(-0.1746940165758133)),(to_sfixed_a(-0.005955874919891357)),(to_sfixed_a(0.00045844350825063884)),(to_sfixed_a(8.555433305446059e-05)),(to_sfixed_a(0.0002489033213350922)),(to_sfixed_a(0.00014403133536688983)),(to_sfixed_a(-5.565236642723903e-05)),(to_sfixed_a(-3.21338557114359e-05)),(to_sfixed_a(6.127417145762593e-05)),(to_sfixed_a(-0.029583698138594627)),(to_sfixed_a(-0.00946820992976427)),(to_sfixed_a(-0.03499195724725723)),(to_sfixed_a(-0.03610072284936905)),(to_sfixed_a(0.11527960002422333)),(to_sfixed_a(0.12147944420576096)),(to_sfixed_a(0.03424306586384773)),(to_sfixed_a(-0.11662568151950836)),(to_sfixed_a(-0.048810750246047974)),(to_sfixed_a(0.07063447684049606)),(to_sfixed_a(0.3134717643260956)),(to_sfixed_a(0.04199019819498062)),(to_sfixed_a(0.13110989332199097)),(to_sfixed_a(0.04347928985953331)),(to_sfixed_a(0.008465904742479324)),(to_sfixed_a(-0.0317060612142086)),(to_sfixed_a(-0.32235196232795715)),(to_sfixed_a(-0.07232104241847992)),(to_sfixed_a(0.044763799756765366)),(to_sfixed_a(-0.09217216074466705)),(to_sfixed_a(-0.06538510322570801)),(to_sfixed_a(0.00015407183673232794)),(to_sfixed_a(-1.7343393210467184e-07)),(to_sfixed_a(7.469718548236415e-05)),(to_sfixed_a(0.00031914535793475807)),(to_sfixed_a(-7.197829836513847e-05)),(to_sfixed_a(-7.366644422290847e-05)),(to_sfixed_a(0.0006876631523482502)),(to_sfixed_a(-0.04136122390627861)),(to_sfixed_a(0.06939348578453064)),(to_sfixed_a(0.09410711377859116)),(to_sfixed_a(-0.0916588082909584)),(to_sfixed_a(0.04077325761318207)),(to_sfixed_a(0.13789135217666626)),(to_sfixed_a(0.12995684146881104)),(to_sfixed_a(0.34944188594818115)),(to_sfixed_a(0.23229162395000458)),(to_sfixed_a(0.12144459038972855)),(to_sfixed_a(0.03510760888457298)),(to_sfixed_a(0.012507162988185883)),(to_sfixed_a(0.12204281985759735)),(to_sfixed_a(0.06873692572116852)),(to_sfixed_a(0.07486354559659958)),(to_sfixed_a(-0.21091768145561218)),(to_sfixed_a(-0.5204569101333618)),(to_sfixed_a(0.0025739704724401236)),(to_sfixed_a(-0.09358549118041992)),(to_sfixed_a(0.0499739870429039)),(to_sfixed_a(-0.04327015578746796)),(to_sfixed_a(-0.010522586293518543)),(to_sfixed_a(0.00011266724322922528)),(to_sfixed_a(-0.00015159128815867007)),(to_sfixed_a(6.289011798799038e-05)),(to_sfixed_a(0.00017305449000559747)),(to_sfixed_a(0.0007256733952090144)),(to_sfixed_a(0.0008053512428887188)),(to_sfixed_a(0.04465043917298317)),(to_sfixed_a(0.03669056296348572)),(to_sfixed_a(0.01259776670485735)),(to_sfixed_a(0.09483347088098526)),(to_sfixed_a(0.1356746256351471)),(to_sfixed_a(0.16482502222061157)),(to_sfixed_a(0.4569224715232849)),(to_sfixed_a(0.22519497573375702)),(to_sfixed_a(0.01349696610122919)),(to_sfixed_a(-0.07698123902082443)),(to_sfixed_a(-0.08794842660427094)),(to_sfixed_a(0.16041520237922668)),(to_sfixed_a(0.1518973559141159)),(to_sfixed_a(0.12358413636684418)),(to_sfixed_a(0.0630841851234436)),(to_sfixed_a(-0.10439164191484451)),(to_sfixed_a(-0.36949780583381653)),(to_sfixed_a(-0.13432885706424713)),(to_sfixed_a(-0.30724331736564636)),(to_sfixed_a(-0.019284743815660477)),(to_sfixed_a(-5.210647577769123e-05)),(to_sfixed_a(2.2596905182581395e-05)),(to_sfixed_a(0.00026811595307663083)),(to_sfixed_a(0.00032510593882761896)),(to_sfixed_a(-0.00018147507216781378)),(to_sfixed_a(0.0001280872238567099)),(to_sfixed_a(0.000317530328175053)),(to_sfixed_a(0.026213163509964943)),(to_sfixed_a(-0.027477959170937538)),(to_sfixed_a(-0.16384483873844147)),(to_sfixed_a(-0.08090198040008545)),(to_sfixed_a(0.03719954937696457)),(to_sfixed_a(0.06615559011697769)),(to_sfixed_a(0.035326868295669556)),(to_sfixed_a(0.16059863567352295)),(to_sfixed_a(0.24201075732707977)),(to_sfixed_a(-0.04983896389603615)),(to_sfixed_a(0.1669536679983139)),(to_sfixed_a(0.08840806782245636)),(to_sfixed_a(0.13014918565750122)),(to_sfixed_a(0.10767149925231934)),(to_sfixed_a(0.16411492228507996)),(to_sfixed_a(-0.11438430100679398)),(to_sfixed_a(-0.0943465605378151)),(to_sfixed_a(-0.10676519572734833)),(to_sfixed_a(-0.4683811068534851)),(to_sfixed_a(-0.0916210263967514)),(to_sfixed_a(-0.04020664468407631)),(to_sfixed_a(-0.004293912090361118)),(to_sfixed_a(0.00014430185547098517)),(to_sfixed_a(-3.917693538824096e-05)),(to_sfixed_a(0.00019756000256165862)),(to_sfixed_a(7.68805475672707e-05)),(to_sfixed_a(0.00012824279838241637)),(to_sfixed_a(-7.031495624687523e-05)),(to_sfixed_a(-0.056117404252290726)),(to_sfixed_a(0.0015416996320709586)),(to_sfixed_a(0.0005622218013741076)),(to_sfixed_a(-0.02763138711452484)),(to_sfixed_a(-0.1574217826128006)),(to_sfixed_a(-0.27757972478866577)),(to_sfixed_a(-0.21206936240196228)),(to_sfixed_a(-0.11814286559820175)),(to_sfixed_a(-0.07519955188035965)),(to_sfixed_a(-0.16998539865016937)),(to_sfixed_a(-0.048207223415374756)),(to_sfixed_a(0.1203199177980423)),(to_sfixed_a(0.015041577629745007)),(to_sfixed_a(-0.029417164623737335)),(to_sfixed_a(0.10642988979816437)),(to_sfixed_a(-0.048209305852651596)),(to_sfixed_a(0.0015209827106446028)),(to_sfixed_a(-0.10648325085639954)),(to_sfixed_a(-0.1726040244102478)),(to_sfixed_a(-0.12488718330860138)),(to_sfixed_a(-0.15863114595413208)),(to_sfixed_a(0.0001322549069300294)),(to_sfixed_a(-0.00013467943063005805)),(to_sfixed_a(0.00012008997873635963)),(to_sfixed_a(-3.3168831578223035e-05)),(to_sfixed_a(-9.596122981747612e-05)),(to_sfixed_a(-0.00019309007620904595)),(to_sfixed_a(4.5862834667786956e-05)),(to_sfixed_a(-8.323565270984545e-05)),(to_sfixed_a(-0.0076998146250844)),(to_sfixed_a(-0.052750032395124435)),(to_sfixed_a(0.015501749701797962)),(to_sfixed_a(-0.1594611257314682)),(to_sfixed_a(0.05982198938727379)),(to_sfixed_a(-0.1090826764702797)),(to_sfixed_a(0.03399135172367096)),(to_sfixed_a(-0.191840261220932)),(to_sfixed_a(-0.2013935148715973)),(to_sfixed_a(-0.2592604160308838)),(to_sfixed_a(-0.09158999472856522)),(to_sfixed_a(0.041802383959293365)),(to_sfixed_a(0.05940045788884163)),(to_sfixed_a(0.09135983884334564)),(to_sfixed_a(0.009680072776973248)),(to_sfixed_a(-0.05017872154712677)),(to_sfixed_a(-0.453713059425354)),(to_sfixed_a(-0.13648952543735504)),(to_sfixed_a(-0.1983257532119751)),(to_sfixed_a(-0.1537737250328064)),(to_sfixed_a(-0.0359644778072834)),(to_sfixed_a(0.00018305022967979312)),(to_sfixed_a(-6.6524458816275e-05)),(to_sfixed_a(-0.00011229654046474025)),(to_sfixed_a(-7.334447582252324e-05)),(to_sfixed_a(-0.00014009176811669022)),(to_sfixed_a(0.0002498575486242771)),(to_sfixed_a(-0.0001415717852069065)),(to_sfixed_a(0.002968207001686096)),(to_sfixed_a(0.0005305776139721274)),(to_sfixed_a(-0.0028404018376022577)),(to_sfixed_a(-0.12368322908878326)),(to_sfixed_a(0.07910935580730438)),(to_sfixed_a(-0.019819313660264015)),(to_sfixed_a(-0.08505800366401672)),(to_sfixed_a(-0.018618924543261528)),(to_sfixed_a(-0.09231053292751312)),(to_sfixed_a(-0.04537350684404373)),(to_sfixed_a(-0.03451048955321312)),(to_sfixed_a(0.00436413986608386)),(to_sfixed_a(0.023704934865236282)),(to_sfixed_a(0.24598783254623413)),(to_sfixed_a(-0.24002207815647125)),(to_sfixed_a(-0.22237350046634674)),(to_sfixed_a(-0.3339601159095764)),(to_sfixed_a(-0.0003688481810968369)),(to_sfixed_a(-0.022214598953723907)),(to_sfixed_a(-0.0012152758426964283)),(to_sfixed_a(0.05153168737888336)),(to_sfixed_a(-9.413436782779172e-05)),(to_sfixed_a(0.00022740884742233902)),(to_sfixed_a(-0.0001232763461302966)),(to_sfixed_a(-0.0001663704460952431)),(to_sfixed_a(0.0002267705713165924)),(to_sfixed_a(9.117391164181754e-05)),(to_sfixed_a(4.7503115638392046e-05)),(to_sfixed_a(-0.0002782245574053377)),(to_sfixed_a(0.1316303312778473)),(to_sfixed_a(0.1001499742269516)),(to_sfixed_a(0.18163204193115234)),(to_sfixed_a(0.03578004986047745)),(to_sfixed_a(0.015748273581266403)),(to_sfixed_a(-0.044744037091732025)),(to_sfixed_a(-0.028091592714190483)),(to_sfixed_a(-0.24323709309101105)),(to_sfixed_a(-0.14240242540836334)),(to_sfixed_a(0.012938432395458221)),(to_sfixed_a(0.013092405162751675)),(to_sfixed_a(0.01960095949470997)),(to_sfixed_a(0.04718029871582985)),(to_sfixed_a(-0.20778214931488037)),(to_sfixed_a(0.01440434716641903)),(to_sfixed_a(-0.004514646250754595)),(to_sfixed_a(-0.004177687224000692)),(to_sfixed_a(0.053358208388090134)),(to_sfixed_a(-0.015699181705713272)),(to_sfixed_a(-9.294936171500012e-05)),(to_sfixed_a(-5.971877908450551e-05)),(to_sfixed_a(-0.0001780217426130548)),(to_sfixed_a(8.744633669266477e-05)),(to_sfixed_a(2.7155178031534888e-05)),(to_sfixed_a(6.639361527049914e-05)),(to_sfixed_a(0.0002551469951868057)),(to_sfixed_a(-0.00015306621207855642)),(to_sfixed_a(-0.0002597257262095809)),(to_sfixed_a(-0.02033628337085247)),(to_sfixed_a(-0.04583612084388733)),(to_sfixed_a(-0.07971954345703125)),(to_sfixed_a(0.1388530135154724)),(to_sfixed_a(-0.048602163791656494)),(to_sfixed_a(-0.05714200437068939)),(to_sfixed_a(-0.057362984865903854)),(to_sfixed_a(0.06955586373806)),(to_sfixed_a(-0.09292343258857727)),(to_sfixed_a(-0.17089833319187164)),(to_sfixed_a(-0.06651807576417923)),(to_sfixed_a(-0.20964333415031433)),(to_sfixed_a(0.11745090782642365)),(to_sfixed_a(-0.06830383837223053)),(to_sfixed_a(-0.10346271097660065)),(to_sfixed_a(0.02163298800587654)),(to_sfixed_a(-0.03561844304203987)),(to_sfixed_a(-0.023555658757686615)),(to_sfixed_a(-0.014997203834354877)),(to_sfixed_a(8.491482003591955e-05)),(to_sfixed_a(-0.00011710340913850814)),(to_sfixed_a(-0.00012836474343203008)),(to_sfixed_a(3.862825542455539e-05)),(to_sfixed_a(0.00011403297685319558)),(to_sfixed_a(-0.00023406711989082396)),(to_sfixed_a(-0.00016768675413914025)),(to_sfixed_a(6.534824933623895e-06)),(to_sfixed_a(0.015626797452569008)),(to_sfixed_a(-0.04646258056163788)),(to_sfixed_a(0.06323013454675674)),(to_sfixed_a(0.12643493711948395)),(to_sfixed_a(0.07080457359552383)),(to_sfixed_a(0.06438720971345901)),(to_sfixed_a(-0.005435371771454811)),(to_sfixed_a(-0.12958240509033203)),(to_sfixed_a(0.03467962518334389)),(to_sfixed_a(0.377470999956131)),(to_sfixed_a(-0.05885619670152664)),(to_sfixed_a(-0.12356103211641312)),(to_sfixed_a(0.5172322392463684)),(to_sfixed_a(-0.09946370869874954)),(to_sfixed_a(-0.00526512460783124)),(to_sfixed_a(-0.07753122597932816)),(to_sfixed_a(-0.0035348657984286547)),(to_sfixed_a(-0.053210582584142685)),(to_sfixed_a(-0.02010534144937992)),(to_sfixed_a(-0.015352039597928524)),(to_sfixed_a(-9.091597894439474e-05)),(to_sfixed_a(0.0001389072131132707)),(to_sfixed_a(0.00020667216449510306)),(to_sfixed_a(-1.951133344846312e-05)),(to_sfixed_a(0.00020073264022357762)),(to_sfixed_a(-5.357979262043955e-06)),(to_sfixed_a(4.188643288216554e-06)),(to_sfixed_a(4.004788934253156e-05)),(to_sfixed_a(-0.00014592136722058058)),(to_sfixed_a(0.012496710754930973)),(to_sfixed_a(0.03918332979083061)),(to_sfixed_a(-0.02317887544631958)),(to_sfixed_a(0.1156831905245781)),(to_sfixed_a(0.18753942847251892)),(to_sfixed_a(0.005777359940111637)),(to_sfixed_a(-0.06895571947097778)),(to_sfixed_a(0.27515795826911926)),(to_sfixed_a(0.10948913544416428)),(to_sfixed_a(0.019009679555892944)),(to_sfixed_a(0.010653679259121418)),(to_sfixed_a(0.14852343499660492)),(to_sfixed_a(-0.022330624982714653)),(to_sfixed_a(0.005410529673099518)),(to_sfixed_a(-0.1371769905090332)),(to_sfixed_a(-0.1440647542476654)),(to_sfixed_a(-0.0010427817469462752)),(to_sfixed_a(-0.007309229113161564)),(to_sfixed_a(-0.008001943118870258)),(to_sfixed_a(2.0827857952099293e-05)),(to_sfixed_a(0.00021928545902483165)),(to_sfixed_a(-2.50889115704922e-06)),(to_sfixed_a(0.00020596012473106384)),(to_sfixed_a(9.107612277148291e-05)),(to_sfixed_a(-0.00010932428995147347)),(to_sfixed_a(0.0003486895002424717)),(to_sfixed_a(-2.398617289145477e-05)),(to_sfixed_a(3.211599323549308e-05)),(to_sfixed_a(0.0009958143346011639)),(to_sfixed_a(0.0012331744655966759)),(to_sfixed_a(-5.450525713968091e-05)),(to_sfixed_a(-0.00010477631440153345)),(to_sfixed_a(0.0003338469541631639)),(to_sfixed_a(-0.10234922170639038)),(to_sfixed_a(-0.009198720566928387)),(to_sfixed_a(-0.002799786627292633)),(to_sfixed_a(-0.06659755110740662)),(to_sfixed_a(-0.0160544253885746)),(to_sfixed_a(0.0041877212934195995)),(to_sfixed_a(-0.020825175568461418)),(to_sfixed_a(-0.07464548945426941)),(to_sfixed_a(-0.09453482180833817)),(to_sfixed_a(0.002638374688103795)),(to_sfixed_a(0.0019320901483297348)),(to_sfixed_a(0.00016374941333197057)),(to_sfixed_a(-0.00011520255793584511)),(to_sfixed_a(0.00041929809958674014)),(to_sfixed_a(-0.00021956702403258532)),(to_sfixed_a(-4.1486007830826566e-05)),(to_sfixed_a(7.872922287788242e-05)),(to_sfixed_a(-5.747355680796318e-05)),(to_sfixed_a(0.00018612494750414044)),(to_sfixed_a(-8.391847950406373e-05)),(to_sfixed_a(-6.352089712891029e-06)),(to_sfixed_a(9.547465197101701e-06)),(to_sfixed_a(-0.00011383341188775375)),(to_sfixed_a(-2.761333053058479e-05)),(to_sfixed_a(-3.151834607706405e-05)),(to_sfixed_a(5.747585601056926e-05)),(to_sfixed_a(0.000358532095560804)),(to_sfixed_a(6.512308755191043e-05)),(to_sfixed_a(-6.027623385307379e-05)),(to_sfixed_a(2.6211886506644078e-05)),(to_sfixed_a(-4.284727765480056e-06)),(to_sfixed_a(3.149025360471569e-05)),(to_sfixed_a(0.00016695783415343612)),(to_sfixed_a(0.0003030298976227641)),(to_sfixed_a(0.00016882986528798938)),(to_sfixed_a(-9.794743164093234e-06)),(to_sfixed_a(-0.0002209107333328575)),(to_sfixed_a(0.00019517213513609022)),(to_sfixed_a(0.00016326822515111417)),(to_sfixed_a(-0.00011823919339803979)),(to_sfixed_a(-7.536691555287689e-05)),(to_sfixed_a(-0.00021482535521499813)),(to_sfixed_a(6.190495332702994e-05)),(to_sfixed_a(7.505776011385024e-05)),(to_sfixed_a(-5.688165401807055e-05)),(to_sfixed_a(-0.00021984221530146897)));

    constant weight_n0_10 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-4.297447594581172e-05)),(to_sfixed_a(-0.00016281200805678964)),(to_sfixed_a(3.3862049804156413e-06)),(to_sfixed_a(1.998576226469595e-05)),(to_sfixed_a(0.00012631421850528568)),(to_sfixed_a(-0.00022523972438648343)),(to_sfixed_a(-6.728381413267925e-05)),(to_sfixed_a(0.0003499386366456747)),(to_sfixed_a(-4.3311800254741684e-05)),(to_sfixed_a(-3.679687870317139e-05)),(to_sfixed_a(1.2593084647960495e-05)),(to_sfixed_a(-0.00023391643480863422)),(to_sfixed_a(-9.853363735601306e-05)),(to_sfixed_a(0.00014073388592805713)),(to_sfixed_a(4.934025855618529e-05)),(to_sfixed_a(0.00013777973072137684)),(to_sfixed_a(1.1874743904627394e-05)),(to_sfixed_a(-2.321982719877269e-05)),(to_sfixed_a(8.937173697631806e-05)),(to_sfixed_a(7.342650496866554e-05)),(to_sfixed_a(-0.00014357856707647443)),(to_sfixed_a(0.0001557389769004658)),(to_sfixed_a(3.6704626836581156e-05)),(to_sfixed_a(0.0001875455491244793)),(to_sfixed_a(-3.034900510101579e-05)),(to_sfixed_a(5.917190355830826e-05)),(to_sfixed_a(7.950825965963304e-05)),(to_sfixed_a(-0.00023417834017891437)),(to_sfixed_a(-0.0002659414312802255)),(to_sfixed_a(4.671363740271772e-08)),(to_sfixed_a(-0.00011345365783199668)),(to_sfixed_a(-0.00014974076475482434)),(to_sfixed_a(-1.3817463695886545e-05)),(to_sfixed_a(-1.6819854863570072e-05)),(to_sfixed_a(7.000956975389272e-05)),(to_sfixed_a(0.0002949096087832004)),(to_sfixed_a(0.00013385874626692384)),(to_sfixed_a(2.3634062017663382e-05)),(to_sfixed_a(0.00030003790743649006)),(to_sfixed_a(0.00020815478637814522)),(to_sfixed_a(-0.0001992308971239254)),(to_sfixed_a(0.00025313792866654694)),(to_sfixed_a(3.2245818147202954e-05)),(to_sfixed_a(4.012220597360283e-05)),(to_sfixed_a(0.0001524726685602218)),(to_sfixed_a(7.130822723411256e-07)),(to_sfixed_a(-0.0001843834324972704)),(to_sfixed_a(-0.0002306762180523947)),(to_sfixed_a(-0.00041899376083165407)),(to_sfixed_a(-0.00032720222952775657)),(to_sfixed_a(-2.951811438833829e-05)),(to_sfixed_a(-1.1587195558604435e-06)),(to_sfixed_a(-0.00010885895608225837)),(to_sfixed_a(9.458002750761807e-05)),(to_sfixed_a(-3.109588215011172e-05)),(to_sfixed_a(-0.00017939847020898014)),(to_sfixed_a(0.00011748525139410049)),(to_sfixed_a(-0.00013628252781927586)),(to_sfixed_a(0.00019370550580788404)),(to_sfixed_a(0.00016803662583697587)),(to_sfixed_a(-5.439528831630014e-05)),(to_sfixed_a(2.0210814909660257e-05)),(to_sfixed_a(1.0063828312922851e-06)),(to_sfixed_a(-0.0002620044397190213)),(to_sfixed_a(0.00012155356671428308)),(to_sfixed_a(-0.00027204988873563707)),(to_sfixed_a(5.305300510372035e-05)),(to_sfixed_a(8.00157431513071e-06)),(to_sfixed_a(-6.194313755258918e-05)),(to_sfixed_a(-0.004541747272014618)),(to_sfixed_a(0.0002506681194063276)),(to_sfixed_a(3.921150346286595e-05)),(to_sfixed_a(4.296178667573258e-05)),(to_sfixed_a(-3.358931644470431e-05)),(to_sfixed_a(8.809034625301138e-05)),(to_sfixed_a(-3.479816950857639e-05)),(to_sfixed_a(-0.00011172605445608497)),(to_sfixed_a(-4.013714351458475e-05)),(to_sfixed_a(9.036117262439802e-06)),(to_sfixed_a(3.102168420809903e-06)),(to_sfixed_a(-0.0003226312401238829)),(to_sfixed_a(1.966153649846092e-05)),(to_sfixed_a(-7.893113797763363e-05)),(to_sfixed_a(-0.00012804906873498112)),(to_sfixed_a(-0.00020559396944008768)),(to_sfixed_a(0.0001444461231585592)),(to_sfixed_a(-0.00012453633826225996)),(to_sfixed_a(-2.358466008445248e-05)),(to_sfixed_a(-2.284038782818243e-05)),(to_sfixed_a(0.00018355327483732253)),(to_sfixed_a(9.164315270027146e-05)),(to_sfixed_a(0.0001837313175201416)),(to_sfixed_a(-0.01072793547064066)),(to_sfixed_a(-1.0042194844572805e-06)),(to_sfixed_a(-0.01215147040784359)),(to_sfixed_a(0.18509887158870697)),(to_sfixed_a(0.01114640012383461)),(to_sfixed_a(0.03652597963809967)),(to_sfixed_a(-0.01752380281686783)),(to_sfixed_a(-0.026069924235343933)),(to_sfixed_a(0.016353001818060875)),(to_sfixed_a(0.03186805173754692)),(to_sfixed_a(-0.11658255010843277)),(to_sfixed_a(-0.012390071526169777)),(to_sfixed_a(-0.0023376846220344305)),(to_sfixed_a(-0.004615224432200193)),(to_sfixed_a(-3.5652181395562366e-05)),(to_sfixed_a(0.00016437149315606803)),(to_sfixed_a(8.680569590069354e-05)),(to_sfixed_a(5.8341847761766985e-05)),(to_sfixed_a(-6.968440720811486e-05)),(to_sfixed_a(-0.00024383034906350076)),(to_sfixed_a(-0.0001951883314177394)),(to_sfixed_a(2.1773596017737873e-05)),(to_sfixed_a(-1.881954631244298e-05)),(to_sfixed_a(-5.4280986660160124e-05)),(to_sfixed_a(-8.375367906410247e-05)),(to_sfixed_a(8.869491284713149e-05)),(to_sfixed_a(0.001362777897156775)),(to_sfixed_a(0.073882095515728)),(to_sfixed_a(-0.025117849931120872)),(to_sfixed_a(-0.016935059800744057)),(to_sfixed_a(0.3007625341415405)),(to_sfixed_a(0.06011374667286873)),(to_sfixed_a(0.19796936213970184)),(to_sfixed_a(0.02719319611787796)),(to_sfixed_a(-0.042224809527397156)),(to_sfixed_a(-0.03315719962120056)),(to_sfixed_a(0.15340864658355713)),(to_sfixed_a(0.05120796710252762)),(to_sfixed_a(0.09276055544614792)),(to_sfixed_a(0.014995056204497814)),(to_sfixed_a(-0.022996455430984497)),(to_sfixed_a(-0.02755420096218586)),(to_sfixed_a(0.012949904426932335)),(to_sfixed_a(0.000386086932849139)),(to_sfixed_a(-0.00011086117592640221)),(to_sfixed_a(0.000144283301779069)),(to_sfixed_a(0.00016030104598030448)),(to_sfixed_a(-0.00013990139996167272)),(to_sfixed_a(0.00025947566609829664)),(to_sfixed_a(-1.902381336549297e-05)),(to_sfixed_a(0.00013659692194778472)),(to_sfixed_a(-0.00031305814627557993)),(to_sfixed_a(0.0013510960852727294)),(to_sfixed_a(0.1184445470571518)),(to_sfixed_a(0.014553649351000786)),(to_sfixed_a(0.1992177963256836)),(to_sfixed_a(0.26710671186447144)),(to_sfixed_a(-0.0022546290419995785)),(to_sfixed_a(0.01676136627793312)),(to_sfixed_a(0.1984689086675644)),(to_sfixed_a(0.20497733354568481)),(to_sfixed_a(0.2542862594127655)),(to_sfixed_a(0.006738625932484865)),(to_sfixed_a(0.11193665117025375)),(to_sfixed_a(0.028550228103995323)),(to_sfixed_a(0.2388506680727005)),(to_sfixed_a(0.2108619064092636)),(to_sfixed_a(-0.11329279094934464)),(to_sfixed_a(-0.07787320017814636)),(to_sfixed_a(-0.11922785639762878)),(to_sfixed_a(-9.10688831936568e-05)),(to_sfixed_a(-0.057923708111047745)),(to_sfixed_a(-0.0007715413812547922)),(to_sfixed_a(0.0006285937852226198)),(to_sfixed_a(0.00019852645345963538)),(to_sfixed_a(-6.970936738071032e-06)),(to_sfixed_a(5.898932067793794e-05)),(to_sfixed_a(-0.00012631277786567807)),(to_sfixed_a(0.00023391525610350072)),(to_sfixed_a(-0.00023958575911819935)),(to_sfixed_a(-0.0003009771171491593)),(to_sfixed_a(0.11397410929203033)),(to_sfixed_a(0.14119671285152435)),(to_sfixed_a(0.13940925896167755)),(to_sfixed_a(0.12271236628293991)),(to_sfixed_a(-0.020586326718330383)),(to_sfixed_a(0.3012748956680298)),(to_sfixed_a(0.28905513882637024)),(to_sfixed_a(0.18922163546085358)),(to_sfixed_a(0.1837908923625946)),(to_sfixed_a(0.21347220242023468)),(to_sfixed_a(0.3072132468223572)),(to_sfixed_a(0.322043776512146)),(to_sfixed_a(0.11467946320772171)),(to_sfixed_a(0.10392126441001892)),(to_sfixed_a(-0.09759433567523956)),(to_sfixed_a(-0.18450325727462769)),(to_sfixed_a(0.05819331109523773)),(to_sfixed_a(-0.21676237881183624)),(to_sfixed_a(-0.2197655439376831)),(to_sfixed_a(0.000613926153164357)),(to_sfixed_a(0.00020940722606610507)),(to_sfixed_a(0.0026118867099285126)),(to_sfixed_a(4.9945974751608446e-05)),(to_sfixed_a(0.00018771963368635625)),(to_sfixed_a(-0.0002494349901098758)),(to_sfixed_a(0.0001343407784588635)),(to_sfixed_a(2.9780730983475223e-05)),(to_sfixed_a(7.743777678115293e-05)),(to_sfixed_a(0.09665442258119583)),(to_sfixed_a(0.11358211934566498)),(to_sfixed_a(-0.08224848657846451)),(to_sfixed_a(-0.16823774576187134)),(to_sfixed_a(0.021415334194898605)),(to_sfixed_a(0.08562655001878738)),(to_sfixed_a(0.0511452741920948)),(to_sfixed_a(-0.07481652498245239)),(to_sfixed_a(0.1208721473813057)),(to_sfixed_a(0.11203332245349884)),(to_sfixed_a(0.1434236466884613)),(to_sfixed_a(0.22446158528327942)),(to_sfixed_a(0.12421824038028717)),(to_sfixed_a(-0.07308397442102432)),(to_sfixed_a(0.2307470589876175)),(to_sfixed_a(-0.34272003173828125)),(to_sfixed_a(-0.10034695267677307)),(to_sfixed_a(-0.28466764092445374)),(to_sfixed_a(-0.3788537085056305)),(to_sfixed_a(-0.08869198709726334)),(to_sfixed_a(-0.009419985115528107)),(to_sfixed_a(5.598584903054871e-05)),(to_sfixed_a(0.0002069144247798249)),(to_sfixed_a(-2.6261777748004533e-05)),(to_sfixed_a(-0.00023741595214232802)),(to_sfixed_a(-0.00020728247181978077)),(to_sfixed_a(-0.0001257482945220545)),(to_sfixed_a(-0.011215128935873508)),(to_sfixed_a(-0.03146544471383095)),(to_sfixed_a(0.09220939129590988)),(to_sfixed_a(0.021276889368891716)),(to_sfixed_a(0.02659309282898903)),(to_sfixed_a(0.09842333942651749)),(to_sfixed_a(0.20168712735176086)),(to_sfixed_a(0.007405559532344341)),(to_sfixed_a(-0.08927887678146362)),(to_sfixed_a(0.02459682524204254)),(to_sfixed_a(0.12471982836723328)),(to_sfixed_a(0.1609063595533371)),(to_sfixed_a(0.11966577917337418)),(to_sfixed_a(-0.09924198687076569)),(to_sfixed_a(-0.3122320771217346)),(to_sfixed_a(-0.3668588697910309)),(to_sfixed_a(-0.18096701800823212)),(to_sfixed_a(-0.2426202893257141)),(to_sfixed_a(0.06412094831466675)),(to_sfixed_a(-0.2754180431365967)),(to_sfixed_a(-0.39229434728622437)),(to_sfixed_a(-0.0814318135380745)),(to_sfixed_a(4.5343487727222964e-05)),(to_sfixed_a(-3.020941448994563e-06)),(to_sfixed_a(3.112245030933991e-05)),(to_sfixed_a(-0.00028990779537707567)),(to_sfixed_a(-4.337075733928941e-05)),(to_sfixed_a(2.9062402973067947e-05)),(to_sfixed_a(0.0005202781176194549)),(to_sfixed_a(0.03975210338830948)),(to_sfixed_a(-0.061360448598861694)),(to_sfixed_a(-0.049143966287374496)),(to_sfixed_a(0.12924417853355408)),(to_sfixed_a(-0.08309505134820938)),(to_sfixed_a(-0.3661157786846161)),(to_sfixed_a(-0.1058179959654808)),(to_sfixed_a(0.11011696606874466)),(to_sfixed_a(-0.16542834043502808)),(to_sfixed_a(-0.068648561835289)),(to_sfixed_a(0.15492479503154755)),(to_sfixed_a(0.22452779114246368)),(to_sfixed_a(0.1623641699552536)),(to_sfixed_a(-0.06808115541934967)),(to_sfixed_a(-0.13906358182430267)),(to_sfixed_a(-0.2517532706260681)),(to_sfixed_a(-0.023012034595012665)),(to_sfixed_a(0.10742446035146713)),(to_sfixed_a(-0.2054091840982437)),(to_sfixed_a(-0.2092403918504715)),(to_sfixed_a(5.839437653776258e-05)),(to_sfixed_a(-6.750811007805169e-05)),(to_sfixed_a(2.9878630812163465e-05)),(to_sfixed_a(-6.820294220233336e-05)),(to_sfixed_a(-0.00010959966311929747)),(to_sfixed_a(-0.00036400178214535117)),(to_sfixed_a(0.00018447621550876647)),(to_sfixed_a(0.003525668289512396)),(to_sfixed_a(0.08109543472528458)),(to_sfixed_a(-0.04613010212779045)),(to_sfixed_a(-0.16115467250347137)),(to_sfixed_a(-0.2789328694343567)),(to_sfixed_a(-0.4983294904232025)),(to_sfixed_a(-0.10030924528837204)),(to_sfixed_a(0.06460723280906677)),(to_sfixed_a(-0.06967322528362274)),(to_sfixed_a(0.2660297751426697)),(to_sfixed_a(0.027532868087291718)),(to_sfixed_a(0.17492744326591492)),(to_sfixed_a(0.40786510705947876)),(to_sfixed_a(0.4206216037273407)),(to_sfixed_a(0.26848235726356506)),(to_sfixed_a(0.09223833680152893)),(to_sfixed_a(-0.12261465936899185)),(to_sfixed_a(-0.11355134099721909)),(to_sfixed_a(0.34827831387519836)),(to_sfixed_a(0.023314645513892174)),(to_sfixed_a(0.08540191501379013)),(to_sfixed_a(-0.02151365950703621)),(to_sfixed_a(-4.180415999144316e-05)),(to_sfixed_a(7.835552969481796e-05)),(to_sfixed_a(-3.49611509591341e-05)),(to_sfixed_a(0.00018759415252134204)),(to_sfixed_a(-1.8100105080520734e-05)),(to_sfixed_a(0.02337261289358139)),(to_sfixed_a(-0.012659704312682152)),(to_sfixed_a(-0.16619780659675598)),(to_sfixed_a(-0.1560676097869873)),(to_sfixed_a(-0.22267790138721466)),(to_sfixed_a(0.0031570231076329947)),(to_sfixed_a(-0.085208460688591)),(to_sfixed_a(-0.09527513384819031)),(to_sfixed_a(0.03883766010403633)),(to_sfixed_a(0.03213806450366974)),(to_sfixed_a(0.01661089062690735)),(to_sfixed_a(0.11963694542646408)),(to_sfixed_a(0.32846227288246155)),(to_sfixed_a(0.27720946073532104)),(to_sfixed_a(0.25360339879989624)),(to_sfixed_a(0.5361509919166565)),(to_sfixed_a(0.4890347719192505)),(to_sfixed_a(0.2392318844795227)),(to_sfixed_a(0.19851334393024445)),(to_sfixed_a(0.030693652108311653)),(to_sfixed_a(-5.686914664693177e-05)),(to_sfixed_a(0.24028408527374268)),(to_sfixed_a(9.873896487988532e-05)),(to_sfixed_a(-0.00017142476281151175)),(to_sfixed_a(-0.00013964055688120425)),(to_sfixed_a(9.401312854606658e-05)),(to_sfixed_a(-3.6186331271892413e-05)),(to_sfixed_a(3.164510053466074e-05)),(to_sfixed_a(-0.00018271533190272748)),(to_sfixed_a(-0.025356071069836617)),(to_sfixed_a(-0.23697049915790558)),(to_sfixed_a(-0.20489706099033356)),(to_sfixed_a(-0.12461453676223755)),(to_sfixed_a(-0.17620591819286346)),(to_sfixed_a(-0.275727778673172)),(to_sfixed_a(-0.12951835989952087)),(to_sfixed_a(-0.3455590009689331)),(to_sfixed_a(-0.5915112495422363)),(to_sfixed_a(-0.5079598426818848)),(to_sfixed_a(0.18929773569107056)),(to_sfixed_a(0.7399762272834778)),(to_sfixed_a(0.3419119715690613)),(to_sfixed_a(0.2180803120136261)),(to_sfixed_a(0.019417356699705124)),(to_sfixed_a(0.17310896515846252)),(to_sfixed_a(0.2598206102848053)),(to_sfixed_a(0.2982492446899414)),(to_sfixed_a(0.19164247810840607)),(to_sfixed_a(-0.03938603773713112)),(to_sfixed_a(0.16232995688915253)),(to_sfixed_a(-7.13979679858312e-05)),(to_sfixed_a(5.5895099649205804e-05)),(to_sfixed_a(-9.696120832813904e-05)),(to_sfixed_a(0.00021864048903807998)),(to_sfixed_a(2.1901105355937034e-06)),(to_sfixed_a(0.00017069578461814672)),(to_sfixed_a(6.960669270483777e-05)),(to_sfixed_a(-0.10014916956424713)),(to_sfixed_a(-0.47902438044548035)),(to_sfixed_a(-0.08283527195453644)),(to_sfixed_a(-0.22569966316223145)),(to_sfixed_a(0.053723305463790894)),(to_sfixed_a(-0.3458028733730316)),(to_sfixed_a(-0.029144737869501114)),(to_sfixed_a(-0.30866146087646484)),(to_sfixed_a(-0.18958339095115662)),(to_sfixed_a(-0.0815143883228302)),(to_sfixed_a(-0.008310407400131226)),(to_sfixed_a(0.13827931880950928)),(to_sfixed_a(0.18219000101089478)),(to_sfixed_a(0.11134251207113266)),(to_sfixed_a(0.02384689263999462)),(to_sfixed_a(-0.2093045860528946)),(to_sfixed_a(0.042722221463918686)),(to_sfixed_a(-0.03887008875608444)),(to_sfixed_a(-0.05685801804065704)),(to_sfixed_a(0.4285283386707306)),(to_sfixed_a(-0.012127967551350594)),(to_sfixed_a(0.0015686952974647284)),(to_sfixed_a(0.0013265236048027873)),(to_sfixed_a(-3.483811815385707e-05)),(to_sfixed_a(0.00023666773631703109)),(to_sfixed_a(-0.0001311791129410267)),(to_sfixed_a(-0.00014504353748634458)),(to_sfixed_a(0.00017847462731879205)),(to_sfixed_a(-0.001602568314410746)),(to_sfixed_a(-0.29970812797546387)),(to_sfixed_a(-0.11493642628192902)),(to_sfixed_a(-0.2758142054080963)),(to_sfixed_a(-0.36902233958244324)),(to_sfixed_a(-0.26896703243255615)),(to_sfixed_a(-0.5562105178833008)),(to_sfixed_a(-0.4026503264904022)),(to_sfixed_a(-0.337704062461853)),(to_sfixed_a(-0.32687291502952576)),(to_sfixed_a(0.14584395289421082)),(to_sfixed_a(0.20597374439239502)),(to_sfixed_a(0.061606213450431824)),(to_sfixed_a(-0.03222605586051941)),(to_sfixed_a(-0.17083904147148132)),(to_sfixed_a(-0.3205157220363617)),(to_sfixed_a(-0.15781736373901367)),(to_sfixed_a(-0.16694849729537964)),(to_sfixed_a(0.016567682847380638)),(to_sfixed_a(-0.04557286575436592)),(to_sfixed_a(0.060465119779109955)),(to_sfixed_a(6.065821708034491e-06)),(to_sfixed_a(-0.00013739749556407332)),(to_sfixed_a(7.305650797206908e-05)),(to_sfixed_a(6.690960435662419e-05)),(to_sfixed_a(6.534688145620748e-05)),(to_sfixed_a(-0.00035148393362760544)),(to_sfixed_a(-0.00016641250113025308)),(to_sfixed_a(-0.05705615505576134)),(to_sfixed_a(-0.3223954737186432)),(to_sfixed_a(-0.1345294862985611)),(to_sfixed_a(-0.2390681803226471)),(to_sfixed_a(-0.14509855210781097)),(to_sfixed_a(-0.05465469881892204)),(to_sfixed_a(-0.2524271011352539)),(to_sfixed_a(-0.32860445976257324)),(to_sfixed_a(-0.5108137726783752)),(to_sfixed_a(-0.14068129658699036)),(to_sfixed_a(-0.0449930876493454)),(to_sfixed_a(0.21069638431072235)),(to_sfixed_a(0.2016306221485138)),(to_sfixed_a(-0.12138165533542633)),(to_sfixed_a(-0.3333042562007904)),(to_sfixed_a(-0.5153123736381531)),(to_sfixed_a(0.057018302381038666)),(to_sfixed_a(0.028440413996577263)),(to_sfixed_a(0.04122160002589226)),(to_sfixed_a(0.11803392320871353)),(to_sfixed_a(-0.01870104670524597)),(to_sfixed_a(0.00033692005672492087)),(to_sfixed_a(-2.6469009753782302e-05)),(to_sfixed_a(5.838916422362672e-06)),(to_sfixed_a(0.0002407038991805166)),(to_sfixed_a(2.6847681510844268e-05)),(to_sfixed_a(-0.0002174340042984113)),(to_sfixed_a(-0.004452084191143513)),(to_sfixed_a(-0.09956725686788559)),(to_sfixed_a(0.12155462801456451)),(to_sfixed_a(0.22434672713279724)),(to_sfixed_a(0.12099859863519669)),(to_sfixed_a(0.11015186458826065)),(to_sfixed_a(0.23044127225875854)),(to_sfixed_a(-0.026856545358896255)),(to_sfixed_a(-0.33442550897598267)),(to_sfixed_a(-0.07090672105550766)),(to_sfixed_a(0.005522916559129953)),(to_sfixed_a(-0.018389441072940826)),(to_sfixed_a(0.07197503745555878)),(to_sfixed_a(0.07823104411363602)),(to_sfixed_a(-0.07010603696107864)),(to_sfixed_a(-0.2087823897600174)),(to_sfixed_a(-0.1257363259792328)),(to_sfixed_a(-0.03577783331274986)),(to_sfixed_a(0.05319301411509514)),(to_sfixed_a(-0.07369501888751984)),(to_sfixed_a(0.23870053887367249)),(to_sfixed_a(-0.03394101560115814)),(to_sfixed_a(0.004329859744757414)),(to_sfixed_a(-0.00015775237989146262)),(to_sfixed_a(0.0002669051755219698)),(to_sfixed_a(-4.6271816245280206e-05)),(to_sfixed_a(-8.842279203236103e-05)),(to_sfixed_a(-0.0027142066974192858)),(to_sfixed_a(-0.004570807330310345)),(to_sfixed_a(0.15836335718631744)),(to_sfixed_a(0.08730781078338623)),(to_sfixed_a(0.16276349127292633)),(to_sfixed_a(0.1052875965833664)),(to_sfixed_a(0.3161596953868866)),(to_sfixed_a(0.2672007083892822)),(to_sfixed_a(0.448758065700531)),(to_sfixed_a(0.24491626024246216)),(to_sfixed_a(-0.09537429362535477)),(to_sfixed_a(0.24304106831550598)),(to_sfixed_a(-0.08239489793777466)),(to_sfixed_a(0.12505429983139038)),(to_sfixed_a(-0.2457713931798935)),(to_sfixed_a(-0.21121688187122345)),(to_sfixed_a(-0.32893550395965576)),(to_sfixed_a(-0.04649488627910614)),(to_sfixed_a(-0.17157389223575592)),(to_sfixed_a(-0.12602262198925018)),(to_sfixed_a(-0.030120372772216797)),(to_sfixed_a(0.004822169430553913)),(to_sfixed_a(0.00016328693891409785)),(to_sfixed_a(-1.2623051588889211e-05)),(to_sfixed_a(4.984019687981345e-05)),(to_sfixed_a(5.0509268476162106e-05)),(to_sfixed_a(-8.714348950888962e-05)),(to_sfixed_a(-0.00016680323460604995)),(to_sfixed_a(-0.00010719527199398726)),(to_sfixed_a(0.024581868201494217)),(to_sfixed_a(0.01114635169506073)),(to_sfixed_a(-0.16231794655323029)),(to_sfixed_a(0.00919139850884676)),(to_sfixed_a(0.18236549198627472)),(to_sfixed_a(0.03941556438803673)),(to_sfixed_a(0.2765389084815979)),(to_sfixed_a(0.09491149336099625)),(to_sfixed_a(-0.21263033151626587)),(to_sfixed_a(-0.028215711936354637)),(to_sfixed_a(-0.06854789704084396)),(to_sfixed_a(-0.06572580337524414)),(to_sfixed_a(-0.09080249071121216)),(to_sfixed_a(-0.2361806035041809)),(to_sfixed_a(-0.1418938785791397)),(to_sfixed_a(-0.05707226321101189)),(to_sfixed_a(-0.1998283565044403)),(to_sfixed_a(-0.08142240345478058)),(to_sfixed_a(-0.25817689299583435)),(to_sfixed_a(0.15423612296581268)),(to_sfixed_a(-0.05890420079231262)),(to_sfixed_a(-0.014440242201089859)),(to_sfixed_a(0.00013421390030998737)),(to_sfixed_a(-0.0003725705901160836)),(to_sfixed_a(0.00021349287999328226)),(to_sfixed_a(-0.00021453054796438664)),(to_sfixed_a(0.0002149628271581605)),(to_sfixed_a(-6.243725692911539e-06)),(to_sfixed_a(0.006495187990367413)),(to_sfixed_a(-0.0031310804188251495)),(to_sfixed_a(0.19144907593727112)),(to_sfixed_a(-0.015241959132254124)),(to_sfixed_a(0.09849805384874344)),(to_sfixed_a(-0.06545736640691757)),(to_sfixed_a(-0.17449520528316498)),(to_sfixed_a(-0.553677499294281)),(to_sfixed_a(-0.4505259096622467)),(to_sfixed_a(-0.4847719073295593)),(to_sfixed_a(0.09724097698926926)),(to_sfixed_a(-0.15627340972423553)),(to_sfixed_a(-0.22783350944519043)),(to_sfixed_a(-0.15933063626289368)),(to_sfixed_a(-0.230991929769516)),(to_sfixed_a(-0.23082499206066132)),(to_sfixed_a(-0.09813534468412399)),(to_sfixed_a(-0.025278214365243912)),(to_sfixed_a(-0.22917059063911438)),(to_sfixed_a(0.19258376955986023)),(to_sfixed_a(-0.07153378427028656)),(to_sfixed_a(-1.5096059541974682e-05)),(to_sfixed_a(-0.0001290059444727376)),(to_sfixed_a(0.00023522638366557658)),(to_sfixed_a(-5.125450843479484e-05)),(to_sfixed_a(-0.00017975996888708323)),(to_sfixed_a(-0.0003044414333999157)),(to_sfixed_a(-0.00010379187733633444)),(to_sfixed_a(-0.0002647076325956732)),(to_sfixed_a(-0.012326112948358059)),(to_sfixed_a(-0.02034158818423748)),(to_sfixed_a(0.052363816648721695)),(to_sfixed_a(0.039202164858579636)),(to_sfixed_a(0.02671804651618004)),(to_sfixed_a(-0.3471090495586395)),(to_sfixed_a(-0.08128216862678528)),(to_sfixed_a(-0.3235185444355011)),(to_sfixed_a(-0.36562579870224)),(to_sfixed_a(0.021685177460312843)),(to_sfixed_a(0.017838919535279274)),(to_sfixed_a(-0.12154186517000198)),(to_sfixed_a(0.04606316611170769)),(to_sfixed_a(-0.22629477083683014)),(to_sfixed_a(0.030002783983945847)),(to_sfixed_a(-0.34623512625694275)),(to_sfixed_a(-0.23934222757816315)),(to_sfixed_a(0.10239679366350174)),(to_sfixed_a(-0.07339555770158768)),(to_sfixed_a(-0.037491895258426666)),(to_sfixed_a(0.03429222106933594)),(to_sfixed_a(0.00010677784302970394)),(to_sfixed_a(-1.2126964975323062e-05)),(to_sfixed_a(-0.0002809001598507166)),(to_sfixed_a(7.126888522179797e-05)),(to_sfixed_a(9.86468730843626e-05)),(to_sfixed_a(2.9983712011016905e-05)),(to_sfixed_a(-3.0116182188066887e-06)),(to_sfixed_a(0.0625111311674118)),(to_sfixed_a(-0.001057189074344933)),(to_sfixed_a(-0.10213903337717056)),(to_sfixed_a(0.11160045862197876)),(to_sfixed_a(-0.13885602355003357)),(to_sfixed_a(0.18615804612636566)),(to_sfixed_a(0.12880705296993256)),(to_sfixed_a(0.25197935104370117)),(to_sfixed_a(-0.08155199140310287)),(to_sfixed_a(-0.008497685194015503)),(to_sfixed_a(-0.029970617964863777)),(to_sfixed_a(0.06021936982870102)),(to_sfixed_a(-0.06610007584095001)),(to_sfixed_a(-0.2508569359779358)),(to_sfixed_a(-0.17695176601409912)),(to_sfixed_a(-0.14443492889404297)),(to_sfixed_a(-0.1460527926683426)),(to_sfixed_a(-0.029088696464896202)),(to_sfixed_a(-0.10332787781953812)),(to_sfixed_a(0.0005012984620407224)),(to_sfixed_a(-0.02998819388449192)),(to_sfixed_a(-4.342643478594255e-06)),(to_sfixed_a(1.693060767138377e-05)),(to_sfixed_a(-3.1110950658330694e-05)),(to_sfixed_a(4.136443749302998e-05)),(to_sfixed_a(3.496568388072774e-05)),(to_sfixed_a(5.225828499533236e-05)),(to_sfixed_a(0.00010037973697762936)),(to_sfixed_a(-0.0005605676560662687)),(to_sfixed_a(-0.004884702619165182)),(to_sfixed_a(0.1737411767244339)),(to_sfixed_a(0.1688733696937561)),(to_sfixed_a(0.022624703124165535)),(to_sfixed_a(0.06254857778549194)),(to_sfixed_a(0.08468496799468994)),(to_sfixed_a(0.048461224883794785)),(to_sfixed_a(-0.04384274780750275)),(to_sfixed_a(0.056306224316358566)),(to_sfixed_a(-0.03419864922761917)),(to_sfixed_a(-0.17371971905231476)),(to_sfixed_a(-0.19322188198566437)),(to_sfixed_a(-0.20153072476387024)),(to_sfixed_a(-0.3388338088989258)),(to_sfixed_a(0.0037159149069339037)),(to_sfixed_a(-0.05891774594783783)),(to_sfixed_a(-0.022718753665685654)),(to_sfixed_a(-0.05806327983736992)),(to_sfixed_a(-0.003004610538482666)),(to_sfixed_a(-0.00013621982361655682)),(to_sfixed_a(0.00015252416778821498)),(to_sfixed_a(-0.00011742733477149159)),(to_sfixed_a(-9.67882588156499e-05)),(to_sfixed_a(-5.076466186437756e-05)),(to_sfixed_a(-0.00018848977924790233)),(to_sfixed_a(6.725703860865906e-05)),(to_sfixed_a(-0.00020802489598281682)),(to_sfixed_a(-0.0006169034750200808)),(to_sfixed_a(0.011820276267826557)),(to_sfixed_a(0.06944781541824341)),(to_sfixed_a(-0.12405460327863693)),(to_sfixed_a(0.09436886012554169)),(to_sfixed_a(0.02962745539844036)),(to_sfixed_a(0.0019084407249465585)),(to_sfixed_a(0.058328233659267426)),(to_sfixed_a(-0.07025711238384247)),(to_sfixed_a(-0.005459066480398178)),(to_sfixed_a(0.09119510650634766)),(to_sfixed_a(-0.01266274694353342)),(to_sfixed_a(-0.26310214400291443)),(to_sfixed_a(0.032705117017030716)),(to_sfixed_a(0.0770130306482315)),(to_sfixed_a(0.016026299446821213)),(to_sfixed_a(0.03568808361887932)),(to_sfixed_a(-0.12035377323627472)),(to_sfixed_a(-0.007234077900648117)),(to_sfixed_a(-0.09138180315494537)),(to_sfixed_a(-3.901421951013617e-05)),(to_sfixed_a(-2.4125434720190242e-05)),(to_sfixed_a(-0.000255434715654701)),(to_sfixed_a(-2.4710830984986387e-05)),(to_sfixed_a(-6.75902483635582e-05)),(to_sfixed_a(0.0003987850795965642)),(to_sfixed_a(1.690170211077202e-05)),(to_sfixed_a(-0.00014275670400820673)),(to_sfixed_a(0.00289850402623415)),(to_sfixed_a(0.0335904136300087)),(to_sfixed_a(0.014501137658953667)),(to_sfixed_a(0.12774521112442017)),(to_sfixed_a(0.3013298809528351)),(to_sfixed_a(0.2508205771446228)),(to_sfixed_a(-0.1154237687587738)),(to_sfixed_a(-0.2412710189819336)),(to_sfixed_a(-0.1913839876651764)),(to_sfixed_a(-0.07134509086608887)),(to_sfixed_a(-0.03377072513103485)),(to_sfixed_a(-0.09056265652179718)),(to_sfixed_a(-0.49385783076286316)),(to_sfixed_a(-0.13895316421985626)),(to_sfixed_a(-0.06009430065751076)),(to_sfixed_a(-0.05208365619182587)),(to_sfixed_a(0.012332948856055737)),(to_sfixed_a(-0.051722850650548935)),(to_sfixed_a(-0.04348897933959961)),(to_sfixed_a(-0.0020673843100667)),(to_sfixed_a(-0.00027593536651693285)),(to_sfixed_a(9.711735765449703e-05)),(to_sfixed_a(-1.993745900108479e-05)),(to_sfixed_a(3.86596548196394e-05)),(to_sfixed_a(0.0002902160631492734)),(to_sfixed_a(-6.934713019290939e-05)),(to_sfixed_a(-8.93011165317148e-05)),(to_sfixed_a(7.180088869063184e-05)),(to_sfixed_a(6.415294774342328e-05)),(to_sfixed_a(0.0480944998562336)),(to_sfixed_a(0.007300259079784155)),(to_sfixed_a(0.05281481146812439)),(to_sfixed_a(0.09317556768655777)),(to_sfixed_a(0.020718686282634735)),(to_sfixed_a(0.044335026293992996)),(to_sfixed_a(-0.0037131954450160265)),(to_sfixed_a(0.1299261748790741)),(to_sfixed_a(0.057446908205747604)),(to_sfixed_a(0.06923219561576843)),(to_sfixed_a(0.009381985291838646)),(to_sfixed_a(-0.0037051152903586626)),(to_sfixed_a(-0.09135013073682785)),(to_sfixed_a(0.009300153702497482)),(to_sfixed_a(0.05500422418117523)),(to_sfixed_a(0.023921815678477287)),(to_sfixed_a(-0.0010981064988300204)),(to_sfixed_a(-0.004361848812550306)),(to_sfixed_a(-0.004883086308836937)),(to_sfixed_a(3.684419425553642e-05)),(to_sfixed_a(0.00028222467517480254)),(to_sfixed_a(2.4753397156018764e-05)),(to_sfixed_a(0.0001939620851771906)),(to_sfixed_a(-0.0002570188953541219)),(to_sfixed_a(0.0002536717802286148)),(to_sfixed_a(-0.0001716477272566408)),(to_sfixed_a(-0.00012663770758081228)),(to_sfixed_a(-0.00013419362949207425)),(to_sfixed_a(0.004053795710206032)),(to_sfixed_a(0.003912505693733692)),(to_sfixed_a(-6.718134682159871e-05)),(to_sfixed_a(-0.00011066511797253042)),(to_sfixed_a(7.182000990724191e-05)),(to_sfixed_a(-0.019666435196995735)),(to_sfixed_a(-9.92704663076438e-05)),(to_sfixed_a(0.0008118503028526902)),(to_sfixed_a(-0.022821009159088135)),(to_sfixed_a(0.011692252941429615)),(to_sfixed_a(-0.008102277293801308)),(to_sfixed_a(-0.0016053528524935246)),(to_sfixed_a(-0.016716018319129944)),(to_sfixed_a(-0.019626857712864876)),(to_sfixed_a(0.0063676671124994755)),(to_sfixed_a(0.0013218133244663477)),(to_sfixed_a(0.00023194191453512758)),(to_sfixed_a(0.0001037477923091501)),(to_sfixed_a(-2.6617661205818877e-05)),(to_sfixed_a(3.179223131155595e-05)),(to_sfixed_a(-0.00011108813487226143)),(to_sfixed_a(-0.0002444279962219298)),(to_sfixed_a(5.851749301655218e-05)),(to_sfixed_a(-1.5491539670620114e-05)),(to_sfixed_a(-0.00018132815603166819)),(to_sfixed_a(0.00018473285308573395)),(to_sfixed_a(-5.285516454023309e-05)),(to_sfixed_a(-0.0002113042864948511)),(to_sfixed_a(0.0001361458853352815)),(to_sfixed_a(0.00012064223847119138)),(to_sfixed_a(2.1526919226744212e-05)),(to_sfixed_a(0.00012985059584025294)),(to_sfixed_a(8.556085958844051e-05)),(to_sfixed_a(-4.118205470149405e-05)),(to_sfixed_a(7.048965926514938e-05)),(to_sfixed_a(-0.0002593253448139876)),(to_sfixed_a(-0.0002202901232521981)),(to_sfixed_a(0.00017904562992043793)),(to_sfixed_a(-2.1121402824064717e-05)),(to_sfixed_a(1.6710211639292538e-05)),(to_sfixed_a(-0.00013929454144090414)),(to_sfixed_a(0.00034093804424628615)),(to_sfixed_a(-0.00011198910215171054)),(to_sfixed_a(0.00010821832256624475)),(to_sfixed_a(8.433286711806431e-05)),(to_sfixed_a(2.1177769667701796e-05)),(to_sfixed_a(-4.3878757423954085e-05)),(to_sfixed_a(7.630157779203728e-05)),(to_sfixed_a(0.00011627909407252446)),(to_sfixed_a(-3.961663242080249e-05)),(to_sfixed_a(6.997044692980126e-05)));

    constant weight_n0_11 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(6.703292456222698e-05)),(to_sfixed_a(0.00013236847007647157)),(to_sfixed_a(-0.00015358341624960303)),(to_sfixed_a(1.988246185646858e-05)),(to_sfixed_a(6.447784835472703e-05)),(to_sfixed_a(6.59689394524321e-05)),(to_sfixed_a(-5.3440442570718005e-05)),(to_sfixed_a(-5.1180166337871924e-05)),(to_sfixed_a(-9.841524297371507e-05)),(to_sfixed_a(-1.724901630950626e-05)),(to_sfixed_a(-0.00016116799088194966)),(to_sfixed_a(-0.000164201992447488)),(to_sfixed_a(-1.6274645531666465e-05)),(to_sfixed_a(-6.232161831576377e-05)),(to_sfixed_a(-5.205855268286541e-05)),(to_sfixed_a(0.00021066378394607455)),(to_sfixed_a(-0.00037186365807428956)),(to_sfixed_a(1.8155040379497223e-05)),(to_sfixed_a(2.946914355561603e-05)),(to_sfixed_a(4.390818503452465e-05)),(to_sfixed_a(0.00017772780847735703)),(to_sfixed_a(0.00012215215247124434)),(to_sfixed_a(-1.57401282194769e-05)),(to_sfixed_a(-8.137107943184674e-05)),(to_sfixed_a(-0.00016722279542591423)),(to_sfixed_a(9.635537571739405e-05)),(to_sfixed_a(-0.00018413906218484044)),(to_sfixed_a(-0.00013380507880356163)),(to_sfixed_a(3.7368819903349504e-05)),(to_sfixed_a(0.00021396417287178338)),(to_sfixed_a(0.00011107585305580869)),(to_sfixed_a(-4.276941763237119e-05)),(to_sfixed_a(-0.00040116862510330975)),(to_sfixed_a(-6.640081119257957e-05)),(to_sfixed_a(0.000119886921311263)),(to_sfixed_a(-7.035119779175147e-05)),(to_sfixed_a(0.00014807205297984183)),(to_sfixed_a(0.00013334036339074373)),(to_sfixed_a(8.039919339353219e-05)),(to_sfixed_a(-0.00022677840024698526)),(to_sfixed_a(-9.975793363992125e-05)),(to_sfixed_a(-2.332269650651142e-05)),(to_sfixed_a(-7.773618563078344e-05)),(to_sfixed_a(-8.31343641038984e-05)),(to_sfixed_a(3.502862819004804e-05)),(to_sfixed_a(-3.4304587188671576e-06)),(to_sfixed_a(3.2848962291609496e-05)),(to_sfixed_a(-6.703105464112014e-05)),(to_sfixed_a(0.0003603707591537386)),(to_sfixed_a(4.052164149470627e-05)),(to_sfixed_a(-5.7667461078381166e-05)),(to_sfixed_a(-1.7135766938736197e-06)),(to_sfixed_a(-9.279757796321064e-05)),(to_sfixed_a(-0.00010561929229879752)),(to_sfixed_a(9.178018081001937e-05)),(to_sfixed_a(-0.0001141806787927635)),(to_sfixed_a(-0.00015011581126600504)),(to_sfixed_a(-3.724509952007793e-05)),(to_sfixed_a(0.00021549088705796748)),(to_sfixed_a(0.00020513722847681493)),(to_sfixed_a(-0.00017847541312221438)),(to_sfixed_a(2.909327668021433e-05)),(to_sfixed_a(3.8314086850732565e-05)),(to_sfixed_a(-0.00011489225289551541)),(to_sfixed_a(2.2543642899108818e-06)),(to_sfixed_a(-0.0001659437984926626)),(to_sfixed_a(7.859797187848017e-05)),(to_sfixed_a(6.131864938652143e-05)),(to_sfixed_a(7.411876867990941e-05)),(to_sfixed_a(0.020306773483753204)),(to_sfixed_a(-3.265105624450371e-05)),(to_sfixed_a(0.00013258644321467727)),(to_sfixed_a(-7.301336154341698e-05)),(to_sfixed_a(7.99205809016712e-05)),(to_sfixed_a(7.983885734574869e-05)),(to_sfixed_a(-0.00021458785340655595)),(to_sfixed_a(2.578912244644016e-05)),(to_sfixed_a(-0.00010306940384907648)),(to_sfixed_a(-0.00017343081708531827)),(to_sfixed_a(0.0001618058158783242)),(to_sfixed_a(-1.969275763258338e-05)),(to_sfixed_a(0.00017051948816515505)),(to_sfixed_a(1.6964946553343907e-05)),(to_sfixed_a(0.00011104207078460604)),(to_sfixed_a(-9.629760461393744e-05)),(to_sfixed_a(0.00027848940226249397)),(to_sfixed_a(-2.7669309929478914e-05)),(to_sfixed_a(-0.00013442919589579105)),(to_sfixed_a(-0.00016335835971403867)),(to_sfixed_a(-9.557720477459952e-05)),(to_sfixed_a(0.00010799035953823477)),(to_sfixed_a(1.5704226825619116e-05)),(to_sfixed_a(0.0647682473063469)),(to_sfixed_a(-0.00010798352741403505)),(to_sfixed_a(0.07321856170892715)),(to_sfixed_a(0.05462300777435303)),(to_sfixed_a(0.12690916657447815)),(to_sfixed_a(-0.019230082631111145)),(to_sfixed_a(0.11438996344804764)),(to_sfixed_a(-0.11327061057090759)),(to_sfixed_a(-0.009814241901040077)),(to_sfixed_a(-0.04849432408809662)),(to_sfixed_a(-0.005415941122919321)),(to_sfixed_a(0.021056871861219406)),(to_sfixed_a(-0.01036064326763153)),(to_sfixed_a(-0.021450962871313095)),(to_sfixed_a(3.752634074771777e-05)),(to_sfixed_a(-3.128215030301362e-05)),(to_sfixed_a(0.0001151998876594007)),(to_sfixed_a(3.293605914223008e-05)),(to_sfixed_a(0.00010556426423136145)),(to_sfixed_a(3.769346221815795e-05)),(to_sfixed_a(-0.00015124735364224762)),(to_sfixed_a(9.270329610444605e-05)),(to_sfixed_a(0.00011633073154371232)),(to_sfixed_a(0.00013963511446490884)),(to_sfixed_a(-0.0002444522688165307)),(to_sfixed_a(6.1017999541945755e-06)),(to_sfixed_a(-0.0003171116695739329)),(to_sfixed_a(0.017818670719861984)),(to_sfixed_a(0.058501385152339935)),(to_sfixed_a(0.09116803109645844)),(to_sfixed_a(0.16754750907421112)),(to_sfixed_a(0.11481811851263046)),(to_sfixed_a(0.11035217344760895)),(to_sfixed_a(0.08177780359983444)),(to_sfixed_a(-0.01100747101008892)),(to_sfixed_a(-0.3692876696586609)),(to_sfixed_a(-0.11116470396518707)),(to_sfixed_a(-0.19133014976978302)),(to_sfixed_a(-0.17302720248699188)),(to_sfixed_a(0.04673213139176369)),(to_sfixed_a(0.003987249452620745)),(to_sfixed_a(0.019680721685290337)),(to_sfixed_a(-0.04970656707882881)),(to_sfixed_a(-9.836866229306906e-05)),(to_sfixed_a(0.0008227492799051106)),(to_sfixed_a(0.00015865822206251323)),(to_sfixed_a(8.526205056114122e-05)),(to_sfixed_a(-0.00012969778617843986)),(to_sfixed_a(0.00013436787412501872)),(to_sfixed_a(-1.3365124686970375e-06)),(to_sfixed_a(8.09061987183668e-07)),(to_sfixed_a(-0.0001279782154597342)),(to_sfixed_a(-0.0011861745733767748)),(to_sfixed_a(0.01943226158618927)),(to_sfixed_a(-0.011106463149189949)),(to_sfixed_a(0.10644108802080154)),(to_sfixed_a(0.038785215467214584)),(to_sfixed_a(0.0253800880163908)),(to_sfixed_a(0.05643896386027336)),(to_sfixed_a(-0.056052278727293015)),(to_sfixed_a(0.13788145780563354)),(to_sfixed_a(-0.008151471614837646)),(to_sfixed_a(0.0045862952247262)),(to_sfixed_a(0.0464305616915226)),(to_sfixed_a(-0.044038549065589905)),(to_sfixed_a(-0.11691080033779144)),(to_sfixed_a(-0.43188774585723877)),(to_sfixed_a(0.07246813178062439)),(to_sfixed_a(-0.10721521079540253)),(to_sfixed_a(-0.08698198944330215)),(to_sfixed_a(0.004153075627982616)),(to_sfixed_a(-0.032037317752838135)),(to_sfixed_a(-0.002651739865541458)),(to_sfixed_a(-0.0006875052931718528)),(to_sfixed_a(-6.476537964772433e-05)),(to_sfixed_a(7.088028360158205e-05)),(to_sfixed_a(-1.5018906196928583e-05)),(to_sfixed_a(0.00017214119725394994)),(to_sfixed_a(3.7164434615988284e-05)),(to_sfixed_a(-0.0001328714279225096)),(to_sfixed_a(0.000349697977071628)),(to_sfixed_a(0.02036404237151146)),(to_sfixed_a(-0.05383874848484993)),(to_sfixed_a(0.045564159750938416)),(to_sfixed_a(0.001581484917551279)),(to_sfixed_a(0.11181525141000748)),(to_sfixed_a(0.04333137348294258)),(to_sfixed_a(0.019368642941117287)),(to_sfixed_a(0.1842288225889206)),(to_sfixed_a(-0.030585335567593575)),(to_sfixed_a(0.042792193591594696)),(to_sfixed_a(-0.16364815831184387)),(to_sfixed_a(-0.1566053032875061)),(to_sfixed_a(-0.1480056494474411)),(to_sfixed_a(-0.2051960974931717)),(to_sfixed_a(-0.2808215320110321)),(to_sfixed_a(-0.19870483875274658)),(to_sfixed_a(-0.0464489683508873)),(to_sfixed_a(-0.01647358015179634)),(to_sfixed_a(0.1973370760679245)),(to_sfixed_a(-0.0002621005696710199)),(to_sfixed_a(0.00022704659204464406)),(to_sfixed_a(0.0002564621390774846)),(to_sfixed_a(-7.215799996629357e-05)),(to_sfixed_a(-0.00014630799705628306)),(to_sfixed_a(-0.00023647338093724102)),(to_sfixed_a(0.00034318052348680794)),(to_sfixed_a(0.00010242026473861188)),(to_sfixed_a(-0.00011750005796784535)),(to_sfixed_a(0.01115400530397892)),(to_sfixed_a(-0.050814274698495865)),(to_sfixed_a(0.19203554093837738)),(to_sfixed_a(-0.08302269130945206)),(to_sfixed_a(-0.05693327635526657)),(to_sfixed_a(0.16635379195213318)),(to_sfixed_a(0.2403600960969925)),(to_sfixed_a(0.11671086400747299)),(to_sfixed_a(0.08353859931230545)),(to_sfixed_a(-0.02080114372074604)),(to_sfixed_a(0.043176375329494476)),(to_sfixed_a(-0.07348379492759705)),(to_sfixed_a(-0.12756215035915375)),(to_sfixed_a(-0.16353733837604523)),(to_sfixed_a(-0.28994831442832947)),(to_sfixed_a(0.14168789982795715)),(to_sfixed_a(-0.1787661612033844)),(to_sfixed_a(0.2162739783525467)),(to_sfixed_a(0.0440739281475544)),(to_sfixed_a(0.10977941751480103)),(to_sfixed_a(0.006740146782249212)),(to_sfixed_a(-3.1736450182506815e-05)),(to_sfixed_a(1.3896941709390376e-05)),(to_sfixed_a(-3.304715210106224e-05)),(to_sfixed_a(0.00011163028102600947)),(to_sfixed_a(-2.613678589113988e-05)),(to_sfixed_a(7.262463441293221e-06)),(to_sfixed_a(0.030198566615581512)),(to_sfixed_a(0.018498588353395462)),(to_sfixed_a(0.05592908337712288)),(to_sfixed_a(-0.11518460512161255)),(to_sfixed_a(0.07462962716817856)),(to_sfixed_a(-0.010263331234455109)),(to_sfixed_a(-0.011938032694160938)),(to_sfixed_a(-0.014211450703442097)),(to_sfixed_a(-0.016066091135144234)),(to_sfixed_a(0.06979876756668091)),(to_sfixed_a(0.016692494973540306)),(to_sfixed_a(0.22407743334770203)),(to_sfixed_a(0.09120912849903107)),(to_sfixed_a(-0.06515047699213028)),(to_sfixed_a(-0.064290352165699)),(to_sfixed_a(-0.03726911172270775)),(to_sfixed_a(0.3203711211681366)),(to_sfixed_a(0.14770261943340302)),(to_sfixed_a(-0.12186412513256073)),(to_sfixed_a(0.08187846094369888)),(to_sfixed_a(0.22178059816360474)),(to_sfixed_a(0.08278214931488037)),(to_sfixed_a(6.286461575655267e-05)),(to_sfixed_a(-1.0378938242183722e-07)),(to_sfixed_a(7.862596976337954e-05)),(to_sfixed_a(0.00010497659241082147)),(to_sfixed_a(8.977533434517682e-05)),(to_sfixed_a(-0.0002060595143120736)),(to_sfixed_a(0.002836767351254821)),(to_sfixed_a(0.057141367346048355)),(to_sfixed_a(-0.05709734186530113)),(to_sfixed_a(0.14981333911418915)),(to_sfixed_a(-0.07306580245494843)),(to_sfixed_a(0.03568732738494873)),(to_sfixed_a(0.08897527307271957)),(to_sfixed_a(-0.04133202135562897)),(to_sfixed_a(-0.10969473421573639)),(to_sfixed_a(-0.11483973264694214)),(to_sfixed_a(0.042761776596307755)),(to_sfixed_a(0.06319583207368851)),(to_sfixed_a(-0.1887047290802002)),(to_sfixed_a(-0.1350478082895279)),(to_sfixed_a(-0.06877636164426804)),(to_sfixed_a(-0.12398234009742737)),(to_sfixed_a(-0.13076816499233246)),(to_sfixed_a(0.01236043218523264)),(to_sfixed_a(0.03798854723572731)),(to_sfixed_a(0.2709287106990814)),(to_sfixed_a(0.23087111115455627)),(to_sfixed_a(-4.6254106564447284e-05)),(to_sfixed_a(-0.00012813002103939652)),(to_sfixed_a(5.722166315536015e-05)),(to_sfixed_a(2.567105730122421e-05)),(to_sfixed_a(0.0001157042570412159)),(to_sfixed_a(7.654057299077976e-06)),(to_sfixed_a(-7.461729546776041e-05)),(to_sfixed_a(0.00011092412023572251)),(to_sfixed_a(-0.007947871461510658)),(to_sfixed_a(0.08578720688819885)),(to_sfixed_a(-0.03894553333520889)),(to_sfixed_a(-0.07229649275541306)),(to_sfixed_a(-0.05902962386608124)),(to_sfixed_a(-0.014823062345385551)),(to_sfixed_a(-0.1081462949514389)),(to_sfixed_a(-0.19224824011325836)),(to_sfixed_a(-0.19286060333251953)),(to_sfixed_a(-0.5789056420326233)),(to_sfixed_a(-0.2806614339351654)),(to_sfixed_a(-0.4445139765739441)),(to_sfixed_a(-0.2321346253156662)),(to_sfixed_a(-0.21038833260536194)),(to_sfixed_a(-0.13678331673145294)),(to_sfixed_a(0.2339680790901184)),(to_sfixed_a(0.24519474804401398)),(to_sfixed_a(-0.13846077024936676)),(to_sfixed_a(0.024320807307958603)),(to_sfixed_a(0.05869666114449501)),(to_sfixed_a(0.012722214683890343)),(to_sfixed_a(-0.0002058198006125167)),(to_sfixed_a(2.4840204787324183e-05)),(to_sfixed_a(-3.540503166732378e-05)),(to_sfixed_a(-0.00013361574383452535)),(to_sfixed_a(-8.51655422593467e-05)),(to_sfixed_a(-0.0348338708281517)),(to_sfixed_a(0.039021480828523636)),(to_sfixed_a(-0.15145480632781982)),(to_sfixed_a(0.04444853216409683)),(to_sfixed_a(0.025942819193005562)),(to_sfixed_a(-0.009920959360897541)),(to_sfixed_a(-0.0041197072714567184)),(to_sfixed_a(-0.07484022527933121)),(to_sfixed_a(-0.03183968737721443)),(to_sfixed_a(-0.30739012360572815)),(to_sfixed_a(-0.3973948657512665)),(to_sfixed_a(-0.48653122782707214)),(to_sfixed_a(-0.3972632586956024)),(to_sfixed_a(-0.23149394989013672)),(to_sfixed_a(-0.3526701331138611)),(to_sfixed_a(-0.24244074523448944)),(to_sfixed_a(-0.13885289430618286)),(to_sfixed_a(-0.008440311998128891)),(to_sfixed_a(-0.1263372302055359)),(to_sfixed_a(0.013247225433588028)),(to_sfixed_a(-0.11089513450860977)),(to_sfixed_a(-0.07827761769294739)),(to_sfixed_a(-0.0001239192788489163)),(to_sfixed_a(4.022594657726586e-05)),(to_sfixed_a(-0.00042335165198892355)),(to_sfixed_a(0.0001151276082964614)),(to_sfixed_a(2.5139908757410012e-05)),(to_sfixed_a(-0.00021310560987330973)),(to_sfixed_a(-0.0002749450213741511)),(to_sfixed_a(-0.1598832607269287)),(to_sfixed_a(-0.17524220049381256)),(to_sfixed_a(-0.08079210668802261)),(to_sfixed_a(0.12921005487442017)),(to_sfixed_a(-0.04998861998319626)),(to_sfixed_a(0.12352200597524643)),(to_sfixed_a(-0.039511408656835556)),(to_sfixed_a(-0.2868057191371918)),(to_sfixed_a(-0.39728137850761414)),(to_sfixed_a(-0.7894819974899292)),(to_sfixed_a(-0.16102807223796844)),(to_sfixed_a(-0.03474639356136322)),(to_sfixed_a(-0.09781577438116074)),(to_sfixed_a(-0.09114661812782288)),(to_sfixed_a(-0.03409635275602341)),(to_sfixed_a(0.15154586732387543)),(to_sfixed_a(-0.13833162188529968)),(to_sfixed_a(-0.08842732757329941)),(to_sfixed_a(-0.036779891699552536)),(to_sfixed_a(-0.14752623438835144)),(to_sfixed_a(-0.258957177400589)),(to_sfixed_a(-8.22983281523193e-07)),(to_sfixed_a(-0.0003442050365265459)),(to_sfixed_a(0.00023588904878124595)),(to_sfixed_a(8.617124694865197e-05)),(to_sfixed_a(5.914382199989632e-05)),(to_sfixed_a(0.0003648996935226023)),(to_sfixed_a(-0.00018820317927747965)),(to_sfixed_a(-0.10550110787153244)),(to_sfixed_a(-0.09019511193037033)),(to_sfixed_a(0.2471553087234497)),(to_sfixed_a(0.0781632661819458)),(to_sfixed_a(0.35438618063926697)),(to_sfixed_a(0.10124225914478302)),(to_sfixed_a(-0.10307753831148148)),(to_sfixed_a(-0.4944632053375244)),(to_sfixed_a(-0.35787543654441833)),(to_sfixed_a(-0.33261728286743164)),(to_sfixed_a(-0.08271774649620056)),(to_sfixed_a(0.0893745869398117)),(to_sfixed_a(0.09724169224500656)),(to_sfixed_a(-0.03184376657009125)),(to_sfixed_a(0.022719785571098328)),(to_sfixed_a(0.09028726816177368)),(to_sfixed_a(-0.1119123324751854)),(to_sfixed_a(-0.1220019981265068)),(to_sfixed_a(-0.02365339919924736)),(to_sfixed_a(-0.1022903248667717)),(to_sfixed_a(0.08070658892393112)),(to_sfixed_a(-0.001951283193193376)),(to_sfixed_a(-0.0014353691367432475)),(to_sfixed_a(5.1090275519527495e-05)),(to_sfixed_a(-0.00017231536912731826)),(to_sfixed_a(-0.00012463118764571846)),(to_sfixed_a(-0.0002638647856656462)),(to_sfixed_a(-0.0001445080852136016)),(to_sfixed_a(-0.00014563863805960864)),(to_sfixed_a(0.2801639437675476)),(to_sfixed_a(0.17342111468315125)),(to_sfixed_a(0.15456527471542358)),(to_sfixed_a(-0.08930253237485886)),(to_sfixed_a(0.13499686121940613)),(to_sfixed_a(-0.34800267219543457)),(to_sfixed_a(-0.27190226316452026)),(to_sfixed_a(-0.644034206867218)),(to_sfixed_a(-0.0833592563867569)),(to_sfixed_a(0.37743356823921204)),(to_sfixed_a(0.17277997732162476)),(to_sfixed_a(0.29446732997894287)),(to_sfixed_a(-0.01984400488436222)),(to_sfixed_a(-0.01656242087483406)),(to_sfixed_a(-0.026091886684298515)),(to_sfixed_a(-0.17498071491718292)),(to_sfixed_a(-0.13771013915538788)),(to_sfixed_a(0.15690378844738007)),(to_sfixed_a(0.13094890117645264)),(to_sfixed_a(-0.10377217084169388)),(to_sfixed_a(-0.00037622355739586055)),(to_sfixed_a(-0.00012452503142412752)),(to_sfixed_a(1.6550176951568574e-05)),(to_sfixed_a(-0.00010856542940018699)),(to_sfixed_a(5.236043580225669e-05)),(to_sfixed_a(-1.5078084288688842e-05)),(to_sfixed_a(-1.5099353731784504e-05)),(to_sfixed_a(0.019976062700152397)),(to_sfixed_a(-0.007283024489879608)),(to_sfixed_a(0.028963444754481316)),(to_sfixed_a(0.12818647921085358)),(to_sfixed_a(0.056437768042087555)),(to_sfixed_a(-0.10858757048845291)),(to_sfixed_a(-0.19871564209461212)),(to_sfixed_a(-0.21547625958919525)),(to_sfixed_a(-0.3836258351802826)),(to_sfixed_a(0.3631053566932678)),(to_sfixed_a(0.2600094974040985)),(to_sfixed_a(0.1318366527557373)),(to_sfixed_a(-0.005347905680537224)),(to_sfixed_a(-0.10623374581336975)),(to_sfixed_a(0.08319926261901855)),(to_sfixed_a(-0.33406174182891846)),(to_sfixed_a(-0.3710283041000366)),(to_sfixed_a(-0.13402396440505981)),(to_sfixed_a(0.05593673139810562)),(to_sfixed_a(0.14250829815864563)),(to_sfixed_a(0.16484007239341736)),(to_sfixed_a(-0.00016781067824922502)),(to_sfixed_a(0.00017197290435433388)),(to_sfixed_a(0.00023841179790906608)),(to_sfixed_a(0.00020665896590799093)),(to_sfixed_a(0.00020007988496217877)),(to_sfixed_a(-0.00012062871974194422)),(to_sfixed_a(-0.001505560358054936)),(to_sfixed_a(-0.17195233702659607)),(to_sfixed_a(-0.2775539457798004)),(to_sfixed_a(-0.1261977106332779)),(to_sfixed_a(0.06438707560300827)),(to_sfixed_a(0.03780142590403557)),(to_sfixed_a(-0.07445657253265381)),(to_sfixed_a(-0.1417328417301178)),(to_sfixed_a(0.00509722949936986)),(to_sfixed_a(0.26037928462028503)),(to_sfixed_a(0.6071804165840149)),(to_sfixed_a(0.1441268026828766)),(to_sfixed_a(0.2833947539329529)),(to_sfixed_a(0.05672907456755638)),(to_sfixed_a(0.14467285573482513)),(to_sfixed_a(-0.258968323469162)),(to_sfixed_a(-0.5233184695243835)),(to_sfixed_a(-0.5129058957099915)),(to_sfixed_a(-0.26592394709587097)),(to_sfixed_a(-0.18015417456626892)),(to_sfixed_a(-0.0659533217549324)),(to_sfixed_a(0.14042644202709198)),(to_sfixed_a(0.020991230383515358)),(to_sfixed_a(-7.436464511556551e-05)),(to_sfixed_a(-0.00012087780487490818)),(to_sfixed_a(5.27523152413778e-05)),(to_sfixed_a(0.00026060501113533974)),(to_sfixed_a(-0.0009075241978280246)),(to_sfixed_a(-0.0019158812938258052)),(to_sfixed_a(-0.016111643984913826)),(to_sfixed_a(-0.022696686908602715)),(to_sfixed_a(0.13814669847488403)),(to_sfixed_a(-0.20767663419246674)),(to_sfixed_a(-0.0004793170664925128)),(to_sfixed_a(-0.17501524090766907)),(to_sfixed_a(-0.12042620033025742)),(to_sfixed_a(0.34112945199012756)),(to_sfixed_a(0.5807918906211853)),(to_sfixed_a(0.3852315843105316)),(to_sfixed_a(0.17292112112045288)),(to_sfixed_a(0.33319881558418274)),(to_sfixed_a(0.12472528964281082)),(to_sfixed_a(-0.1074962466955185)),(to_sfixed_a(-0.12946853041648865)),(to_sfixed_a(-0.09589410573244095)),(to_sfixed_a(0.01343740988522768)),(to_sfixed_a(0.08598475158214569)),(to_sfixed_a(0.01860337145626545)),(to_sfixed_a(0.008675464428961277)),(to_sfixed_a(1.2854237866122276e-05)),(to_sfixed_a(-6.443688471335918e-05)),(to_sfixed_a(-3.0150275051710196e-05)),(to_sfixed_a(-1.0784275218611583e-05)),(to_sfixed_a(-5.874927592230961e-05)),(to_sfixed_a(3.441819717409089e-05)),(to_sfixed_a(-3.185277819284238e-05)),(to_sfixed_a(-0.019278965890407562)),(to_sfixed_a(0.12508006393909454)),(to_sfixed_a(0.08130098134279251)),(to_sfixed_a(-0.11983219534158707)),(to_sfixed_a(-0.06344064325094223)),(to_sfixed_a(-0.15329979360103607)),(to_sfixed_a(-0.09371259063482285)),(to_sfixed_a(0.2270938754081726)),(to_sfixed_a(0.21518082916736603)),(to_sfixed_a(0.47422337532043457)),(to_sfixed_a(0.5497372150421143)),(to_sfixed_a(0.22920574247837067)),(to_sfixed_a(0.0781046599149704)),(to_sfixed_a(0.22721825540065765)),(to_sfixed_a(-0.052024245262145996)),(to_sfixed_a(-0.18069623410701752)),(to_sfixed_a(-0.3830210268497467)),(to_sfixed_a(-0.15345898270606995)),(to_sfixed_a(-0.07849694788455963)),(to_sfixed_a(0.029115106910467148)),(to_sfixed_a(0.12202061712741852)),(to_sfixed_a(0.038202930241823196)),(to_sfixed_a(-9.004570165416226e-05)),(to_sfixed_a(5.435609637061134e-05)),(to_sfixed_a(-0.00017319750622846186)),(to_sfixed_a(0.00045110913924872875)),(to_sfixed_a(0.000311816023895517)),(to_sfixed_a(-0.00018705583352129906)),(to_sfixed_a(-0.09336014091968536)),(to_sfixed_a(-0.004206148907542229)),(to_sfixed_a(-0.15611816942691803)),(to_sfixed_a(-0.07102347910404205)),(to_sfixed_a(-0.20167817175388336)),(to_sfixed_a(-0.33802857995033264)),(to_sfixed_a(-0.19971801340579987)),(to_sfixed_a(0.15716294944286346)),(to_sfixed_a(0.43328657746315)),(to_sfixed_a(0.2977750599384308)),(to_sfixed_a(0.35763901472091675)),(to_sfixed_a(0.533473551273346)),(to_sfixed_a(0.21084094047546387)),(to_sfixed_a(0.015117869712412357)),(to_sfixed_a(0.025822091847658157)),(to_sfixed_a(-0.12157543003559113)),(to_sfixed_a(0.05910778045654297)),(to_sfixed_a(0.12357475608587265)),(to_sfixed_a(0.1161157637834549)),(to_sfixed_a(0.09173659980297089)),(to_sfixed_a(0.025347460061311722)),(to_sfixed_a(0.00014280292089097202)),(to_sfixed_a(0.00014784271479584277)),(to_sfixed_a(3.283515980001539e-05)),(to_sfixed_a(-4.202771742711775e-05)),(to_sfixed_a(-0.00012554459681268781)),(to_sfixed_a(-0.00011546174937393516)),(to_sfixed_a(0.0001493857562309131)),(to_sfixed_a(-9.235337347490713e-05)),(to_sfixed_a(-0.018770700320601463)),(to_sfixed_a(-0.01817285642027855)),(to_sfixed_a(-0.3253028988838196)),(to_sfixed_a(-0.26362666487693787)),(to_sfixed_a(0.04740552976727486)),(to_sfixed_a(-0.021243009716272354)),(to_sfixed_a(0.027279485017061234)),(to_sfixed_a(0.20779599249362946)),(to_sfixed_a(0.16925588250160217)),(to_sfixed_a(0.16076281666755676)),(to_sfixed_a(0.3422617018222809)),(to_sfixed_a(0.11969736218452454)),(to_sfixed_a(0.05285540968179703)),(to_sfixed_a(-0.04520072042942047)),(to_sfixed_a(-0.2569199204444885)),(to_sfixed_a(0.17958992719650269)),(to_sfixed_a(0.012035537511110306)),(to_sfixed_a(-0.13464975357055664)),(to_sfixed_a(-0.022436505183577538)),(to_sfixed_a(0.14916476607322693)),(to_sfixed_a(0.08963516354560852)),(to_sfixed_a(0.00012916956620756537)),(to_sfixed_a(-3.120779729215428e-05)),(to_sfixed_a(-0.00020486248831730336)),(to_sfixed_a(0.00014300504699349403)),(to_sfixed_a(9.686580597190186e-05)),(to_sfixed_a(0.00011265480861766264)),(to_sfixed_a(-0.00019192487525288016)),(to_sfixed_a(0.005575473420321941)),(to_sfixed_a(-0.0010178042575716972)),(to_sfixed_a(-0.2015335112810135)),(to_sfixed_a(-0.176333487033844)),(to_sfixed_a(0.01111865695565939)),(to_sfixed_a(-0.03969307616353035)),(to_sfixed_a(0.11844862997531891)),(to_sfixed_a(0.228862464427948)),(to_sfixed_a(0.08513885736465454)),(to_sfixed_a(0.0010369842639192939)),(to_sfixed_a(-0.12757661938667297)),(to_sfixed_a(0.03435681015253067)),(to_sfixed_a(-0.047979287803173065)),(to_sfixed_a(-0.14973540604114532)),(to_sfixed_a(-0.1123218685388565)),(to_sfixed_a(-0.10634281486272812)),(to_sfixed_a(-0.010401817969977856)),(to_sfixed_a(-0.00399735989049077)),(to_sfixed_a(0.0751107856631279)),(to_sfixed_a(-0.0007241012062877417)),(to_sfixed_a(0.022771185263991356)),(to_sfixed_a(0.00011002661631209776)),(to_sfixed_a(0.00020342539937701076)),(to_sfixed_a(9.182263602269813e-05)),(to_sfixed_a(-0.00026431685546413064)),(to_sfixed_a(-0.0001287884806515649)),(to_sfixed_a(0.00011893431656062603)),(to_sfixed_a(8.964361040852964e-05)),(to_sfixed_a(0.00012131199036957696)),(to_sfixed_a(0.03535859286785126)),(to_sfixed_a(-0.031319376081228256)),(to_sfixed_a(-0.0962207019329071)),(to_sfixed_a(0.14355091750621796)),(to_sfixed_a(0.0017964949365705252)),(to_sfixed_a(0.06071952357888222)),(to_sfixed_a(0.10114956647157669)),(to_sfixed_a(0.04614420235157013)),(to_sfixed_a(0.06133975088596344)),(to_sfixed_a(-0.018733028322458267)),(to_sfixed_a(-0.0505700521171093)),(to_sfixed_a(-0.3757592737674713)),(to_sfixed_a(-0.13067597150802612)),(to_sfixed_a(-0.04053855314850807)),(to_sfixed_a(-0.003644123673439026)),(to_sfixed_a(-0.03250717744231224)),(to_sfixed_a(0.035385068506002426)),(to_sfixed_a(0.07034853845834732)),(to_sfixed_a(0.006103897467255592)),(to_sfixed_a(-0.0001450333365937695)),(to_sfixed_a(0.00022498144244309515)),(to_sfixed_a(-2.8997928893659264e-05)),(to_sfixed_a(-7.426966476486996e-05)),(to_sfixed_a(-6.225582910701632e-05)),(to_sfixed_a(5.59984655410517e-05)),(to_sfixed_a(4.376814467832446e-05)),(to_sfixed_a(-7.656412344658747e-05)),(to_sfixed_a(0.00042307464173063636)),(to_sfixed_a(-0.0011287882225587964)),(to_sfixed_a(0.0946907252073288)),(to_sfixed_a(0.04943099245429039)),(to_sfixed_a(-0.17834000289440155)),(to_sfixed_a(0.169269859790802)),(to_sfixed_a(-0.005543238017708063)),(to_sfixed_a(-0.2254108041524887)),(to_sfixed_a(-0.06272945553064346)),(to_sfixed_a(-0.012903690338134766)),(to_sfixed_a(-0.11944825947284698)),(to_sfixed_a(-0.10070837289094925)),(to_sfixed_a(-0.21558628976345062)),(to_sfixed_a(-0.4525824189186096)),(to_sfixed_a(-0.015896592289209366)),(to_sfixed_a(0.07129982858896255)),(to_sfixed_a(-0.1313546597957611)),(to_sfixed_a(0.13017967343330383)),(to_sfixed_a(0.015059389173984528)),(to_sfixed_a(0.09057288616895676)),(to_sfixed_a(0.00018598638416733593)),(to_sfixed_a(9.92765199043788e-05)),(to_sfixed_a(0.0001839486649259925)),(to_sfixed_a(-4.2615785787347704e-05)),(to_sfixed_a(9.481388406129554e-05)),(to_sfixed_a(-2.8570188987941947e-06)),(to_sfixed_a(1.921594957821071e-06)),(to_sfixed_a(-1.48194260418677e-06)),(to_sfixed_a(-0.023916032165288925)),(to_sfixed_a(-0.005057742353528738)),(to_sfixed_a(-0.10043633729219437)),(to_sfixed_a(-0.17341294884681702)),(to_sfixed_a(0.16092896461486816)),(to_sfixed_a(-0.057149093598127365)),(to_sfixed_a(-0.03106255829334259)),(to_sfixed_a(0.1320662945508957)),(to_sfixed_a(-0.14857518672943115)),(to_sfixed_a(-0.2698337435722351)),(to_sfixed_a(-0.11527981609106064)),(to_sfixed_a(-0.004181308671832085)),(to_sfixed_a(-0.5426103472709656)),(to_sfixed_a(-0.30782797932624817)),(to_sfixed_a(-0.14534616470336914)),(to_sfixed_a(-0.054519493132829666)),(to_sfixed_a(-0.007052022032439709)),(to_sfixed_a(0.12272224575281143)),(to_sfixed_a(0.052716728299856186)),(to_sfixed_a(0.007929109036922455)),(to_sfixed_a(0.00012772373156622052)),(to_sfixed_a(2.0722459339594934e-06)),(to_sfixed_a(0.0002482403360772878)),(to_sfixed_a(7.550695590907708e-05)),(to_sfixed_a(-0.00015352378250099719)),(to_sfixed_a(0.00015115660789888352)),(to_sfixed_a(-2.8512675271485932e-05)),(to_sfixed_a(-6.938957812963054e-05)),(to_sfixed_a(0.00020401008077897131)),(to_sfixed_a(-0.06460591405630112)),(to_sfixed_a(-0.05996307358145714)),(to_sfixed_a(-0.08043655753135681)),(to_sfixed_a(-0.299101859331131)),(to_sfixed_a(-0.09665792435407639)),(to_sfixed_a(-0.12889701128005981)),(to_sfixed_a(-0.010797332040965557)),(to_sfixed_a(0.10268425941467285)),(to_sfixed_a(-0.018986184149980545)),(to_sfixed_a(-0.10281452536582947)),(to_sfixed_a(-0.026198141276836395)),(to_sfixed_a(-0.11624689400196075)),(to_sfixed_a(-0.04708048328757286)),(to_sfixed_a(-0.0008613948011770844)),(to_sfixed_a(-0.02195163443684578)),(to_sfixed_a(-0.08667594194412231)),(to_sfixed_a(-4.2753697925945744e-05)),(to_sfixed_a(0.0016177009092643857)),(to_sfixed_a(0.0026862628292292356)),(to_sfixed_a(2.2600142983719707e-06)),(to_sfixed_a(-0.0001499909267295152)),(to_sfixed_a(0.00023235751723404974)),(to_sfixed_a(0.00019930208509322256)),(to_sfixed_a(0.00011933049972867593)),(to_sfixed_a(2.1708538042730652e-05)),(to_sfixed_a(-3.105566793237813e-05)),(to_sfixed_a(-9.587044041836634e-05)),(to_sfixed_a(-7.87419849075377e-05)),(to_sfixed_a(-0.0017507692100480199)),(to_sfixed_a(-0.0014863808173686266)),(to_sfixed_a(0.00010798466246342286)),(to_sfixed_a(0.00018526522035244852)),(to_sfixed_a(0.00014423874381463975)),(to_sfixed_a(-0.06688462197780609)),(to_sfixed_a(-0.006152601446956396)),(to_sfixed_a(-0.0010779885342344642)),(to_sfixed_a(-0.04332846775650978)),(to_sfixed_a(0.06458227336406708)),(to_sfixed_a(0.009721898473799229)),(to_sfixed_a(0.0019014952704310417)),(to_sfixed_a(-0.04883652552962303)),(to_sfixed_a(-0.06569210439920425)),(to_sfixed_a(0.0015404880978167057)),(to_sfixed_a(0.002039461862295866)),(to_sfixed_a(5.5159805924631655e-05)),(to_sfixed_a(-0.0001306843914790079)),(to_sfixed_a(3.902593380189501e-05)),(to_sfixed_a(8.61001099110581e-05)),(to_sfixed_a(0.00012470848741941154)),(to_sfixed_a(-0.0001121236928156577)),(to_sfixed_a(5.524785228772089e-05)),(to_sfixed_a(-0.00026179192354902625)),(to_sfixed_a(-0.000177179099409841)),(to_sfixed_a(-0.0001586285070516169)),(to_sfixed_a(-0.00017120626580435783)),(to_sfixed_a(-0.00022143698879517615)),(to_sfixed_a(-0.00021620336337946355)),(to_sfixed_a(0.00016464508371427655)),(to_sfixed_a(-0.00023238352150656283)),(to_sfixed_a(-0.00012439835700206459)),(to_sfixed_a(-0.00010093766468344256)),(to_sfixed_a(-2.6294626877643168e-05)),(to_sfixed_a(-0.0003077676519751549)),(to_sfixed_a(0.0001477215118939057)),(to_sfixed_a(-5.7572747209633235e-06)),(to_sfixed_a(-0.00032691951491869986)),(to_sfixed_a(-0.00017904059495776892)),(to_sfixed_a(0.00014127118629403412)),(to_sfixed_a(-5.556117685046047e-05)),(to_sfixed_a(0.0001249009947059676)),(to_sfixed_a(-9.102515832637437e-06)),(to_sfixed_a(-0.00011692672705976292)),(to_sfixed_a(-6.997038872214034e-05)),(to_sfixed_a(0.0001801229373086244)),(to_sfixed_a(0.0001753254618961364)),(to_sfixed_a(-6.166264029161539e-06)),(to_sfixed_a(0.00011116552195744589)),(to_sfixed_a(-6.275809573708102e-05)),(to_sfixed_a(-0.00011627922503976151)));

    constant weight_n0_12 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(3.184497109032236e-05)),(to_sfixed_a(4.6054199628997594e-05)),(to_sfixed_a(-7.755085243843496e-05)),(to_sfixed_a(-1.7451384337618947e-05)),(to_sfixed_a(-0.00023367578978650272)),(to_sfixed_a(-0.0001021123316604644)),(to_sfixed_a(-0.00017064860730897635)),(to_sfixed_a(-0.00012605448137037456)),(to_sfixed_a(-4.2140567529713735e-05)),(to_sfixed_a(8.718227036297321e-05)),(to_sfixed_a(6.711813330184668e-05)),(to_sfixed_a(0.0002707754902075976)),(to_sfixed_a(0.0002445914433337748)),(to_sfixed_a(6.941916944924742e-05)),(to_sfixed_a(0.0001503652601968497)),(to_sfixed_a(0.00010145197302335873)),(to_sfixed_a(1.3618257980851922e-05)),(to_sfixed_a(0.00017054274212568998)),(to_sfixed_a(-0.00018005151650868356)),(to_sfixed_a(-0.00010102202941197902)),(to_sfixed_a(-0.00017212766397278756)),(to_sfixed_a(5.039839743403718e-05)),(to_sfixed_a(0.00027206269442103803)),(to_sfixed_a(0.00016944206436164677)),(to_sfixed_a(8.304674702230841e-05)),(to_sfixed_a(5.4376956541091204e-05)),(to_sfixed_a(-0.0001316638954449445)),(to_sfixed_a(0.0003545984218362719)),(to_sfixed_a(9.802910062717274e-05)),(to_sfixed_a(0.00014994780940469354)),(to_sfixed_a(0.00015099297161214054)),(to_sfixed_a(-9.096010762732476e-05)),(to_sfixed_a(4.455732778296806e-06)),(to_sfixed_a(-0.0001084717659978196)),(to_sfixed_a(0.00024094354012049735)),(to_sfixed_a(1.651609636610374e-05)),(to_sfixed_a(0.0001595791254658252)),(to_sfixed_a(0.00016293727094307542)),(to_sfixed_a(2.2624257326242514e-05)),(to_sfixed_a(-0.00012951424287166446)),(to_sfixed_a(0.00013797671999782324)),(to_sfixed_a(3.695849591167644e-05)),(to_sfixed_a(-5.4389438446378335e-05)),(to_sfixed_a(-0.0001828258828027174)),(to_sfixed_a(2.7581574613577686e-05)),(to_sfixed_a(-0.00011144113523187116)),(to_sfixed_a(0.00016211633919738233)),(to_sfixed_a(-0.00039731673314236104)),(to_sfixed_a(-9.934236004482955e-05)),(to_sfixed_a(-1.9549406715668738e-05)),(to_sfixed_a(0.00022697969689033926)),(to_sfixed_a(6.567200762219727e-05)),(to_sfixed_a(-0.0005248560337349772)),(to_sfixed_a(-0.00015294666809495538)),(to_sfixed_a(-0.0001002134958980605)),(to_sfixed_a(0.00036806819844059646)),(to_sfixed_a(-4.6625224058516324e-05)),(to_sfixed_a(-4.887974137091078e-05)),(to_sfixed_a(6.598023173864931e-05)),(to_sfixed_a(-9.211754513671622e-05)),(to_sfixed_a(0.00011427720892243087)),(to_sfixed_a(-0.00014384396490640938)),(to_sfixed_a(2.987917287100572e-05)),(to_sfixed_a(-9.72207635641098e-05)),(to_sfixed_a(0.0002961610443890095)),(to_sfixed_a(-0.0001605077850399539)),(to_sfixed_a(-1.529419569124002e-05)),(to_sfixed_a(0.00015617730969097465)),(to_sfixed_a(-0.00019638589583337307)),(to_sfixed_a(-0.012816805392503738)),(to_sfixed_a(-1.227029861183837e-05)),(to_sfixed_a(-0.0001867350219981745)),(to_sfixed_a(3.621227006078698e-05)),(to_sfixed_a(1.730908297759015e-05)),(to_sfixed_a(-2.6624662496033125e-05)),(to_sfixed_a(-6.42220038571395e-05)),(to_sfixed_a(-0.00014037937216926366)),(to_sfixed_a(-6.174472946440801e-05)),(to_sfixed_a(-0.00023420536308549345)),(to_sfixed_a(-0.00024496056721545756)),(to_sfixed_a(-0.00013977628259453923)),(to_sfixed_a(0.00014693367120344192)),(to_sfixed_a(-3.802856326728943e-06)),(to_sfixed_a(-4.888753028353676e-05)),(to_sfixed_a(-8.870509918779135e-05)),(to_sfixed_a(-0.00024317298084497452)),(to_sfixed_a(-9.915485861711204e-05)),(to_sfixed_a(-1.51133053805097e-05)),(to_sfixed_a(-0.0001012053107842803)),(to_sfixed_a(8.36075414554216e-05)),(to_sfixed_a(-9.304851846536621e-05)),(to_sfixed_a(0.00016252617933787405)),(to_sfixed_a(0.01588832214474678)),(to_sfixed_a(0.00021949065558146685)),(to_sfixed_a(0.017847156152129173)),(to_sfixed_a(-0.12213881313800812)),(to_sfixed_a(-0.00026820850325748324)),(to_sfixed_a(-0.026700925081968307)),(to_sfixed_a(0.03169422224164009)),(to_sfixed_a(0.18210147321224213)),(to_sfixed_a(0.020042553544044495)),(to_sfixed_a(0.005510933697223663)),(to_sfixed_a(0.1710052341222763)),(to_sfixed_a(0.004687483422458172)),(to_sfixed_a(0.01656351238489151)),(to_sfixed_a(0.03342106193304062)),(to_sfixed_a(6.693774776067585e-05)),(to_sfixed_a(-0.00033065464231185615)),(to_sfixed_a(0.0002077193494187668)),(to_sfixed_a(0.00022034170979168266)),(to_sfixed_a(0.00022342149168252945)),(to_sfixed_a(6.0311602283036336e-05)),(to_sfixed_a(3.4244865219079657e-06)),(to_sfixed_a(4.9266498535871506e-05)),(to_sfixed_a(9.182167559629306e-05)),(to_sfixed_a(-0.00027503358433023095)),(to_sfixed_a(-0.00020000043150503188)),(to_sfixed_a(-0.00013584447151515633)),(to_sfixed_a(0.002063910709694028)),(to_sfixed_a(-0.060906361788511276)),(to_sfixed_a(0.032088879495859146)),(to_sfixed_a(0.022524749860167503)),(to_sfixed_a(-0.14970369637012482)),(to_sfixed_a(-0.0717422366142273)),(to_sfixed_a(0.10451149195432663)),(to_sfixed_a(0.23633430898189545)),(to_sfixed_a(0.20011471211910248)),(to_sfixed_a(0.024480868130922318)),(to_sfixed_a(0.2297038733959198)),(to_sfixed_a(-0.13705888390541077)),(to_sfixed_a(0.0694216638803482)),(to_sfixed_a(0.052919503301382065)),(to_sfixed_a(0.017762821167707443)),(to_sfixed_a(-0.0039193411357700825)),(to_sfixed_a(-0.03227551653981209)),(to_sfixed_a(0.0003225031541660428)),(to_sfixed_a(0.0005095448577776551)),(to_sfixed_a(5.086556120659225e-05)),(to_sfixed_a(-2.7882269932888448e-05)),(to_sfixed_a(0.00011076775990659371)),(to_sfixed_a(2.4310076696565375e-05)),(to_sfixed_a(-0.00024238227342721075)),(to_sfixed_a(8.714079740457237e-05)),(to_sfixed_a(3.363639552844688e-05)),(to_sfixed_a(0.00031311606289818883)),(to_sfixed_a(-0.07625837624073029)),(to_sfixed_a(0.019719399511814117)),(to_sfixed_a(-0.19850295782089233)),(to_sfixed_a(-0.07456929981708527)),(to_sfixed_a(-0.042409125715494156)),(to_sfixed_a(0.005700299050658941)),(to_sfixed_a(-0.08684897422790527)),(to_sfixed_a(-0.26028433442115784)),(to_sfixed_a(-0.26230472326278687)),(to_sfixed_a(0.004843317437916994)),(to_sfixed_a(0.10324103385210037)),(to_sfixed_a(0.18253789842128754)),(to_sfixed_a(-0.24034839868545532)),(to_sfixed_a(0.20872275531291962)),(to_sfixed_a(-0.025960320606827736)),(to_sfixed_a(0.0834888368844986)),(to_sfixed_a(0.2725892663002014)),(to_sfixed_a(0.004996501374989748)),(to_sfixed_a(0.050530076026916504)),(to_sfixed_a(6.211355503182858e-05)),(to_sfixed_a(0.0007616515504196286)),(to_sfixed_a(0.0001068413257598877)),(to_sfixed_a(0.00011876572534674779)),(to_sfixed_a(-0.0002335235185455531)),(to_sfixed_a(8.962166612036526e-05)),(to_sfixed_a(-0.0001809345412766561)),(to_sfixed_a(0.0001272465306101367)),(to_sfixed_a(0.00010430852853460237)),(to_sfixed_a(-0.07477691024541855)),(to_sfixed_a(-0.052253853529691696)),(to_sfixed_a(-0.14029905200004578)),(to_sfixed_a(-0.030018962919712067)),(to_sfixed_a(-0.15971457958221436)),(to_sfixed_a(-0.33755922317504883)),(to_sfixed_a(-0.11331360787153244)),(to_sfixed_a(-0.05916731804609299)),(to_sfixed_a(-0.09217320382595062)),(to_sfixed_a(-0.03657850995659828)),(to_sfixed_a(-0.22651077806949615)),(to_sfixed_a(-0.16710759699344635)),(to_sfixed_a(-0.21208080649375916)),(to_sfixed_a(0.13159886002540588)),(to_sfixed_a(0.017182832583785057)),(to_sfixed_a(0.1527140885591507)),(to_sfixed_a(0.05676623061299324)),(to_sfixed_a(0.13405457139015198)),(to_sfixed_a(0.07288393378257751)),(to_sfixed_a(-0.0038857797626405954)),(to_sfixed_a(-0.005267731845378876)),(to_sfixed_a(-0.0014526300365105271)),(to_sfixed_a(-0.0002447694423608482)),(to_sfixed_a(-3.113201091764495e-05)),(to_sfixed_a(-2.7443800718174316e-05)),(to_sfixed_a(7.85297597758472e-05)),(to_sfixed_a(-6.349379691528156e-05)),(to_sfixed_a(-0.0002702803467400372)),(to_sfixed_a(-0.05444428324699402)),(to_sfixed_a(-0.2673787772655487)),(to_sfixed_a(-0.07076428085565567)),(to_sfixed_a(-0.03259846568107605)),(to_sfixed_a(-0.16721998155117035)),(to_sfixed_a(-0.3239089548587799)),(to_sfixed_a(-0.19265899062156677)),(to_sfixed_a(0.09720275551080704)),(to_sfixed_a(0.18668615818023682)),(to_sfixed_a(-0.024596678093075752)),(to_sfixed_a(-0.07764153182506561)),(to_sfixed_a(-0.2739226222038269)),(to_sfixed_a(-0.14670482277870178)),(to_sfixed_a(-0.11895114183425903)),(to_sfixed_a(0.08634635806083679)),(to_sfixed_a(-0.11989489942789078)),(to_sfixed_a(0.02952556498348713)),(to_sfixed_a(-0.5101600289344788)),(to_sfixed_a(-0.10113821178674698)),(to_sfixed_a(-0.1345292627811432)),(to_sfixed_a(-0.004925938788801432)),(to_sfixed_a(0.00019820919260382652)),(to_sfixed_a(1.2170147783763241e-05)),(to_sfixed_a(6.922279862919822e-05)),(to_sfixed_a(-0.00011111618368886411)),(to_sfixed_a(2.3959612008184195e-05)),(to_sfixed_a(-1.0733432645793073e-05)),(to_sfixed_a(0.03397425636649132)),(to_sfixed_a(-0.015090669505298138)),(to_sfixed_a(-0.10382430255413055)),(to_sfixed_a(-0.06641001254320145)),(to_sfixed_a(-0.37105679512023926)),(to_sfixed_a(-0.03198741003870964)),(to_sfixed_a(0.037301745265722275)),(to_sfixed_a(0.11356799304485321)),(to_sfixed_a(0.10845421254634857)),(to_sfixed_a(0.14625906944274902)),(to_sfixed_a(-0.1504909247159958)),(to_sfixed_a(-0.2979778051376343)),(to_sfixed_a(-0.37029972672462463)),(to_sfixed_a(0.015660008415579796)),(to_sfixed_a(0.1321360319852829)),(to_sfixed_a(0.035433996468782425)),(to_sfixed_a(-0.0692228227853775)),(to_sfixed_a(-0.1266755908727646)),(to_sfixed_a(-0.13971014320850372)),(to_sfixed_a(-0.1214340329170227)),(to_sfixed_a(-0.3804381489753723)),(to_sfixed_a(0.015770776197314262)),(to_sfixed_a(9.892298112390563e-05)),(to_sfixed_a(0.0001909415441332385)),(to_sfixed_a(7.431695848936215e-05)),(to_sfixed_a(-0.00010030068369815126)),(to_sfixed_a(2.7256395696895197e-05)),(to_sfixed_a(8.530234481440857e-05)),(to_sfixed_a(8.352585427928716e-05)),(to_sfixed_a(0.061291664838790894)),(to_sfixed_a(-0.04703535512089729)),(to_sfixed_a(0.05060352385044098)),(to_sfixed_a(-0.12531974911689758)),(to_sfixed_a(0.004506988450884819)),(to_sfixed_a(0.13237431645393372)),(to_sfixed_a(0.011523270048201084)),(to_sfixed_a(0.09294319152832031)),(to_sfixed_a(0.17123086750507355)),(to_sfixed_a(-0.20382478833198547)),(to_sfixed_a(-0.03051619790494442)),(to_sfixed_a(-0.04151766002178192)),(to_sfixed_a(0.1258283406496048)),(to_sfixed_a(0.23231661319732666)),(to_sfixed_a(0.08976313471794128)),(to_sfixed_a(-0.10123168677091599)),(to_sfixed_a(-0.12069365382194519)),(to_sfixed_a(-0.07377833873033524)),(to_sfixed_a(-0.20322595536708832)),(to_sfixed_a(0.018582504242658615)),(to_sfixed_a(9.509021765552461e-05)),(to_sfixed_a(1.568802872498054e-05)),(to_sfixed_a(-3.2362149795517325e-05)),(to_sfixed_a(-7.958588685141876e-05)),(to_sfixed_a(0.00011816956975962967)),(to_sfixed_a(-1.8143777197110467e-05)),(to_sfixed_a(-0.00018092499522026628)),(to_sfixed_a(-0.001278283423744142)),(to_sfixed_a(-0.030186230316758156)),(to_sfixed_a(0.11989691108465195)),(to_sfixed_a(0.182334303855896)),(to_sfixed_a(0.23040752112865448)),(to_sfixed_a(0.4012407958507538)),(to_sfixed_a(0.10185208916664124)),(to_sfixed_a(0.10129429399967194)),(to_sfixed_a(0.06962356716394424)),(to_sfixed_a(0.12570816278457642)),(to_sfixed_a(0.16418898105621338)),(to_sfixed_a(-0.04705038666725159)),(to_sfixed_a(0.43526095151901245)),(to_sfixed_a(0.20832796394824982)),(to_sfixed_a(0.30499038100242615)),(to_sfixed_a(0.051985953003168106)),(to_sfixed_a(-0.6469767689704895)),(to_sfixed_a(-0.24911534786224365)),(to_sfixed_a(-0.006619917694479227)),(to_sfixed_a(-0.2602119445800781)),(to_sfixed_a(-0.026386091485619545)),(to_sfixed_a(0.005927866790443659)),(to_sfixed_a(-2.4432629288639873e-05)),(to_sfixed_a(2.7020158086088486e-05)),(to_sfixed_a(-0.000222233182284981)),(to_sfixed_a(-1.846033046604134e-05)),(to_sfixed_a(-6.739650416420773e-05)),(to_sfixed_a(0.017187731340527534)),(to_sfixed_a(0.060086894780397415)),(to_sfixed_a(0.07717692852020264)),(to_sfixed_a(0.1518293172121048)),(to_sfixed_a(-0.03687189146876335)),(to_sfixed_a(-0.11913526803255081)),(to_sfixed_a(0.10293038934469223)),(to_sfixed_a(-0.07097255438566208)),(to_sfixed_a(0.23524440824985504)),(to_sfixed_a(-0.2431449592113495)),(to_sfixed_a(-0.1432860642671585)),(to_sfixed_a(-0.29225024580955505)),(to_sfixed_a(0.1436811238527298)),(to_sfixed_a(0.527442455291748)),(to_sfixed_a(0.38729506731033325)),(to_sfixed_a(0.5521292090415955)),(to_sfixed_a(0.033986303955316544)),(to_sfixed_a(-0.22556430101394653)),(to_sfixed_a(0.0378725491464138)),(to_sfixed_a(-0.21087953448295593)),(to_sfixed_a(-0.09756134450435638)),(to_sfixed_a(-0.007596250623464584)),(to_sfixed_a(0.00013497521285898983)),(to_sfixed_a(-1.4988270777394064e-05)),(to_sfixed_a(0.00015319713565986603)),(to_sfixed_a(-0.00024394792853854597)),(to_sfixed_a(-3.275486596976407e-05)),(to_sfixed_a(-7.084045500960201e-05)),(to_sfixed_a(0.00018649360572453588)),(to_sfixed_a(-0.1566351354122162)),(to_sfixed_a(-0.1450907438993454)),(to_sfixed_a(0.07511389255523682)),(to_sfixed_a(-0.1811651587486267)),(to_sfixed_a(-0.22404736280441284)),(to_sfixed_a(-0.06359156221151352)),(to_sfixed_a(-0.07254922389984131)),(to_sfixed_a(-0.05507969856262207)),(to_sfixed_a(0.2640509009361267)),(to_sfixed_a(-0.20922857522964478)),(to_sfixed_a(-0.09908109903335571)),(to_sfixed_a(0.1393015831708908)),(to_sfixed_a(0.7070276737213135)),(to_sfixed_a(0.39893651008605957)),(to_sfixed_a(0.0524291954934597)),(to_sfixed_a(-0.3158084452152252)),(to_sfixed_a(-0.5584902763366699)),(to_sfixed_a(0.08277702331542969)),(to_sfixed_a(0.007687387987971306)),(to_sfixed_a(-0.15579502284526825)),(to_sfixed_a(-0.05712289735674858)),(to_sfixed_a(4.1041690565180033e-05)),(to_sfixed_a(8.94877957762219e-05)),(to_sfixed_a(-0.00018840926350094378)),(to_sfixed_a(0.00023133723880164325)),(to_sfixed_a(0.00018141961481887847)),(to_sfixed_a(-7.259858102770522e-05)),(to_sfixed_a(-0.0001455843885196373)),(to_sfixed_a(-0.051651597023010254)),(to_sfixed_a(0.10736440122127533)),(to_sfixed_a(0.12237890064716339)),(to_sfixed_a(-0.022655321285128593)),(to_sfixed_a(0.036550331860780716)),(to_sfixed_a(0.16862113773822784)),(to_sfixed_a(0.072484090924263)),(to_sfixed_a(0.03626310080289841)),(to_sfixed_a(0.1530391126871109)),(to_sfixed_a(-0.1023101732134819)),(to_sfixed_a(-0.12289757281541824)),(to_sfixed_a(0.09182725101709366)),(to_sfixed_a(0.28713852167129517)),(to_sfixed_a(-0.01209914032369852)),(to_sfixed_a(-0.10154219716787338)),(to_sfixed_a(-0.789475679397583)),(to_sfixed_a(-0.21206238865852356)),(to_sfixed_a(-0.2144189178943634)),(to_sfixed_a(-0.02316860668361187)),(to_sfixed_a(0.1753126084804535)),(to_sfixed_a(0.017917444929480553)),(to_sfixed_a(-0.002548472722992301)),(to_sfixed_a(-0.0019072226714342833)),(to_sfixed_a(-0.00022839101438876241)),(to_sfixed_a(-0.00023626461916137487)),(to_sfixed_a(-0.00018969253869727254)),(to_sfixed_a(-0.000133760942844674)),(to_sfixed_a(0.0002085952874040231)),(to_sfixed_a(0.0019799857400357723)),(to_sfixed_a(0.19372080266475677)),(to_sfixed_a(0.08021236211061478)),(to_sfixed_a(0.21284419298171997)),(to_sfixed_a(0.22375193238258362)),(to_sfixed_a(0.213922381401062)),(to_sfixed_a(0.13184645771980286)),(to_sfixed_a(0.26211053133010864)),(to_sfixed_a(-0.18952959775924683)),(to_sfixed_a(-0.01383822038769722)),(to_sfixed_a(0.08297622203826904)),(to_sfixed_a(-0.027197223156690598)),(to_sfixed_a(0.08497047424316406)),(to_sfixed_a(-0.009446422569453716)),(to_sfixed_a(-0.13789638876914978)),(to_sfixed_a(-0.657177746295929)),(to_sfixed_a(-0.5202957987785339)),(to_sfixed_a(-0.2506701350212097)),(to_sfixed_a(0.027035661041736603)),(to_sfixed_a(0.1015537828207016)),(to_sfixed_a(0.02074017934501171)),(to_sfixed_a(1.6563509461775539e-06)),(to_sfixed_a(-1.5094194168341346e-05)),(to_sfixed_a(0.0002322903455933556)),(to_sfixed_a(0.00011610231013037264)),(to_sfixed_a(-0.00025885619106702507)),(to_sfixed_a(6.795363151468337e-05)),(to_sfixed_a(-8.590766083216295e-05)),(to_sfixed_a(-0.053687628358602524)),(to_sfixed_a(0.16955877840518951)),(to_sfixed_a(0.05458668991923332)),(to_sfixed_a(0.19758759438991547)),(to_sfixed_a(0.16421669721603394)),(to_sfixed_a(0.21163137257099152)),(to_sfixed_a(0.2992863655090332)),(to_sfixed_a(0.004721911624073982)),(to_sfixed_a(-0.09611328691244125)),(to_sfixed_a(0.20661719143390656)),(to_sfixed_a(0.1575343906879425)),(to_sfixed_a(0.10908378660678864)),(to_sfixed_a(0.013583304360508919)),(to_sfixed_a(-0.11170732975006104)),(to_sfixed_a(-0.41984447836875916)),(to_sfixed_a(-0.3762512505054474)),(to_sfixed_a(-0.37762972712516785)),(to_sfixed_a(-0.1482638567686081)),(to_sfixed_a(-0.21412688493728638)),(to_sfixed_a(0.009562053717672825)),(to_sfixed_a(0.18150605261325836)),(to_sfixed_a(-0.00012773237540386617)),(to_sfixed_a(0.00024342328833881766)),(to_sfixed_a(4.2169413063675165e-06)),(to_sfixed_a(-0.0001549380976939574)),(to_sfixed_a(0.0002074908697977662)),(to_sfixed_a(0.00022746722970623523)),(to_sfixed_a(0.002881500869989395)),(to_sfixed_a(0.11031481623649597)),(to_sfixed_a(0.037923749536275864)),(to_sfixed_a(0.11448956280946732)),(to_sfixed_a(0.3701696991920471)),(to_sfixed_a(0.1773553341627121)),(to_sfixed_a(-0.06431572884321213)),(to_sfixed_a(-0.07296835631132126)),(to_sfixed_a(-0.28256455063819885)),(to_sfixed_a(-0.1282424032688141)),(to_sfixed_a(-0.0922466516494751)),(to_sfixed_a(0.12752175331115723)),(to_sfixed_a(0.15874187648296356)),(to_sfixed_a(-0.050096798688173294)),(to_sfixed_a(-0.11901618540287018)),(to_sfixed_a(-0.5633772015571594)),(to_sfixed_a(-0.10026562213897705)),(to_sfixed_a(-0.25295737385749817)),(to_sfixed_a(0.008331915363669395)),(to_sfixed_a(0.002606438472867012)),(to_sfixed_a(0.11735046654939651)),(to_sfixed_a(0.07010538876056671)),(to_sfixed_a(0.009494717232882977)),(to_sfixed_a(6.440255674533546e-05)),(to_sfixed_a(3.661389200715348e-05)),(to_sfixed_a(-0.0001009968327707611)),(to_sfixed_a(4.748253559228033e-05)),(to_sfixed_a(0.0025994463358074427)),(to_sfixed_a(0.002972498070448637)),(to_sfixed_a(-0.028662998229265213)),(to_sfixed_a(0.14471586048603058)),(to_sfixed_a(0.03487369418144226)),(to_sfixed_a(-0.18592092394828796)),(to_sfixed_a(0.0649469718337059)),(to_sfixed_a(-0.06916488707065582)),(to_sfixed_a(-0.27588871121406555)),(to_sfixed_a(-0.24582451581954956)),(to_sfixed_a(-0.1372670829296112)),(to_sfixed_a(-0.12981151044368744)),(to_sfixed_a(0.17145764827728271)),(to_sfixed_a(-0.09935284405946732)),(to_sfixed_a(-0.42439401149749756)),(to_sfixed_a(-0.26669368147850037)),(to_sfixed_a(-0.18430837988853455)),(to_sfixed_a(-0.020421810448169708)),(to_sfixed_a(-0.09299121797084808)),(to_sfixed_a(0.04491817578673363)),(to_sfixed_a(-0.12193615734577179)),(to_sfixed_a(0.024583106860518456)),(to_sfixed_a(-0.0001388231903547421)),(to_sfixed_a(-2.665934334800113e-05)),(to_sfixed_a(0.0002411511813988909)),(to_sfixed_a(0.00010263417061651126)),(to_sfixed_a(-0.0001905307435663417)),(to_sfixed_a(2.9082035325700417e-05)),(to_sfixed_a(-0.0005587564082816243)),(to_sfixed_a(0.0047693075612187386)),(to_sfixed_a(0.16633237898349762)),(to_sfixed_a(0.24725624918937683)),(to_sfixed_a(-0.010050841607153416)),(to_sfixed_a(-0.16452442109584808)),(to_sfixed_a(-0.15921704471111298)),(to_sfixed_a(-0.006329106632620096)),(to_sfixed_a(-0.06403066962957382)),(to_sfixed_a(-0.250624418258667)),(to_sfixed_a(0.007313376758247614)),(to_sfixed_a(0.16235266625881195)),(to_sfixed_a(0.09878745675086975)),(to_sfixed_a(-0.1987912952899933)),(to_sfixed_a(-0.20087914168834686)),(to_sfixed_a(-0.32777610421180725)),(to_sfixed_a(0.0024010157212615013)),(to_sfixed_a(0.1179766058921814)),(to_sfixed_a(0.05835999175906181)),(to_sfixed_a(0.12998028099536896)),(to_sfixed_a(-0.1421419233083725)),(to_sfixed_a(0.049428317695856094)),(to_sfixed_a(0.011921546421945095)),(to_sfixed_a(0.00017935372306965292)),(to_sfixed_a(0.00019453157437965274)),(to_sfixed_a(1.4591755643778015e-05)),(to_sfixed_a(-4.416634328663349e-05)),(to_sfixed_a(0.0002837352512869984)),(to_sfixed_a(-4.758226714329794e-05)),(to_sfixed_a(-0.0235200934112072)),(to_sfixed_a(-0.0037123742513358593)),(to_sfixed_a(0.10996945947408676)),(to_sfixed_a(0.01680741086602211)),(to_sfixed_a(-0.03605475276708603)),(to_sfixed_a(-0.22377558052539825)),(to_sfixed_a(-0.030158961191773415)),(to_sfixed_a(0.1349818855524063)),(to_sfixed_a(0.0809808224439621)),(to_sfixed_a(-0.03565197065472603)),(to_sfixed_a(0.2356966882944107)),(to_sfixed_a(-0.011494050733745098)),(to_sfixed_a(-0.04321760684251785)),(to_sfixed_a(0.13829761743545532)),(to_sfixed_a(0.05456603318452835)),(to_sfixed_a(0.030021509155631065)),(to_sfixed_a(0.06959749013185501)),(to_sfixed_a(0.09307791292667389)),(to_sfixed_a(0.07333024591207504)),(to_sfixed_a(-0.019332867115736008)),(to_sfixed_a(0.43297430872917175)),(to_sfixed_a(-7.477496637875447e-06)),(to_sfixed_a(4.0304355934495106e-05)),(to_sfixed_a(0.0002262953348690644)),(to_sfixed_a(0.00015720483497716486)),(to_sfixed_a(-0.00010841203038580716)),(to_sfixed_a(-2.7279869755147956e-05)),(to_sfixed_a(-0.0001983141846721992)),(to_sfixed_a(2.561527480793302e-06)),(to_sfixed_a(-0.037559136748313904)),(to_sfixed_a(0.0358072891831398)),(to_sfixed_a(0.15049345791339874)),(to_sfixed_a(-0.19342480599880219)),(to_sfixed_a(-0.20622368156909943)),(to_sfixed_a(-0.013652143068611622)),(to_sfixed_a(-0.00868391152471304)),(to_sfixed_a(0.13465537130832672)),(to_sfixed_a(0.35394445061683655)),(to_sfixed_a(0.07444439083337784)),(to_sfixed_a(0.08262985944747925)),(to_sfixed_a(0.06527497619390488)),(to_sfixed_a(0.12170694023370743)),(to_sfixed_a(-0.05474585294723511)),(to_sfixed_a(0.2393776923418045)),(to_sfixed_a(0.3448875844478607)),(to_sfixed_a(0.26697802543640137)),(to_sfixed_a(0.07619775831699371)),(to_sfixed_a(0.2447553426027298)),(to_sfixed_a(0.2699684798717499)),(to_sfixed_a(0.06969040632247925)),(to_sfixed_a(-0.00013175445201341063)),(to_sfixed_a(-0.00015524166519753635)),(to_sfixed_a(8.417361823376268e-05)),(to_sfixed_a(0.00020344437507446855)),(to_sfixed_a(4.288614491088083e-06)),(to_sfixed_a(-6.566870433744043e-05)),(to_sfixed_a(4.492964581004344e-05)),(to_sfixed_a(-0.021624261513352394)),(to_sfixed_a(-0.0004004981310572475)),(to_sfixed_a(-0.007617947179824114)),(to_sfixed_a(-0.18342648446559906)),(to_sfixed_a(-0.05492814630270004)),(to_sfixed_a(-0.04269302263855934)),(to_sfixed_a(0.0360836423933506)),(to_sfixed_a(-0.033643126487731934)),(to_sfixed_a(0.031157556921243668)),(to_sfixed_a(0.1555243879556656)),(to_sfixed_a(-0.09451412409543991)),(to_sfixed_a(0.10579542070627213)),(to_sfixed_a(0.05800137668848038)),(to_sfixed_a(0.26031070947647095)),(to_sfixed_a(0.28947949409484863)),(to_sfixed_a(0.10007523000240326)),(to_sfixed_a(0.568105936050415)),(to_sfixed_a(0.11206721514463425)),(to_sfixed_a(0.18370620906352997)),(to_sfixed_a(0.0009678289643488824)),(to_sfixed_a(-0.006699030753225088)),(to_sfixed_a(-2.6249492293572985e-05)),(to_sfixed_a(-0.00017830207070801407)),(to_sfixed_a(0.00019068922847509384)),(to_sfixed_a(-9.591333218850195e-05)),(to_sfixed_a(0.0001396796724293381)),(to_sfixed_a(0.00021421696874313056)),(to_sfixed_a(-0.00010119482612935826)),(to_sfixed_a(-4.653067207982531e-06)),(to_sfixed_a(0.12855972349643707)),(to_sfixed_a(0.012305008247494698)),(to_sfixed_a(-0.05280124023556709)),(to_sfixed_a(-0.0487922802567482)),(to_sfixed_a(0.01154358685016632)),(to_sfixed_a(-0.16348634660243988)),(to_sfixed_a(-0.04768873751163483)),(to_sfixed_a(-0.09955019503831863)),(to_sfixed_a(-0.00048226318904198706)),(to_sfixed_a(-0.08328429609537125)),(to_sfixed_a(-0.048692844808101654)),(to_sfixed_a(-0.143588587641716)),(to_sfixed_a(0.18481498956680298)),(to_sfixed_a(0.23546558618545532)),(to_sfixed_a(0.022008761763572693)),(to_sfixed_a(-0.011276421137154102)),(to_sfixed_a(0.012609708122909069)),(to_sfixed_a(-0.017232133075594902)),(to_sfixed_a(-0.009598709642887115)),(to_sfixed_a(6.37771881883964e-05)),(to_sfixed_a(0.0001030671555781737)),(to_sfixed_a(-8.458834054181352e-05)),(to_sfixed_a(-3.0253790100687183e-05)),(to_sfixed_a(0.00016400442109443247)),(to_sfixed_a(-0.0002379479119554162)),(to_sfixed_a(-5.547336331801489e-05)),(to_sfixed_a(-1.5289613656932488e-05)),(to_sfixed_a(1.1715907021425664e-05)),(to_sfixed_a(0.003789349226281047)),(to_sfixed_a(-0.04281904920935631)),(to_sfixed_a(0.04885931313037872)),(to_sfixed_a(-0.1323145627975464)),(to_sfixed_a(0.08002283424139023)),(to_sfixed_a(-0.019732395187020302)),(to_sfixed_a(-0.1717015504837036)),(to_sfixed_a(-0.19159989058971405)),(to_sfixed_a(-0.054156966507434845)),(to_sfixed_a(0.01813851296901703)),(to_sfixed_a(-0.041704997420310974)),(to_sfixed_a(0.048678409308195114)),(to_sfixed_a(-0.059138767421245575)),(to_sfixed_a(0.09508362412452698)),(to_sfixed_a(0.07044059038162231)),(to_sfixed_a(-0.06638342887163162)),(to_sfixed_a(-0.020341923460364342)),(to_sfixed_a(-0.01782444305717945)),(to_sfixed_a(-0.009623712860047817)),(to_sfixed_a(0.00018850626656785607)),(to_sfixed_a(-8.417100616497919e-05)),(to_sfixed_a(-1.7595883036847226e-05)),(to_sfixed_a(-3.317181835882366e-05)),(to_sfixed_a(-8.588621858507395e-05)),(to_sfixed_a(0.00011115975212305784)),(to_sfixed_a(0.000175905748619698)),(to_sfixed_a(4.268202246748842e-05)),(to_sfixed_a(-0.03381986916065216)),(to_sfixed_a(-0.006847281474620104)),(to_sfixed_a(-0.14218223094940186)),(to_sfixed_a(-0.27254918217658997)),(to_sfixed_a(-0.12444262206554413)),(to_sfixed_a(-0.012036656960844994)),(to_sfixed_a(-0.17547354102134705)),(to_sfixed_a(-0.012872970663011074)),(to_sfixed_a(-0.2836179733276367)),(to_sfixed_a(-0.3015495240688324)),(to_sfixed_a(-0.10444275289773941)),(to_sfixed_a(0.03499210998415947)),(to_sfixed_a(0.1613401472568512)),(to_sfixed_a(0.08330332487821579)),(to_sfixed_a(0.04400763288140297)),(to_sfixed_a(0.02170022390782833)),(to_sfixed_a(0.01055844221264124)),(to_sfixed_a(0.0019433830166235566)),(to_sfixed_a(-0.005059629678726196)),(to_sfixed_a(-0.007702550385147333)),(to_sfixed_a(-7.242120045702904e-05)),(to_sfixed_a(-0.0001030739804264158)),(to_sfixed_a(0.00014628730423282832)),(to_sfixed_a(-0.0002669066598173231)),(to_sfixed_a(0.00013285037130117416)),(to_sfixed_a(-1.3504664821084589e-05)),(to_sfixed_a(-0.00032281968742609024)),(to_sfixed_a(-4.929819169774419e-06)),(to_sfixed_a(1.228260543939541e-06)),(to_sfixed_a(0.004090879578143358)),(to_sfixed_a(-0.08526909351348877)),(to_sfixed_a(-0.11335878074169159)),(to_sfixed_a(-0.2432858794927597)),(to_sfixed_a(-0.13597925007343292)),(to_sfixed_a(-0.17031821608543396)),(to_sfixed_a(0.04627181589603424)),(to_sfixed_a(-0.06766273081302643)),(to_sfixed_a(-0.2601335346698761)),(to_sfixed_a(-0.1058860719203949)),(to_sfixed_a(-0.06440457701683044)),(to_sfixed_a(0.18861277401447296)),(to_sfixed_a(-0.0349624902009964)),(to_sfixed_a(-0.00722148222848773)),(to_sfixed_a(0.054481390863657)),(to_sfixed_a(0.09085678309202194)),(to_sfixed_a(8.129000343615189e-05)),(to_sfixed_a(-0.0029789460822939873)),(to_sfixed_a(-0.003824302228167653)),(to_sfixed_a(0.00013541730004362762)),(to_sfixed_a(0.00014278660819400102)),(to_sfixed_a(2.553419108153321e-05)),(to_sfixed_a(8.740847988519818e-05)),(to_sfixed_a(-7.446168456226587e-05)),(to_sfixed_a(-0.00012660025095101446)),(to_sfixed_a(8.533748768968508e-05)),(to_sfixed_a(0.00019009463721886277)),(to_sfixed_a(-0.00012827319733332843)),(to_sfixed_a(0.001898718299344182)),(to_sfixed_a(0.0017261991742998362)),(to_sfixed_a(3.972681224695407e-05)),(to_sfixed_a(0.00013889378169551492)),(to_sfixed_a(0.00041975677595473826)),(to_sfixed_a(0.07754429429769516)),(to_sfixed_a(-0.0007722733425907791)),(to_sfixed_a(-0.0018944048788398504)),(to_sfixed_a(0.05489601939916611)),(to_sfixed_a(-0.13776490092277527)),(to_sfixed_a(-0.012195540592074394)),(to_sfixed_a(0.0015262877568602562)),(to_sfixed_a(0.06469884514808655)),(to_sfixed_a(0.086422398686409)),(to_sfixed_a(0.003243133658543229)),(to_sfixed_a(0.0036429029423743486)),(to_sfixed_a(-8.50625383463921e-06)),(to_sfixed_a(-5.467768005473772e-06)),(to_sfixed_a(-7.068587729008868e-05)),(to_sfixed_a(-0.0004120173689443618)),(to_sfixed_a(-0.00012120231986045837)),(to_sfixed_a(3.50458976754453e-05)),(to_sfixed_a(0.00023414882889483124)),(to_sfixed_a(0.00010834060230990872)),(to_sfixed_a(-7.809055387042463e-05)),(to_sfixed_a(0.00025753575027920306)),(to_sfixed_a(0.00019606665591709316)),(to_sfixed_a(8.097020327113569e-05)),(to_sfixed_a(-4.338413418736309e-05)),(to_sfixed_a(0.00028450574609450996)),(to_sfixed_a(0.0002197681023972109)),(to_sfixed_a(-0.00021433350048027933)),(to_sfixed_a(7.405199994536815e-06)),(to_sfixed_a(8.332319703185931e-05)),(to_sfixed_a(4.470067142392509e-05)),(to_sfixed_a(-0.00013864597713109106)),(to_sfixed_a(3.698213185998611e-05)),(to_sfixed_a(7.311886292882264e-05)),(to_sfixed_a(3.561324774636887e-05)),(to_sfixed_a(5.551857248065062e-05)),(to_sfixed_a(-0.00012213800800964236)),(to_sfixed_a(0.00016186069115065038)),(to_sfixed_a(-0.000140848831506446)),(to_sfixed_a(-4.127131978748366e-05)),(to_sfixed_a(-7.16609283699654e-05)),(to_sfixed_a(0.00021502291201613843)),(to_sfixed_a(3.13831719722657e-06)),(to_sfixed_a(-7.061255746521056e-05)),(to_sfixed_a(-4.637422080122633e-06)),(to_sfixed_a(-0.00023513822816312313)),(to_sfixed_a(-0.00020649937505368143)));

    constant weight_n0_13 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(0.00010981001105392352)),(to_sfixed_a(-0.00014526004088111222)),(to_sfixed_a(-9.642725444791722e-07)),(to_sfixed_a(1.5247676856233738e-05)),(to_sfixed_a(0.00035046739503741264)),(to_sfixed_a(0.0002513656218070537)),(to_sfixed_a(-0.00013220912660472095)),(to_sfixed_a(0.0001857506576925516)),(to_sfixed_a(-0.00010156175267184153)),(to_sfixed_a(0.000237374086282216)),(to_sfixed_a(9.418415720574558e-05)),(to_sfixed_a(0.00016205591964535415)),(to_sfixed_a(0.00013814817066304386)),(to_sfixed_a(5.557193799177185e-05)),(to_sfixed_a(1.7338797988486476e-05)),(to_sfixed_a(2.2570928194909357e-05)),(to_sfixed_a(3.774967262870632e-05)),(to_sfixed_a(2.3870838958828244e-06)),(to_sfixed_a(-7.570019806735218e-05)),(to_sfixed_a(0.00020882616809103638)),(to_sfixed_a(-3.604055746109225e-05)),(to_sfixed_a(-9.85189326456748e-05)),(to_sfixed_a(-0.00016329440404661)),(to_sfixed_a(6.245248368941247e-05)),(to_sfixed_a(7.772774551995099e-05)),(to_sfixed_a(-8.54355821502395e-05)),(to_sfixed_a(-0.00022160577645990998)),(to_sfixed_a(0.00016052454884629697)),(to_sfixed_a(-7.258350524352863e-05)),(to_sfixed_a(-9.399525151820853e-05)),(to_sfixed_a(1.8243574231746607e-05)),(to_sfixed_a(-7.098763308022171e-05)),(to_sfixed_a(6.770032632630318e-05)),(to_sfixed_a(7.71780323702842e-05)),(to_sfixed_a(0.0003165476373396814)),(to_sfixed_a(0.0001546815619803965)),(to_sfixed_a(-8.884403359843418e-05)),(to_sfixed_a(-4.479144990909845e-06)),(to_sfixed_a(-0.0001929731370182708)),(to_sfixed_a(-0.00015980425814632326)),(to_sfixed_a(-8.617796265752986e-05)),(to_sfixed_a(-7.476921746274456e-05)),(to_sfixed_a(-0.0001428890391252935)),(to_sfixed_a(-5.588281783275306e-05)),(to_sfixed_a(-0.00025099844788201153)),(to_sfixed_a(1.495189826528076e-05)),(to_sfixed_a(-1.291499847866362e-05)),(to_sfixed_a(4.3416497646830976e-05)),(to_sfixed_a(-0.0003341663395985961)),(to_sfixed_a(2.8147331249783747e-05)),(to_sfixed_a(0.00012414288357831538)),(to_sfixed_a(-7.270877540577203e-05)),(to_sfixed_a(0.0002725869126152247)),(to_sfixed_a(-1.5592375348205678e-05)),(to_sfixed_a(9.182640496874228e-05)),(to_sfixed_a(-4.4654341763816774e-05)),(to_sfixed_a(5.404587500379421e-05)),(to_sfixed_a(-4.2647043301258236e-05)),(to_sfixed_a(0.0002110775385517627)),(to_sfixed_a(-0.00018150679534301162)),(to_sfixed_a(8.20888380985707e-05)),(to_sfixed_a(-0.00032178458059206605)),(to_sfixed_a(7.780483429087326e-05)),(to_sfixed_a(0.00033865985460579395)),(to_sfixed_a(0.00016014106222428381)),(to_sfixed_a(0.00036519611603580415)),(to_sfixed_a(-7.516928599216044e-05)),(to_sfixed_a(-3.6661960621131584e-05)),(to_sfixed_a(-0.0001441578206140548)),(to_sfixed_a(0.00029747403459623456)),(to_sfixed_a(2.5498142349533737e-05)),(to_sfixed_a(-3.334037319291383e-05)),(to_sfixed_a(0.00011138319678138942)),(to_sfixed_a(-3.771771662286483e-05)),(to_sfixed_a(1.1826025001937523e-05)),(to_sfixed_a(0.00014630235091317445)),(to_sfixed_a(-0.00013833257253281772)),(to_sfixed_a(-5.045552097726613e-05)),(to_sfixed_a(0.00021341822866816074)),(to_sfixed_a(-0.00017362374637741596)),(to_sfixed_a(0.00018446148897055537)),(to_sfixed_a(3.731166725629009e-05)),(to_sfixed_a(6.199935887707397e-05)),(to_sfixed_a(0.00012825783051084727)),(to_sfixed_a(9.78193711489439e-05)),(to_sfixed_a(-0.00011940578406210989)),(to_sfixed_a(-2.8686108635156415e-06)),(to_sfixed_a(0.00024563600891269743)),(to_sfixed_a(7.252940849866718e-05)),(to_sfixed_a(0.0002216446737293154)),(to_sfixed_a(5.79608058615122e-05)),(to_sfixed_a(-0.00012453181261662394)),(to_sfixed_a(0.020230691879987717)),(to_sfixed_a(-0.00017786752141546458)),(to_sfixed_a(0.0229190681129694)),(to_sfixed_a(-0.04499530419707298)),(to_sfixed_a(-0.0899813175201416)),(to_sfixed_a(-0.31209734082221985)),(to_sfixed_a(0.04838506132364273)),(to_sfixed_a(0.06454475969076157)),(to_sfixed_a(0.003210717812180519)),(to_sfixed_a(0.002948295557871461)),(to_sfixed_a(0.08588619530200958)),(to_sfixed_a(0.1548806130886078)),(to_sfixed_a(0.08522292971611023)),(to_sfixed_a(0.17281918227672577)),(to_sfixed_a(2.836003841366619e-05)),(to_sfixed_a(-0.0001786989305401221)),(to_sfixed_a(-0.00012944739137310535)),(to_sfixed_a(0.0003132927231490612)),(to_sfixed_a(-3.2878484489629045e-05)),(to_sfixed_a(0.00010120169463334605)),(to_sfixed_a(-5.8242287195753306e-05)),(to_sfixed_a(-0.0001035617824527435)),(to_sfixed_a(-0.00017886624846141785)),(to_sfixed_a(-8.851019811118022e-05)),(to_sfixed_a(-9.113962732953951e-05)),(to_sfixed_a(-5.476131627801806e-05)),(to_sfixed_a(-0.0009118674206547439)),(to_sfixed_a(-0.01529041025787592)),(to_sfixed_a(-0.11397378891706467)),(to_sfixed_a(0.025368204340338707)),(to_sfixed_a(-0.4035642445087433)),(to_sfixed_a(-0.1194004938006401)),(to_sfixed_a(-0.3816867470741272)),(to_sfixed_a(-0.2611847519874573)),(to_sfixed_a(-0.006550045683979988)),(to_sfixed_a(-0.05254373699426651)),(to_sfixed_a(-0.14042632281780243)),(to_sfixed_a(-0.22665190696716309)),(to_sfixed_a(-0.01822352036833763)),(to_sfixed_a(0.06205083057284355)),(to_sfixed_a(-0.006250882986932993)),(to_sfixed_a(-0.021420162171125412)),(to_sfixed_a(0.031061885878443718)),(to_sfixed_a(0.0001351906976196915)),(to_sfixed_a(-0.0029434040188789368)),(to_sfixed_a(-1.8269422071170993e-05)),(to_sfixed_a(0.00031344956369139254)),(to_sfixed_a(1.5987228835001588e-05)),(to_sfixed_a(-0.00017488165758550167)),(to_sfixed_a(-8.982345025287941e-05)),(to_sfixed_a(6.91748209646903e-05)),(to_sfixed_a(5.0050362915499136e-05)),(to_sfixed_a(0.0010875168954953551)),(to_sfixed_a(-0.02590855583548546)),(to_sfixed_a(-0.005601902492344379)),(to_sfixed_a(-0.06902816891670227)),(to_sfixed_a(-0.032942935824394226)),(to_sfixed_a(-0.05506670102477074)),(to_sfixed_a(-0.0007818284211680293)),(to_sfixed_a(-0.06145956739783287)),(to_sfixed_a(-0.3883011043071747)),(to_sfixed_a(-0.3903485834598541)),(to_sfixed_a(-0.21061749756336212)),(to_sfixed_a(-0.3336053788661957)),(to_sfixed_a(-0.45574951171875)),(to_sfixed_a(-0.32226672768592834)),(to_sfixed_a(-0.14706049859523773)),(to_sfixed_a(-0.17316918075084686)),(to_sfixed_a(0.0164189413189888)),(to_sfixed_a(0.016234133392572403)),(to_sfixed_a(-0.005020593758672476)),(to_sfixed_a(0.1378908008337021)),(to_sfixed_a(-0.0042116679251194)),(to_sfixed_a(-8.460052049485967e-05)),(to_sfixed_a(0.00014592622756026685)),(to_sfixed_a(-0.00010374465637141839)),(to_sfixed_a(6.56507836538367e-05)),(to_sfixed_a(-0.00020575083908624947)),(to_sfixed_a(0.00026796883321367204)),(to_sfixed_a(6.57660566503182e-05)),(to_sfixed_a(0.00010579218360362574)),(to_sfixed_a(-0.02429901249706745)),(to_sfixed_a(-0.032346561551094055)),(to_sfixed_a(-0.20457452535629272)),(to_sfixed_a(-0.0833168625831604)),(to_sfixed_a(-0.11724884808063507)),(to_sfixed_a(-0.13642112910747528)),(to_sfixed_a(-0.10651054978370667)),(to_sfixed_a(0.08201070874929428)),(to_sfixed_a(0.08631078153848648)),(to_sfixed_a(-0.07578905671834946)),(to_sfixed_a(-0.2727143466472626)),(to_sfixed_a(-0.21438558399677277)),(to_sfixed_a(-0.10479845851659775)),(to_sfixed_a(0.11179054528474808)),(to_sfixed_a(0.02362757734954357)),(to_sfixed_a(0.28602975606918335)),(to_sfixed_a(0.016908753663301468)),(to_sfixed_a(-0.17036600410938263)),(to_sfixed_a(-0.1162588894367218)),(to_sfixed_a(-0.001312532927840948)),(to_sfixed_a(-0.0015270625008270144)),(to_sfixed_a(0.00040382632869295776)),(to_sfixed_a(-0.0002177059359382838)),(to_sfixed_a(3.242299135308713e-05)),(to_sfixed_a(2.506722739781253e-05)),(to_sfixed_a(9.223917004419491e-05)),(to_sfixed_a(9.030261571751907e-05)),(to_sfixed_a(0.00035025691613554955)),(to_sfixed_a(-0.041991233825683594)),(to_sfixed_a(-0.09226153790950775)),(to_sfixed_a(0.07071477174758911)),(to_sfixed_a(0.020688682794570923)),(to_sfixed_a(0.18738791346549988)),(to_sfixed_a(0.08867904543876648)),(to_sfixed_a(0.25885066390037537)),(to_sfixed_a(0.4075358808040619)),(to_sfixed_a(0.4721601605415344)),(to_sfixed_a(0.44801315665245056)),(to_sfixed_a(0.30860772728919983)),(to_sfixed_a(-0.08771812915802002)),(to_sfixed_a(0.40580466389656067)),(to_sfixed_a(-0.10096777975559235)),(to_sfixed_a(-0.17959746718406677)),(to_sfixed_a(-0.020435508340597153)),(to_sfixed_a(0.02779231406748295)),(to_sfixed_a(-0.10680592805147171)),(to_sfixed_a(-0.07147761434316635)),(to_sfixed_a(-0.037469640374183655)),(to_sfixed_a(0.001335764303803444)),(to_sfixed_a(2.1456323793245247e-06)),(to_sfixed_a(2.4422573915217072e-05)),(to_sfixed_a(-5.572912414208986e-05)),(to_sfixed_a(-2.4742896130192094e-05)),(to_sfixed_a(0.0001459425111534074)),(to_sfixed_a(8.506136509822682e-05)),(to_sfixed_a(-0.10551673173904419)),(to_sfixed_a(-0.013175195083022118)),(to_sfixed_a(-0.0033144375775009394)),(to_sfixed_a(-0.1410442292690277)),(to_sfixed_a(0.04267742484807968)),(to_sfixed_a(0.133978471159935)),(to_sfixed_a(0.3373267948627472)),(to_sfixed_a(0.16400104761123657)),(to_sfixed_a(0.2851608991622925)),(to_sfixed_a(0.17075246572494507)),(to_sfixed_a(0.07352933287620544)),(to_sfixed_a(-0.18699504435062408)),(to_sfixed_a(-0.08474733680486679)),(to_sfixed_a(-0.07951144129037857)),(to_sfixed_a(0.1670410931110382)),(to_sfixed_a(-0.08635750412940979)),(to_sfixed_a(-0.08136630058288574)),(to_sfixed_a(-0.17105627059936523)),(to_sfixed_a(-0.1627349704504013)),(to_sfixed_a(0.0813194140791893)),(to_sfixed_a(-0.10542932897806168)),(to_sfixed_a(-0.0005142667796462774)),(to_sfixed_a(-4.9613263399805874e-05)),(to_sfixed_a(-7.512589945690706e-05)),(to_sfixed_a(4.77546636830084e-05)),(to_sfixed_a(6.652584852417931e-05)),(to_sfixed_a(0.0003095594875048846)),(to_sfixed_a(0.0003840607241727412)),(to_sfixed_a(0.0017696238355711102)),(to_sfixed_a(-0.09912802278995514)),(to_sfixed_a(0.009800754487514496)),(to_sfixed_a(0.0010583442635834217)),(to_sfixed_a(-0.04973462596535683)),(to_sfixed_a(-0.018057994544506073)),(to_sfixed_a(0.08554212003946304)),(to_sfixed_a(0.017544133588671684)),(to_sfixed_a(0.024601684883236885)),(to_sfixed_a(0.19791097939014435)),(to_sfixed_a(0.15325818955898285)),(to_sfixed_a(-0.0023288812953978777)),(to_sfixed_a(0.145269975066185)),(to_sfixed_a(0.16585402190685272)),(to_sfixed_a(0.01242161262780428)),(to_sfixed_a(-0.31548115611076355)),(to_sfixed_a(-0.5252559185028076)),(to_sfixed_a(-0.41631069779396057)),(to_sfixed_a(-0.24218185245990753)),(to_sfixed_a(-0.3067370355129242)),(to_sfixed_a(0.11860689520835876)),(to_sfixed_a(-4.575940693030134e-06)),(to_sfixed_a(-0.00013651198241859674)),(to_sfixed_a(4.724238533526659e-05)),(to_sfixed_a(-0.00017066480359062552)),(to_sfixed_a(0.00012398532999213785)),(to_sfixed_a(-9.188399417325854e-05)),(to_sfixed_a(7.514832395827398e-05)),(to_sfixed_a(0.006864119786769152)),(to_sfixed_a(-0.06922049820423126)),(to_sfixed_a(-0.29473191499710083)),(to_sfixed_a(-0.013406302779912949)),(to_sfixed_a(0.02455344796180725)),(to_sfixed_a(0.11829380691051483)),(to_sfixed_a(-0.2347237765789032)),(to_sfixed_a(-0.3527205288410187)),(to_sfixed_a(-0.185048907995224)),(to_sfixed_a(0.029806066304445267)),(to_sfixed_a(-0.16730089485645294)),(to_sfixed_a(0.16179701685905457)),(to_sfixed_a(0.27591583132743835)),(to_sfixed_a(0.2336728423833847)),(to_sfixed_a(0.17066706717014313)),(to_sfixed_a(-0.056880883872509)),(to_sfixed_a(-0.37318727374076843)),(to_sfixed_a(-0.2969059944152832)),(to_sfixed_a(-0.17210276424884796)),(to_sfixed_a(-0.34761783480644226)),(to_sfixed_a(0.013255364261567593)),(to_sfixed_a(0.03912122920155525)),(to_sfixed_a(-8.416779019171372e-05)),(to_sfixed_a(-0.0001963570830412209)),(to_sfixed_a(0.00013766103074885905)),(to_sfixed_a(-0.00013951578876003623)),(to_sfixed_a(5.080747723695822e-05)),(to_sfixed_a(0.014695003628730774)),(to_sfixed_a(-0.2749618589878082)),(to_sfixed_a(-0.1101301833987236)),(to_sfixed_a(-0.029484452679753304)),(to_sfixed_a(-0.011263531632721424)),(to_sfixed_a(-0.1316508799791336)),(to_sfixed_a(-0.029910339042544365)),(to_sfixed_a(-0.0351988784968853)),(to_sfixed_a(0.030119415372610092)),(to_sfixed_a(0.02190285362303257)),(to_sfixed_a(-0.142916738986969)),(to_sfixed_a(-0.12253646552562714)),(to_sfixed_a(-0.10701465606689453)),(to_sfixed_a(0.1408800482749939)),(to_sfixed_a(0.23252953588962555)),(to_sfixed_a(0.35255536437034607)),(to_sfixed_a(0.16836610436439514)),(to_sfixed_a(0.046041954308748245)),(to_sfixed_a(-0.05823912471532822)),(to_sfixed_a(-0.014545424841344357)),(to_sfixed_a(-0.24843209981918335)),(to_sfixed_a(-0.1938142478466034)),(to_sfixed_a(5.146882540429942e-05)),(to_sfixed_a(-4.488430204219185e-05)),(to_sfixed_a(-5.810368384118192e-05)),(to_sfixed_a(-2.2938187612453476e-05)),(to_sfixed_a(6.597866740776226e-05)),(to_sfixed_a(7.03134064679034e-05)),(to_sfixed_a(-0.00019448247621767223)),(to_sfixed_a(-0.04731472581624985)),(to_sfixed_a(0.10775434225797653)),(to_sfixed_a(0.07077918201684952)),(to_sfixed_a(0.11940724402666092)),(to_sfixed_a(0.06651473790407181)),(to_sfixed_a(0.29101860523223877)),(to_sfixed_a(0.17868323624134064)),(to_sfixed_a(0.1405511200428009)),(to_sfixed_a(0.009396367706358433)),(to_sfixed_a(-0.11443426460027695)),(to_sfixed_a(-0.1059880182147026)),(to_sfixed_a(0.17462565004825592)),(to_sfixed_a(0.08896743506193161)),(to_sfixed_a(0.22413323819637299)),(to_sfixed_a(0.16673678159713745)),(to_sfixed_a(-0.0351913757622242)),(to_sfixed_a(0.383561372756958)),(to_sfixed_a(0.1608491986989975)),(to_sfixed_a(0.08634933084249496)),(to_sfixed_a(-0.09701098501682281)),(to_sfixed_a(0.053874410688877106)),(to_sfixed_a(-3.2609452318865806e-05)),(to_sfixed_a(-0.00029923373949714005)),(to_sfixed_a(7.582998659927398e-05)),(to_sfixed_a(1.2196566956390598e-07)),(to_sfixed_a(7.81372727942653e-05)),(to_sfixed_a(2.0667956050601788e-05)),(to_sfixed_a(-3.205037864972837e-05)),(to_sfixed_a(0.041012030094861984)),(to_sfixed_a(0.20482565462589264)),(to_sfixed_a(0.1856841742992401)),(to_sfixed_a(0.2661416232585907)),(to_sfixed_a(0.18237783014774323)),(to_sfixed_a(0.25591495633125305)),(to_sfixed_a(0.29471006989479065)),(to_sfixed_a(-0.14561370015144348)),(to_sfixed_a(-0.13775159418582916)),(to_sfixed_a(-0.2996481955051422)),(to_sfixed_a(-0.23512230813503265)),(to_sfixed_a(-0.010650728829205036)),(to_sfixed_a(0.046842243522405624)),(to_sfixed_a(-0.0051643275655806065)),(to_sfixed_a(-0.047594666481018066)),(to_sfixed_a(-0.2846390902996063)),(to_sfixed_a(-0.11734570562839508)),(to_sfixed_a(-0.12140470743179321)),(to_sfixed_a(0.12881426513195038)),(to_sfixed_a(0.23925523459911346)),(to_sfixed_a(0.024858349934220314)),(to_sfixed_a(0.0008158429991453886)),(to_sfixed_a(-0.0008143715094774961)),(to_sfixed_a(0.0002818356442730874)),(to_sfixed_a(-0.00016305602912325412)),(to_sfixed_a(1.2968312148586847e-05)),(to_sfixed_a(0.00015613794676028192)),(to_sfixed_a(-4.555491977953352e-05)),(to_sfixed_a(-0.00037014903500676155)),(to_sfixed_a(0.08535739779472351)),(to_sfixed_a(0.055333275347948074)),(to_sfixed_a(0.34172314405441284)),(to_sfixed_a(0.19842053949832916)),(to_sfixed_a(0.31881582736968994)),(to_sfixed_a(-0.14772379398345947)),(to_sfixed_a(-0.04349089413881302)),(to_sfixed_a(-0.05059678107500076)),(to_sfixed_a(-0.18458330631256104)),(to_sfixed_a(-0.19436892867088318)),(to_sfixed_a(-0.007802285254001617)),(to_sfixed_a(-0.1093001589179039)),(to_sfixed_a(-0.020607493817806244)),(to_sfixed_a(0.17810586094856262)),(to_sfixed_a(0.25513601303100586)),(to_sfixed_a(0.09079939126968384)),(to_sfixed_a(-0.03630946949124336)),(to_sfixed_a(0.009755539707839489)),(to_sfixed_a(0.13989366590976715)),(to_sfixed_a(-0.00893572997301817)),(to_sfixed_a(-0.00027013837825506926)),(to_sfixed_a(-0.00031079858308658004)),(to_sfixed_a(-0.00020667604985646904)),(to_sfixed_a(0.00017280572501476854)),(to_sfixed_a(-4.9299735110253096e-05)),(to_sfixed_a(0.00022544401872437447)),(to_sfixed_a(0.00013776290870737284)),(to_sfixed_a(0.027808988466858864)),(to_sfixed_a(0.1191827803850174)),(to_sfixed_a(-0.08625125885009766)),(to_sfixed_a(-0.03136901557445526)),(to_sfixed_a(-0.1145220473408699)),(to_sfixed_a(-0.20065303146839142)),(to_sfixed_a(-0.14358700811862946)),(to_sfixed_a(0.10019712895154953)),(to_sfixed_a(0.13876225054264069)),(to_sfixed_a(-0.06128022074699402)),(to_sfixed_a(-0.2676742672920227)),(to_sfixed_a(-0.15846113860607147)),(to_sfixed_a(-0.06504103541374207)),(to_sfixed_a(0.060165368020534515)),(to_sfixed_a(0.14946861565113068)),(to_sfixed_a(0.04193159192800522)),(to_sfixed_a(-0.06443025916814804)),(to_sfixed_a(0.027974793687462807)),(to_sfixed_a(0.32735469937324524)),(to_sfixed_a(0.03433787450194359)),(to_sfixed_a(0.07635772228240967)),(to_sfixed_a(-0.0001836608280427754)),(to_sfixed_a(2.4525183107471094e-05)),(to_sfixed_a(0.00024640237097628415)),(to_sfixed_a(-0.00019052348216064274)),(to_sfixed_a(3.4385971957817674e-05)),(to_sfixed_a(-0.00010145348642254248)),(to_sfixed_a(0.0006026943447068334)),(to_sfixed_a(-0.11668378859758377)),(to_sfixed_a(-0.23956821858882904)),(to_sfixed_a(-0.2603486478328705)),(to_sfixed_a(-0.2742360234260559)),(to_sfixed_a(-0.36219513416290283)),(to_sfixed_a(-0.18307004868984222)),(to_sfixed_a(0.01537819392979145)),(to_sfixed_a(0.7253554463386536)),(to_sfixed_a(-0.08262258023023605)),(to_sfixed_a(-0.0666065514087677)),(to_sfixed_a(-0.33992621302604675)),(to_sfixed_a(-0.10976538062095642)),(to_sfixed_a(-0.3344217538833618)),(to_sfixed_a(0.06581218540668488)),(to_sfixed_a(-0.14132727682590485)),(to_sfixed_a(-0.06776811927556992)),(to_sfixed_a(-0.042656898498535156)),(to_sfixed_a(-0.3364357352256775)),(to_sfixed_a(-0.09488420933485031)),(to_sfixed_a(0.07638061791658401)),(to_sfixed_a(0.07818716764450073)),(to_sfixed_a(-0.00920148566365242)),(to_sfixed_a(0.00047475151950493455)),(to_sfixed_a(-0.00014994227967690676)),(to_sfixed_a(7.602777623105794e-05)),(to_sfixed_a(0.000365199928637594)),(to_sfixed_a(0.0009787364397197962)),(to_sfixed_a(0.0008660160819999874)),(to_sfixed_a(-0.05393523722887039)),(to_sfixed_a(-0.2010486125946045)),(to_sfixed_a(0.009768219664692879)),(to_sfixed_a(-0.19910630583763123)),(to_sfixed_a(-0.3986077308654785)),(to_sfixed_a(-0.0157451294362545)),(to_sfixed_a(0.6549059152603149)),(to_sfixed_a(0.4266999661922455)),(to_sfixed_a(-0.06994543969631195)),(to_sfixed_a(-0.2668473422527313)),(to_sfixed_a(-0.3219478130340576)),(to_sfixed_a(-0.1804269254207611)),(to_sfixed_a(0.011395403183996677)),(to_sfixed_a(0.012945527210831642)),(to_sfixed_a(0.07265973091125488)),(to_sfixed_a(0.0962296724319458)),(to_sfixed_a(0.1477448046207428)),(to_sfixed_a(-0.049663059413433075)),(to_sfixed_a(0.0912739485502243)),(to_sfixed_a(-0.014579487964510918)),(to_sfixed_a(8.240771421696991e-05)),(to_sfixed_a(0.00018982648907694966)),(to_sfixed_a(-8.852838072925806e-05)),(to_sfixed_a(0.00024077897251117975)),(to_sfixed_a(0.00011314231960568577)),(to_sfixed_a(8.165757026290521e-05)),(to_sfixed_a(-4.273305967217311e-05)),(to_sfixed_a(0.008932755328714848)),(to_sfixed_a(0.07813417166471481)),(to_sfixed_a(0.1305086612701416)),(to_sfixed_a(-0.2187996506690979)),(to_sfixed_a(0.07735536247491837)),(to_sfixed_a(0.1368907392024994)),(to_sfixed_a(0.10632581263780594)),(to_sfixed_a(0.11968968063592911)),(to_sfixed_a(0.17175404727458954)),(to_sfixed_a(-0.12945206463336945)),(to_sfixed_a(-0.26011431217193604)),(to_sfixed_a(0.014875062741339207)),(to_sfixed_a(-0.034548815339803696)),(to_sfixed_a(0.08520784974098206)),(to_sfixed_a(-0.19226479530334473)),(to_sfixed_a(0.04773328825831413)),(to_sfixed_a(-0.06441422551870346)),(to_sfixed_a(-0.04057212173938751)),(to_sfixed_a(0.0913177877664566)),(to_sfixed_a(-0.011310463771224022)),(to_sfixed_a(-0.018818197771906853)),(to_sfixed_a(-0.01799510419368744)),(to_sfixed_a(7.436953455908224e-05)),(to_sfixed_a(9.979999049392063e-06)),(to_sfixed_a(9.7016389190685e-05)),(to_sfixed_a(5.712181518902071e-05)),(to_sfixed_a(1.8207674656878226e-05)),(to_sfixed_a(-1.909603270178195e-05)),(to_sfixed_a(-0.0017424003453925252)),(to_sfixed_a(-4.2275765736121684e-05)),(to_sfixed_a(0.03797437623143196)),(to_sfixed_a(-0.040512025356292725)),(to_sfixed_a(-0.06254220008850098)),(to_sfixed_a(0.23207461833953857)),(to_sfixed_a(0.018985921517014503)),(to_sfixed_a(-0.16852609813213348)),(to_sfixed_a(-0.011493240483105183)),(to_sfixed_a(-0.0742889866232872)),(to_sfixed_a(-0.25245824456214905)),(to_sfixed_a(0.06705831736326218)),(to_sfixed_a(0.05263817310333252)),(to_sfixed_a(-0.24254350364208221)),(to_sfixed_a(-0.015001315623521805)),(to_sfixed_a(-0.040848374366760254)),(to_sfixed_a(0.003256944939494133)),(to_sfixed_a(0.06296908855438232)),(to_sfixed_a(-0.052841708064079285)),(to_sfixed_a(-0.011695285327732563)),(to_sfixed_a(-0.5795881748199463)),(to_sfixed_a(-3.862864559778245e-06)),(to_sfixed_a(0.0001786154170986265)),(to_sfixed_a(0.000260477012488991)),(to_sfixed_a(0.00018849861226044595)),(to_sfixed_a(-0.0003635305038187653)),(to_sfixed_a(0.000128881583805196)),(to_sfixed_a(0.00010051229037344456)),(to_sfixed_a(0.00010491936700418591)),(to_sfixed_a(-0.018065836280584335)),(to_sfixed_a(0.18316026031970978)),(to_sfixed_a(-0.3589034378528595)),(to_sfixed_a(-0.14283183217048645)),(to_sfixed_a(-0.03277391567826271)),(to_sfixed_a(-0.010654937475919724)),(to_sfixed_a(0.018302956596016884)),(to_sfixed_a(0.15927568078041077)),(to_sfixed_a(0.09974342584609985)),(to_sfixed_a(-0.2106417417526245)),(to_sfixed_a(-0.15606380999088287)),(to_sfixed_a(-0.21946494281291962)),(to_sfixed_a(-0.27917999029159546)),(to_sfixed_a(-0.015172258950769901)),(to_sfixed_a(-0.26978620886802673)),(to_sfixed_a(-0.10573842376470566)),(to_sfixed_a(-0.3141041696071625)),(to_sfixed_a(-0.23743021488189697)),(to_sfixed_a(-0.36566728353500366)),(to_sfixed_a(-0.24204149842262268)),(to_sfixed_a(0.017048515379428864)),(to_sfixed_a(-1.5928435459500179e-06)),(to_sfixed_a(-0.0001136980572482571)),(to_sfixed_a(-0.00011988139158347622)),(to_sfixed_a(4.6806904720142484e-05)),(to_sfixed_a(-3.138992906315252e-05)),(to_sfixed_a(-0.0002867623115889728)),(to_sfixed_a(6.820897056059039e-07)),(to_sfixed_a(-0.043701257556676865)),(to_sfixed_a(-0.0004929651040583849)),(to_sfixed_a(0.0868135541677475)),(to_sfixed_a(0.003140147775411606)),(to_sfixed_a(-0.0033638481982052326)),(to_sfixed_a(0.09684263169765472)),(to_sfixed_a(0.14160338044166565)),(to_sfixed_a(-0.14844831824302673)),(to_sfixed_a(0.12280025333166122)),(to_sfixed_a(-0.3090701997280121)),(to_sfixed_a(0.09703738242387772)),(to_sfixed_a(-0.03155362606048584)),(to_sfixed_a(-0.04518544301390648)),(to_sfixed_a(-0.1856933981180191)),(to_sfixed_a(-0.2266455590724945)),(to_sfixed_a(-0.08770786970853806)),(to_sfixed_a(-0.5799239277839661)),(to_sfixed_a(-0.16292527318000793)),(to_sfixed_a(-0.3107903301715851)),(to_sfixed_a(0.0004440605698619038)),(to_sfixed_a(-0.06378372013568878)),(to_sfixed_a(-9.671216685092077e-05)),(to_sfixed_a(0.00016920150665100664)),(to_sfixed_a(9.048819629242644e-05)),(to_sfixed_a(-4.312476085033268e-05)),(to_sfixed_a(9.65781364357099e-05)),(to_sfixed_a(-0.0001387222291668877)),(to_sfixed_a(0.00012176438758615404)),(to_sfixed_a(0.0001849218679126352)),(to_sfixed_a(-0.07248087972402573)),(to_sfixed_a(-0.0410938635468483)),(to_sfixed_a(0.0700756162405014)),(to_sfixed_a(-0.03937023878097534)),(to_sfixed_a(-0.010914686135947704)),(to_sfixed_a(0.013452383689582348)),(to_sfixed_a(0.004647971596568823)),(to_sfixed_a(0.0945981964468956)),(to_sfixed_a(0.09329212456941605)),(to_sfixed_a(-0.12064824253320694)),(to_sfixed_a(-0.02337573654949665)),(to_sfixed_a(-0.06495555490255356)),(to_sfixed_a(-0.015109867788851261)),(to_sfixed_a(-0.006140677258372307)),(to_sfixed_a(-0.186460480093956)),(to_sfixed_a(-0.12007458508014679)),(to_sfixed_a(-0.02525663748383522)),(to_sfixed_a(-0.09132129698991776)),(to_sfixed_a(-0.0038099924568086863)),(to_sfixed_a(0.00011581564467633143)),(to_sfixed_a(7.596601790282875e-05)),(to_sfixed_a(6.381914863595739e-05)),(to_sfixed_a(4.1223520383937284e-05)),(to_sfixed_a(8.788794366410002e-05)),(to_sfixed_a(0.0001624774740776047)),(to_sfixed_a(4.805768912774511e-05)),(to_sfixed_a(0.00016633805353194475)),(to_sfixed_a(0.00014824574464000762)),(to_sfixed_a(-0.029752586036920547)),(to_sfixed_a(0.017214994877576828)),(to_sfixed_a(0.2288302630186081)),(to_sfixed_a(-0.08331207931041718)),(to_sfixed_a(0.02430112659931183)),(to_sfixed_a(0.0076349107548594475)),(to_sfixed_a(-0.029275143519043922)),(to_sfixed_a(-0.15385940670967102)),(to_sfixed_a(0.11828333139419556)),(to_sfixed_a(-0.051323749125003815)),(to_sfixed_a(0.017640370875597)),(to_sfixed_a(-0.07452002912759781)),(to_sfixed_a(-0.22515809535980225)),(to_sfixed_a(-0.05718788132071495)),(to_sfixed_a(-0.12804169952869415)),(to_sfixed_a(-0.03959227353334427)),(to_sfixed_a(-0.16763204336166382)),(to_sfixed_a(-0.001314960652962327)),(to_sfixed_a(-0.12293771654367447)),(to_sfixed_a(0.00020181617583148181)),(to_sfixed_a(3.883153112838045e-05)),(to_sfixed_a(-0.00032080590608529747)),(to_sfixed_a(-7.543093670392409e-05)),(to_sfixed_a(0.00024389068130403757)),(to_sfixed_a(0.00016256202070508152)),(to_sfixed_a(9.077805771084968e-06)),(to_sfixed_a(-0.00010687181202229112)),(to_sfixed_a(-0.005861158948391676)),(to_sfixed_a(0.010651668533682823)),(to_sfixed_a(-0.024264339357614517)),(to_sfixed_a(-0.024260330945253372)),(to_sfixed_a(-0.03165422007441521)),(to_sfixed_a(-0.04272136837244034)),(to_sfixed_a(0.1909194141626358)),(to_sfixed_a(0.07100588828325272)),(to_sfixed_a(-0.1984747350215912)),(to_sfixed_a(0.1107010692358017)),(to_sfixed_a(-0.01060784887522459)),(to_sfixed_a(0.04697763919830322)),(to_sfixed_a(0.07321231812238693)),(to_sfixed_a(-0.15655004978179932)),(to_sfixed_a(0.027829790487885475)),(to_sfixed_a(-0.13084374368190765)),(to_sfixed_a(-0.005587409716099501)),(to_sfixed_a(-0.10613838583230972)),(to_sfixed_a(-0.06287290155887604)),(to_sfixed_a(0.001126133487559855)),(to_sfixed_a(-7.962223753565922e-05)),(to_sfixed_a(0.0002678881282918155)),(to_sfixed_a(-0.00024074251996353269)),(to_sfixed_a(8.513093052897602e-05)),(to_sfixed_a(-0.00010358464351156726)),(to_sfixed_a(1.4231331988412421e-05)),(to_sfixed_a(0.000331683928379789)),(to_sfixed_a(-4.563116453937255e-05)),(to_sfixed_a(8.895034989109263e-05)),(to_sfixed_a(-0.009383054450154305)),(to_sfixed_a(-0.014865325763821602)),(to_sfixed_a(-0.04118317738175392)),(to_sfixed_a(-0.09937461465597153)),(to_sfixed_a(0.09096261113882065)),(to_sfixed_a(0.042197685688734055)),(to_sfixed_a(0.14185525476932526)),(to_sfixed_a(0.20604294538497925)),(to_sfixed_a(-0.008855149149894714)),(to_sfixed_a(-0.1156487911939621)),(to_sfixed_a(-0.004729812033474445)),(to_sfixed_a(0.16798120737075806)),(to_sfixed_a(0.0568186491727829)),(to_sfixed_a(-0.001122006680816412)),(to_sfixed_a(0.29687368869781494)),(to_sfixed_a(0.18463942408561707)),(to_sfixed_a(0.00019038189202547073)),(to_sfixed_a(-0.0006724774139001966)),(to_sfixed_a(-0.0017532911151647568)),(to_sfixed_a(-7.287818880286068e-05)),(to_sfixed_a(-2.3156242605182342e-05)),(to_sfixed_a(5.248567958915373e-06)),(to_sfixed_a(0.00014474581985268742)),(to_sfixed_a(-7.545045809820294e-05)),(to_sfixed_a(-0.00011576699034776539)),(to_sfixed_a(-5.55641163373366e-05)),(to_sfixed_a(-0.00023972519556991756)),(to_sfixed_a(-1.9082982305462792e-07)),(to_sfixed_a(0.0014535593800246716)),(to_sfixed_a(0.0014744866639375687)),(to_sfixed_a(0.00011589814675971866)),(to_sfixed_a(0.00018527892825659364)),(to_sfixed_a(-0.00017215957632288337)),(to_sfixed_a(0.1810692995786667)),(to_sfixed_a(-0.0031046057119965553)),(to_sfixed_a(-0.0010333508253097534)),(to_sfixed_a(0.13722579181194305)),(to_sfixed_a(0.18859444558620453)),(to_sfixed_a(0.017209570854902267)),(to_sfixed_a(0.10983897745609283)),(to_sfixed_a(0.14454472064971924)),(to_sfixed_a(0.19488027691841125)),(to_sfixed_a(0.009769309312105179)),(to_sfixed_a(0.004523893352597952)),(to_sfixed_a(1.811198308132589e-05)),(to_sfixed_a(-1.32872655740357e-05)),(to_sfixed_a(1.4331761121866293e-05)),(to_sfixed_a(-2.2236057702684775e-05)),(to_sfixed_a(-0.00011285070650046691)),(to_sfixed_a(0.0002622302854433656)),(to_sfixed_a(-7.767498027533293e-05)),(to_sfixed_a(-2.5246612494811416e-05)),(to_sfixed_a(-0.00011627515777945518)),(to_sfixed_a(-0.00016033051360864192)),(to_sfixed_a(-0.00012029528443235904)),(to_sfixed_a(-0.00041060452349483967)),(to_sfixed_a(3.250305962865241e-05)),(to_sfixed_a(-3.83262631657999e-05)),(to_sfixed_a(-0.0001246944593731314)),(to_sfixed_a(0.00019818710279650986)),(to_sfixed_a(-5.4567830375162885e-05)),(to_sfixed_a(-0.00013070310524199158)),(to_sfixed_a(-0.000267611671006307)),(to_sfixed_a(-0.00017468685109633952)),(to_sfixed_a(0.0002693752176128328)),(to_sfixed_a(5.167966446606442e-05)),(to_sfixed_a(0.00010958877828670666)),(to_sfixed_a(1.4479447600024287e-05)),(to_sfixed_a(7.639583054697141e-05)),(to_sfixed_a(-0.00020619697170332074)),(to_sfixed_a(-0.0002410356537438929)),(to_sfixed_a(0.00030969514045864344)),(to_sfixed_a(-2.740871423156932e-06)),(to_sfixed_a(0.00017129040497820824)),(to_sfixed_a(0.00024967562058009207)),(to_sfixed_a(-1.547303668303357e-06)),(to_sfixed_a(-0.0001541025994811207)),(to_sfixed_a(5.160695582162589e-05)),(to_sfixed_a(0.0004063384549226612)));

    constant weight_n0_14 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(9.232769662048668e-05)),(to_sfixed_a(0.0001061729562934488)),(to_sfixed_a(-0.0003311135806143284)),(to_sfixed_a(0.0002588743227533996)),(to_sfixed_a(4.395955693325959e-05)),(to_sfixed_a(-0.00015326292486861348)),(to_sfixed_a(0.0002266935771331191)),(to_sfixed_a(0.00010878252214752138)),(to_sfixed_a(0.0002495530934538692)),(to_sfixed_a(-0.00014110907795839012)),(to_sfixed_a(-0.0001583208068041131)),(to_sfixed_a(-3.4392123779980466e-05)),(to_sfixed_a(-6.291190948104486e-05)),(to_sfixed_a(0.00016101018991321325)),(to_sfixed_a(0.00015372820780612528)),(to_sfixed_a(-0.0001070583239197731)),(to_sfixed_a(0.0001501278456998989)),(to_sfixed_a(-8.062865163083188e-06)),(to_sfixed_a(0.00010992681927746162)),(to_sfixed_a(-0.000453267217380926)),(to_sfixed_a(-4.7925906983437017e-05)),(to_sfixed_a(1.4274584827944636e-05)),(to_sfixed_a(0.0003037700953427702)),(to_sfixed_a(0.00018522058962844312)),(to_sfixed_a(8.332840479852166e-06)),(to_sfixed_a(-0.00017475703498348594)),(to_sfixed_a(-4.5670232793781906e-05)),(to_sfixed_a(-0.00038455025060102344)),(to_sfixed_a(0.00033410813193768263)),(to_sfixed_a(-0.000277425890089944)),(to_sfixed_a(7.087218546075746e-05)),(to_sfixed_a(-2.7737278287531808e-05)),(to_sfixed_a(-0.0003146457311231643)),(to_sfixed_a(1.2947114555572625e-05)),(to_sfixed_a(-0.0004513444728218019)),(to_sfixed_a(-1.4475363968813326e-05)),(to_sfixed_a(4.104943855054444e-06)),(to_sfixed_a(-0.0002628148649819195)),(to_sfixed_a(-0.00015962179168127477)),(to_sfixed_a(7.098380592651665e-05)),(to_sfixed_a(-3.2116547199478873e-09)),(to_sfixed_a(8.418613288085908e-05)),(to_sfixed_a(0.00011795514001278207)),(to_sfixed_a(0.00017602481239009649)),(to_sfixed_a(-0.000409547210438177)),(to_sfixed_a(1.0322811249352526e-05)),(to_sfixed_a(0.0001630897750146687)),(to_sfixed_a(-0.00016346485062967986)),(to_sfixed_a(3.868638668791391e-05)),(to_sfixed_a(8.840460941428319e-05)),(to_sfixed_a(-0.00016659076209180057)),(to_sfixed_a(-4.258775879861787e-05)),(to_sfixed_a(0.00014273502165451646)),(to_sfixed_a(4.3282616388751194e-05)),(to_sfixed_a(-0.00012863989104516804)),(to_sfixed_a(0.00023801150382496417)),(to_sfixed_a(-1.370223344565602e-05)),(to_sfixed_a(0.00023792409047018737)),(to_sfixed_a(-3.591350468923338e-05)),(to_sfixed_a(5.7659017329569906e-05)),(to_sfixed_a(7.270754576893523e-05)),(to_sfixed_a(-9.211694123223424e-05)),(to_sfixed_a(-2.3958982637850568e-05)),(to_sfixed_a(6.560940528288484e-05)),(to_sfixed_a(-7.115131302271038e-05)),(to_sfixed_a(0.00027380240499041975)),(to_sfixed_a(2.743118238868192e-05)),(to_sfixed_a(2.3352848074864596e-05)),(to_sfixed_a(-5.2506698011711705e-06)),(to_sfixed_a(0.010948159731924534)),(to_sfixed_a(6.875287363072857e-05)),(to_sfixed_a(-8.116806566249579e-05)),(to_sfixed_a(-9.623949154047295e-05)),(to_sfixed_a(0.00016385888739023358)),(to_sfixed_a(-0.00015956444258335978)),(to_sfixed_a(-5.204457920626737e-05)),(to_sfixed_a(-0.00018017133697867393)),(to_sfixed_a(-0.00029935649945400655)),(to_sfixed_a(-1.49620245792903e-05)),(to_sfixed_a(0.000272634148132056)),(to_sfixed_a(-8.82509266375564e-05)),(to_sfixed_a(0.00024201010819524527)),(to_sfixed_a(1.9798578421159618e-07)),(to_sfixed_a(7.199382525868714e-05)),(to_sfixed_a(-6.666884291917086e-05)),(to_sfixed_a(0.00033899329719133675)),(to_sfixed_a(0.000289319985313341)),(to_sfixed_a(1.646786040510051e-05)),(to_sfixed_a(-5.129136116011068e-05)),(to_sfixed_a(-0.00018963679031003267)),(to_sfixed_a(0.0002853711193893105)),(to_sfixed_a(-6.469245272455737e-05)),(to_sfixed_a(-0.014082503505051136)),(to_sfixed_a(-7.668681064387783e-05)),(to_sfixed_a(-0.016058465465903282)),(to_sfixed_a(-0.05142868682742119)),(to_sfixed_a(-0.04830928146839142)),(to_sfixed_a(0.03553503379225731)),(to_sfixed_a(-0.054849524050951004)),(to_sfixed_a(0.0979078933596611)),(to_sfixed_a(-0.009249419905245304)),(to_sfixed_a(-0.018146062269806862)),(to_sfixed_a(0.07211262732744217)),(to_sfixed_a(0.07183884084224701)),(to_sfixed_a(0.028509778901934624)),(to_sfixed_a(0.0576135478913784)),(to_sfixed_a(9.33329138206318e-05)),(to_sfixed_a(-0.00014735784498043358)),(to_sfixed_a(1.2073471225448884e-05)),(to_sfixed_a(-8.748129039304331e-05)),(to_sfixed_a(0.00023577922547701746)),(to_sfixed_a(0.00010503894736757502)),(to_sfixed_a(-1.272697227250319e-05)),(to_sfixed_a(0.0001089817815227434)),(to_sfixed_a(0.0002485634759068489)),(to_sfixed_a(0.00035914353793486953)),(to_sfixed_a(-2.5517603717162274e-05)),(to_sfixed_a(5.630025043501519e-05)),(to_sfixed_a(0.0003054471453651786)),(to_sfixed_a(-0.043707337230443954)),(to_sfixed_a(0.04461784288287163)),(to_sfixed_a(-0.020146239548921585)),(to_sfixed_a(0.22527264058589935)),(to_sfixed_a(-0.023406600579619408)),(to_sfixed_a(0.08061957359313965)),(to_sfixed_a(0.1284884512424469)),(to_sfixed_a(0.06823761761188507)),(to_sfixed_a(0.05382498353719711)),(to_sfixed_a(0.1262834668159485)),(to_sfixed_a(0.10430257767438889)),(to_sfixed_a(-0.012524658814072609)),(to_sfixed_a(0.046232130378484726)),(to_sfixed_a(0.008557282388210297)),(to_sfixed_a(0.02584010735154152)),(to_sfixed_a(0.021691756322979927)),(to_sfixed_a(-2.16008356801467e-06)),(to_sfixed_a(0.0005731232231482863)),(to_sfixed_a(-3.4939919714815915e-05)),(to_sfixed_a(-0.0001920616050483659)),(to_sfixed_a(0.00024042153381742537)),(to_sfixed_a(0.0001038905029417947)),(to_sfixed_a(3.898439172189683e-05)),(to_sfixed_a(3.717430081451312e-05)),(to_sfixed_a(-0.0001345134514849633)),(to_sfixed_a(0.0009085259516723454)),(to_sfixed_a(-0.07891125977039337)),(to_sfixed_a(-0.013319792225956917)),(to_sfixed_a(-0.12625864148139954)),(to_sfixed_a(0.012049213983118534)),(to_sfixed_a(0.039358220994472504)),(to_sfixed_a(0.03019353374838829)),(to_sfixed_a(-0.2183811068534851)),(to_sfixed_a(-0.12569816410541534)),(to_sfixed_a(-0.037901848554611206)),(to_sfixed_a(-0.07939162105321884)),(to_sfixed_a(0.013608548790216446)),(to_sfixed_a(0.02362196147441864)),(to_sfixed_a(0.03771141916513443)),(to_sfixed_a(0.12308614701032639)),(to_sfixed_a(-0.03136010095477104)),(to_sfixed_a(0.07561536878347397)),(to_sfixed_a(-0.013295253738760948)),(to_sfixed_a(0.0018537468276917934)),(to_sfixed_a(0.06581667810678482)),(to_sfixed_a(0.0010287122568115592)),(to_sfixed_a(0.0006853670929558575)),(to_sfixed_a(-6.0526519519044086e-05)),(to_sfixed_a(-0.00010979911166941747)),(to_sfixed_a(-0.00031088004470802844)),(to_sfixed_a(0.00019480461196508259)),(to_sfixed_a(9.612170833861455e-05)),(to_sfixed_a(0.00019063238869421184)),(to_sfixed_a(0.00022378528956323862)),(to_sfixed_a(-0.07485498487949371)),(to_sfixed_a(-0.09246505051851273)),(to_sfixed_a(-0.02632218599319458)),(to_sfixed_a(0.005292609799653292)),(to_sfixed_a(-0.1533142626285553)),(to_sfixed_a(-0.03647048398852348)),(to_sfixed_a(-0.13881216943264008)),(to_sfixed_a(0.0855991467833519)),(to_sfixed_a(0.06673045456409454)),(to_sfixed_a(0.10461888462305069)),(to_sfixed_a(0.1267627477645874)),(to_sfixed_a(0.15397751331329346)),(to_sfixed_a(0.09179557114839554)),(to_sfixed_a(0.3291940689086914)),(to_sfixed_a(0.04200967773795128)),(to_sfixed_a(0.018015870824456215)),(to_sfixed_a(-0.013229801319539547)),(to_sfixed_a(-0.16134071350097656)),(to_sfixed_a(-0.12405059486627579)),(to_sfixed_a(0.0008948705508373678)),(to_sfixed_a(0.0005171378725208342)),(to_sfixed_a(0.0003878589777741581)),(to_sfixed_a(4.1721916204551235e-05)),(to_sfixed_a(0.00019775117107201368)),(to_sfixed_a(-0.000133577806991525)),(to_sfixed_a(0.0002409242297289893)),(to_sfixed_a(0.0001369748351862654)),(to_sfixed_a(0.0001002070857794024)),(to_sfixed_a(-0.03935880959033966)),(to_sfixed_a(-0.03160449489951134)),(to_sfixed_a(0.1471816450357437)),(to_sfixed_a(-0.2546120584011078)),(to_sfixed_a(-0.24365335702896118)),(to_sfixed_a(-0.3556288480758667)),(to_sfixed_a(-0.511868417263031)),(to_sfixed_a(-0.3033379912376404)),(to_sfixed_a(-0.45447033643722534)),(to_sfixed_a(-0.10827812552452087)),(to_sfixed_a(0.04021291807293892)),(to_sfixed_a(0.17356999218463898)),(to_sfixed_a(0.09047159552574158)),(to_sfixed_a(0.13558141887187958)),(to_sfixed_a(0.057201821357011795)),(to_sfixed_a(-0.12861832976341248)),(to_sfixed_a(0.01729321852326393)),(to_sfixed_a(-0.09611120074987411)),(to_sfixed_a(-0.10192450881004333)),(to_sfixed_a(-0.07862136512994766)),(to_sfixed_a(-0.0008460937533527613)),(to_sfixed_a(0.00012523421901278198)),(to_sfixed_a(-4.468468978302553e-05)),(to_sfixed_a(0.00017684561316855252)),(to_sfixed_a(-0.00019673534552566707)),(to_sfixed_a(3.785468652495183e-05)),(to_sfixed_a(-2.01158309209859e-05)),(to_sfixed_a(0.060577455908060074)),(to_sfixed_a(0.006911936216056347)),(to_sfixed_a(0.02645784057676792)),(to_sfixed_a(0.0997220054268837)),(to_sfixed_a(0.04303828999400139)),(to_sfixed_a(-0.18074414134025574)),(to_sfixed_a(-0.31019294261932373)),(to_sfixed_a(-0.1275402456521988)),(to_sfixed_a(-0.15035390853881836)),(to_sfixed_a(0.030143210664391518)),(to_sfixed_a(-0.01373734138906002)),(to_sfixed_a(0.16107779741287231)),(to_sfixed_a(-0.03822813555598259)),(to_sfixed_a(0.020474139600992203)),(to_sfixed_a(0.0010438195895403624)),(to_sfixed_a(-0.06848857551813126)),(to_sfixed_a(-0.12948442995548248)),(to_sfixed_a(-0.015442226082086563)),(to_sfixed_a(0.028705688193440437)),(to_sfixed_a(-0.20068752765655518)),(to_sfixed_a(-0.1015700101852417)),(to_sfixed_a(0.053587667644023895)),(to_sfixed_a(9.438386769033968e-05)),(to_sfixed_a(-0.00021926563931629062)),(to_sfixed_a(-6.143224891275167e-05)),(to_sfixed_a(-3.4600376238813624e-05)),(to_sfixed_a(-0.00014718026795890182)),(to_sfixed_a(-8.148056804202497e-05)),(to_sfixed_a(0.0006581256166100502)),(to_sfixed_a(-0.01599973253905773)),(to_sfixed_a(0.07236602157354355)),(to_sfixed_a(0.16414915025234222)),(to_sfixed_a(0.005945665296167135)),(to_sfixed_a(0.050406284630298615)),(to_sfixed_a(-0.3988519608974457)),(to_sfixed_a(-0.24358367919921875)),(to_sfixed_a(-0.42257630825042725)),(to_sfixed_a(-0.18206463754177094)),(to_sfixed_a(-0.2191552370786667)),(to_sfixed_a(0.016809746623039246)),(to_sfixed_a(0.2609507143497467)),(to_sfixed_a(0.03490271419286728)),(to_sfixed_a(0.09314731508493423)),(to_sfixed_a(-0.04349062219262123)),(to_sfixed_a(-0.03591964393854141)),(to_sfixed_a(-0.15156809985637665)),(to_sfixed_a(-0.150089830160141)),(to_sfixed_a(-0.0699453353881836)),(to_sfixed_a(0.06924623996019363)),(to_sfixed_a(6.140589903225191e-06)),(to_sfixed_a(-3.746795482584275e-05)),(to_sfixed_a(-5.679572495864704e-05)),(to_sfixed_a(-2.5011158868437633e-05)),(to_sfixed_a(1.827175947255455e-05)),(to_sfixed_a(0.0003366720920894295)),(to_sfixed_a(3.1399107683682814e-05)),(to_sfixed_a(-0.005575146060436964)),(to_sfixed_a(0.004551286809146404)),(to_sfixed_a(0.09274805337190628)),(to_sfixed_a(0.10437405109405518)),(to_sfixed_a(0.09952516853809357)),(to_sfixed_a(-0.057991091161966324)),(to_sfixed_a(0.052339326590299606)),(to_sfixed_a(-0.018152939155697823)),(to_sfixed_a(0.0935235321521759)),(to_sfixed_a(0.21746104955673218)),(to_sfixed_a(0.13410566747188568)),(to_sfixed_a(0.4058496952056885)),(to_sfixed_a(0.20795074105262756)),(to_sfixed_a(0.18972225487232208)),(to_sfixed_a(0.16626803576946259)),(to_sfixed_a(0.133169487118721)),(to_sfixed_a(-0.08682587742805481)),(to_sfixed_a(-0.3206895887851715)),(to_sfixed_a(0.11392869055271149)),(to_sfixed_a(-0.029381053522229195)),(to_sfixed_a(0.11636079847812653)),(to_sfixed_a(0.001132803037762642)),(to_sfixed_a(3.344150854900363e-06)),(to_sfixed_a(5.7654415286378935e-05)),(to_sfixed_a(0.00023835331376176327)),(to_sfixed_a(1.0459628356329631e-05)),(to_sfixed_a(-0.00011117885878775269)),(to_sfixed_a(0.03741106018424034)),(to_sfixed_a(0.14567464590072632)),(to_sfixed_a(0.1393055021762848)),(to_sfixed_a(0.053353581577539444)),(to_sfixed_a(0.1939932405948639)),(to_sfixed_a(-0.01078916434198618)),(to_sfixed_a(-0.04593278840184212)),(to_sfixed_a(-0.07117466628551483)),(to_sfixed_a(-0.15138530731201172)),(to_sfixed_a(-0.2268151193857193)),(to_sfixed_a(0.11804036796092987)),(to_sfixed_a(-0.15878655016422272)),(to_sfixed_a(0.3225403130054474)),(to_sfixed_a(0.057910844683647156)),(to_sfixed_a(-0.10039281100034714)),(to_sfixed_a(0.07178319245576859)),(to_sfixed_a(0.22340445220470428)),(to_sfixed_a(0.25692641735076904)),(to_sfixed_a(0.06903987377882004)),(to_sfixed_a(-0.15530607104301453)),(to_sfixed_a(-0.011652148328721523)),(to_sfixed_a(0.1768115907907486)),(to_sfixed_a(0.00013891640992369503)),(to_sfixed_a(-4.02272999053821e-05)),(to_sfixed_a(0.00013472657883539796)),(to_sfixed_a(6.932010728633031e-05)),(to_sfixed_a(0.00019257447274867445)),(to_sfixed_a(-0.00025330751668661833)),(to_sfixed_a(7.004325743764639e-05)),(to_sfixed_a(-0.03325118497014046)),(to_sfixed_a(-0.11257120221853256)),(to_sfixed_a(0.002024225890636444)),(to_sfixed_a(-0.05874723568558693)),(to_sfixed_a(0.06325887888669968)),(to_sfixed_a(-0.2611834704875946)),(to_sfixed_a(-0.3553241491317749)),(to_sfixed_a(-0.33897456526756287)),(to_sfixed_a(-0.31808820366859436)),(to_sfixed_a(0.18270951509475708)),(to_sfixed_a(-0.1339130401611328)),(to_sfixed_a(0.060067202895879745)),(to_sfixed_a(-0.05695130303502083)),(to_sfixed_a(-0.1380373239517212)),(to_sfixed_a(-0.06612478196620941)),(to_sfixed_a(-0.23408474028110504)),(to_sfixed_a(0.4374091923236847)),(to_sfixed_a(0.09864547103643417)),(to_sfixed_a(0.025876492261886597)),(to_sfixed_a(0.25974905490875244)),(to_sfixed_a(-0.2211010605096817)),(to_sfixed_a(-5.254521602182649e-05)),(to_sfixed_a(0.0005670203827321529)),(to_sfixed_a(9.634403141944858e-08)),(to_sfixed_a(-0.00011931782501051202)),(to_sfixed_a(8.994658128358424e-05)),(to_sfixed_a(-1.4925662981113419e-05)),(to_sfixed_a(0.00031955569284036756)),(to_sfixed_a(-0.03714684396982193)),(to_sfixed_a(0.04716816172003746)),(to_sfixed_a(-0.10511825233697891)),(to_sfixed_a(-0.034015554934740067)),(to_sfixed_a(-0.06188059598207474)),(to_sfixed_a(-0.17145253717899323)),(to_sfixed_a(0.013452336192131042)),(to_sfixed_a(-0.052649177610874176)),(to_sfixed_a(-0.29078441858291626)),(to_sfixed_a(-0.24710431694984436)),(to_sfixed_a(-0.5384657979011536)),(to_sfixed_a(-0.48553192615509033)),(to_sfixed_a(-0.20380151271820068)),(to_sfixed_a(-0.32302016019821167)),(to_sfixed_a(-0.14040666818618774)),(to_sfixed_a(0.02535567805171013)),(to_sfixed_a(-0.03260905295610428)),(to_sfixed_a(0.046923618763685226)),(to_sfixed_a(0.1255543977022171)),(to_sfixed_a(-0.0017842577071860433)),(to_sfixed_a(-0.016693616285920143)),(to_sfixed_a(0.0016724570887163281)),(to_sfixed_a(0.0014373058220371604)),(to_sfixed_a(-0.00013805952039547265)),(to_sfixed_a(-0.0002661388134583831)),(to_sfixed_a(-2.907825546571985e-06)),(to_sfixed_a(-1.7564794688951224e-05)),(to_sfixed_a(-0.00010713136725826189)),(to_sfixed_a(-0.0013617066433653235)),(to_sfixed_a(0.2029993087053299)),(to_sfixed_a(0.14049816131591797)),(to_sfixed_a(-0.021006470546126366)),(to_sfixed_a(0.16505374014377594)),(to_sfixed_a(-0.19232042133808136)),(to_sfixed_a(-0.09789638221263885)),(to_sfixed_a(0.09705567359924316)),(to_sfixed_a(-0.028333202004432678)),(to_sfixed_a(0.0498555488884449)),(to_sfixed_a(-0.21793577075004578)),(to_sfixed_a(-0.17523866891860962)),(to_sfixed_a(-0.17799049615859985)),(to_sfixed_a(-0.10700707137584686)),(to_sfixed_a(0.13634636998176575)),(to_sfixed_a(0.1778813600540161)),(to_sfixed_a(0.07395615428686142)),(to_sfixed_a(0.12850800156593323)),(to_sfixed_a(-0.00904749520123005)),(to_sfixed_a(-0.10468897223472595)),(to_sfixed_a(-0.10173749178647995)),(to_sfixed_a(-0.0002251725527457893)),(to_sfixed_a(-0.00024708634009584785)),(to_sfixed_a(1.4878161891829222e-05)),(to_sfixed_a(0.00016791047528386116)),(to_sfixed_a(-0.00019993717432953417)),(to_sfixed_a(-0.0001581064279889688)),(to_sfixed_a(1.1658179573714733e-05)),(to_sfixed_a(0.036452241241931915)),(to_sfixed_a(0.18037134408950806)),(to_sfixed_a(0.2060391902923584)),(to_sfixed_a(0.21154798567295074)),(to_sfixed_a(0.21359804272651672)),(to_sfixed_a(0.22019346058368683)),(to_sfixed_a(0.02854837477207184)),(to_sfixed_a(-0.0627325028181076)),(to_sfixed_a(0.16157205402851105)),(to_sfixed_a(-0.053480446338653564)),(to_sfixed_a(-0.21252773702144623)),(to_sfixed_a(-0.05801694467663765)),(to_sfixed_a(-0.015677355229854584)),(to_sfixed_a(-0.32012271881103516)),(to_sfixed_a(0.012709027156233788)),(to_sfixed_a(-0.023950699716806412)),(to_sfixed_a(-0.14013181626796722)),(to_sfixed_a(-0.02996160089969635)),(to_sfixed_a(0.10687437653541565)),(to_sfixed_a(-0.12031538784503937)),(to_sfixed_a(-0.09885457158088684)),(to_sfixed_a(-0.00014796132745686918)),(to_sfixed_a(5.919790419284254e-05)),(to_sfixed_a(2.0996718376409262e-05)),(to_sfixed_a(6.021236549713649e-05)),(to_sfixed_a(-0.0002368386776652187)),(to_sfixed_a(0.0004759903240483254)),(to_sfixed_a(0.002234991639852524)),(to_sfixed_a(0.04559760168194771)),(to_sfixed_a(0.11065446585416794)),(to_sfixed_a(0.00040377260302193463)),(to_sfixed_a(0.036592934280633926)),(to_sfixed_a(-0.03691554442048073)),(to_sfixed_a(-0.24830223619937897)),(to_sfixed_a(0.04540480300784111)),(to_sfixed_a(0.20014333724975586)),(to_sfixed_a(0.20944324135780334)),(to_sfixed_a(-0.20974324643611908)),(to_sfixed_a(-0.011907982639968395)),(to_sfixed_a(-0.15092997252941132)),(to_sfixed_a(0.058238182216882706)),(to_sfixed_a(-0.08246995508670807)),(to_sfixed_a(0.14913584291934967)),(to_sfixed_a(-0.01291398424655199)),(to_sfixed_a(-0.08396269381046295)),(to_sfixed_a(-0.03704463317990303)),(to_sfixed_a(0.0014804238453507423)),(to_sfixed_a(0.10977691411972046)),(to_sfixed_a(-0.05052518844604492)),(to_sfixed_a(0.018074210733175278)),(to_sfixed_a(9.40040081331972e-06)),(to_sfixed_a(0.00017560728883836418)),(to_sfixed_a(0.00023049353330861777)),(to_sfixed_a(-8.7419779447373e-05)),(to_sfixed_a(0.0015320932725444436)),(to_sfixed_a(0.0019800022710114717)),(to_sfixed_a(0.14896337687969208)),(to_sfixed_a(0.043831948190927505)),(to_sfixed_a(-0.020115403458476067)),(to_sfixed_a(-0.11119549721479416)),(to_sfixed_a(-0.4159241020679474)),(to_sfixed_a(-0.44348469376564026)),(to_sfixed_a(-0.09903470426797867)),(to_sfixed_a(0.19286267459392548)),(to_sfixed_a(0.5809189677238464)),(to_sfixed_a(0.11095483601093292)),(to_sfixed_a(-0.003595733782276511)),(to_sfixed_a(0.1095641478896141)),(to_sfixed_a(0.09294898062944412)),(to_sfixed_a(0.04116327315568924)),(to_sfixed_a(-0.019259992986917496)),(to_sfixed_a(-0.05534438043832779)),(to_sfixed_a(-0.0028541383799165487)),(to_sfixed_a(-0.006142588797956705)),(to_sfixed_a(-0.1585816890001297)),(to_sfixed_a(0.033617399632930756)),(to_sfixed_a(-0.00013413916167337447)),(to_sfixed_a(-0.00011345365783199668)),(to_sfixed_a(-4.843604619964026e-05)),(to_sfixed_a(-0.00028552449657581747)),(to_sfixed_a(-0.00017472232866566628)),(to_sfixed_a(4.1207920730812475e-05)),(to_sfixed_a(0.00035856489557772875)),(to_sfixed_a(-0.08031754940748215)),(to_sfixed_a(-0.18441356718540192)),(to_sfixed_a(0.007129507139325142)),(to_sfixed_a(-0.20863187313079834)),(to_sfixed_a(0.23585297167301178)),(to_sfixed_a(0.007613722234964371)),(to_sfixed_a(-0.2456798106431961)),(to_sfixed_a(-0.257355660200119)),(to_sfixed_a(0.016125788912177086)),(to_sfixed_a(0.3829757273197174)),(to_sfixed_a(0.2559703588485718)),(to_sfixed_a(-0.00797036848962307)),(to_sfixed_a(0.2863008975982666)),(to_sfixed_a(-0.020166737958788872)),(to_sfixed_a(0.04053351655602455)),(to_sfixed_a(0.0980127602815628)),(to_sfixed_a(-0.09813034534454346)),(to_sfixed_a(-0.031974658370018005)),(to_sfixed_a(-0.45042136311531067)),(to_sfixed_a(-0.11741641163825989)),(to_sfixed_a(0.009081867523491383)),(to_sfixed_a(0.023883556947112083)),(to_sfixed_a(1.5053530660225078e-05)),(to_sfixed_a(-0.0003050788654945791)),(to_sfixed_a(-0.0001990404271055013)),(to_sfixed_a(-0.000128591651446186)),(to_sfixed_a(0.00025092693977057934)),(to_sfixed_a(4.4739565055351704e-05)),(to_sfixed_a(-0.1184925064444542)),(to_sfixed_a(0.0028915945440530777)),(to_sfixed_a(0.05867336690425873)),(to_sfixed_a(-0.11372777819633484)),(to_sfixed_a(-0.23249049484729767)),(to_sfixed_a(-0.34682533144950867)),(to_sfixed_a(-0.14133746922016144)),(to_sfixed_a(0.08814242482185364)),(to_sfixed_a(0.0752822607755661)),(to_sfixed_a(0.023160308599472046)),(to_sfixed_a(0.20452040433883667)),(to_sfixed_a(0.2815495431423187)),(to_sfixed_a(0.35640618205070496)),(to_sfixed_a(-0.052338287234306335)),(to_sfixed_a(0.041354089975357056)),(to_sfixed_a(0.0422426275908947)),(to_sfixed_a(-0.0022586355917155743)),(to_sfixed_a(-0.12876783311367035)),(to_sfixed_a(-0.26828494668006897)),(to_sfixed_a(-0.15787142515182495)),(to_sfixed_a(-0.13329249620437622)),(to_sfixed_a(2.9201662982814014e-05)),(to_sfixed_a(-0.00011334118607919663)),(to_sfixed_a(-0.00014531287888530642)),(to_sfixed_a(4.208774771541357e-05)),(to_sfixed_a(-7.133709914342035e-06)),(to_sfixed_a(-8.88223439687863e-05)),(to_sfixed_a(-0.00019166120910085738)),(to_sfixed_a(-0.00010487027611816302)),(to_sfixed_a(0.006510268431156874)),(to_sfixed_a(0.03515185788273811)),(to_sfixed_a(0.006347862537950277)),(to_sfixed_a(0.13705815374851227)),(to_sfixed_a(-0.23634958267211914)),(to_sfixed_a(0.028390390798449516)),(to_sfixed_a(0.17486517131328583)),(to_sfixed_a(0.6813410520553589)),(to_sfixed_a(0.6954467296600342)),(to_sfixed_a(0.08387858420610428)),(to_sfixed_a(0.5553216934204102)),(to_sfixed_a(0.13864393532276154)),(to_sfixed_a(0.04808256775140762)),(to_sfixed_a(0.4287674129009247)),(to_sfixed_a(0.022116325795650482)),(to_sfixed_a(-0.24634769558906555)),(to_sfixed_a(-0.40867576003074646)),(to_sfixed_a(-0.11244337260723114)),(to_sfixed_a(-0.080951988697052)),(to_sfixed_a(-0.02005583420395851)),(to_sfixed_a(0.05199175700545311)),(to_sfixed_a(0.000244193768594414)),(to_sfixed_a(-0.00028079876210540533)),(to_sfixed_a(-0.0001764883636496961)),(to_sfixed_a(2.9383369110291824e-05)),(to_sfixed_a(-7.743113383185118e-05)),(to_sfixed_a(7.625017315149307e-05)),(to_sfixed_a(-7.012456626398489e-05)),(to_sfixed_a(-0.010360865853726864)),(to_sfixed_a(-0.0003066523640882224)),(to_sfixed_a(-0.079582579433918)),(to_sfixed_a(0.05670354887843132)),(to_sfixed_a(0.2653086483478546)),(to_sfixed_a(0.12116225808858871)),(to_sfixed_a(0.15260183811187744)),(to_sfixed_a(0.3218518793582916)),(to_sfixed_a(0.43744122982025146)),(to_sfixed_a(0.3855297863483429)),(to_sfixed_a(0.6474530100822449)),(to_sfixed_a(0.28183501958847046)),(to_sfixed_a(0.17374181747436523)),(to_sfixed_a(0.40694770216941833)),(to_sfixed_a(-0.008381656371057034)),(to_sfixed_a(-0.1356082707643509)),(to_sfixed_a(-0.4043339192867279)),(to_sfixed_a(-0.13509799540042877)),(to_sfixed_a(-0.1285339742898941)),(to_sfixed_a(-0.0006438244599848986)),(to_sfixed_a(-0.08654575794935226)),(to_sfixed_a(-5.048178354627453e-05)),(to_sfixed_a(-9.418228000868112e-05)),(to_sfixed_a(6.736120121786371e-05)),(to_sfixed_a(4.737201743409969e-05)),(to_sfixed_a(-4.358630030765198e-05)),(to_sfixed_a(-9.70600922300946e-06)),(to_sfixed_a(-0.0001260278222616762)),(to_sfixed_a(-0.0001877628092188388)),(to_sfixed_a(0.06748364865779877)),(to_sfixed_a(-0.08751751482486725)),(to_sfixed_a(0.014029237441718578)),(to_sfixed_a(0.025393497198820114)),(to_sfixed_a(0.23807848989963531)),(to_sfixed_a(0.2930627465248108)),(to_sfixed_a(0.21890302002429962)),(to_sfixed_a(0.21483387053012848)),(to_sfixed_a(0.24272038042545319)),(to_sfixed_a(0.14258906245231628)),(to_sfixed_a(0.4590497612953186)),(to_sfixed_a(0.15942151844501495)),(to_sfixed_a(-0.16216160356998444)),(to_sfixed_a(-0.04672866687178612)),(to_sfixed_a(0.09464624524116516)),(to_sfixed_a(-0.04522058740258217)),(to_sfixed_a(-0.018323823809623718)),(to_sfixed_a(-0.09891372174024582)),(to_sfixed_a(0.003149047726765275)),(to_sfixed_a(-3.4504944778745994e-05)),(to_sfixed_a(-0.0003246220585424453)),(to_sfixed_a(-5.2362302085384727e-05)),(to_sfixed_a(-9.370195039082319e-05)),(to_sfixed_a(-9.76968658505939e-05)),(to_sfixed_a(9.619382763048634e-05)),(to_sfixed_a(0.0001309537183260545)),(to_sfixed_a(-7.213079516077414e-05)),(to_sfixed_a(-0.00040734626236371696)),(to_sfixed_a(0.019428687170147896)),(to_sfixed_a(-0.023065289482474327)),(to_sfixed_a(-0.1458478569984436)),(to_sfixed_a(-0.21637572348117828)),(to_sfixed_a(0.18034228682518005)),(to_sfixed_a(0.08755096793174744)),(to_sfixed_a(0.18573816120624542)),(to_sfixed_a(0.046287886798381805)),(to_sfixed_a(0.014926615171134472)),(to_sfixed_a(0.0087524289265275)),(to_sfixed_a(0.24368001520633698)),(to_sfixed_a(0.06195713207125664)),(to_sfixed_a(0.10754060745239258)),(to_sfixed_a(0.027703002095222473)),(to_sfixed_a(-0.03898981958627701)),(to_sfixed_a(0.02792702056467533)),(to_sfixed_a(-0.01897668093442917)),(to_sfixed_a(-0.008638952858746052)),(to_sfixed_a(-0.011494260281324387)),(to_sfixed_a(0.00019917925237677991)),(to_sfixed_a(-0.00014343678776640445)),(to_sfixed_a(7.36266520107165e-05)),(to_sfixed_a(3.27565248881001e-05)),(to_sfixed_a(1.9729541236301884e-05)),(to_sfixed_a(3.8275007682386786e-05)),(to_sfixed_a(0.00011081998673034832)),(to_sfixed_a(-7.292455120477825e-05)),(to_sfixed_a(0.001554455840960145)),(to_sfixed_a(0.00029019592329859734)),(to_sfixed_a(0.005725301802158356)),(to_sfixed_a(0.05440332740545273)),(to_sfixed_a(-0.08520609885454178)),(to_sfixed_a(-0.11624226719141006)),(to_sfixed_a(-0.13927410542964935)),(to_sfixed_a(0.05532694607973099)),(to_sfixed_a(-0.09806004166603088)),(to_sfixed_a(0.11596301198005676)),(to_sfixed_a(-0.1722177416086197)),(to_sfixed_a(0.09307784587144852)),(to_sfixed_a(0.2578706443309784)),(to_sfixed_a(0.4504433870315552)),(to_sfixed_a(-0.01352649461477995)),(to_sfixed_a(-0.016399413347244263)),(to_sfixed_a(-0.006748090032488108)),(to_sfixed_a(-0.03788380324840546)),(to_sfixed_a(-0.031741514801979065)),(to_sfixed_a(-0.02553764171898365)),(to_sfixed_a(-0.00026000174693763256)),(to_sfixed_a(6.443130132538499e-06)),(to_sfixed_a(0.00012600481568370014)),(to_sfixed_a(9.956111171049997e-05)),(to_sfixed_a(0.00010461026977282017)),(to_sfixed_a(-3.1911498808767647e-05)),(to_sfixed_a(8.204477489925921e-05)),(to_sfixed_a(-0.00014283631753642112)),(to_sfixed_a(-0.0003004627942573279)),(to_sfixed_a(-0.028490539640188217)),(to_sfixed_a(0.003809843910858035)),(to_sfixed_a(0.020331745967268944)),(to_sfixed_a(0.05743783339858055)),(to_sfixed_a(0.137782484292984)),(to_sfixed_a(-0.014586293138563633)),(to_sfixed_a(-0.14257676899433136)),(to_sfixed_a(-0.09800813347101212)),(to_sfixed_a(-0.12491209805011749)),(to_sfixed_a(0.06544386595487595)),(to_sfixed_a(0.08741305768489838)),(to_sfixed_a(0.04553770273923874)),(to_sfixed_a(-0.01312924548983574)),(to_sfixed_a(-0.005683894269168377)),(to_sfixed_a(-0.10839243978261948)),(to_sfixed_a(-0.08686794340610504)),(to_sfixed_a(-0.001321339514106512)),(to_sfixed_a(-0.006076856050640345)),(to_sfixed_a(-0.007128952071070671)),(to_sfixed_a(-1.249064825969981e-05)),(to_sfixed_a(-0.00017846217087935656)),(to_sfixed_a(7.289257337106392e-05)),(to_sfixed_a(-4.847560830967268e-06)),(to_sfixed_a(8.051255281316116e-05)),(to_sfixed_a(-3.490430026431568e-05)),(to_sfixed_a(0.00010012416896643117)),(to_sfixed_a(0.0002147964114556089)),(to_sfixed_a(-5.5545959185110405e-05)),(to_sfixed_a(0.001385197159834206)),(to_sfixed_a(0.0013289098860695958)),(to_sfixed_a(-1.467217458639425e-07)),(to_sfixed_a(-3.264922997914255e-05)),(to_sfixed_a(-0.0003547185624483973)),(to_sfixed_a(-0.08122208714485168)),(to_sfixed_a(-0.006902661174535751)),(to_sfixed_a(0.0011183388996869326)),(to_sfixed_a(-0.06313575804233551)),(to_sfixed_a(0.06287454068660736)),(to_sfixed_a(0.006393060088157654)),(to_sfixed_a(-0.022074712440371513)),(to_sfixed_a(-0.0630032941699028)),(to_sfixed_a(-0.08885692059993744)),(to_sfixed_a(-0.006419735960662365)),(to_sfixed_a(-0.004413362592458725)),(to_sfixed_a(0.0001594316854607314)),(to_sfixed_a(-0.0001308991340920329)),(to_sfixed_a(-4.132604590267874e-05)),(to_sfixed_a(-3.6737827031174675e-05)),(to_sfixed_a(-0.00010341274173697457)),(to_sfixed_a(0.00017765947268344462)),(to_sfixed_a(-6.344738358166069e-05)),(to_sfixed_a(-8.377728227060288e-05)),(to_sfixed_a(-0.0004972179303877056)),(to_sfixed_a(6.259678048081696e-05)),(to_sfixed_a(9.886779298540205e-05)),(to_sfixed_a(9.846310422290117e-05)),(to_sfixed_a(0.00028084387304261327)),(to_sfixed_a(7.462932990165427e-05)),(to_sfixed_a(-0.00012789924221578985)),(to_sfixed_a(0.00029862302471883595)),(to_sfixed_a(7.070855644997209e-05)),(to_sfixed_a(-0.0002245232171844691)),(to_sfixed_a(0.0001667510805418715)),(to_sfixed_a(0.00029650269425474107)),(to_sfixed_a(0.0001602252887096256)),(to_sfixed_a(-0.0001487478002673015)),(to_sfixed_a(3.1898915040073916e-05)),(to_sfixed_a(3.9421342080459e-05)),(to_sfixed_a(3.731468314072117e-05)),(to_sfixed_a(2.7523106837179512e-05)),(to_sfixed_a(-1.839235847000964e-05)),(to_sfixed_a(-6.876913539599627e-05)),(to_sfixed_a(-0.000224092771532014)),(to_sfixed_a(-3.471085801720619e-05)),(to_sfixed_a(7.70882106735371e-05)),(to_sfixed_a(-8.435919153271243e-05)),(to_sfixed_a(0.00021264016686473042)),(to_sfixed_a(-3.50285044987686e-05)),(to_sfixed_a(-0.000340430939104408)));

    constant weight_n0_15 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(9.494935511611402e-05)),(to_sfixed_a(-0.0003201631479896605)),(to_sfixed_a(-6.100515747675672e-05)),(to_sfixed_a(0.0005344618111848831)),(to_sfixed_a(-0.00017638245481066406)),(to_sfixed_a(0.0002118901611538604)),(to_sfixed_a(-0.0003509313683025539)),(to_sfixed_a(8.680066093802452e-05)),(to_sfixed_a(-6.336237129289657e-05)),(to_sfixed_a(0.00015700455696787685)),(to_sfixed_a(9.162275091512129e-05)),(to_sfixed_a(-0.00014126941096037626)),(to_sfixed_a(3.974799983552657e-05)),(to_sfixed_a(9.219579806085676e-05)),(to_sfixed_a(2.5993669623858295e-05)),(to_sfixed_a(-4.048399205203168e-05)),(to_sfixed_a(9.247071830031928e-06)),(to_sfixed_a(7.700115929765161e-06)),(to_sfixed_a(-0.00016538859927095473)),(to_sfixed_a(-4.653229552786797e-05)),(to_sfixed_a(0.00037963397335261106)),(to_sfixed_a(3.224477404728532e-05)),(to_sfixed_a(-0.000293643563054502)),(to_sfixed_a(6.31019429420121e-05)),(to_sfixed_a(0.0001508092536823824)),(to_sfixed_a(-0.0003186596732120961)),(to_sfixed_a(0.00019171526946593076)),(to_sfixed_a(5.543352381209843e-05)),(to_sfixed_a(-6.050406227586791e-05)),(to_sfixed_a(6.106174987507984e-05)),(to_sfixed_a(0.00020701884932350367)),(to_sfixed_a(0.00011610157525865361)),(to_sfixed_a(-6.0855043557239696e-05)),(to_sfixed_a(0.00013089952699374408)),(to_sfixed_a(6.498058792203665e-05)),(to_sfixed_a(0.0002640091988723725)),(to_sfixed_a(-0.000169567356351763)),(to_sfixed_a(0.00027659095940180123)),(to_sfixed_a(-0.00033400728716515005)),(to_sfixed_a(-5.753305958933197e-05)),(to_sfixed_a(0.00012960282037965953)),(to_sfixed_a(0.0001804193016141653)),(to_sfixed_a(1.0898391337832436e-05)),(to_sfixed_a(-0.00011213200923521072)),(to_sfixed_a(0.000227013006224297)),(to_sfixed_a(0.00013400113675743341)),(to_sfixed_a(-0.00017602075240574777)),(to_sfixed_a(-3.0035230338398833e-06)),(to_sfixed_a(-0.0002851895696949214)),(to_sfixed_a(-0.00018635104061104357)),(to_sfixed_a(-0.00032917558564804494)),(to_sfixed_a(-0.0001813816634239629)),(to_sfixed_a(-9.457849955651909e-05)),(to_sfixed_a(0.00023115810472518206)),(to_sfixed_a(4.3270982132526115e-05)),(to_sfixed_a(-0.00023211154621094465)),(to_sfixed_a(7.735293183941394e-05)),(to_sfixed_a(-2.3964163119671866e-05)),(to_sfixed_a(7.65684453654103e-05)),(to_sfixed_a(1.1490125871205237e-05)),(to_sfixed_a(0.000334374257363379)),(to_sfixed_a(1.1490410543046892e-05)),(to_sfixed_a(0.00014864314289297909)),(to_sfixed_a(3.091669350396842e-05)),(to_sfixed_a(-0.0004444414225872606)),(to_sfixed_a(0.0002363808307563886)),(to_sfixed_a(0.00016940214845817536)),(to_sfixed_a(0.00016026604862418026)),(to_sfixed_a(0.00022054840519558638)),(to_sfixed_a(-0.004430805332958698)),(to_sfixed_a(-9.119027708948124e-06)),(to_sfixed_a(4.752466702484526e-05)),(to_sfixed_a(0.0002144019235856831)),(to_sfixed_a(-6.359696999425068e-05)),(to_sfixed_a(0.0001942100061569363)),(to_sfixed_a(0.0001739030994940549)),(to_sfixed_a(0.00010377671424066648)),(to_sfixed_a(2.368481546000112e-05)),(to_sfixed_a(-1.4109253925198573e-06)),(to_sfixed_a(1.8909830032498576e-05)),(to_sfixed_a(-0.00026532483752816916)),(to_sfixed_a(7.791584835104004e-07)),(to_sfixed_a(1.278711533814203e-05)),(to_sfixed_a(-1.5807738236617297e-05)),(to_sfixed_a(0.00023398133635055274)),(to_sfixed_a(-7.964544784044847e-05)),(to_sfixed_a(3.890949301421642e-05)),(to_sfixed_a(9.531339310342446e-05)),(to_sfixed_a(-0.0001467960828449577)),(to_sfixed_a(-0.00011972014181083068)),(to_sfixed_a(0.00013444444630295038)),(to_sfixed_a(-2.7305184175929753e-06)),(to_sfixed_a(-0.06628350913524628)),(to_sfixed_a(-8.03021393949166e-05)),(to_sfixed_a(-0.07519406080245972)),(to_sfixed_a(0.02716020494699478)),(to_sfixed_a(-0.14844325184822083)),(to_sfixed_a(-0.06784029304981232)),(to_sfixed_a(-0.13426722586154938)),(to_sfixed_a(-0.22716403007507324)),(to_sfixed_a(-0.001996168401092291)),(to_sfixed_a(-0.18949873745441437)),(to_sfixed_a(-0.1761256903409958)),(to_sfixed_a(0.03986562043428421)),(to_sfixed_a(0.026597188785672188)),(to_sfixed_a(0.05390492081642151)),(to_sfixed_a(3.081826798734255e-05)),(to_sfixed_a(-6.636708712903783e-05)),(to_sfixed_a(0.00013568198482971638)),(to_sfixed_a(0.0001098618158721365)),(to_sfixed_a(3.4300719562452286e-05)),(to_sfixed_a(-7.207546786958119e-06)),(to_sfixed_a(-5.6012420827755705e-05)),(to_sfixed_a(-0.00018308611470274627)),(to_sfixed_a(-9.715613487060182e-06)),(to_sfixed_a(-8.001983951544389e-05)),(to_sfixed_a(-0.00013081527140457183)),(to_sfixed_a(1.2223150406498462e-05)),(to_sfixed_a(0.0004354129487182945)),(to_sfixed_a(0.06710074841976166)),(to_sfixed_a(0.017212051898241043)),(to_sfixed_a(-0.09553533792495728)),(to_sfixed_a(-0.28864479064941406)),(to_sfixed_a(-0.11351576447486877)),(to_sfixed_a(0.03186517208814621)),(to_sfixed_a(-0.011290116235613823)),(to_sfixed_a(-0.04136928915977478)),(to_sfixed_a(-0.22239834070205688)),(to_sfixed_a(-0.2876738905906677)),(to_sfixed_a(-0.21391288936138153)),(to_sfixed_a(-0.18356852233409882)),(to_sfixed_a(0.026877954602241516)),(to_sfixed_a(0.004520428366959095)),(to_sfixed_a(0.1340755969285965)),(to_sfixed_a(-0.028684815391898155)),(to_sfixed_a(2.9053060643491335e-05)),(to_sfixed_a(-0.0017246183706447482)),(to_sfixed_a(-1.3155810847820248e-05)),(to_sfixed_a(-0.00016542896628379822)),(to_sfixed_a(0.0004151111643295735)),(to_sfixed_a(-0.00024844022118486464)),(to_sfixed_a(-3.144993388559669e-05)),(to_sfixed_a(-2.988392225233838e-05)),(to_sfixed_a(-0.00032640082645229995)),(to_sfixed_a(-0.00012483976024668664)),(to_sfixed_a(0.1048799678683281)),(to_sfixed_a(0.00650067487731576)),(to_sfixed_a(0.15263251960277557)),(to_sfixed_a(-0.07836568355560303)),(to_sfixed_a(0.05589871481060982)),(to_sfixed_a(0.03340020775794983)),(to_sfixed_a(0.08673940598964691)),(to_sfixed_a(0.1405058652162552)),(to_sfixed_a(0.01018655113875866)),(to_sfixed_a(-0.19008885324001312)),(to_sfixed_a(-0.15788495540618896)),(to_sfixed_a(-0.02057344652712345)),(to_sfixed_a(-0.17148713767528534)),(to_sfixed_a(0.1717478334903717)),(to_sfixed_a(-0.11781208217144012)),(to_sfixed_a(-0.058880362659692764)),(to_sfixed_a(0.03000294789671898)),(to_sfixed_a(0.00015121788601391017)),(to_sfixed_a(0.03854374215006828)),(to_sfixed_a(0.00020224324543960392)),(to_sfixed_a(-6.86452112859115e-05)),(to_sfixed_a(0.00017151811334770173)),(to_sfixed_a(-0.00011688335507642478)),(to_sfixed_a(-7.395699867629446e-06)),(to_sfixed_a(-4.605237700161524e-05)),(to_sfixed_a(-9.441641304874793e-05)),(to_sfixed_a(-0.00017850750009529293)),(to_sfixed_a(0.0001257225521840155)),(to_sfixed_a(0.09728700667619705)),(to_sfixed_a(0.10161242634057999)),(to_sfixed_a(0.22272536158561707)),(to_sfixed_a(-0.028810255229473114)),(to_sfixed_a(0.28774622082710266)),(to_sfixed_a(0.1847473680973053)),(to_sfixed_a(0.24315230548381805)),(to_sfixed_a(-0.22987061738967896)),(to_sfixed_a(-0.26192787289619446)),(to_sfixed_a(-0.3745204508304596)),(to_sfixed_a(-0.21909105777740479)),(to_sfixed_a(-0.31420424580574036)),(to_sfixed_a(-0.15490375459194183)),(to_sfixed_a(-0.00013269425835460424)),(to_sfixed_a(0.09721539169549942)),(to_sfixed_a(0.1553577482700348)),(to_sfixed_a(-0.007500152103602886)),(to_sfixed_a(0.16053491830825806)),(to_sfixed_a(0.16013756394386292)),(to_sfixed_a(0.005739861633628607)),(to_sfixed_a(0.007314158137887716)),(to_sfixed_a(0.0029196348041296005)),(to_sfixed_a(3.7715035432484e-05)),(to_sfixed_a(-0.00010301032307324931)),(to_sfixed_a(1.767686626408249e-05)),(to_sfixed_a(-4.217536479700357e-05)),(to_sfixed_a(-9.891546505969018e-05)),(to_sfixed_a(-6.257511267904192e-05)),(to_sfixed_a(-0.009722785092890263)),(to_sfixed_a(0.13990312814712524)),(to_sfixed_a(-0.022303622215986252)),(to_sfixed_a(0.14036598801612854)),(to_sfixed_a(0.24167369306087494)),(to_sfixed_a(0.21583634614944458)),(to_sfixed_a(0.20461918413639069)),(to_sfixed_a(0.13321571052074432)),(to_sfixed_a(-0.18215711414813995)),(to_sfixed_a(-0.22624246776103973)),(to_sfixed_a(-0.2857722043991089)),(to_sfixed_a(-0.2515709698200226)),(to_sfixed_a(-0.057545892894268036)),(to_sfixed_a(-0.20052754878997803)),(to_sfixed_a(0.12370068579912186)),(to_sfixed_a(0.0764150321483612)),(to_sfixed_a(0.0994129329919815)),(to_sfixed_a(0.052968189120292664)),(to_sfixed_a(0.2793118953704834)),(to_sfixed_a(0.06802239269018173)),(to_sfixed_a(0.004234161227941513)),(to_sfixed_a(5.856405186932534e-05)),(to_sfixed_a(0.00017830760043580085)),(to_sfixed_a(0.0002457873779349029)),(to_sfixed_a(-0.000348409143043682)),(to_sfixed_a(0.00020054151536896825)),(to_sfixed_a(-7.323230965994298e-05)),(to_sfixed_a(0.022859051823616028)),(to_sfixed_a(0.10046364367008209)),(to_sfixed_a(-0.0672077015042305)),(to_sfixed_a(0.08130229264497757)),(to_sfixed_a(-0.2844485342502594)),(to_sfixed_a(0.32096609473228455)),(to_sfixed_a(0.38172873854637146)),(to_sfixed_a(-0.0117917750030756)),(to_sfixed_a(0.2211613804101944)),(to_sfixed_a(0.09595680236816406)),(to_sfixed_a(-0.21942991018295288)),(to_sfixed_a(-0.0036905757151544094)),(to_sfixed_a(-0.1370994597673416)),(to_sfixed_a(0.03970152884721756)),(to_sfixed_a(-0.0051795486360788345)),(to_sfixed_a(-0.13258036971092224)),(to_sfixed_a(0.012881665490567684)),(to_sfixed_a(-0.023324452340602875)),(to_sfixed_a(0.06695830076932907)),(to_sfixed_a(0.14361321926116943)),(to_sfixed_a(0.03191032260656357)),(to_sfixed_a(-0.004116765223443508)),(to_sfixed_a(-7.965503755258396e-05)),(to_sfixed_a(0.0001073412859113887)),(to_sfixed_a(-0.00010071729775518179)),(to_sfixed_a(-9.273592149838805e-05)),(to_sfixed_a(3.794855729211122e-05)),(to_sfixed_a(-0.0002962905855383724)),(to_sfixed_a(-0.0017632225062698126)),(to_sfixed_a(0.04173463210463524)),(to_sfixed_a(-0.003938326146453619)),(to_sfixed_a(0.219354048371315)),(to_sfixed_a(-0.08269061893224716)),(to_sfixed_a(0.05721672251820564)),(to_sfixed_a(0.18412624299526215)),(to_sfixed_a(0.43393170833587646)),(to_sfixed_a(0.0651182234287262)),(to_sfixed_a(-0.008093860000371933)),(to_sfixed_a(0.17825809121131897)),(to_sfixed_a(0.1572074443101883)),(to_sfixed_a(0.19417934119701385)),(to_sfixed_a(0.10684636235237122)),(to_sfixed_a(0.010338437743484974)),(to_sfixed_a(-0.5132634043693542)),(to_sfixed_a(-0.47977325320243835)),(to_sfixed_a(-0.11582665145397186)),(to_sfixed_a(0.14948689937591553)),(to_sfixed_a(-0.13118577003479004)),(to_sfixed_a(-0.11421211063861847)),(to_sfixed_a(-0.0002702937927097082)),(to_sfixed_a(-0.0001246201863978058)),(to_sfixed_a(0.00019931643328163773)),(to_sfixed_a(0.00016335588588844985)),(to_sfixed_a(-0.00017691087850835174)),(to_sfixed_a(-0.00023424097162205726)),(to_sfixed_a(0.00011964895384153351)),(to_sfixed_a(-0.009232636541128159)),(to_sfixed_a(-0.03653270751237869)),(to_sfixed_a(-0.334222674369812)),(to_sfixed_a(-0.13756412267684937)),(to_sfixed_a(-0.16610881686210632)),(to_sfixed_a(0.0655151978135109)),(to_sfixed_a(0.2676258683204651)),(to_sfixed_a(0.2861197590827942)),(to_sfixed_a(0.13366861641407013)),(to_sfixed_a(0.22553741931915283)),(to_sfixed_a(0.15472331643104553)),(to_sfixed_a(0.6115001440048218)),(to_sfixed_a(0.1747683733701706)),(to_sfixed_a(-0.005017354618757963)),(to_sfixed_a(-0.0738881304860115)),(to_sfixed_a(0.01524563878774643)),(to_sfixed_a(-0.07460997253656387)),(to_sfixed_a(-0.014751598238945007)),(to_sfixed_a(-0.2553575932979584)),(to_sfixed_a(0.058139268308877945)),(to_sfixed_a(-0.03552105650305748)),(to_sfixed_a(0.004499774891883135)),(to_sfixed_a(3.825437670457177e-05)),(to_sfixed_a(-7.582108810311183e-05)),(to_sfixed_a(2.7935358957620338e-05)),(to_sfixed_a(-0.00014776209718547761)),(to_sfixed_a(-0.00025930022820830345)),(to_sfixed_a(0.002585100941359997)),(to_sfixed_a(0.011875614523887634)),(to_sfixed_a(-0.19025765359401703)),(to_sfixed_a(-0.13188768923282623)),(to_sfixed_a(-0.21994644403457642)),(to_sfixed_a(-0.2019820511341095)),(to_sfixed_a(-0.2559976577758789)),(to_sfixed_a(-0.03522372618317604)),(to_sfixed_a(0.01225259155035019)),(to_sfixed_a(0.2858317792415619)),(to_sfixed_a(0.32732445001602173)),(to_sfixed_a(0.033076707273721695)),(to_sfixed_a(0.16743114590644836)),(to_sfixed_a(0.08252071589231491)),(to_sfixed_a(-0.06817495822906494)),(to_sfixed_a(-0.09100460261106491)),(to_sfixed_a(0.08247554302215576)),(to_sfixed_a(0.047383859753608704)),(to_sfixed_a(-0.06118317320942879)),(to_sfixed_a(-0.05484267696738243)),(to_sfixed_a(-0.1016397625207901)),(to_sfixed_a(-0.13048849999904633)),(to_sfixed_a(5.074434284324525e-06)),(to_sfixed_a(9.515867714071646e-05)),(to_sfixed_a(-0.00029239131254144013)),(to_sfixed_a(5.821839749842184e-06)),(to_sfixed_a(4.490706851356663e-05)),(to_sfixed_a(-0.000203198374947533)),(to_sfixed_a(0.00038326423964463174)),(to_sfixed_a(0.030787639319896698)),(to_sfixed_a(-0.12338947504758835)),(to_sfixed_a(-0.25267601013183594)),(to_sfixed_a(-0.21268367767333984)),(to_sfixed_a(-0.1598798632621765)),(to_sfixed_a(-0.22805388271808624)),(to_sfixed_a(0.016458362340927124)),(to_sfixed_a(0.5730329155921936)),(to_sfixed_a(0.7484021782875061)),(to_sfixed_a(0.252060204744339)),(to_sfixed_a(0.14754757285118103)),(to_sfixed_a(0.4641721546649933)),(to_sfixed_a(-0.18546873331069946)),(to_sfixed_a(0.12029232084751129)),(to_sfixed_a(0.07617378979921341)),(to_sfixed_a(0.24736982583999634)),(to_sfixed_a(0.18676066398620605)),(to_sfixed_a(-0.07808005809783936)),(to_sfixed_a(-0.03432377055287361)),(to_sfixed_a(0.015449500642716885)),(to_sfixed_a(-0.26924630999565125)),(to_sfixed_a(1.0609850505716167e-05)),(to_sfixed_a(-0.00017844045942183584)),(to_sfixed_a(-7.066460239002481e-05)),(to_sfixed_a(-0.0001594577042851597)),(to_sfixed_a(-1.313404573011212e-05)),(to_sfixed_a(-9.927220162353478e-06)),(to_sfixed_a(-0.00012856628745794296)),(to_sfixed_a(-0.055832043290138245)),(to_sfixed_a(-0.1352829784154892)),(to_sfixed_a(-0.21340225636959076)),(to_sfixed_a(-0.24742832779884338)),(to_sfixed_a(-0.1553952991962433)),(to_sfixed_a(0.07094339281320572)),(to_sfixed_a(0.16340309381484985)),(to_sfixed_a(0.3377993702888489)),(to_sfixed_a(0.18695074319839478)),(to_sfixed_a(0.07199787348508835)),(to_sfixed_a(-0.25044533610343933)),(to_sfixed_a(0.04077170044183731)),(to_sfixed_a(0.09824378043413162)),(to_sfixed_a(0.1720060557126999)),(to_sfixed_a(0.16424858570098877)),(to_sfixed_a(0.2881369888782501)),(to_sfixed_a(0.1390152871608734)),(to_sfixed_a(-0.2051832377910614)),(to_sfixed_a(-0.06589248031377792)),(to_sfixed_a(-0.5295949578285217)),(to_sfixed_a(-0.08259282261133194)),(to_sfixed_a(0.0012682428350672126)),(to_sfixed_a(-0.0005890766624361277)),(to_sfixed_a(4.834908395423554e-05)),(to_sfixed_a(0.00013099968782626092)),(to_sfixed_a(-5.8378547691972926e-05)),(to_sfixed_a(-0.00025679171085357666)),(to_sfixed_a(-5.971292921458371e-05)),(to_sfixed_a(-0.00038278003921732306)),(to_sfixed_a(-0.05668637901544571)),(to_sfixed_a(-0.00922379270195961)),(to_sfixed_a(-0.07137603312730789)),(to_sfixed_a(-0.23005187511444092)),(to_sfixed_a(-0.076291024684906)),(to_sfixed_a(-0.04828176274895668)),(to_sfixed_a(-0.032992515712976456)),(to_sfixed_a(-0.005786743480712175)),(to_sfixed_a(-0.2237757444381714)),(to_sfixed_a(0.11780238896608353)),(to_sfixed_a(0.1839960217475891)),(to_sfixed_a(-0.0009790584444999695)),(to_sfixed_a(0.060652509331703186)),(to_sfixed_a(0.05983293429017067)),(to_sfixed_a(-0.008571195416152477)),(to_sfixed_a(0.00857485830783844)),(to_sfixed_a(-0.08436943590641022)),(to_sfixed_a(-0.18458260595798492)),(to_sfixed_a(-0.20834627747535706)),(to_sfixed_a(0.07888149470090866)),(to_sfixed_a(0.0010505671380087733)),(to_sfixed_a(9.554539701639442e-07)),(to_sfixed_a(0.00024211895652115345)),(to_sfixed_a(0.00018890960200224072)),(to_sfixed_a(0.0002851221652235836)),(to_sfixed_a(-5.5535360843350645e-06)),(to_sfixed_a(-1.7247542928089388e-05)),(to_sfixed_a(-0.06738971173763275)),(to_sfixed_a(-0.08262936770915985)),(to_sfixed_a(0.07567203044891357)),(to_sfixed_a(-0.1622130423784256)),(to_sfixed_a(-0.2882448136806488)),(to_sfixed_a(-0.00144993606954813)),(to_sfixed_a(-0.230687215924263)),(to_sfixed_a(-0.09004874527454376)),(to_sfixed_a(-0.05527316778898239)),(to_sfixed_a(-0.08797747641801834)),(to_sfixed_a(0.13366778194904327)),(to_sfixed_a(0.07574272155761719)),(to_sfixed_a(0.28406408429145813)),(to_sfixed_a(-0.24424853920936584)),(to_sfixed_a(-0.07208602130413055)),(to_sfixed_a(0.008527683094143867)),(to_sfixed_a(-0.11830053478479385)),(to_sfixed_a(-0.019780246540904045)),(to_sfixed_a(-0.11691741645336151)),(to_sfixed_a(-0.03370356932282448)),(to_sfixed_a(-0.1115521788597107)),(to_sfixed_a(0.0011288393288850784)),(to_sfixed_a(0.0001512879243819043)),(to_sfixed_a(0.00027637151652015746)),(to_sfixed_a(-2.4491866497555748e-05)),(to_sfixed_a(-0.0001023057266138494)),(to_sfixed_a(3.659549474832602e-05)),(to_sfixed_a(-0.003943756688386202)),(to_sfixed_a(0.1422075629234314)),(to_sfixed_a(0.17193035781383514)),(to_sfixed_a(0.40021923184394836)),(to_sfixed_a(-0.0650620386004448)),(to_sfixed_a(0.14553841948509216)),(to_sfixed_a(-0.2852266728878021)),(to_sfixed_a(-0.09368076175451279)),(to_sfixed_a(-0.10973310470581055)),(to_sfixed_a(0.08694259822368622)),(to_sfixed_a(0.0018107234500348568)),(to_sfixed_a(-0.04816266894340515)),(to_sfixed_a(0.0338122732937336)),(to_sfixed_a(0.21867839992046356)),(to_sfixed_a(-0.02403610199689865)),(to_sfixed_a(-0.21442586183547974)),(to_sfixed_a(-0.08481840789318085)),(to_sfixed_a(0.06375360488891602)),(to_sfixed_a(0.22953161597251892)),(to_sfixed_a(0.042314622551202774)),(to_sfixed_a(-0.012859736569225788)),(to_sfixed_a(-0.10652262717485428)),(to_sfixed_a(-0.011145119555294514)),(to_sfixed_a(-0.00012113878619857132)),(to_sfixed_a(-5.79071493120864e-05)),(to_sfixed_a(7.097137859091163e-05)),(to_sfixed_a(-7.923951670818496e-06)),(to_sfixed_a(-0.0030577434226870537)),(to_sfixed_a(-0.003928746562451124)),(to_sfixed_a(-0.09335244446992874)),(to_sfixed_a(0.16769008338451385)),(to_sfixed_a(0.14026705920696259)),(to_sfixed_a(-0.06951839476823807)),(to_sfixed_a(-0.18776780366897583)),(to_sfixed_a(-0.08519066870212555)),(to_sfixed_a(0.014190074056386948)),(to_sfixed_a(0.116803839802742)),(to_sfixed_a(0.3084527552127838)),(to_sfixed_a(0.06805213540792465)),(to_sfixed_a(0.09779108315706253)),(to_sfixed_a(0.48380813002586365)),(to_sfixed_a(-0.07348808646202087)),(to_sfixed_a(0.003223937703296542)),(to_sfixed_a(-0.06099072843790054)),(to_sfixed_a(-0.1785462200641632)),(to_sfixed_a(0.1549682766199112)),(to_sfixed_a(-0.1176946610212326)),(to_sfixed_a(-0.06080075353384018)),(to_sfixed_a(0.05064665153622627)),(to_sfixed_a(0.0001499462523497641)),(to_sfixed_a(-9.834732736635488e-06)),(to_sfixed_a(-0.00010247150203213096)),(to_sfixed_a(0.00011283477215329185)),(to_sfixed_a(2.7475158276502043e-05)),(to_sfixed_a(-0.00013413088163360953)),(to_sfixed_a(0.00025503928191028535)),(to_sfixed_a(-0.016237106174230576)),(to_sfixed_a(-0.11888085305690765)),(to_sfixed_a(-0.0931512862443924)),(to_sfixed_a(-0.17848174273967743)),(to_sfixed_a(-0.008449180983006954)),(to_sfixed_a(-0.11761193722486496)),(to_sfixed_a(-0.2138538807630539)),(to_sfixed_a(-0.07267707586288452)),(to_sfixed_a(0.3281041383743286)),(to_sfixed_a(0.6330446600914001)),(to_sfixed_a(0.16337649524211884)),(to_sfixed_a(0.19462719559669495)),(to_sfixed_a(0.05443895608186722)),(to_sfixed_a(-0.02296900935471058)),(to_sfixed_a(-0.30186179280281067)),(to_sfixed_a(-0.024714410305023193)),(to_sfixed_a(-0.13666628301143646)),(to_sfixed_a(0.025072887539863586)),(to_sfixed_a(0.19573339819908142)),(to_sfixed_a(0.13958074152469635)),(to_sfixed_a(-0.10532449185848236)),(to_sfixed_a(0.0017350066918879747)),(to_sfixed_a(7.859921606723219e-05)),(to_sfixed_a(2.7977600893791532e-06)),(to_sfixed_a(0.00025615940103307366)),(to_sfixed_a(-3.303156699985266e-05)),(to_sfixed_a(-0.0001739698345772922)),(to_sfixed_a(0.00035927107091993093)),(to_sfixed_a(0.03775791823863983)),(to_sfixed_a(0.0004069598508067429)),(to_sfixed_a(0.1129334419965744)),(to_sfixed_a(-0.10186667740345001)),(to_sfixed_a(-0.15386953949928284)),(to_sfixed_a(-0.309194952249527)),(to_sfixed_a(-0.1966647505760193)),(to_sfixed_a(-0.07531904429197311)),(to_sfixed_a(0.08784741163253784)),(to_sfixed_a(0.25093960762023926)),(to_sfixed_a(0.2734586298465729)),(to_sfixed_a(0.10694007575511932)),(to_sfixed_a(0.027129851281642914)),(to_sfixed_a(-0.20935742557048798)),(to_sfixed_a(-0.3796011507511139)),(to_sfixed_a(-0.10172347724437714)),(to_sfixed_a(0.10304161161184311)),(to_sfixed_a(-0.03652633726596832)),(to_sfixed_a(0.06414084136486053)),(to_sfixed_a(0.16291171312332153)),(to_sfixed_a(0.09946173429489136)),(to_sfixed_a(5.443831469165161e-05)),(to_sfixed_a(2.7724456231226213e-05)),(to_sfixed_a(0.0001438419276382774)),(to_sfixed_a(-9.599774784874171e-05)),(to_sfixed_a(1.897261790873017e-05)),(to_sfixed_a(0.00012951232201885432)),(to_sfixed_a(0.00018367846496403217)),(to_sfixed_a(0.00013815093552693725)),(to_sfixed_a(-0.009696213528513908)),(to_sfixed_a(0.026735816150903702)),(to_sfixed_a(0.15930664539337158)),(to_sfixed_a(-0.4013141095638275)),(to_sfixed_a(-0.068287692964077)),(to_sfixed_a(-0.2165970355272293)),(to_sfixed_a(-0.15541404485702515)),(to_sfixed_a(0.14361342787742615)),(to_sfixed_a(0.48401695489883423)),(to_sfixed_a(-0.03748002275824547)),(to_sfixed_a(-0.03626241907477379)),(to_sfixed_a(-0.05129125341773033)),(to_sfixed_a(0.029741613194346428)),(to_sfixed_a(-0.04457923769950867)),(to_sfixed_a(0.10857369005680084)),(to_sfixed_a(0.14514006674289703)),(to_sfixed_a(0.22748129069805145)),(to_sfixed_a(0.14792633056640625)),(to_sfixed_a(-0.02079327590763569)),(to_sfixed_a(-0.028390413150191307)),(to_sfixed_a(0.020506905391812325)),(to_sfixed_a(-0.0001082267626770772)),(to_sfixed_a(-0.00016725943714845926)),(to_sfixed_a(-0.00030942645389586687)),(to_sfixed_a(-0.000279218889772892)),(to_sfixed_a(0.0001658398687141016)),(to_sfixed_a(-4.9436759582022205e-05)),(to_sfixed_a(-0.0003161186177749187)),(to_sfixed_a(-0.03873346745967865)),(to_sfixed_a(-0.0009004962048493326)),(to_sfixed_a(-0.21115736663341522)),(to_sfixed_a(-0.2397466003894806)),(to_sfixed_a(-0.25571727752685547)),(to_sfixed_a(-0.10637222230434418)),(to_sfixed_a(-0.01548463199287653)),(to_sfixed_a(-0.007687679026275873)),(to_sfixed_a(-0.018894903361797333)),(to_sfixed_a(-0.0751664787530899)),(to_sfixed_a(0.15423651039600372)),(to_sfixed_a(-0.05049661174416542)),(to_sfixed_a(-0.14310164749622345)),(to_sfixed_a(-0.23335060477256775)),(to_sfixed_a(0.14083698391914368)),(to_sfixed_a(0.015188725665211678)),(to_sfixed_a(-0.1055726632475853)),(to_sfixed_a(-0.03246096894145012)),(to_sfixed_a(0.024204622954130173)),(to_sfixed_a(-0.0005629210500046611)),(to_sfixed_a(-0.0916208028793335)),(to_sfixed_a(0.00022017092851456255)),(to_sfixed_a(0.0001813996786950156)),(to_sfixed_a(4.054534656461328e-05)),(to_sfixed_a(-6.641964137088507e-05)),(to_sfixed_a(-0.00017114220827352256)),(to_sfixed_a(-4.890747004537843e-05)),(to_sfixed_a(-4.2068040784215555e-05)),(to_sfixed_a(0.0003577310126274824)),(to_sfixed_a(-0.010447410866618156)),(to_sfixed_a(-0.029529057443141937)),(to_sfixed_a(0.105067677795887)),(to_sfixed_a(0.04301841929554939)),(to_sfixed_a(0.12890473008155823)),(to_sfixed_a(-0.041807107627391815)),(to_sfixed_a(0.09293638914823532)),(to_sfixed_a(0.0831177830696106)),(to_sfixed_a(0.1268927901983261)),(to_sfixed_a(0.23137551546096802)),(to_sfixed_a(0.17466139793395996)),(to_sfixed_a(-0.025936361402273178)),(to_sfixed_a(-0.02516341395676136)),(to_sfixed_a(0.10796858370304108)),(to_sfixed_a(0.08572211861610413)),(to_sfixed_a(-0.06466878950595856)),(to_sfixed_a(-0.021852383390069008)),(to_sfixed_a(-0.1355714350938797)),(to_sfixed_a(0.004769318737089634)),(to_sfixed_a(5.1893730415031314e-05)),(to_sfixed_a(-1.3802139619656373e-05)),(to_sfixed_a(5.160936416359618e-05)),(to_sfixed_a(1.0574569387244992e-05)),(to_sfixed_a(0.00018993399862665683)),(to_sfixed_a(-4.081437873537652e-05)),(to_sfixed_a(0.0003084289492107928)),(to_sfixed_a(3.682590613607317e-05)),(to_sfixed_a(0.00046937758452259004)),(to_sfixed_a(0.00487591652199626)),(to_sfixed_a(-0.033422693610191345)),(to_sfixed_a(0.17183592915534973)),(to_sfixed_a(0.15789954364299774)),(to_sfixed_a(0.07514937222003937)),(to_sfixed_a(0.01517408899962902)),(to_sfixed_a(0.05848877504467964)),(to_sfixed_a(0.25366103649139404)),(to_sfixed_a(0.023850610479712486)),(to_sfixed_a(0.3324345350265503)),(to_sfixed_a(0.25718238949775696)),(to_sfixed_a(0.3937578499317169)),(to_sfixed_a(0.26201164722442627)),(to_sfixed_a(0.02612266130745411)),(to_sfixed_a(0.0894404873251915)),(to_sfixed_a(0.1160254254937172)),(to_sfixed_a(-0.06781678646802902)),(to_sfixed_a(0.008586962707340717)),(to_sfixed_a(-0.051740966737270355)),(to_sfixed_a(-9.6799289167393e-05)),(to_sfixed_a(-0.0003100686299148947)),(to_sfixed_a(-0.0001646825548959896)),(to_sfixed_a(-8.60646614455618e-05)),(to_sfixed_a(0.00014570220082532614)),(to_sfixed_a(6.706963904434815e-05)),(to_sfixed_a(-5.556788528338075e-05)),(to_sfixed_a(4.727095802081749e-05)),(to_sfixed_a(-0.010754546150565147)),(to_sfixed_a(0.007517751771956682)),(to_sfixed_a(-0.04553305730223656)),(to_sfixed_a(0.05512438714504242)),(to_sfixed_a(0.10820744186639786)),(to_sfixed_a(0.013822878710925579)),(to_sfixed_a(0.1680297702550888)),(to_sfixed_a(0.07695210725069046)),(to_sfixed_a(0.11786060035228729)),(to_sfixed_a(0.552239179611206)),(to_sfixed_a(0.2754490375518799)),(to_sfixed_a(0.11531971395015717)),(to_sfixed_a(0.006594976410269737)),(to_sfixed_a(-0.13996466994285583)),(to_sfixed_a(0.003925208002328873)),(to_sfixed_a(0.030274417251348495)),(to_sfixed_a(0.005913387052714825)),(to_sfixed_a(-0.07617270946502686)),(to_sfixed_a(-0.022258970886468887)),(to_sfixed_a(0.006059560924768448)),(to_sfixed_a(-5.395602056523785e-05)),(to_sfixed_a(0.0002177284623030573)),(to_sfixed_a(9.732862235978246e-05)),(to_sfixed_a(0.00015539587184321135)),(to_sfixed_a(6.247369310585782e-05)),(to_sfixed_a(9.128200326813385e-05)),(to_sfixed_a(-0.00021428077889140695)),(to_sfixed_a(7.006759551586583e-05)),(to_sfixed_a(0.00011313112918287516)),(to_sfixed_a(0.023806998506188393)),(to_sfixed_a(-0.026578206568956375)),(to_sfixed_a(-0.06479146331548691)),(to_sfixed_a(0.11733387410640717)),(to_sfixed_a(0.007128132041543722)),(to_sfixed_a(-0.07861928641796112)),(to_sfixed_a(0.028717726469039917)),(to_sfixed_a(-0.054030731320381165)),(to_sfixed_a(-0.07508984208106995)),(to_sfixed_a(0.10900504887104034)),(to_sfixed_a(0.09480427205562592)),(to_sfixed_a(-0.002267414005473256)),(to_sfixed_a(-0.03520909324288368)),(to_sfixed_a(-0.00319239916279912)),(to_sfixed_a(-0.019060330465435982)),(to_sfixed_a(-0.12710873782634735)),(to_sfixed_a(-0.0003943062329199165)),(to_sfixed_a(-0.00047904462553560734)),(to_sfixed_a(-0.00020921842951793224)),(to_sfixed_a(-9.137974120676517e-05)),(to_sfixed_a(8.491324479109608e-07)),(to_sfixed_a(-0.00013502055662684143)),(to_sfixed_a(0.00024205366207752377)),(to_sfixed_a(-5.424918344942853e-05)),(to_sfixed_a(7.813535921741277e-05)),(to_sfixed_a(-0.00012794385838788003)),(to_sfixed_a(4.392234041006304e-05)),(to_sfixed_a(4.8465848522027954e-05)),(to_sfixed_a(-0.0002327391557628289)),(to_sfixed_a(3.6898265534546226e-05)),(to_sfixed_a(-1.0545018085394986e-05)),(to_sfixed_a(0.00013784883776679635)),(to_sfixed_a(0.0005431267782114446)),(to_sfixed_a(0.020850377157330513)),(to_sfixed_a(-0.0040346295572817326)),(to_sfixed_a(-0.0027432593051344156)),(to_sfixed_a(0.013308536261320114)),(to_sfixed_a(-0.08174148201942444)),(to_sfixed_a(0.002498057670891285)),(to_sfixed_a(-0.04173076152801514)),(to_sfixed_a(0.019984368234872818)),(to_sfixed_a(0.017360424622893333)),(to_sfixed_a(-0.011884892359375954)),(to_sfixed_a(-0.006150494795292616)),(to_sfixed_a(0.00014856822963338345)),(to_sfixed_a(0.0001040742572513409)),(to_sfixed_a(-8.652321412228048e-05)),(to_sfixed_a(0.00015366001753136516)),(to_sfixed_a(0.0001796973228920251)),(to_sfixed_a(6.483001925516874e-05)),(to_sfixed_a(-0.0001707014162093401)),(to_sfixed_a(-0.00014953433128539473)),(to_sfixed_a(-0.0001298821734962985)),(to_sfixed_a(8.39170825202018e-05)),(to_sfixed_a(4.655838347389363e-05)),(to_sfixed_a(-1.983973561436869e-06)),(to_sfixed_a(-8.716784213902429e-05)),(to_sfixed_a(-1.5068077118485235e-05)),(to_sfixed_a(0.00033884719596244395)),(to_sfixed_a(5.9327758208382875e-06)),(to_sfixed_a(-0.00017667561769485474)),(to_sfixed_a(0.0002629747032187879)),(to_sfixed_a(-2.4088598365779035e-05)),(to_sfixed_a(9.814702207222581e-05)),(to_sfixed_a(0.00027933728415519)),(to_sfixed_a(0.0003751229669433087)),(to_sfixed_a(-0.00015544284542556852)),(to_sfixed_a(-4.867911047767848e-05)),(to_sfixed_a(-1.3511137694877107e-05)),(to_sfixed_a(0.0001522799429949373)),(to_sfixed_a(-4.722238008980639e-05)),(to_sfixed_a(-0.00014972723147366196)),(to_sfixed_a(-0.0003722121473401785)),(to_sfixed_a(-0.00020469834271352738)),(to_sfixed_a(-4.707526386482641e-05)),(to_sfixed_a(2.599554500193335e-05)),(to_sfixed_a(0.0002984464808832854)),(to_sfixed_a(4.081410224898718e-05)),(to_sfixed_a(-0.00022382871247828007)));

    constant weight_n0_16 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(6.254162144614384e-05)),(to_sfixed_a(0.00019014028657693416)),(to_sfixed_a(-4.364584128779825e-06)),(to_sfixed_a(-1.4251058018999174e-05)),(to_sfixed_a(0.0001811254769563675)),(to_sfixed_a(1.5980047010089038e-06)),(to_sfixed_a(-4.9276255595032126e-05)),(to_sfixed_a(-0.00024418835528194904)),(to_sfixed_a(0.0001832517154980451)),(to_sfixed_a(-0.0001691002253210172)),(to_sfixed_a(7.326577906496823e-05)),(to_sfixed_a(9.869493806036189e-05)),(to_sfixed_a(-4.806050128536299e-06)),(to_sfixed_a(-0.00013347227650228888)),(to_sfixed_a(6.651288913417375e-06)),(to_sfixed_a(-4.749946674564853e-05)),(to_sfixed_a(-0.00021584464411716908)),(to_sfixed_a(-0.00023632991360500455)),(to_sfixed_a(0.00023353211872745305)),(to_sfixed_a(4.3330488551873714e-05)),(to_sfixed_a(0.00019163724209647626)),(to_sfixed_a(0.0002027191367233172)),(to_sfixed_a(-2.1495048713404685e-05)),(to_sfixed_a(-4.1280349250882864e-05)),(to_sfixed_a(-9.530180250294507e-05)),(to_sfixed_a(-4.338304279372096e-05)),(to_sfixed_a(1.0500746611796785e-05)),(to_sfixed_a(-0.00026539916871115565)),(to_sfixed_a(-6.629528070334345e-05)),(to_sfixed_a(-8.791632717475295e-05)),(to_sfixed_a(6.565712828887627e-05)),(to_sfixed_a(-0.0002065422886516899)),(to_sfixed_a(-8.268922101706266e-06)),(to_sfixed_a(7.233724318211898e-05)),(to_sfixed_a(-0.00020153980585746467)),(to_sfixed_a(6.293781916610897e-05)),(to_sfixed_a(5.3219744586385787e-05)),(to_sfixed_a(0.0001130243472289294)),(to_sfixed_a(0.00018292640743311495)),(to_sfixed_a(-0.00012025002797599882)),(to_sfixed_a(1.969633376575075e-05)),(to_sfixed_a(-0.00012553493434097618)),(to_sfixed_a(-2.7304917239234783e-05)),(to_sfixed_a(-0.00024358794325962663)),(to_sfixed_a(6.194857996888459e-05)),(to_sfixed_a(-6.273754115682095e-05)),(to_sfixed_a(-0.0001049892307491973)),(to_sfixed_a(0.0002832365280482918)),(to_sfixed_a(0.0001235345407621935)),(to_sfixed_a(-0.00014165241736918688)),(to_sfixed_a(8.640961459605023e-05)),(to_sfixed_a(-7.257259130710736e-05)),(to_sfixed_a(0.00010086205293191597)),(to_sfixed_a(0.0001510808215243742)),(to_sfixed_a(8.607663767179474e-05)),(to_sfixed_a(-0.00020969223987776786)),(to_sfixed_a(-3.478656435618177e-05)),(to_sfixed_a(-3.359696620464092e-06)),(to_sfixed_a(-9.949019840860274e-06)),(to_sfixed_a(5.698594031855464e-05)),(to_sfixed_a(-5.625392077490687e-06)),(to_sfixed_a(-9.442429291084409e-05)),(to_sfixed_a(6.837724504293874e-05)),(to_sfixed_a(-2.505264319552225e-06)),(to_sfixed_a(-0.0001950692676473409)),(to_sfixed_a(0.00016776513075456023)),(to_sfixed_a(-6.735949864378199e-05)),(to_sfixed_a(-4.411000190884806e-05)),(to_sfixed_a(7.862699931138195e-06)),(to_sfixed_a(-0.006433446425944567)),(to_sfixed_a(3.03573197015794e-05)),(to_sfixed_a(5.030279862694442e-05)),(to_sfixed_a(0.00011524741421453655)),(to_sfixed_a(-2.5736662792041898e-05)),(to_sfixed_a(0.0001454704615753144)),(to_sfixed_a(-7.28668601368554e-05)),(to_sfixed_a(0.0001923637028085068)),(to_sfixed_a(0.00020141751156188548)),(to_sfixed_a(0.0001270719658350572)),(to_sfixed_a(0.00017555523663759232)),(to_sfixed_a(-0.0002738412586040795)),(to_sfixed_a(-1.847199564508628e-05)),(to_sfixed_a(-1.2320864698267542e-05)),(to_sfixed_a(-0.0002792907471302897)),(to_sfixed_a(0.00010389649105491117)),(to_sfixed_a(-0.0002087840111926198)),(to_sfixed_a(0.00010633826605044305)),(to_sfixed_a(-6.67239601170877e-06)),(to_sfixed_a(8.212629472836852e-05)),(to_sfixed_a(-3.693962571560405e-05)),(to_sfixed_a(-2.537027648941148e-05)),(to_sfixed_a(-0.0002837029460351914)),(to_sfixed_a(-0.023449242115020752)),(to_sfixed_a(-3.806845052167773e-05)),(to_sfixed_a(-0.02673826925456524)),(to_sfixed_a(-0.07687930762767792)),(to_sfixed_a(-0.050772882997989655)),(to_sfixed_a(-0.09612124413251877)),(to_sfixed_a(-0.07260142266750336)),(to_sfixed_a(-0.1441880315542221)),(to_sfixed_a(-0.007106977980583906)),(to_sfixed_a(-0.14823904633522034)),(to_sfixed_a(-0.09972860664129257)),(to_sfixed_a(0.035803891718387604)),(to_sfixed_a(0.027070187032222748)),(to_sfixed_a(0.05481398478150368)),(to_sfixed_a(1.3949444337413297e-06)),(to_sfixed_a(0.00012584605428855866)),(to_sfixed_a(2.1973459297441877e-05)),(to_sfixed_a(-0.00013649981701746583)),(to_sfixed_a(0.0002362007217016071)),(to_sfixed_a(0.0001719989813864231)),(to_sfixed_a(0.0001106414056266658)),(to_sfixed_a(-8.068107126746327e-05)),(to_sfixed_a(0.00016857561422511935)),(to_sfixed_a(4.7765024646651e-05)),(to_sfixed_a(0.00012995324505027384)),(to_sfixed_a(3.2507516152691096e-05)),(to_sfixed_a(-0.0012365368893370032)),(to_sfixed_a(-0.025502804666757584)),(to_sfixed_a(-0.08012399822473526)),(to_sfixed_a(-0.03300488367676735)),(to_sfixed_a(-0.04623265191912651)),(to_sfixed_a(-0.1644248217344284)),(to_sfixed_a(-0.14543013274669647)),(to_sfixed_a(-0.26804402470588684)),(to_sfixed_a(-0.03884771093726158)),(to_sfixed_a(-0.052609823644161224)),(to_sfixed_a(0.07007487118244171)),(to_sfixed_a(0.27536797523498535)),(to_sfixed_a(-0.01770796999335289)),(to_sfixed_a(0.029459098353981972)),(to_sfixed_a(0.0010701996507123113)),(to_sfixed_a(0.19263765215873718)),(to_sfixed_a(0.0011966059682890773)),(to_sfixed_a(-0.00011631631787167862)),(to_sfixed_a(-0.0017513877246528864)),(to_sfixed_a(-1.5892890132818138e-06)),(to_sfixed_a(0.00012569595128297806)),(to_sfixed_a(-0.0002387201093370095)),(to_sfixed_a(-0.0004165805294178426)),(to_sfixed_a(6.355662480928004e-05)),(to_sfixed_a(-7.072980224620551e-05)),(to_sfixed_a(-0.00014603356248699129)),(to_sfixed_a(0.0012621113564819098)),(to_sfixed_a(-0.0067915357649326324)),(to_sfixed_a(0.02208859845995903)),(to_sfixed_a(0.000820688612293452)),(to_sfixed_a(-0.09034483134746552)),(to_sfixed_a(0.08492932468652725)),(to_sfixed_a(0.14571094512939453)),(to_sfixed_a(-0.10964136570692062)),(to_sfixed_a(-0.3465203642845154)),(to_sfixed_a(-0.1304212361574173)),(to_sfixed_a(-0.11239432543516159)),(to_sfixed_a(-0.1524820327758789)),(to_sfixed_a(0.20755434036254883)),(to_sfixed_a(0.1816985160112381)),(to_sfixed_a(0.2951647937297821)),(to_sfixed_a(-0.1428321748971939)),(to_sfixed_a(-0.06943289190530777)),(to_sfixed_a(0.12886199355125427)),(to_sfixed_a(-0.006946744862943888)),(to_sfixed_a(0.04776662960648537)),(to_sfixed_a(-0.005157326813787222)),(to_sfixed_a(-0.0006053042598068714)),(to_sfixed_a(4.331310265115462e-05)),(to_sfixed_a(0.00022903541685082018)),(to_sfixed_a(-1.261086708836956e-05)),(to_sfixed_a(-8.247227378888056e-05)),(to_sfixed_a(4.0847447962732986e-05)),(to_sfixed_a(-0.00010466740786796436)),(to_sfixed_a(-0.00012489722575992346)),(to_sfixed_a(-0.013695843517780304)),(to_sfixed_a(-0.058792658150196075)),(to_sfixed_a(0.1884448528289795)),(to_sfixed_a(0.23214952647686005)),(to_sfixed_a(-0.015219037421047688)),(to_sfixed_a(-0.0287304874509573)),(to_sfixed_a(-0.0020186484325677156)),(to_sfixed_a(-0.012356508523225784)),(to_sfixed_a(-0.19274353981018066)),(to_sfixed_a(-0.15098749101161957)),(to_sfixed_a(-0.21622464060783386)),(to_sfixed_a(-0.135801300406456)),(to_sfixed_a(0.05090642347931862)),(to_sfixed_a(0.2233435958623886)),(to_sfixed_a(0.20112960040569305)),(to_sfixed_a(0.2160213142633438)),(to_sfixed_a(0.09643924981355667)),(to_sfixed_a(0.2385159432888031)),(to_sfixed_a(0.23930546641349792)),(to_sfixed_a(-0.0004875557206105441)),(to_sfixed_a(-0.0008382605155929923)),(to_sfixed_a(0.002592592965811491)),(to_sfixed_a(0.0002063932770397514)),(to_sfixed_a(0.00032952456967905164)),(to_sfixed_a(-0.0002923810970969498)),(to_sfixed_a(5.012888664168713e-07)),(to_sfixed_a(0.00010322596062906086)),(to_sfixed_a(-0.00029158475808799267)),(to_sfixed_a(-0.042704831808805466)),(to_sfixed_a(0.021626895293593407)),(to_sfixed_a(-0.23852023482322693)),(to_sfixed_a(0.07893447577953339)),(to_sfixed_a(0.15217141807079315)),(to_sfixed_a(0.42820268869400024)),(to_sfixed_a(0.04863078519701958)),(to_sfixed_a(0.006448162253946066)),(to_sfixed_a(-0.4056808054447174)),(to_sfixed_a(-0.1984526515007019)),(to_sfixed_a(-0.08337754011154175)),(to_sfixed_a(0.16867852210998535)),(to_sfixed_a(-0.07382237166166306)),(to_sfixed_a(0.02740524336695671)),(to_sfixed_a(0.19150301814079285)),(to_sfixed_a(-0.26122307777404785)),(to_sfixed_a(0.16391950845718384)),(to_sfixed_a(0.14835944771766663)),(to_sfixed_a(-0.04402891919016838)),(to_sfixed_a(0.10509628802537918)),(to_sfixed_a(0.00357057130895555)),(to_sfixed_a(0.00021893304074183106)),(to_sfixed_a(-1.3655620932695456e-05)),(to_sfixed_a(0.00015881411673035473)),(to_sfixed_a(1.2000780770904385e-05)),(to_sfixed_a(-6.387002031260636e-06)),(to_sfixed_a(-0.00010173172631766647)),(to_sfixed_a(-0.06825251132249832)),(to_sfixed_a(0.07019972056150436)),(to_sfixed_a(-0.17161215841770172)),(to_sfixed_a(0.08336413651704788)),(to_sfixed_a(-0.09626500308513641)),(to_sfixed_a(0.2108408510684967)),(to_sfixed_a(-0.013530408963561058)),(to_sfixed_a(-0.02347925491631031)),(to_sfixed_a(0.01683058775961399)),(to_sfixed_a(-0.1493266224861145)),(to_sfixed_a(-0.2854035198688507)),(to_sfixed_a(0.20698010921478271)),(to_sfixed_a(0.4029029607772827)),(to_sfixed_a(-0.0013120152289047837)),(to_sfixed_a(0.03443126007914543)),(to_sfixed_a(0.13170939683914185)),(to_sfixed_a(0.038612812757492065)),(to_sfixed_a(0.06754381954669952)),(to_sfixed_a(0.2696104645729065)),(to_sfixed_a(0.11258304119110107)),(to_sfixed_a(0.15122656524181366)),(to_sfixed_a(0.030095456168055534)),(to_sfixed_a(-2.0115003280807287e-05)),(to_sfixed_a(-0.00016222029807977378)),(to_sfixed_a(-8.404100663028657e-05)),(to_sfixed_a(4.868013638770208e-05)),(to_sfixed_a(-0.00010181470861425623)),(to_sfixed_a(0.00019229270401410758)),(to_sfixed_a(-0.004867029841989279)),(to_sfixed_a(-0.05127264931797981)),(to_sfixed_a(0.04846614599227905)),(to_sfixed_a(-0.1723778396844864)),(to_sfixed_a(0.014932665973901749)),(to_sfixed_a(0.10701299458742142)),(to_sfixed_a(0.321929931640625)),(to_sfixed_a(0.3506610095500946)),(to_sfixed_a(0.0599031038582325)),(to_sfixed_a(-0.2020895928144455)),(to_sfixed_a(-0.1655554473400116)),(to_sfixed_a(0.02787637524306774)),(to_sfixed_a(-0.09205053746700287)),(to_sfixed_a(-0.25605228543281555)),(to_sfixed_a(-0.3506280779838562)),(to_sfixed_a(-0.20513829588890076)),(to_sfixed_a(-0.13659898936748505)),(to_sfixed_a(-0.2179570198059082)),(to_sfixed_a(-0.1510998159646988)),(to_sfixed_a(0.1614064872264862)),(to_sfixed_a(0.08802419155836105)),(to_sfixed_a(-0.00011481085675768554)),(to_sfixed_a(0.00021848878532182425)),(to_sfixed_a(-0.0001724567118799314)),(to_sfixed_a(0.0001620595285203308)),(to_sfixed_a(-5.657790461555123e-05)),(to_sfixed_a(0.0002292256394866854)),(to_sfixed_a(0.00031672525801695883)),(to_sfixed_a(-0.005600782111287117)),(to_sfixed_a(-0.04838748648762703)),(to_sfixed_a(-0.16437546908855438)),(to_sfixed_a(0.06380093842744827)),(to_sfixed_a(0.1654929667711258)),(to_sfixed_a(0.1823481172323227)),(to_sfixed_a(0.39901790022850037)),(to_sfixed_a(0.11395376175642014)),(to_sfixed_a(0.009414269588887691)),(to_sfixed_a(0.03757896274328232)),(to_sfixed_a(-0.07087370753288269)),(to_sfixed_a(0.26988866925239563)),(to_sfixed_a(0.06790397316217422)),(to_sfixed_a(-0.11545339226722717)),(to_sfixed_a(0.006972258910536766)),(to_sfixed_a(-0.046501513570547104)),(to_sfixed_a(0.3169284462928772)),(to_sfixed_a(0.06272581964731216)),(to_sfixed_a(-0.059488147497177124)),(to_sfixed_a(0.07469470053911209)),(to_sfixed_a(0.1421063095331192)),(to_sfixed_a(0.027603795751929283)),(to_sfixed_a(-0.000224838440772146)),(to_sfixed_a(3.3949319913517684e-05)),(to_sfixed_a(-0.00029419356724247336)),(to_sfixed_a(5.040970063419081e-05)),(to_sfixed_a(0.00012377604434732348)),(to_sfixed_a(0.04292941093444824)),(to_sfixed_a(-0.15689297020435333)),(to_sfixed_a(-0.0033701732754707336)),(to_sfixed_a(0.12266375124454498)),(to_sfixed_a(0.02216632105410099)),(to_sfixed_a(0.03625527769327164)),(to_sfixed_a(0.11077804118394852)),(to_sfixed_a(-0.05616181716322899)),(to_sfixed_a(-0.013692514970898628)),(to_sfixed_a(-0.015814587473869324)),(to_sfixed_a(-0.08825556933879852)),(to_sfixed_a(0.1433335840702057)),(to_sfixed_a(0.021155240014195442)),(to_sfixed_a(-0.15643998980522156)),(to_sfixed_a(-0.24936750531196594)),(to_sfixed_a(-0.038333047181367874)),(to_sfixed_a(0.24423179030418396)),(to_sfixed_a(0.3394358456134796)),(to_sfixed_a(0.26388072967529297)),(to_sfixed_a(0.3188132643699646)),(to_sfixed_a(0.1191796287894249)),(to_sfixed_a(0.13480882346630096)),(to_sfixed_a(3.988598837167956e-05)),(to_sfixed_a(8.85228073457256e-05)),(to_sfixed_a(-0.00012041769514326006)),(to_sfixed_a(0.00011619205179158598)),(to_sfixed_a(-0.0002157737035304308)),(to_sfixed_a(-0.00017286068759858608)),(to_sfixed_a(-7.06261198502034e-05)),(to_sfixed_a(-0.04533980414271355)),(to_sfixed_a(0.11809472739696503)),(to_sfixed_a(0.03665967658162117)),(to_sfixed_a(-0.017084935680031776)),(to_sfixed_a(0.0622231662273407)),(to_sfixed_a(0.11941903829574585)),(to_sfixed_a(0.018259096890687943)),(to_sfixed_a(-0.07282271236181259)),(to_sfixed_a(-0.04466252401471138)),(to_sfixed_a(-0.019785316661000252)),(to_sfixed_a(0.08330681174993515)),(to_sfixed_a(-0.15876145660877228)),(to_sfixed_a(-0.23540066182613373)),(to_sfixed_a(-0.2920338213443756)),(to_sfixed_a(-0.1310334950685501)),(to_sfixed_a(0.19839933514595032)),(to_sfixed_a(0.11539816111326218)),(to_sfixed_a(0.15468381345272064)),(to_sfixed_a(0.1571059674024582)),(to_sfixed_a(0.1498965322971344)),(to_sfixed_a(0.2630402743816376)),(to_sfixed_a(0.00010279787238687277)),(to_sfixed_a(-8.114362572086975e-05)),(to_sfixed_a(-0.00011301283666398376)),(to_sfixed_a(6.431460496969521e-05)),(to_sfixed_a(5.632550528389402e-05)),(to_sfixed_a(-6.944923370610923e-05)),(to_sfixed_a(-0.00011409933358663693)),(to_sfixed_a(-0.029656175523996353)),(to_sfixed_a(0.12146678566932678)),(to_sfixed_a(0.23277264833450317)),(to_sfixed_a(0.1456064134836197)),(to_sfixed_a(0.07672671973705292)),(to_sfixed_a(0.06275990605354309)),(to_sfixed_a(0.09229637682437897)),(to_sfixed_a(0.05772995576262474)),(to_sfixed_a(0.3033319115638733)),(to_sfixed_a(0.0609903447329998)),(to_sfixed_a(-0.05884364992380142)),(to_sfixed_a(-0.14691029489040375)),(to_sfixed_a(-0.26183006167411804)),(to_sfixed_a(-0.31677815318107605)),(to_sfixed_a(-0.07381648570299149)),(to_sfixed_a(0.10848596692085266)),(to_sfixed_a(0.00042053734068758786)),(to_sfixed_a(-0.005001178476959467)),(to_sfixed_a(0.05060647800564766)),(to_sfixed_a(0.3226812481880188)),(to_sfixed_a(-0.03254147619009018)),(to_sfixed_a(-0.0031375864055007696)),(to_sfixed_a(-0.004569192882627249)),(to_sfixed_a(-0.0002607674105092883)),(to_sfixed_a(0.00013123831013217568)),(to_sfixed_a(0.0002085841551888734)),(to_sfixed_a(-0.0005694815190508962)),(to_sfixed_a(-2.1151887267478742e-05)),(to_sfixed_a(0.0019732164219021797)),(to_sfixed_a(0.23002709448337555)),(to_sfixed_a(0.06720487028360367)),(to_sfixed_a(0.2694205641746521)),(to_sfixed_a(0.16287240386009216)),(to_sfixed_a(0.22126004099845886)),(to_sfixed_a(0.26688167452812195)),(to_sfixed_a(0.15192922949790955)),(to_sfixed_a(0.10883065313100815)),(to_sfixed_a(-0.02639545127749443)),(to_sfixed_a(-0.12276288121938705)),(to_sfixed_a(-0.051721785217523575)),(to_sfixed_a(-0.1545034945011139)),(to_sfixed_a(-0.30398982763290405)),(to_sfixed_a(-0.2524118721485138)),(to_sfixed_a(-0.2614399790763855)),(to_sfixed_a(0.06590277701616287)),(to_sfixed_a(-0.008273203857243061)),(to_sfixed_a(-0.06298305839300156)),(to_sfixed_a(0.10178549587726593)),(to_sfixed_a(-0.06205132231116295)),(to_sfixed_a(-7.792375981807709e-05)),(to_sfixed_a(5.950725244474597e-05)),(to_sfixed_a(0.0001284301542909816)),(to_sfixed_a(-0.00019839245942421257)),(to_sfixed_a(0.00020884518744423985)),(to_sfixed_a(0.0002003788686124608)),(to_sfixed_a(0.00017247095820493996)),(to_sfixed_a(0.050501372665166855)),(to_sfixed_a(0.26923519372940063)),(to_sfixed_a(0.12049289047718048)),(to_sfixed_a(0.20876388251781464)),(to_sfixed_a(0.1499122530221939)),(to_sfixed_a(0.16896654665470123)),(to_sfixed_a(0.2663005292415619)),(to_sfixed_a(-0.13866733014583588)),(to_sfixed_a(0.007850429974496365)),(to_sfixed_a(-0.06234490126371384)),(to_sfixed_a(-0.2854788899421692)),(to_sfixed_a(-0.038566358387470245)),(to_sfixed_a(-0.3028291165828705)),(to_sfixed_a(-0.19733862578868866)),(to_sfixed_a(-0.06351689249277115)),(to_sfixed_a(-0.28450652956962585)),(to_sfixed_a(0.1691819131374359)),(to_sfixed_a(0.012011880986392498)),(to_sfixed_a(-0.16506733000278473)),(to_sfixed_a(0.010127894580364227)),(to_sfixed_a(0.05133608728647232)),(to_sfixed_a(-0.0003965049982070923)),(to_sfixed_a(-7.812050898792222e-05)),(to_sfixed_a(-0.0002427232393529266)),(to_sfixed_a(0.00019751381478272378)),(to_sfixed_a(-2.2043665012461133e-05)),(to_sfixed_a(5.088644684292376e-05)),(to_sfixed_a(0.0007391144754365087)),(to_sfixed_a(0.07790869474411011)),(to_sfixed_a(0.055102989077568054)),(to_sfixed_a(-0.1987132877111435)),(to_sfixed_a(0.03755122423171997)),(to_sfixed_a(0.0027049388736486435)),(to_sfixed_a(-0.06330397725105286)),(to_sfixed_a(-0.02078341506421566)),(to_sfixed_a(-0.13830284774303436)),(to_sfixed_a(-0.015569265931844711)),(to_sfixed_a(-0.30944502353668213)),(to_sfixed_a(-0.020877182483673096)),(to_sfixed_a(0.1035861000418663)),(to_sfixed_a(-0.4040375053882599)),(to_sfixed_a(-0.15825670957565308)),(to_sfixed_a(-0.018250877037644386)),(to_sfixed_a(-0.20473934710025787)),(to_sfixed_a(-0.11737487465143204)),(to_sfixed_a(-0.2689417004585266)),(to_sfixed_a(-0.08434370160102844)),(to_sfixed_a(0.024712054058909416)),(to_sfixed_a(-0.01922784186899662)),(to_sfixed_a(-0.007708998396992683)),(to_sfixed_a(-0.0001157090300694108)),(to_sfixed_a(4.440778138814494e-05)),(to_sfixed_a(-7.34377681510523e-06)),(to_sfixed_a(0.0002937757526524365)),(to_sfixed_a(0.0014502134872600436)),(to_sfixed_a(0.0005594157264567912)),(to_sfixed_a(0.07922215014696121)),(to_sfixed_a(0.04130180925130844)),(to_sfixed_a(-0.0693494975566864)),(to_sfixed_a(-0.3682754635810852)),(to_sfixed_a(-0.06520821154117584)),(to_sfixed_a(0.022747278213500977)),(to_sfixed_a(0.02230245992541313)),(to_sfixed_a(-0.07498642802238464)),(to_sfixed_a(-0.17733973264694214)),(to_sfixed_a(-0.23127034306526184)),(to_sfixed_a(-0.07107380777597427)),(to_sfixed_a(0.02878105267882347)),(to_sfixed_a(-0.37385839223861694)),(to_sfixed_a(-0.24711637198925018)),(to_sfixed_a(-0.2693248987197876)),(to_sfixed_a(-0.06505946815013885)),(to_sfixed_a(-0.02293277345597744)),(to_sfixed_a(-0.1646798849105835)),(to_sfixed_a(-0.01876010186970234)),(to_sfixed_a(0.02042052522301674)),(to_sfixed_a(-6.659892096649855e-05)),(to_sfixed_a(4.970835107087623e-06)),(to_sfixed_a(-6.122255581431091e-05)),(to_sfixed_a(4.413682108861394e-05)),(to_sfixed_a(-6.808416947023943e-05)),(to_sfixed_a(0.00024725706316530704)),(to_sfixed_a(-4.717383853858337e-05)),(to_sfixed_a(-0.026281027123332024)),(to_sfixed_a(0.012914675287902355)),(to_sfixed_a(0.1944779008626938)),(to_sfixed_a(0.14745791256427765)),(to_sfixed_a(0.10783512145280838)),(to_sfixed_a(0.054224953055381775)),(to_sfixed_a(0.16526131331920624)),(to_sfixed_a(-0.0819719061255455)),(to_sfixed_a(-0.21466240286827087)),(to_sfixed_a(-0.23707924783229828)),(to_sfixed_a(-0.07756198197603226)),(to_sfixed_a(0.08364565670490265)),(to_sfixed_a(-0.09218687564134598)),(to_sfixed_a(-0.14480438828468323)),(to_sfixed_a(-0.19259291887283325)),(to_sfixed_a(-0.2664877474308014)),(to_sfixed_a(-0.3701084554195404)),(to_sfixed_a(-0.177725687623024)),(to_sfixed_a(-0.2987736165523529)),(to_sfixed_a(0.017695607617497444)),(to_sfixed_a(0.020649611949920654)),(to_sfixed_a(0.0015231013530865312)),(to_sfixed_a(8.550031634513289e-05)),(to_sfixed_a(-0.00012891917140223086)),(to_sfixed_a(-0.00015576838632114232)),(to_sfixed_a(7.023759098956361e-05)),(to_sfixed_a(-0.00015641615027561784)),(to_sfixed_a(4.363276457297616e-05)),(to_sfixed_a(-0.01890798844397068)),(to_sfixed_a(-0.002362085971981287)),(to_sfixed_a(0.0187800582498312)),(to_sfixed_a(0.0587579719722271)),(to_sfixed_a(0.05343618988990784)),(to_sfixed_a(0.32509735226631165)),(to_sfixed_a(0.12079261243343353)),(to_sfixed_a(0.19284634292125702)),(to_sfixed_a(0.05427195131778717)),(to_sfixed_a(-0.06739789247512817)),(to_sfixed_a(0.05879608169198036)),(to_sfixed_a(0.0332111157476902)),(to_sfixed_a(-0.38762167096138)),(to_sfixed_a(-0.04349112883210182)),(to_sfixed_a(-0.1464628279209137)),(to_sfixed_a(-0.17685571312904358)),(to_sfixed_a(-0.1264524757862091)),(to_sfixed_a(-0.024518253281712532)),(to_sfixed_a(-0.2499603033065796)),(to_sfixed_a(0.03752799704670906)),(to_sfixed_a(0.39270538091659546)),(to_sfixed_a(0.00021584522619377822)),(to_sfixed_a(7.570093293907121e-05)),(to_sfixed_a(-0.00013397066504694521)),(to_sfixed_a(0.00013972941087558866)),(to_sfixed_a(0.00028096334426663816)),(to_sfixed_a(4.3356507376302034e-05)),(to_sfixed_a(4.5405144192045555e-05)),(to_sfixed_a(-0.00014109440962783992)),(to_sfixed_a(0.02371126599609852)),(to_sfixed_a(0.08025285601615906)),(to_sfixed_a(0.2803483009338379)),(to_sfixed_a(-0.00531577505171299)),(to_sfixed_a(0.14786286652088165)),(to_sfixed_a(0.28799429535865784)),(to_sfixed_a(0.06944429129362106)),(to_sfixed_a(0.4192543625831604)),(to_sfixed_a(0.2502637803554535)),(to_sfixed_a(0.06833834946155548)),(to_sfixed_a(-0.25227823853492737)),(to_sfixed_a(-0.27820831537246704)),(to_sfixed_a(-0.1639855057001114)),(to_sfixed_a(-0.18627828359603882)),(to_sfixed_a(-0.49711430072784424)),(to_sfixed_a(-0.28382760286331177)),(to_sfixed_a(-0.028159277513623238)),(to_sfixed_a(0.3612375557422638)),(to_sfixed_a(0.08440449833869934)),(to_sfixed_a(0.07057793438434601)),(to_sfixed_a(0.019617898389697075)),(to_sfixed_a(9.682211384642869e-05)),(to_sfixed_a(0.00011822285887319595)),(to_sfixed_a(-4.259970228304155e-05)),(to_sfixed_a(-0.0003010470827575773)),(to_sfixed_a(0.0003329607716295868)),(to_sfixed_a(-0.00012311719183344394)),(to_sfixed_a(0.00013757146371062845)),(to_sfixed_a(-0.056242313235998154)),(to_sfixed_a(-0.00030861294362694025)),(to_sfixed_a(0.26315510272979736)),(to_sfixed_a(0.12010455876588821)),(to_sfixed_a(0.10485557466745377)),(to_sfixed_a(0.2234242558479309)),(to_sfixed_a(0.2697382867336273)),(to_sfixed_a(0.2970341145992279)),(to_sfixed_a(0.14274847507476807)),(to_sfixed_a(0.14130179584026337)),(to_sfixed_a(-0.053287114948034286)),(to_sfixed_a(0.054272882640361786)),(to_sfixed_a(-0.17261438071727753)),(to_sfixed_a(-0.5573079586029053)),(to_sfixed_a(-0.3304480314254761)),(to_sfixed_a(-0.13825955986976624)),(to_sfixed_a(0.4746472239494324)),(to_sfixed_a(0.18263521790504456)),(to_sfixed_a(0.3061147630214691)),(to_sfixed_a(-0.0009321183897554874)),(to_sfixed_a(0.03400935232639313)),(to_sfixed_a(-0.00013492272410076112)),(to_sfixed_a(-0.00010783641482703388)),(to_sfixed_a(0.00011306535452604294)),(to_sfixed_a(5.275104922475293e-05)),(to_sfixed_a(-0.00024458402185700834)),(to_sfixed_a(0.00016012116975616664)),(to_sfixed_a(0.00013501527428161353)),(to_sfixed_a(6.0389735153876245e-05)),(to_sfixed_a(-0.08072184771299362)),(to_sfixed_a(0.015959925949573517)),(to_sfixed_a(0.20719410479068756)),(to_sfixed_a(0.11198902875185013)),(to_sfixed_a(0.07407404482364655)),(to_sfixed_a(0.19159413874149323)),(to_sfixed_a(0.06363984197378159)),(to_sfixed_a(0.12713877856731415)),(to_sfixed_a(0.050041019916534424)),(to_sfixed_a(-0.10070950537919998)),(to_sfixed_a(-0.03781343251466751)),(to_sfixed_a(-0.16611891984939575)),(to_sfixed_a(-0.2303011417388916)),(to_sfixed_a(-0.3151310682296753)),(to_sfixed_a(-0.13560084998607635)),(to_sfixed_a(0.08335509896278381)),(to_sfixed_a(0.031884532421827316)),(to_sfixed_a(0.03647420182824135)),(to_sfixed_a(0.00140235701110214)),(to_sfixed_a(-7.226104207802564e-05)),(to_sfixed_a(0.00014833372551947832)),(to_sfixed_a(-0.00011938879470108077)),(to_sfixed_a(2.72340571427776e-06)),(to_sfixed_a(0.00011795174214057624)),(to_sfixed_a(-1.3905719242757186e-05)),(to_sfixed_a(-0.00025568969431333244)),(to_sfixed_a(0.0002262815396534279)),(to_sfixed_a(0.00018909428035840392)),(to_sfixed_a(-0.007511096075177193)),(to_sfixed_a(0.1902589648962021)),(to_sfixed_a(-0.14431820809841156)),(to_sfixed_a(0.11962808668613434)),(to_sfixed_a(0.14519579708576202)),(to_sfixed_a(0.061974652111530304)),(to_sfixed_a(0.05761103704571724)),(to_sfixed_a(0.24366916716098785)),(to_sfixed_a(-0.08341260999441147)),(to_sfixed_a(-0.09565415233373642)),(to_sfixed_a(-0.09323764592409134)),(to_sfixed_a(-0.43125051259994507)),(to_sfixed_a(-0.046527199447155)),(to_sfixed_a(-0.017505813390016556)),(to_sfixed_a(-0.008006369695067406)),(to_sfixed_a(0.03470799699425697)),(to_sfixed_a(0.11993084102869034)),(to_sfixed_a(0.001342038856819272)),(to_sfixed_a(0.07928785681724548)),(to_sfixed_a(-3.9719259802950546e-05)),(to_sfixed_a(1.7000032812575228e-06)),(to_sfixed_a(0.0003055882116314024)),(to_sfixed_a(8.987384353531525e-05)),(to_sfixed_a(5.938165122643113e-05)),(to_sfixed_a(-0.00010097766789840534)),(to_sfixed_a(0.00010379763989476487)),(to_sfixed_a(-3.577728057280183e-05)),(to_sfixed_a(-0.003199870465323329)),(to_sfixed_a(0.031185006722807884)),(to_sfixed_a(-0.011273008771240711)),(to_sfixed_a(-0.13069483637809753)),(to_sfixed_a(0.09925319254398346)),(to_sfixed_a(0.13308432698249817)),(to_sfixed_a(-0.10568558424711227)),(to_sfixed_a(-0.02816612459719181)),(to_sfixed_a(-0.14033161103725433)),(to_sfixed_a(0.14378416538238525)),(to_sfixed_a(-0.046665892004966736)),(to_sfixed_a(-0.07164227217435837)),(to_sfixed_a(-0.416202574968338)),(to_sfixed_a(-0.346132755279541)),(to_sfixed_a(-0.1292562186717987)),(to_sfixed_a(-0.012664485722780228)),(to_sfixed_a(0.018393943086266518)),(to_sfixed_a(0.10465370118618011)),(to_sfixed_a(0.04449792951345444)),(to_sfixed_a(-0.004832453094422817)),(to_sfixed_a(-8.67251874296926e-05)),(to_sfixed_a(-0.00016407026851084083)),(to_sfixed_a(-6.951074465177953e-05)),(to_sfixed_a(0.00011950764746870846)),(to_sfixed_a(0.0001018230541376397)),(to_sfixed_a(-0.0001020242998492904)),(to_sfixed_a(0.0002543179434724152)),(to_sfixed_a(-0.0001178826205432415)),(to_sfixed_a(-8.14979721326381e-05)),(to_sfixed_a(-0.044726841151714325)),(to_sfixed_a(-0.0076781874522566795)),(to_sfixed_a(0.026473332196474075)),(to_sfixed_a(-0.11346922814846039)),(to_sfixed_a(-0.10646115988492966)),(to_sfixed_a(-0.006089663133025169)),(to_sfixed_a(0.024719513952732086)),(to_sfixed_a(-0.19312669336795807)),(to_sfixed_a(-0.06508142501115799)),(to_sfixed_a(-0.017534883692860603)),(to_sfixed_a(-0.019948197528719902)),(to_sfixed_a(0.013311718590557575)),(to_sfixed_a(0.011841796338558197)),(to_sfixed_a(0.004027070477604866)),(to_sfixed_a(0.03427113965153694)),(to_sfixed_a(-0.1200828105211258)),(to_sfixed_a(-0.000613601878285408)),(to_sfixed_a(-0.0033799600787460804)),(to_sfixed_a(-0.0035111468750983477)),(to_sfixed_a(-9.660687646828592e-05)),(to_sfixed_a(0.0001711505465209484)),(to_sfixed_a(-0.00010243673023069277)),(to_sfixed_a(-0.0002002661203732714)),(to_sfixed_a(-2.4777034923317842e-05)),(to_sfixed_a(-4.998477015760727e-05)),(to_sfixed_a(-0.00013021539780311286)),(to_sfixed_a(0.00015342261758632958)),(to_sfixed_a(-2.4463195586577058e-05)),(to_sfixed_a(0.0006157382158562541)),(to_sfixed_a(0.000682758807670325)),(to_sfixed_a(-7.50554318074137e-05)),(to_sfixed_a(-0.00012370676267892122)),(to_sfixed_a(0.00036160016315989196)),(to_sfixed_a(0.026760714128613472)),(to_sfixed_a(-0.004949756897985935)),(to_sfixed_a(-0.0009957881411537528)),(to_sfixed_a(0.011810239404439926)),(to_sfixed_a(-0.17898592352867126)),(to_sfixed_a(0.0037721474654972553)),(to_sfixed_a(-0.0014981355052441359)),(to_sfixed_a(0.024502750486135483)),(to_sfixed_a(0.03143102675676346)),(to_sfixed_a(-0.003992937970906496)),(to_sfixed_a(0.00035921556991524994)),(to_sfixed_a(0.00013591187598649412)),(to_sfixed_a(0.00011558774713193998)),(to_sfixed_a(-0.00026041455566883087)),(to_sfixed_a(6.394466618075967e-05)),(to_sfixed_a(-0.0003088129451498389)),(to_sfixed_a(5.124882954987697e-05)),(to_sfixed_a(4.980747326044366e-05)),(to_sfixed_a(-0.00011609394277911633)),(to_sfixed_a(-1.5480237607334857e-06)),(to_sfixed_a(0.0002784702810458839)),(to_sfixed_a(-0.00020521173428278416)),(to_sfixed_a(0.0003220803337171674)),(to_sfixed_a(-0.00016906566452234983)),(to_sfixed_a(-0.0001252263755304739)),(to_sfixed_a(-6.085454060666962e-06)),(to_sfixed_a(-3.069519152631983e-05)),(to_sfixed_a(-0.00013613556802738458)),(to_sfixed_a(2.611765239635133e-06)),(to_sfixed_a(2.866360046027694e-05)),(to_sfixed_a(0.00017586983449291438)),(to_sfixed_a(-0.00018288346473127604)),(to_sfixed_a(-0.00015245037502609193)),(to_sfixed_a(0.00013015736476518214)),(to_sfixed_a(-4.24107420258224e-05)),(to_sfixed_a(3.017937342519872e-05)),(to_sfixed_a(-6.415363168343902e-05)),(to_sfixed_a(-1.2956157661392353e-05)),(to_sfixed_a(-7.867711974540725e-05)),(to_sfixed_a(3.916594141628593e-05)),(to_sfixed_a(4.315137630328536e-05)),(to_sfixed_a(4.7214278311003e-05)),(to_sfixed_a(-0.0002479685063008219)),(to_sfixed_a(0.00027004245202988386)),(to_sfixed_a(-0.0003058520669583231)),(to_sfixed_a(0.00011994731175946072)));

    constant weight_n0_17 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-0.00013584221596829593)),(to_sfixed_a(-0.00011153803643537685)),(to_sfixed_a(0.00019465557124931365)),(to_sfixed_a(9.947286889655516e-05)),(to_sfixed_a(3.995343286078423e-05)),(to_sfixed_a(2.838357431755867e-05)),(to_sfixed_a(9.807009519136045e-06)),(to_sfixed_a(2.8590517104021274e-05)),(to_sfixed_a(-3.993365680798888e-05)),(to_sfixed_a(-7.709843339398503e-05)),(to_sfixed_a(-0.00020889889856334776)),(to_sfixed_a(0.0002004380658036098)),(to_sfixed_a(0.000122519995784387)),(to_sfixed_a(-3.2658139389241114e-05)),(to_sfixed_a(6.383705112966709e-06)),(to_sfixed_a(-0.00012566072109621018)),(to_sfixed_a(-3.175912206643261e-05)),(to_sfixed_a(-0.00010420633770991117)),(to_sfixed_a(-0.00022591606830246747)),(to_sfixed_a(-0.00014720053877681494)),(to_sfixed_a(4.171834370936267e-05)),(to_sfixed_a(9.83017889666371e-06)),(to_sfixed_a(6.0830676375189796e-05)),(to_sfixed_a(1.7640020814724267e-05)),(to_sfixed_a(0.00029403576627373695)),(to_sfixed_a(-4.979319783160463e-05)),(to_sfixed_a(0.00023478176444768906)),(to_sfixed_a(2.4429977202089503e-05)),(to_sfixed_a(-0.0001197907404275611)),(to_sfixed_a(1.1221930435567629e-05)),(to_sfixed_a(3.85191997338552e-05)),(to_sfixed_a(1.711879349386436e-08)),(to_sfixed_a(0.00022678716049995273)),(to_sfixed_a(0.0002726704115048051)),(to_sfixed_a(0.00034521499765105546)),(to_sfixed_a(-0.00010525083780521527)),(to_sfixed_a(0.00019294711819384247)),(to_sfixed_a(-3.163045403198339e-05)),(to_sfixed_a(4.2528020571808156e-07)),(to_sfixed_a(4.224869189783931e-05)),(to_sfixed_a(-3.516477590892464e-05)),(to_sfixed_a(-7.879280019551516e-05)),(to_sfixed_a(4.215574881527573e-05)),(to_sfixed_a(-6.573663267772645e-05)),(to_sfixed_a(-0.00011656647257041186)),(to_sfixed_a(-7.168369484134018e-05)),(to_sfixed_a(5.7127635955112055e-05)),(to_sfixed_a(0.00014102086424827576)),(to_sfixed_a(0.0001599844399606809)),(to_sfixed_a(-3.91702342312783e-05)),(to_sfixed_a(-4.101619197172113e-05)),(to_sfixed_a(-6.637074693571776e-05)),(to_sfixed_a(-8.319811604451388e-05)),(to_sfixed_a(-0.00012243584205862135)),(to_sfixed_a(-0.0001889461709652096)),(to_sfixed_a(4.049062408739701e-05)),(to_sfixed_a(-0.0001593652123119682)),(to_sfixed_a(0.0004225815355312079)),(to_sfixed_a(-8.054743375396356e-05)),(to_sfixed_a(0.00011293307761661708)),(to_sfixed_a(-5.101052738609724e-05)),(to_sfixed_a(-0.00024066826154012233)),(to_sfixed_a(-0.00022967193217482418)),(to_sfixed_a(0.00015806133160367608)),(to_sfixed_a(4.4526223064167425e-05)),(to_sfixed_a(-6.998373282840475e-05)),(to_sfixed_a(-8.683577107149176e-06)),(to_sfixed_a(-0.00017662438040133566)),(to_sfixed_a(8.130168862408027e-05)),(to_sfixed_a(0.01126146875321865)),(to_sfixed_a(-0.00011185489711351693)),(to_sfixed_a(-3.014587491634302e-05)),(to_sfixed_a(0.00012385461013764143)),(to_sfixed_a(-1.8074999388772994e-05)),(to_sfixed_a(-0.00020266987849026918)),(to_sfixed_a(-6.43932389721158e-06)),(to_sfixed_a(7.924795500002801e-05)),(to_sfixed_a(0.00023158638214226812)),(to_sfixed_a(-0.00015180707850959152)),(to_sfixed_a(0.0002771683211904019)),(to_sfixed_a(0.00018038069538306445)),(to_sfixed_a(8.816396439215168e-05)),(to_sfixed_a(-0.00019676687952596694)),(to_sfixed_a(5.543522274820134e-05)),(to_sfixed_a(-0.00018908013589680195)),(to_sfixed_a(-0.000267323775915429)),(to_sfixed_a(-0.0003037108399439603)),(to_sfixed_a(0.00013792861136607826)),(to_sfixed_a(5.857830910827033e-05)),(to_sfixed_a(-0.0002481121919117868)),(to_sfixed_a(5.68617622320744e-07)),(to_sfixed_a(0.00016885316290427)),(to_sfixed_a(0.014888448640704155)),(to_sfixed_a(-5.411518486653222e-06)),(to_sfixed_a(0.01692182756960392)),(to_sfixed_a(0.00970859918743372)),(to_sfixed_a(-0.016000283882021904)),(to_sfixed_a(0.08885487914085388)),(to_sfixed_a(0.03826112300157547)),(to_sfixed_a(-0.030890844762325287)),(to_sfixed_a(-0.020001066848635674)),(to_sfixed_a(0.04948688670992851)),(to_sfixed_a(0.06126834824681282)),(to_sfixed_a(0.0185032207518816)),(to_sfixed_a(-0.0022032565902918577)),(to_sfixed_a(-0.004312028642743826)),(to_sfixed_a(-0.00015191000420600176)),(to_sfixed_a(-4.7388348320964724e-05)),(to_sfixed_a(8.485838770866394e-05)),(to_sfixed_a(-0.0002149590291082859)),(to_sfixed_a(-1.140451422543265e-05)),(to_sfixed_a(9.341466648038477e-05)),(to_sfixed_a(0.000319914921419695)),(to_sfixed_a(-5.99784470978193e-06)),(to_sfixed_a(-7.95952928456245e-07)),(to_sfixed_a(5.2161685744067654e-05)),(to_sfixed_a(0.00030174441053532064)),(to_sfixed_a(1.3778623724647332e-05)),(to_sfixed_a(-0.0001968753058463335)),(to_sfixed_a(0.012988993898034096)),(to_sfixed_a(-0.11776509881019592)),(to_sfixed_a(0.023425955325365067)),(to_sfixed_a(0.2737351059913635)),(to_sfixed_a(-0.0018136491999030113)),(to_sfixed_a(0.1945931315422058)),(to_sfixed_a(0.06964287161827087)),(to_sfixed_a(0.02676430158317089)),(to_sfixed_a(0.2544576823711395)),(to_sfixed_a(0.08193168044090271)),(to_sfixed_a(0.22429583966732025)),(to_sfixed_a(0.0228115227073431)),(to_sfixed_a(0.06574497371912003)),(to_sfixed_a(-0.018431363627314568)),(to_sfixed_a(-0.0031047493685036898)),(to_sfixed_a(0.050082866102457047)),(to_sfixed_a(0.00022765800531487912)),(to_sfixed_a(-0.0028905323706567287)),(to_sfixed_a(-3.844550155918114e-05)),(to_sfixed_a(-0.00013336408301256597)),(to_sfixed_a(0.00015040063590276986)),(to_sfixed_a(0.00030652686837129295)),(to_sfixed_a(2.744292578427121e-05)),(to_sfixed_a(0.00017135441885329783)),(to_sfixed_a(-4.893497680313885e-05)),(to_sfixed_a(-0.0002998052223119885)),(to_sfixed_a(0.0420365184545517)),(to_sfixed_a(0.017383785918354988)),(to_sfixed_a(0.030439775437116623)),(to_sfixed_a(-0.009887928143143654)),(to_sfixed_a(-0.03305337205529213)),(to_sfixed_a(-0.05306268855929375)),(to_sfixed_a(0.019608795642852783)),(to_sfixed_a(0.11159343272447586)),(to_sfixed_a(0.15975835919380188)),(to_sfixed_a(0.09304823726415634)),(to_sfixed_a(0.15086033940315247)),(to_sfixed_a(0.15575307607650757)),(to_sfixed_a(0.2283327430486679)),(to_sfixed_a(0.14794375002384186)),(to_sfixed_a(-0.14287517964839935)),(to_sfixed_a(0.05987746641039848)),(to_sfixed_a(0.015440806746482849)),(to_sfixed_a(-0.0067076776176691055)),(to_sfixed_a(0.005830790847539902)),(to_sfixed_a(0.00029729187372140586)),(to_sfixed_a(4.4534272092278115e-07)),(to_sfixed_a(-0.00015020798309706151)),(to_sfixed_a(-5.962555587757379e-05)),(to_sfixed_a(0.00034013547701761127)),(to_sfixed_a(0.00015562574844807386)),(to_sfixed_a(-0.0001592335756868124)),(to_sfixed_a(8.846295531839132e-05)),(to_sfixed_a(-1.4251233551476616e-05)),(to_sfixed_a(0.036164525896310806)),(to_sfixed_a(-0.004620353225618601)),(to_sfixed_a(0.06796596199274063)),(to_sfixed_a(-0.015714609995484352)),(to_sfixed_a(0.1658674031496048)),(to_sfixed_a(-0.21315360069274902)),(to_sfixed_a(-0.2671733796596527)),(to_sfixed_a(-0.11337128281593323)),(to_sfixed_a(0.0696743056178093)),(to_sfixed_a(-0.03838749974966049)),(to_sfixed_a(0.09346622973680496)),(to_sfixed_a(0.09967755526304245)),(to_sfixed_a(0.2108083814382553)),(to_sfixed_a(0.06228596717119217)),(to_sfixed_a(0.018771491944789886)),(to_sfixed_a(0.08775204420089722)),(to_sfixed_a(-0.08537913858890533)),(to_sfixed_a(-0.04217459261417389)),(to_sfixed_a(0.0830899178981781)),(to_sfixed_a(0.004223901778459549)),(to_sfixed_a(0.005795177072286606)),(to_sfixed_a(0.002182627795264125)),(to_sfixed_a(0.0002861101529560983)),(to_sfixed_a(-3.197044861735776e-05)),(to_sfixed_a(3.635351458797231e-05)),(to_sfixed_a(-0.0002156140108127147)),(to_sfixed_a(0.00018988497322425246)),(to_sfixed_a(-3.3183086998178624e-06)),(to_sfixed_a(0.04576247185468674)),(to_sfixed_a(0.0044902232475578785)),(to_sfixed_a(-0.09139984846115112)),(to_sfixed_a(0.1485775113105774)),(to_sfixed_a(-0.12905408442020416)),(to_sfixed_a(-0.30223095417022705)),(to_sfixed_a(-0.10066742449998856)),(to_sfixed_a(-0.10104671865701675)),(to_sfixed_a(-0.2733927071094513)),(to_sfixed_a(-0.049909621477127075)),(to_sfixed_a(0.006516674999147654)),(to_sfixed_a(0.10460933297872543)),(to_sfixed_a(0.15997926890850067)),(to_sfixed_a(-0.0520700141787529)),(to_sfixed_a(-0.021590810269117355)),(to_sfixed_a(0.1627195030450821)),(to_sfixed_a(-0.029737439006567)),(to_sfixed_a(0.07897290587425232)),(to_sfixed_a(-0.07398343086242676)),(to_sfixed_a(0.03094143234193325)),(to_sfixed_a(0.003447264665737748)),(to_sfixed_a(-3.0440673072007485e-05)),(to_sfixed_a(-6.296533683780581e-06)),(to_sfixed_a(-0.00012805958976969123)),(to_sfixed_a(0.00011859304504469037)),(to_sfixed_a(0.00014711200492456555)),(to_sfixed_a(0.0001168401722679846)),(to_sfixed_a(-0.11964458227157593)),(to_sfixed_a(0.005542748142033815)),(to_sfixed_a(-0.015420977026224136)),(to_sfixed_a(-0.10363399237394333)),(to_sfixed_a(-0.08592282235622406)),(to_sfixed_a(-0.05462590977549553)),(to_sfixed_a(0.05263352021574974)),(to_sfixed_a(-0.05189184844493866)),(to_sfixed_a(-0.022005656734108925)),(to_sfixed_a(0.03379858285188675)),(to_sfixed_a(0.12428361177444458)),(to_sfixed_a(0.22130565345287323)),(to_sfixed_a(0.2910867929458618)),(to_sfixed_a(-0.050503022968769073)),(to_sfixed_a(0.010539657436311245)),(to_sfixed_a(0.029324529692530632)),(to_sfixed_a(0.12581370770931244)),(to_sfixed_a(0.03936208412051201)),(to_sfixed_a(-0.09727325290441513)),(to_sfixed_a(0.04825182259082794)),(to_sfixed_a(0.04571690037846565)),(to_sfixed_a(0.0648464635014534)),(to_sfixed_a(0.000107666572148446)),(to_sfixed_a(0.00012397214595694095)),(to_sfixed_a(9.416727698408067e-05)),(to_sfixed_a(-7.919164636405185e-05)),(to_sfixed_a(-9.795978985494003e-05)),(to_sfixed_a(0.0002606296620797366)),(to_sfixed_a(-0.0017692047404125333)),(to_sfixed_a(-0.20590773224830627)),(to_sfixed_a(-0.07175389677286148)),(to_sfixed_a(-0.16650164127349854)),(to_sfixed_a(-0.022521881386637688)),(to_sfixed_a(-0.0438067764043808)),(to_sfixed_a(0.027116214856505394)),(to_sfixed_a(0.17802885174751282)),(to_sfixed_a(0.12740078568458557)),(to_sfixed_a(0.21352936327457428)),(to_sfixed_a(0.22878675162792206)),(to_sfixed_a(0.1222810447216034)),(to_sfixed_a(0.09380082786083221)),(to_sfixed_a(-0.12252160161733627)),(to_sfixed_a(-0.034252192825078964)),(to_sfixed_a(0.15940873324871063)),(to_sfixed_a(-0.04188301041722298)),(to_sfixed_a(-0.04901625216007233)),(to_sfixed_a(0.0717020183801651)),(to_sfixed_a(0.2494397908449173)),(to_sfixed_a(0.15497788786888123)),(to_sfixed_a(-1.4405570254893973e-05)),(to_sfixed_a(6.78760334267281e-05)),(to_sfixed_a(-8.494437497574836e-05)),(to_sfixed_a(3.475357880233787e-05)),(to_sfixed_a(-5.271102418191731e-05)),(to_sfixed_a(4.7887006076052785e-05)),(to_sfixed_a(0.00010848061356227845)),(to_sfixed_a(-0.0018383347196504474)),(to_sfixed_a(0.05550146475434303)),(to_sfixed_a(-0.06708208471536636)),(to_sfixed_a(0.006539229769259691)),(to_sfixed_a(-0.05687861889600754)),(to_sfixed_a(0.024629822000861168)),(to_sfixed_a(-0.02899269573390484)),(to_sfixed_a(0.2632381319999695)),(to_sfixed_a(0.21566982567310333)),(to_sfixed_a(0.18199053406715393)),(to_sfixed_a(0.06325056403875351)),(to_sfixed_a(-0.12046562135219574)),(to_sfixed_a(-0.17187504470348358)),(to_sfixed_a(-0.07898956537246704)),(to_sfixed_a(0.0013401401229202747)),(to_sfixed_a(-0.02525162138044834)),(to_sfixed_a(-0.04510875418782234)),(to_sfixed_a(0.10023726522922516)),(to_sfixed_a(-0.1501256376504898)),(to_sfixed_a(-0.07139863073825836)),(to_sfixed_a(-0.061539120972156525)),(to_sfixed_a(0.021638553589582443)),(to_sfixed_a(0.0001898693008115515)),(to_sfixed_a(-0.00027266007964499295)),(to_sfixed_a(0.0002970920177176595)),(to_sfixed_a(-0.00017703694174997509)),(to_sfixed_a(-0.00022996759798843414)),(to_sfixed_a(0.0008178958669304848)),(to_sfixed_a(-0.1176287978887558)),(to_sfixed_a(-0.10547126084566116)),(to_sfixed_a(-0.05499682575464249)),(to_sfixed_a(-0.07123760879039764)),(to_sfixed_a(-0.15826308727264404)),(to_sfixed_a(-0.26284506916999817)),(to_sfixed_a(-0.05399726703763008)),(to_sfixed_a(0.0312763936817646)),(to_sfixed_a(-0.07948427647352219)),(to_sfixed_a(0.09179854393005371)),(to_sfixed_a(-0.18506252765655518)),(to_sfixed_a(-0.30992186069488525)),(to_sfixed_a(-0.1976054161787033)),(to_sfixed_a(-0.19718413054943085)),(to_sfixed_a(-0.11555908620357513)),(to_sfixed_a(0.23296085000038147)),(to_sfixed_a(0.11043143272399902)),(to_sfixed_a(-0.008929984644055367)),(to_sfixed_a(0.03947897255420685)),(to_sfixed_a(0.03159784898161888)),(to_sfixed_a(-0.14893381297588348)),(to_sfixed_a(-8.062046981649473e-05)),(to_sfixed_a(-0.00010673090582713485)),(to_sfixed_a(5.625517587759532e-05)),(to_sfixed_a(-0.00019823815091513097)),(to_sfixed_a(2.9597158572869375e-05)),(to_sfixed_a(-4.5261313061928377e-05)),(to_sfixed_a(0.00021526234922930598)),(to_sfixed_a(-0.23693175613880157)),(to_sfixed_a(-0.3587653636932373)),(to_sfixed_a(-0.25438445806503296)),(to_sfixed_a(-0.07664696127176285)),(to_sfixed_a(-0.21215875446796417)),(to_sfixed_a(-0.25506314635276794)),(to_sfixed_a(-0.2423751950263977)),(to_sfixed_a(0.3780880570411682)),(to_sfixed_a(0.40202629566192627)),(to_sfixed_a(-0.19391703605651855)),(to_sfixed_a(-0.21312502026557922)),(to_sfixed_a(-0.5227583646774292)),(to_sfixed_a(-0.10946954041719437)),(to_sfixed_a(-0.3514547646045685)),(to_sfixed_a(-0.11356639862060547)),(to_sfixed_a(-0.0507768951356411)),(to_sfixed_a(0.0879158228635788)),(to_sfixed_a(-0.10020021349191666)),(to_sfixed_a(-0.129414364695549)),(to_sfixed_a(-0.42205050587654114)),(to_sfixed_a(0.1925230473279953)),(to_sfixed_a(-2.9297334549482912e-05)),(to_sfixed_a(0.00017162262520287186)),(to_sfixed_a(0.00016190386668313295)),(to_sfixed_a(-0.00014149505295790732)),(to_sfixed_a(2.7314034014125355e-05)),(to_sfixed_a(0.00019844439520966262)),(to_sfixed_a(0.00012334460916463286)),(to_sfixed_a(-0.07930382341146469)),(to_sfixed_a(-0.20369811356067657)),(to_sfixed_a(-0.2542906701564789)),(to_sfixed_a(-0.34223127365112305)),(to_sfixed_a(-0.18937966227531433)),(to_sfixed_a(-0.0764489620923996)),(to_sfixed_a(-0.2250647246837616)),(to_sfixed_a(0.1897677630186081)),(to_sfixed_a(0.32733264565467834)),(to_sfixed_a(-0.09442432969808578)),(to_sfixed_a(-0.4621049463748932)),(to_sfixed_a(-0.02108151465654373)),(to_sfixed_a(0.06445326656103134)),(to_sfixed_a(-0.22373706102371216)),(to_sfixed_a(0.047759559005498886)),(to_sfixed_a(-0.3363235294818878)),(to_sfixed_a(-0.11435192078351974)),(to_sfixed_a(-0.19101402163505554)),(to_sfixed_a(-0.21002039313316345)),(to_sfixed_a(-0.07821938395500183)),(to_sfixed_a(0.017151212319731712)),(to_sfixed_a(-0.0026079609524458647)),(to_sfixed_a(-0.002254500752314925)),(to_sfixed_a(0.00014387708506546915)),(to_sfixed_a(-3.3551218621141743e-06)),(to_sfixed_a(9.471458906773478e-05)),(to_sfixed_a(8.25617607915774e-05)),(to_sfixed_a(5.95433812122792e-05)),(to_sfixed_a(-0.000862944289110601)),(to_sfixed_a(-0.5298068523406982)),(to_sfixed_a(-0.03043566271662712)),(to_sfixed_a(-0.02425343170762062)),(to_sfixed_a(-0.26140615344047546)),(to_sfixed_a(-0.241013303399086)),(to_sfixed_a(0.03411255031824112)),(to_sfixed_a(0.10912537574768066)),(to_sfixed_a(0.11157529056072235)),(to_sfixed_a(-0.18597349524497986)),(to_sfixed_a(-0.018200291320681572)),(to_sfixed_a(-0.10665438324213028)),(to_sfixed_a(-0.04034379869699478)),(to_sfixed_a(-0.08123183250427246)),(to_sfixed_a(-0.1379241794347763)),(to_sfixed_a(-0.2576906979084015)),(to_sfixed_a(-0.22000445425510406)),(to_sfixed_a(-0.11863567680120468)),(to_sfixed_a(-0.022424932569265366)),(to_sfixed_a(0.12120246887207031)),(to_sfixed_a(-0.07804933190345764)),(to_sfixed_a(0.00022458478633780032)),(to_sfixed_a(9.05754859559238e-05)),(to_sfixed_a(0.000139310272061266)),(to_sfixed_a(-0.0003745304129552096)),(to_sfixed_a(2.883972592826467e-05)),(to_sfixed_a(-0.00018061380251310766)),(to_sfixed_a(-0.00013462465722113848)),(to_sfixed_a(-0.06590920686721802)),(to_sfixed_a(-0.2715076208114624)),(to_sfixed_a(-0.1612958461046219)),(to_sfixed_a(-0.2861280143260956)),(to_sfixed_a(-0.24037808179855347)),(to_sfixed_a(0.021292289718985558)),(to_sfixed_a(-0.016024185344576836)),(to_sfixed_a(0.2111433744430542)),(to_sfixed_a(0.11579544097185135)),(to_sfixed_a(-0.13547846674919128)),(to_sfixed_a(-0.13220642507076263)),(to_sfixed_a(-0.09629713743925095)),(to_sfixed_a(0.0063707600347697735)),(to_sfixed_a(-0.20739871263504028)),(to_sfixed_a(-0.015502242371439934)),(to_sfixed_a(-0.3169917166233063)),(to_sfixed_a(-0.1761089414358139)),(to_sfixed_a(-0.08359307050704956)),(to_sfixed_a(-0.06654607504606247)),(to_sfixed_a(0.058033186942338943)),(to_sfixed_a(0.2802501916885376)),(to_sfixed_a(-1.1629544133029412e-05)),(to_sfixed_a(-0.0001893956505227834)),(to_sfixed_a(3.174980156472884e-05)),(to_sfixed_a(-3.631991785368882e-05)),(to_sfixed_a(-4.69828701170627e-05)),(to_sfixed_a(-0.00015706574777141213)),(to_sfixed_a(-0.0014833708992227912)),(to_sfixed_a(-0.032647423446178436)),(to_sfixed_a(-0.2188737988471985)),(to_sfixed_a(-0.0643918588757515)),(to_sfixed_a(-0.17128100991249084)),(to_sfixed_a(-0.36804261803627014)),(to_sfixed_a(-0.00767596485093236)),(to_sfixed_a(-0.019706353545188904)),(to_sfixed_a(0.48810893297195435)),(to_sfixed_a(0.03681546077132225)),(to_sfixed_a(-0.2312328964471817)),(to_sfixed_a(-0.10126235336065292)),(to_sfixed_a(0.10087919980287552)),(to_sfixed_a(-0.02715328149497509)),(to_sfixed_a(0.0007275156094692647)),(to_sfixed_a(-0.12268061190843582)),(to_sfixed_a(-0.14974187314510345)),(to_sfixed_a(-0.10698059946298599)),(to_sfixed_a(0.049632806330919266)),(to_sfixed_a(0.06102645397186279)),(to_sfixed_a(0.005458198953419924)),(to_sfixed_a(0.11375253647565842)),(to_sfixed_a(0.004044783301651478)),(to_sfixed_a(0.00021633283176925033)),(to_sfixed_a(0.00018734965124167502)),(to_sfixed_a(-0.0003810665803030133)),(to_sfixed_a(0.0003691662277560681)),(to_sfixed_a(-0.00010483829828444868)),(to_sfixed_a(-0.0011083156568929553)),(to_sfixed_a(-0.13844366371631622)),(to_sfixed_a(-0.08157704770565033)),(to_sfixed_a(-0.07091313600540161)),(to_sfixed_a(-0.06737511605024338)),(to_sfixed_a(-0.08803393691778183)),(to_sfixed_a(-0.025648219510912895)),(to_sfixed_a(0.5388931632041931)),(to_sfixed_a(0.4178816080093384)),(to_sfixed_a(-0.33748528361320496)),(to_sfixed_a(-0.29303741455078125)),(to_sfixed_a(0.09794038534164429)),(to_sfixed_a(0.1408233493566513)),(to_sfixed_a(0.12836116552352905)),(to_sfixed_a(0.15054838359355927)),(to_sfixed_a(0.05492695793509483)),(to_sfixed_a(-0.05959991738200188)),(to_sfixed_a(-0.17122958600521088)),(to_sfixed_a(0.18659572303295135)),(to_sfixed_a(-0.0737842470407486)),(to_sfixed_a(0.007300824858248234)),(to_sfixed_a(0.00013113624299876392)),(to_sfixed_a(3.540153556969017e-05)),(to_sfixed_a(-0.00017258884327020496)),(to_sfixed_a(-0.0001052966108545661)),(to_sfixed_a(0.00014917201770003885)),(to_sfixed_a(-0.00012606554082594812)),(to_sfixed_a(-0.00037051516119390726)),(to_sfixed_a(-0.030728435143828392)),(to_sfixed_a(0.21342472732067108)),(to_sfixed_a(0.00815459992736578)),(to_sfixed_a(-0.12280898541212082)),(to_sfixed_a(0.033752404153347015)),(to_sfixed_a(0.17186802625656128)),(to_sfixed_a(0.22634673118591309)),(to_sfixed_a(0.17981590330600739)),(to_sfixed_a(-0.14918121695518494)),(to_sfixed_a(-0.05173066258430481)),(to_sfixed_a(-0.2587861716747284)),(to_sfixed_a(0.13616099953651428)),(to_sfixed_a(0.03891398757696152)),(to_sfixed_a(0.22204385697841644)),(to_sfixed_a(-0.2704767882823944)),(to_sfixed_a(0.08747927099466324)),(to_sfixed_a(-0.044250261038541794)),(to_sfixed_a(0.13448596000671387)),(to_sfixed_a(0.24371473491191864)),(to_sfixed_a(0.05768685042858124)),(to_sfixed_a(0.10864879190921783)),(to_sfixed_a(0.01910378970205784)),(to_sfixed_a(-0.0001800694881239906)),(to_sfixed_a(-0.00016349439101759344)),(to_sfixed_a(-0.00031388079514726996)),(to_sfixed_a(8.694858843227848e-05)),(to_sfixed_a(5.739698463003151e-05)),(to_sfixed_a(0.0002500567934475839)),(to_sfixed_a(0.0894043818116188)),(to_sfixed_a(-0.006746968720108271)),(to_sfixed_a(0.16227740049362183)),(to_sfixed_a(-0.07351767271757126)),(to_sfixed_a(0.12893052399158478)),(to_sfixed_a(0.23518356680870056)),(to_sfixed_a(0.020952468737959862)),(to_sfixed_a(-0.2750716805458069)),(to_sfixed_a(-0.3144437074661255)),(to_sfixed_a(-0.19451139867305756)),(to_sfixed_a(-0.21461671590805054)),(to_sfixed_a(0.3668938875198364)),(to_sfixed_a(0.756160318851471)),(to_sfixed_a(0.2101086676120758)),(to_sfixed_a(0.1580881029367447)),(to_sfixed_a(0.018169013783335686)),(to_sfixed_a(-0.03774334862828255)),(to_sfixed_a(0.03181303292512894)),(to_sfixed_a(0.21589277684688568)),(to_sfixed_a(0.051326096057891846)),(to_sfixed_a(0.019808296114206314)),(to_sfixed_a(-7.613520665472606e-06)),(to_sfixed_a(7.031505083432421e-05)),(to_sfixed_a(-5.301924466039054e-05)),(to_sfixed_a(0.00018684571841731668)),(to_sfixed_a(4.607573828252498e-06)),(to_sfixed_a(-3.0261235224315897e-05)),(to_sfixed_a(-9.292030154028907e-05)),(to_sfixed_a(-5.8062909374712035e-05)),(to_sfixed_a(-0.002416193252429366)),(to_sfixed_a(0.028217315673828125)),(to_sfixed_a(0.05299413204193115)),(to_sfixed_a(0.25516611337661743)),(to_sfixed_a(0.24369241297245026)),(to_sfixed_a(0.004293885547667742)),(to_sfixed_a(-0.0825834795832634)),(to_sfixed_a(0.057695422321558)),(to_sfixed_a(-0.05922180786728859)),(to_sfixed_a(0.009409132413566113)),(to_sfixed_a(0.28752145171165466)),(to_sfixed_a(0.1111779436469078)),(to_sfixed_a(0.07617012411355972)),(to_sfixed_a(-0.17222654819488525)),(to_sfixed_a(0.2592545449733734)),(to_sfixed_a(0.39945533871650696)),(to_sfixed_a(0.17582322657108307)),(to_sfixed_a(0.057563066482543945)),(to_sfixed_a(-0.040771838277578354)),(to_sfixed_a(0.054672569036483765)),(to_sfixed_a(0.1158294677734375)),(to_sfixed_a(4.279269705875777e-05)),(to_sfixed_a(0.0001231827773153782)),(to_sfixed_a(-3.5399276384850964e-05)),(to_sfixed_a(0.00023728428641334176)),(to_sfixed_a(0.00014850535080768168)),(to_sfixed_a(0.0003101486654486507)),(to_sfixed_a(0.0003071025130338967)),(to_sfixed_a(0.047635409981012344)),(to_sfixed_a(-0.0009059527073986828)),(to_sfixed_a(0.14308686554431915)),(to_sfixed_a(0.3124163746833801)),(to_sfixed_a(0.19367516040802002)),(to_sfixed_a(0.23082362115383148)),(to_sfixed_a(0.04601246118545532)),(to_sfixed_a(0.08142058551311493)),(to_sfixed_a(0.2990611493587494)),(to_sfixed_a(-0.04802998527884483)),(to_sfixed_a(0.003225217340514064)),(to_sfixed_a(0.27020856738090515)),(to_sfixed_a(0.06319290399551392)),(to_sfixed_a(0.0662543848156929)),(to_sfixed_a(0.050691794604063034)),(to_sfixed_a(0.20332379639148712)),(to_sfixed_a(0.011294681578874588)),(to_sfixed_a(0.08978643268346786)),(to_sfixed_a(0.09332656115293503)),(to_sfixed_a(-0.00042652583215385675)),(to_sfixed_a(0.08686570078134537)),(to_sfixed_a(-2.7247144316788763e-05)),(to_sfixed_a(5.863655678695068e-05)),(to_sfixed_a(1.2722657629637979e-05)),(to_sfixed_a(-0.00026199896819889545)),(to_sfixed_a(-0.00012262279051356018)),(to_sfixed_a(0.00018472182273399085)),(to_sfixed_a(0.0001741239393595606)),(to_sfixed_a(0.00021675755851902068)),(to_sfixed_a(0.07094763219356537)),(to_sfixed_a(0.15589365363121033)),(to_sfixed_a(0.24111966788768768)),(to_sfixed_a(0.10959069430828094)),(to_sfixed_a(0.1823153793811798)),(to_sfixed_a(0.3833235800266266)),(to_sfixed_a(0.15397927165031433)),(to_sfixed_a(0.1015777587890625)),(to_sfixed_a(0.028808949515223503)),(to_sfixed_a(-0.22240018844604492)),(to_sfixed_a(-0.010153520852327347)),(to_sfixed_a(-0.1530027687549591)),(to_sfixed_a(0.2005954533815384)),(to_sfixed_a(0.3085747957229614)),(to_sfixed_a(-0.048343054950237274)),(to_sfixed_a(0.1327214539051056)),(to_sfixed_a(0.027438385412096977)),(to_sfixed_a(0.10672654211521149)),(to_sfixed_a(0.003760252147912979)),(to_sfixed_a(0.00018476371769793332)),(to_sfixed_a(1.3483213479048572e-05)),(to_sfixed_a(0.00013174180639907718)),(to_sfixed_a(0.00019983641686849296)),(to_sfixed_a(0.0001453140430385247)),(to_sfixed_a(4.239277041051537e-05)),(to_sfixed_a(0.0002706707746256143)),(to_sfixed_a(0.00012119076563976705)),(to_sfixed_a(0.00019786180928349495)),(to_sfixed_a(0.02773360162973404)),(to_sfixed_a(-0.08054888248443604)),(to_sfixed_a(0.22224459052085876)),(to_sfixed_a(0.29793983697891235)),(to_sfixed_a(0.22019197046756744)),(to_sfixed_a(0.09426150470972061)),(to_sfixed_a(0.19146116077899933)),(to_sfixed_a(0.1020229309797287)),(to_sfixed_a(-0.1301874816417694)),(to_sfixed_a(-0.14816470444202423)),(to_sfixed_a(0.01979791186749935)),(to_sfixed_a(0.0005849472945556045)),(to_sfixed_a(-0.20958808064460754)),(to_sfixed_a(-0.16377735137939453)),(to_sfixed_a(-0.050815775990486145)),(to_sfixed_a(-0.0698978453874588)),(to_sfixed_a(0.029812905937433243)),(to_sfixed_a(0.0052328286692500114)),(to_sfixed_a(0.016616079956293106)),(to_sfixed_a(-1.3356570889300201e-06)),(to_sfixed_a(-5.6278135161846876e-05)),(to_sfixed_a(0.00020075486099813133)),(to_sfixed_a(-0.00013168003351893276)),(to_sfixed_a(-8.55769121699268e-06)),(to_sfixed_a(-0.000295473902951926)),(to_sfixed_a(0.0003887325874529779)),(to_sfixed_a(-6.615422898903489e-05)),(to_sfixed_a(-0.013184072449803352)),(to_sfixed_a(-0.0712476298213005)),(to_sfixed_a(-0.051932428032159805)),(to_sfixed_a(0.006244229152798653)),(to_sfixed_a(0.17485782504081726)),(to_sfixed_a(0.10087443888187408)),(to_sfixed_a(0.3733340799808502)),(to_sfixed_a(0.2537907063961029)),(to_sfixed_a(-0.34603509306907654)),(to_sfixed_a(-0.18836069107055664)),(to_sfixed_a(0.09282767027616501)),(to_sfixed_a(0.06712095439434052)),(to_sfixed_a(-0.009742776863276958)),(to_sfixed_a(0.3036579489707947)),(to_sfixed_a(-0.01959482952952385)),(to_sfixed_a(-0.04342379793524742)),(to_sfixed_a(0.012473798356950283)),(to_sfixed_a(0.018606994301080704)),(to_sfixed_a(0.011011305265128613)),(to_sfixed_a(0.0017819245113059878)),(to_sfixed_a(-5.968545792711666e-06)),(to_sfixed_a(7.861172343837097e-05)),(to_sfixed_a(2.165725345548708e-05)),(to_sfixed_a(0.00016522292571607977)),(to_sfixed_a(2.753716216830071e-05)),(to_sfixed_a(4.531348167802207e-05)),(to_sfixed_a(9.576133379596286e-06)),(to_sfixed_a(0.0002599830331746489)),(to_sfixed_a(7.061076757963747e-05)),(to_sfixed_a(-0.03165000304579735)),(to_sfixed_a(-0.03248807415366173)),(to_sfixed_a(-0.0043996055610477924)),(to_sfixed_a(-0.3377513587474823)),(to_sfixed_a(-0.14914950728416443)),(to_sfixed_a(0.07762279361486435)),(to_sfixed_a(-0.05242540314793587)),(to_sfixed_a(0.106300950050354)),(to_sfixed_a(0.06904994696378708)),(to_sfixed_a(-0.13016390800476074)),(to_sfixed_a(-0.16735821962356567)),(to_sfixed_a(0.035420551896095276)),(to_sfixed_a(-0.04737760126590729)),(to_sfixed_a(-0.01289138663560152)),(to_sfixed_a(-0.14020030200481415)),(to_sfixed_a(-0.06974051147699356)),(to_sfixed_a(-0.000548133160918951)),(to_sfixed_a(-0.00042167652281932533)),(to_sfixed_a(0.0001254135713679716)),(to_sfixed_a(-4.3761083361459896e-05)),(to_sfixed_a(0.0003141329507343471)),(to_sfixed_a(-0.00022994093887973577)),(to_sfixed_a(-0.00017638782446738333)),(to_sfixed_a(-8.89177099452354e-05)),(to_sfixed_a(-2.785242031677626e-05)),(to_sfixed_a(-5.015060378354974e-05)),(to_sfixed_a(-0.00028742002905346453)),(to_sfixed_a(1.090240493795136e-05)),(to_sfixed_a(-7.142903632484376e-05)),(to_sfixed_a(-6.663436215603724e-05)),(to_sfixed_a(0.00024347196449525654)),(to_sfixed_a(0.00011791151337092742)),(to_sfixed_a(0.0008296800660900772)),(to_sfixed_a(-0.08391176164150238)),(to_sfixed_a(0.0005524176522158086)),(to_sfixed_a(-0.00048804463585838675)),(to_sfixed_a(-0.06439611315727234)),(to_sfixed_a(-0.06678769737482071)),(to_sfixed_a(-0.005072818603366613)),(to_sfixed_a(-0.04698231816291809)),(to_sfixed_a(-0.06597322970628738)),(to_sfixed_a(-0.08731404691934586)),(to_sfixed_a(0.002182522090151906)),(to_sfixed_a(0.00014250889944378287)),(to_sfixed_a(0.0001151472024503164)),(to_sfixed_a(-6.546660733874887e-05)),(to_sfixed_a(-0.00010516562178963795)),(to_sfixed_a(-0.00013584730913862586)),(to_sfixed_a(0.00015576693112961948)),(to_sfixed_a(6.284578557824716e-05)),(to_sfixed_a(7.866094529163092e-05)),(to_sfixed_a(2.4705504984012805e-05)),(to_sfixed_a(-0.00019666059233713895)),(to_sfixed_a(-0.0003572080167941749)),(to_sfixed_a(-0.00018646343960426748)),(to_sfixed_a(-8.651513053337112e-05)),(to_sfixed_a(9.430647332919762e-05)),(to_sfixed_a(-8.732209971640259e-05)),(to_sfixed_a(-2.2814076146460138e-05)),(to_sfixed_a(0.0001032911823131144)),(to_sfixed_a(0.0001607670565135777)),(to_sfixed_a(0.00013769393262919039)),(to_sfixed_a(-0.00010043574729934335)),(to_sfixed_a(-5.868360312888399e-05)),(to_sfixed_a(8.780907228356227e-05)),(to_sfixed_a(2.7924526875722222e-05)),(to_sfixed_a(-3.038633440155536e-05)),(to_sfixed_a(6.163139914860949e-05)),(to_sfixed_a(2.0852092347922735e-05)),(to_sfixed_a(-2.4743329049670137e-05)),(to_sfixed_a(-1.905432691273745e-05)),(to_sfixed_a(-0.00017731636762619019)),(to_sfixed_a(-0.0003132343990728259)),(to_sfixed_a(-2.0540514015010558e-05)),(to_sfixed_a(-0.0001315821282332763)),(to_sfixed_a(-0.00038543681148439646)),(to_sfixed_a(0.00011958016693824902)),(to_sfixed_a(8.375260222237557e-05)),(to_sfixed_a(0.0002215387939941138)));

    constant weight_n0_18 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-0.0004131252062506974)),(to_sfixed_a(-5.9689169574994594e-05)),(to_sfixed_a(-1.0034118531621061e-05)),(to_sfixed_a(6.989094981690869e-05)),(to_sfixed_a(-0.00021854968508705497)),(to_sfixed_a(0.00014341663336381316)),(to_sfixed_a(0.0003567337989807129)),(to_sfixed_a(0.0001624298165552318)),(to_sfixed_a(5.625849371426739e-05)),(to_sfixed_a(-2.5765255486476235e-05)),(to_sfixed_a(-8.525962039129809e-05)),(to_sfixed_a(-0.00011791804718086496)),(to_sfixed_a(4.838125823880546e-05)),(to_sfixed_a(-0.00021095392003189772)),(to_sfixed_a(0.00022724394511897117)),(to_sfixed_a(-8.380604413105175e-05)),(to_sfixed_a(-0.00013967056293040514)),(to_sfixed_a(-0.0001587651640875265)),(to_sfixed_a(3.3700125641189516e-05)),(to_sfixed_a(-0.00012768726446665823)),(to_sfixed_a(0.00010952126467600465)),(to_sfixed_a(0.0002678142045624554)),(to_sfixed_a(-0.0002458615635987371)),(to_sfixed_a(-0.00018101828754879534)),(to_sfixed_a(5.0622802518773824e-05)),(to_sfixed_a(8.244071068475023e-05)),(to_sfixed_a(5.7777589972829446e-05)),(to_sfixed_a(-5.580649303738028e-05)),(to_sfixed_a(-4.8387653805548325e-05)),(to_sfixed_a(-7.03157638781704e-05)),(to_sfixed_a(1.0010814548877534e-05)),(to_sfixed_a(0.00010593482875265181)),(to_sfixed_a(0.00010271898645441979)),(to_sfixed_a(-0.00011189474753336981)),(to_sfixed_a(0.00021171553817112)),(to_sfixed_a(-0.00012885684554930776)),(to_sfixed_a(4.984725819667801e-05)),(to_sfixed_a(-0.00015364520368166268)),(to_sfixed_a(-0.00016243525897152722)),(to_sfixed_a(-4.6742925974285754e-07)),(to_sfixed_a(1.518897624919191e-05)),(to_sfixed_a(0.0001582190889166668)),(to_sfixed_a(0.00027082572341896594)),(to_sfixed_a(8.793703455012292e-05)),(to_sfixed_a(7.378263399004936e-05)),(to_sfixed_a(4.624000212061219e-05)),(to_sfixed_a(9.376127127325162e-05)),(to_sfixed_a(-7.574972551083192e-05)),(to_sfixed_a(0.00020264825434423983)),(to_sfixed_a(0.00014486582949757576)),(to_sfixed_a(-6.047455099178478e-05)),(to_sfixed_a(-0.00018411071505397558)),(to_sfixed_a(-2.7588837838266045e-05)),(to_sfixed_a(-1.9917932149837725e-05)),(to_sfixed_a(0.00030585535569116473)),(to_sfixed_a(-6.761452095815912e-05)),(to_sfixed_a(2.4002943973755464e-05)),(to_sfixed_a(-7.57966045057401e-05)),(to_sfixed_a(3.576207745936699e-05)),(to_sfixed_a(0.00022899277973920107)),(to_sfixed_a(-0.0003620931238401681)),(to_sfixed_a(-0.00023421058722306043)),(to_sfixed_a(-0.0002395711198914796)),(to_sfixed_a(-5.7695244322530925e-05)),(to_sfixed_a(0.0002489352773409337)),(to_sfixed_a(5.048268212703988e-05)),(to_sfixed_a(-7.651200576219708e-05)),(to_sfixed_a(-0.00021910987561568618)),(to_sfixed_a(0.0002042827836703509)),(to_sfixed_a(0.03181326016783714)),(to_sfixed_a(-0.00012214973685331643)),(to_sfixed_a(4.5525754103437066e-05)),(to_sfixed_a(-0.0001417432795278728)),(to_sfixed_a(-0.00019011908443644643)),(to_sfixed_a(5.778607737738639e-05)),(to_sfixed_a(8.450807945337147e-05)),(to_sfixed_a(-6.469843356171623e-05)),(to_sfixed_a(3.4760989365167916e-05)),(to_sfixed_a(-6.321219552773982e-05)),(to_sfixed_a(-9.40486861509271e-05)),(to_sfixed_a(3.38151803589426e-05)),(to_sfixed_a(-0.0002356330369366333)),(to_sfixed_a(-0.00018666553660295904)),(to_sfixed_a(0.00010828206723090261)),(to_sfixed_a(1.6197984223254025e-05)),(to_sfixed_a(6.914266850799322e-05)),(to_sfixed_a(-0.0003587957180570811)),(to_sfixed_a(6.906013823027024e-06)),(to_sfixed_a(0.000158658716827631)),(to_sfixed_a(-7.211300544440746e-05)),(to_sfixed_a(7.09240703145042e-05)),(to_sfixed_a(-4.4902455556439236e-05)),(to_sfixed_a(0.05823671072721481)),(to_sfixed_a(-6.442479934776202e-05)),(to_sfixed_a(0.06626903265714645)),(to_sfixed_a(-0.007027315441519022)),(to_sfixed_a(0.16503717005252838)),(to_sfixed_a(0.15498754382133484)),(to_sfixed_a(0.08740902692079544)),(to_sfixed_a(-0.13801363110542297)),(to_sfixed_a(0.03735456243157387)),(to_sfixed_a(-0.12815925478935242)),(to_sfixed_a(0.1175212413072586)),(to_sfixed_a(-0.02544279582798481)),(to_sfixed_a(-0.04884316027164459)),(to_sfixed_a(-0.09927663207054138)),(to_sfixed_a(0.00013803470938000828)),(to_sfixed_a(-0.00011264226486673579)),(to_sfixed_a(1.5327900655393023e-06)),(to_sfixed_a(3.520843165460974e-05)),(to_sfixed_a(1.6059950212365948e-05)),(to_sfixed_a(-0.00015270750736817718)),(to_sfixed_a(-0.00032838163315318525)),(to_sfixed_a(-0.0001648114703129977)),(to_sfixed_a(-0.000235585801419802)),(to_sfixed_a(4.797062501893379e-05)),(to_sfixed_a(-7.2007474045676645e-06)),(to_sfixed_a(-1.6466334272990935e-05)),(to_sfixed_a(0.001311873784288764)),(to_sfixed_a(-0.0028522040229290724)),(to_sfixed_a(-0.06531447172164917)),(to_sfixed_a(0.08128337562084198)),(to_sfixed_a(0.3733212351799011)),(to_sfixed_a(0.17523455619812012)),(to_sfixed_a(0.25703829526901245)),(to_sfixed_a(0.21018055081367493)),(to_sfixed_a(0.14025135338306427)),(to_sfixed_a(-0.083006851375103)),(to_sfixed_a(-0.24334922432899475)),(to_sfixed_a(0.03099038638174534)),(to_sfixed_a(-0.15020370483398438)),(to_sfixed_a(-0.015006509609520435)),(to_sfixed_a(-0.0054026031866669655)),(to_sfixed_a(0.17759327590465546)),(to_sfixed_a(-0.0003608802508097142)),(to_sfixed_a(0.0008580653229728341)),(to_sfixed_a(-0.0020674520637840033)),(to_sfixed_a(6.477983697550371e-05)),(to_sfixed_a(-0.00016677696839906275)),(to_sfixed_a(3.67972970707342e-05)),(to_sfixed_a(-6.280008528847247e-05)),(to_sfixed_a(-5.556895848712884e-05)),(to_sfixed_a(0.00016216868243645877)),(to_sfixed_a(3.70551242667716e-05)),(to_sfixed_a(0.0012106855865567923)),(to_sfixed_a(-0.009476471692323685)),(to_sfixed_a(-0.0053803701885044575)),(to_sfixed_a(0.06832887977361679)),(to_sfixed_a(-0.023495933040976524)),(to_sfixed_a(0.09118068963289261)),(to_sfixed_a(0.15477976202964783)),(to_sfixed_a(0.03807070851325989)),(to_sfixed_a(0.04829883202910423)),(to_sfixed_a(0.04515216127038002)),(to_sfixed_a(0.04328940436244011)),(to_sfixed_a(-0.0816582515835762)),(to_sfixed_a(0.07753048092126846)),(to_sfixed_a(0.09561952203512192)),(to_sfixed_a(-0.45534875988960266)),(to_sfixed_a(-0.17819467186927795)),(to_sfixed_a(-0.07007931172847748)),(to_sfixed_a(-0.2020823210477829)),(to_sfixed_a(-0.0019062302308157086)),(to_sfixed_a(-0.07768338173627853)),(to_sfixed_a(-0.00036055201780982316)),(to_sfixed_a(-7.897846808191389e-05)),(to_sfixed_a(-0.0002536489046178758)),(to_sfixed_a(0.00021131712128408253)),(to_sfixed_a(-0.00020277200383134186)),(to_sfixed_a(-0.00012010436330456287)),(to_sfixed_a(-8.22033325675875e-05)),(to_sfixed_a(2.4114469852065668e-05)),(to_sfixed_a(0.0004554619954433292)),(to_sfixed_a(-0.008888855576515198)),(to_sfixed_a(-0.020891154184937477)),(to_sfixed_a(0.1180809736251831)),(to_sfixed_a(0.04287772625684738)),(to_sfixed_a(0.019469408318400383)),(to_sfixed_a(0.17734242975711823)),(to_sfixed_a(0.17184068262577057)),(to_sfixed_a(-0.0734642893075943)),(to_sfixed_a(-0.16900628805160522)),(to_sfixed_a(-0.1709882915019989)),(to_sfixed_a(-0.21929898858070374)),(to_sfixed_a(-0.15070675313472748)),(to_sfixed_a(-0.1565386950969696)),(to_sfixed_a(-0.19829262793064117)),(to_sfixed_a(-0.3564956486225128)),(to_sfixed_a(-0.3600179851055145)),(to_sfixed_a(-0.15184219181537628)),(to_sfixed_a(-0.08147913217544556)),(to_sfixed_a(0.03766552358865738)),(to_sfixed_a(0.0006464689504355192)),(to_sfixed_a(0.0001495715550845489)),(to_sfixed_a(-0.0008446324500255287)),(to_sfixed_a(-3.8374131690943614e-05)),(to_sfixed_a(9.133133426075801e-05)),(to_sfixed_a(-0.0002510701597202569)),(to_sfixed_a(-0.00010295533138560131)),(to_sfixed_a(2.322804539289791e-05)),(to_sfixed_a(9.140264592133462e-05)),(to_sfixed_a(-0.019625267013907433)),(to_sfixed_a(-0.02794182114303112)),(to_sfixed_a(0.13876959681510925)),(to_sfixed_a(-0.2409633994102478)),(to_sfixed_a(-0.13695304095745087)),(to_sfixed_a(0.3384736180305481)),(to_sfixed_a(-0.024137135595083237)),(to_sfixed_a(-0.11912595480680466)),(to_sfixed_a(-0.046850331127643585)),(to_sfixed_a(-0.1768280416727066)),(to_sfixed_a(-0.24733518064022064)),(to_sfixed_a(0.051835160702466965)),(to_sfixed_a(-0.014528801664710045)),(to_sfixed_a(-0.21436463296413422)),(to_sfixed_a(-0.5152084231376648)),(to_sfixed_a(-0.02866542711853981)),(to_sfixed_a(-0.2567073702812195)),(to_sfixed_a(0.006200065370649099)),(to_sfixed_a(-0.019338587298989296)),(to_sfixed_a(0.11135293543338776)),(to_sfixed_a(0.004897229839116335)),(to_sfixed_a(0.00010825737263076007)),(to_sfixed_a(0.0001411461125826463)),(to_sfixed_a(1.0315573490515817e-05)),(to_sfixed_a(-9.934024274116382e-05)),(to_sfixed_a(-1.1451879800006282e-05)),(to_sfixed_a(7.938370254123583e-05)),(to_sfixed_a(-0.07043550163507462)),(to_sfixed_a(0.06489542871713638)),(to_sfixed_a(0.0033281929790973663)),(to_sfixed_a(0.14404529333114624)),(to_sfixed_a(0.12377727031707764)),(to_sfixed_a(0.09289529174566269)),(to_sfixed_a(0.4001569151878357)),(to_sfixed_a(0.11238215118646622)),(to_sfixed_a(0.025736959651112556)),(to_sfixed_a(-0.27040454745292664)),(to_sfixed_a(-0.006799250841140747)),(to_sfixed_a(0.04864473268389702)),(to_sfixed_a(-0.06294435262680054)),(to_sfixed_a(-0.22947539389133453)),(to_sfixed_a(-0.19357895851135254)),(to_sfixed_a(-0.15056651830673218)),(to_sfixed_a(0.0014042105758562684)),(to_sfixed_a(0.09851650148630142)),(to_sfixed_a(-0.1114882081747055)),(to_sfixed_a(0.02005680277943611)),(to_sfixed_a(0.1590748131275177)),(to_sfixed_a(0.010692440904676914)),(to_sfixed_a(-0.00011480885586934164)),(to_sfixed_a(7.497121987398714e-05)),(to_sfixed_a(-0.00034253785270266235)),(to_sfixed_a(-0.0002004448906518519)),(to_sfixed_a(7.16063950676471e-05)),(to_sfixed_a(2.202674477302935e-05)),(to_sfixed_a(0.003043955657631159)),(to_sfixed_a(-0.004986136220395565)),(to_sfixed_a(0.04636291787028313)),(to_sfixed_a(0.081695057451725)),(to_sfixed_a(0.06150677427649498)),(to_sfixed_a(0.09199657291173935)),(to_sfixed_a(0.2754685580730438)),(to_sfixed_a(0.1562040150165558)),(to_sfixed_a(0.10407701134681702)),(to_sfixed_a(-0.25771111249923706)),(to_sfixed_a(-0.03702719509601593)),(to_sfixed_a(-0.25432077050209045)),(to_sfixed_a(-0.5307989716529846)),(to_sfixed_a(-0.2147616446018219)),(to_sfixed_a(-0.3258790373802185)),(to_sfixed_a(0.08149135857820511)),(to_sfixed_a(0.22775700688362122)),(to_sfixed_a(0.003557795425876975)),(to_sfixed_a(-0.017999034374952316)),(to_sfixed_a(0.3954789340496063)),(to_sfixed_a(0.2599736750125885)),(to_sfixed_a(-0.0002181049931095913)),(to_sfixed_a(0.00010240300616715103)),(to_sfixed_a(5.180769949220121e-05)),(to_sfixed_a(-1.3887733985029627e-05)),(to_sfixed_a(-3.427842239034362e-05)),(to_sfixed_a(0.0001925620890688151)),(to_sfixed_a(-0.0002571591467130929)),(to_sfixed_a(0.004057872574776411)),(to_sfixed_a(0.0014597260160371661)),(to_sfixed_a(-0.0840248391032219)),(to_sfixed_a(0.01864033006131649)),(to_sfixed_a(-0.02461829036474228)),(to_sfixed_a(0.09020224958658218)),(to_sfixed_a(0.16361011564731598)),(to_sfixed_a(0.2151932567358017)),(to_sfixed_a(-0.02692609280347824)),(to_sfixed_a(0.02036348730325699)),(to_sfixed_a(-0.10604701191186905)),(to_sfixed_a(-0.22793696820735931)),(to_sfixed_a(-0.21652202308177948)),(to_sfixed_a(-0.31780412793159485)),(to_sfixed_a(-0.3122817277908325)),(to_sfixed_a(-0.26581835746765137)),(to_sfixed_a(0.0156408604234457)),(to_sfixed_a(0.24659891426563263)),(to_sfixed_a(0.018188998103141785)),(to_sfixed_a(0.18877725303173065)),(to_sfixed_a(0.1272488236427307)),(to_sfixed_a(0.05493567883968353)),(to_sfixed_a(4.9868318455992267e-05)),(to_sfixed_a(-1.16658575279871e-05)),(to_sfixed_a(-0.0002544928574934602)),(to_sfixed_a(-0.00030825036810711026)),(to_sfixed_a(0.00025206603459082544)),(to_sfixed_a(0.00012136580335209146)),(to_sfixed_a(-0.034631673246622086)),(to_sfixed_a(0.04084921255707741)),(to_sfixed_a(-0.05651887133717537)),(to_sfixed_a(0.05194410681724548)),(to_sfixed_a(-0.09364677220582962)),(to_sfixed_a(0.09090033918619156)),(to_sfixed_a(-0.0316266193985939)),(to_sfixed_a(0.13945545256137848)),(to_sfixed_a(0.008327987976372242)),(to_sfixed_a(0.3944523334503174)),(to_sfixed_a(-0.035707987844944)),(to_sfixed_a(0.33694344758987427)),(to_sfixed_a(0.17595848441123962)),(to_sfixed_a(-0.020067157223820686)),(to_sfixed_a(-0.0411575548350811)),(to_sfixed_a(-0.21821458637714386)),(to_sfixed_a(-0.29413971304893494)),(to_sfixed_a(-0.05594580993056297)),(to_sfixed_a(0.16242165863513947)),(to_sfixed_a(0.1373887062072754)),(to_sfixed_a(0.12757085263729095)),(to_sfixed_a(-0.0001238896802533418)),(to_sfixed_a(4.4857009925181046e-05)),(to_sfixed_a(-7.013927097432315e-05)),(to_sfixed_a(-4.4884094677399844e-05)),(to_sfixed_a(1.1185019502590876e-05)),(to_sfixed_a(-7.3125320341205224e-06)),(to_sfixed_a(2.43985286942916e-05)),(to_sfixed_a(0.05854853615164757)),(to_sfixed_a(-0.2139746993780136)),(to_sfixed_a(-0.0027188907843083143)),(to_sfixed_a(-0.08367915451526642)),(to_sfixed_a(-0.07202144712209702)),(to_sfixed_a(-0.11979462951421738)),(to_sfixed_a(0.14303253591060638)),(to_sfixed_a(0.01673109643161297)),(to_sfixed_a(0.024137208238244057)),(to_sfixed_a(0.1816164255142212)),(to_sfixed_a(0.2717079520225525)),(to_sfixed_a(0.731560230255127)),(to_sfixed_a(0.36397838592529297)),(to_sfixed_a(-0.15091249346733093)),(to_sfixed_a(-0.16000232100486755)),(to_sfixed_a(-0.04496913030743599)),(to_sfixed_a(-0.25178200006484985)),(to_sfixed_a(-0.06809017062187195)),(to_sfixed_a(-0.10668903589248657)),(to_sfixed_a(0.272137314081192)),(to_sfixed_a(0.08803273737430573)),(to_sfixed_a(2.8779970307368785e-05)),(to_sfixed_a(0.0003110539400950074)),(to_sfixed_a(3.685984847834334e-05)),(to_sfixed_a(0.00023691763635724783)),(to_sfixed_a(0.00011883345723617822)),(to_sfixed_a(0.00010503120574867353)),(to_sfixed_a(3.1703602871857584e-06)),(to_sfixed_a(-0.03464128449559212)),(to_sfixed_a(0.055792659521102905)),(to_sfixed_a(0.03175193816423416)),(to_sfixed_a(0.057873062789440155)),(to_sfixed_a(0.05640048161149025)),(to_sfixed_a(0.045033734291791916)),(to_sfixed_a(0.04907778277993202)),(to_sfixed_a(0.18220682442188263)),(to_sfixed_a(0.029834622517228127)),(to_sfixed_a(-0.09577307105064392)),(to_sfixed_a(0.08725549280643463)),(to_sfixed_a(0.15999986231327057)),(to_sfixed_a(0.018771246075630188)),(to_sfixed_a(-0.06935649365186691)),(to_sfixed_a(-0.12103331834077835)),(to_sfixed_a(-0.4493255913257599)),(to_sfixed_a(0.020221032202243805)),(to_sfixed_a(0.1096939966082573)),(to_sfixed_a(0.1304701864719391)),(to_sfixed_a(0.1470734030008316)),(to_sfixed_a(0.07496669143438339)),(to_sfixed_a(0.001195334130898118)),(to_sfixed_a(0.002060066210106015)),(to_sfixed_a(-9.308962762588635e-05)),(to_sfixed_a(-0.00012326051364652812)),(to_sfixed_a(-0.00027555596898309886)),(to_sfixed_a(-0.0001904335367726162)),(to_sfixed_a(0.00023328869428951293)),(to_sfixed_a(-2.9270864615682513e-05)),(to_sfixed_a(0.04849721118807793)),(to_sfixed_a(-0.007599144242703915)),(to_sfixed_a(-0.08632059395313263)),(to_sfixed_a(-0.09271770715713501)),(to_sfixed_a(0.08959075063467026)),(to_sfixed_a(0.1267978549003601)),(to_sfixed_a(0.26352718472480774)),(to_sfixed_a(0.026563052088022232)),(to_sfixed_a(0.02021712437272072)),(to_sfixed_a(-0.10815601795911789)),(to_sfixed_a(0.09939311444759369)),(to_sfixed_a(-0.2880970239639282)),(to_sfixed_a(-0.10483840852975845)),(to_sfixed_a(0.03431880101561546)),(to_sfixed_a(-0.3380584716796875)),(to_sfixed_a(-0.18409807980060577)),(to_sfixed_a(-0.011538345366716385)),(to_sfixed_a(0.1371624916791916)),(to_sfixed_a(-0.19507300853729248)),(to_sfixed_a(0.020540833473205566)),(to_sfixed_a(-0.0003830795467365533)),(to_sfixed_a(-7.269137859111652e-05)),(to_sfixed_a(0.0001547423016745597)),(to_sfixed_a(-0.00029002930386923254)),(to_sfixed_a(4.8398852925402025e-08)),(to_sfixed_a(-0.00015653081936761737)),(to_sfixed_a(-9.548707021167502e-05)),(to_sfixed_a(-0.03971020132303238)),(to_sfixed_a(0.07470588386058807)),(to_sfixed_a(0.08645115792751312)),(to_sfixed_a(0.13049226999282837)),(to_sfixed_a(0.1294269859790802)),(to_sfixed_a(0.1844547539949417)),(to_sfixed_a(0.25296929478645325)),(to_sfixed_a(-0.07400110363960266)),(to_sfixed_a(-0.14155136048793793)),(to_sfixed_a(-0.020645873621106148)),(to_sfixed_a(0.030373279005289078)),(to_sfixed_a(0.05199764296412468)),(to_sfixed_a(-0.0696137398481369)),(to_sfixed_a(-0.052064523100852966)),(to_sfixed_a(-0.2601368725299835)),(to_sfixed_a(-0.28140363097190857)),(to_sfixed_a(-0.3238056004047394)),(to_sfixed_a(-0.00971432775259018)),(to_sfixed_a(0.17084769904613495)),(to_sfixed_a(-0.07042552530765533)),(to_sfixed_a(-0.18725666403770447)),(to_sfixed_a(-0.0004904379020445049)),(to_sfixed_a(0.00038529557059518993)),(to_sfixed_a(0.0002168565260944888)),(to_sfixed_a(-5.5181873904075474e-05)),(to_sfixed_a(0.00018721510423347354)),(to_sfixed_a(0.00017895811470225453)),(to_sfixed_a(9.718840738059953e-05)),(to_sfixed_a(0.16617806255817413)),(to_sfixed_a(0.1628653109073639)),(to_sfixed_a(0.11971018463373184)),(to_sfixed_a(-0.153485506772995)),(to_sfixed_a(0.09740856289863586)),(to_sfixed_a(-0.04952499270439148)),(to_sfixed_a(0.020983979105949402)),(to_sfixed_a(0.13742350041866302)),(to_sfixed_a(-0.3376990556716919)),(to_sfixed_a(-0.37469202280044556)),(to_sfixed_a(-0.18355083465576172)),(to_sfixed_a(-0.17781753838062286)),(to_sfixed_a(-0.15034279227256775)),(to_sfixed_a(-0.268667608499527)),(to_sfixed_a(-0.2318749725818634)),(to_sfixed_a(-0.09377237409353256)),(to_sfixed_a(-0.33318081498146057)),(to_sfixed_a(-0.23612938821315765)),(to_sfixed_a(0.0034202421084046364)),(to_sfixed_a(-0.07322259992361069)),(to_sfixed_a(-0.017695961520075798)),(to_sfixed_a(0.0019565674010664225)),(to_sfixed_a(-8.753530710237101e-05)),(to_sfixed_a(-0.00014666907372884452)),(to_sfixed_a(0.0002702728961594403)),(to_sfixed_a(-5.235395292402245e-05)),(to_sfixed_a(-0.0004950827569700778)),(to_sfixed_a(-6.272680911934003e-05)),(to_sfixed_a(0.037360645830631256)),(to_sfixed_a(0.10263147950172424)),(to_sfixed_a(-0.04984329268336296)),(to_sfixed_a(0.014868772588670254)),(to_sfixed_a(-0.1312323659658432)),(to_sfixed_a(0.05704505369067192)),(to_sfixed_a(0.21541157364845276)),(to_sfixed_a(0.01781802996993065)),(to_sfixed_a(-0.327210396528244)),(to_sfixed_a(-0.062049299478530884)),(to_sfixed_a(-0.13164456188678741)),(to_sfixed_a(-0.23454906046390533)),(to_sfixed_a(-0.046952761709690094)),(to_sfixed_a(-0.18839997053146362)),(to_sfixed_a(-0.01873418129980564)),(to_sfixed_a(-0.18371756374835968)),(to_sfixed_a(0.11167198419570923)),(to_sfixed_a(0.06878509372472763)),(to_sfixed_a(-0.03651316836476326)),(to_sfixed_a(-0.018659980967640877)),(to_sfixed_a(4.633648495655507e-05)),(to_sfixed_a(0.0001382543268846348)),(to_sfixed_a(-7.735039253020659e-05)),(to_sfixed_a(0.0002205640630563721)),(to_sfixed_a(0.00012190996494609863)),(to_sfixed_a(0.00013962865341454744)),(to_sfixed_a(0.000133552064653486)),(to_sfixed_a(-0.017239771783351898)),(to_sfixed_a(-0.18740934133529663)),(to_sfixed_a(-0.2782876193523407)),(to_sfixed_a(-0.09300174564123154)),(to_sfixed_a(0.1906493902206421)),(to_sfixed_a(0.21012653410434723)),(to_sfixed_a(0.05374467372894287)),(to_sfixed_a(0.08949653059244156)),(to_sfixed_a(-0.13394103944301605)),(to_sfixed_a(-0.2776736319065094)),(to_sfixed_a(-0.46591341495513916)),(to_sfixed_a(-0.2684456706047058)),(to_sfixed_a(-0.03147425130009651)),(to_sfixed_a(-0.24052582681179047)),(to_sfixed_a(-0.11655811965465546)),(to_sfixed_a(0.13304415345191956)),(to_sfixed_a(0.06369564682245255)),(to_sfixed_a(0.0440450944006443)),(to_sfixed_a(-0.0850302129983902)),(to_sfixed_a(-0.0932779461145401)),(to_sfixed_a(0.10214343667030334)),(to_sfixed_a(0.0046907635405659676)),(to_sfixed_a(9.659615170676261e-05)),(to_sfixed_a(-0.00027983865584246814)),(to_sfixed_a(0.0005055329529568553)),(to_sfixed_a(0.00010738449054770172)),(to_sfixed_a(-5.274544491840061e-06)),(to_sfixed_a(-0.00018365372670814395)),(to_sfixed_a(0.003117811167612672)),(to_sfixed_a(0.003427959978580475)),(to_sfixed_a(-0.06440409272909164)),(to_sfixed_a(0.01770549640059471)),(to_sfixed_a(0.011785120703279972)),(to_sfixed_a(0.07617304474115372)),(to_sfixed_a(0.11261752247810364)),(to_sfixed_a(0.15177087485790253)),(to_sfixed_a(0.13697932660579681)),(to_sfixed_a(0.07218125462532043)),(to_sfixed_a(-0.21903695166110992)),(to_sfixed_a(0.12084904313087463)),(to_sfixed_a(0.02138531766831875)),(to_sfixed_a(-0.2582319974899292)),(to_sfixed_a(0.2135435938835144)),(to_sfixed_a(-0.05952683091163635)),(to_sfixed_a(0.000921096361707896)),(to_sfixed_a(0.06205308064818382)),(to_sfixed_a(-0.026343975216150284)),(to_sfixed_a(-0.06817691028118134)),(to_sfixed_a(-0.4240042269229889)),(to_sfixed_a(-6.66356718284078e-05)),(to_sfixed_a(-0.0001269378699362278)),(to_sfixed_a(-0.0002196403656853363)),(to_sfixed_a(-1.6693897123332135e-05)),(to_sfixed_a(0.00019474417786113918)),(to_sfixed_a(-4.115708179597277e-06)),(to_sfixed_a(-6.844331801403314e-05)),(to_sfixed_a(2.3725344362901524e-05)),(to_sfixed_a(0.010197421535849571)),(to_sfixed_a(-0.15856893360614777)),(to_sfixed_a(-0.09960183501243591)),(to_sfixed_a(0.01687815599143505)),(to_sfixed_a(0.026555094867944717)),(to_sfixed_a(0.12449384480714798)),(to_sfixed_a(0.06100361794233322)),(to_sfixed_a(0.11050879210233688)),(to_sfixed_a(0.23673802614212036)),(to_sfixed_a(0.028025150299072266)),(to_sfixed_a(0.21367791295051575)),(to_sfixed_a(0.15638750791549683)),(to_sfixed_a(0.033806633204221725)),(to_sfixed_a(0.05254141986370087)),(to_sfixed_a(0.15219846367835999)),(to_sfixed_a(0.05572221800684929)),(to_sfixed_a(-0.23525190353393555)),(to_sfixed_a(-0.17577923834323883)),(to_sfixed_a(-0.17313139140605927)),(to_sfixed_a(-0.06203993782401085)),(to_sfixed_a(0.031209591776132584)),(to_sfixed_a(3.018835195689462e-05)),(to_sfixed_a(-7.2199932219518814e-06)),(to_sfixed_a(-0.0002073112118523568)),(to_sfixed_a(4.74029548058752e-05)),(to_sfixed_a(-0.00014318038302008063)),(to_sfixed_a(-8.429805893683806e-05)),(to_sfixed_a(6.731789471814409e-05)),(to_sfixed_a(-0.012949884869158268)),(to_sfixed_a(0.0007884571678005159)),(to_sfixed_a(0.0783449038863182)),(to_sfixed_a(0.027084510773420334)),(to_sfixed_a(-0.012770374305546284)),(to_sfixed_a(0.02146962843835354)),(to_sfixed_a(-0.09978703409433365)),(to_sfixed_a(0.17189234495162964)),(to_sfixed_a(0.041610367596149445)),(to_sfixed_a(-0.18782781064510345)),(to_sfixed_a(-0.05052778497338295)),(to_sfixed_a(0.1966944932937622)),(to_sfixed_a(0.06046630069613457)),(to_sfixed_a(0.20339833199977875)),(to_sfixed_a(-0.04428783804178238)),(to_sfixed_a(0.055971890687942505)),(to_sfixed_a(-0.35041481256484985)),(to_sfixed_a(-0.16120725870132446)),(to_sfixed_a(-0.36228564381599426)),(to_sfixed_a(-0.00026872099260799587)),(to_sfixed_a(-0.09412194788455963)),(to_sfixed_a(7.038180046947673e-05)),(to_sfixed_a(-1.4144272427074611e-05)),(to_sfixed_a(0.00017449381994083524)),(to_sfixed_a(0.0001708869094727561)),(to_sfixed_a(-0.00019626939320005476)),(to_sfixed_a(0.00014866082346998155)),(to_sfixed_a(0.00011671978427330032)),(to_sfixed_a(0.00022377407003659755)),(to_sfixed_a(0.09716561436653137)),(to_sfixed_a(0.06473558396100998)),(to_sfixed_a(-0.016777843236923218)),(to_sfixed_a(0.024899397045373917)),(to_sfixed_a(-0.08838710188865662)),(to_sfixed_a(-0.12253454327583313)),(to_sfixed_a(0.05638495460152626)),(to_sfixed_a(0.08841218054294586)),(to_sfixed_a(0.09169120341539383)),(to_sfixed_a(0.07597211003303528)),(to_sfixed_a(0.201967254281044)),(to_sfixed_a(0.0237031988799572)),(to_sfixed_a(0.06461972743272781)),(to_sfixed_a(-0.006414005998522043)),(to_sfixed_a(-0.24441644549369812)),(to_sfixed_a(-0.13152247667312622)),(to_sfixed_a(0.04152602329850197)),(to_sfixed_a(-0.028962187469005585)),(to_sfixed_a(0.011323791928589344)),(to_sfixed_a(-4.685799285653047e-05)),(to_sfixed_a(-6.479943112935871e-05)),(to_sfixed_a(6.31892544333823e-05)),(to_sfixed_a(-3.180851126671769e-05)),(to_sfixed_a(-0.0001723224122542888)),(to_sfixed_a(9.252641757484525e-05)),(to_sfixed_a(0.00021817712695337832)),(to_sfixed_a(-8.917511149775237e-05)),(to_sfixed_a(0.00047250385978259146)),(to_sfixed_a(-0.007329369895160198)),(to_sfixed_a(-0.05809818580746651)),(to_sfixed_a(0.1489141434431076)),(to_sfixed_a(0.16220985352993011)),(to_sfixed_a(0.06405331194400787)),(to_sfixed_a(0.05256761983036995)),(to_sfixed_a(-0.1936284899711609)),(to_sfixed_a(0.09384171664714813)),(to_sfixed_a(0.18362468481063843)),(to_sfixed_a(-0.029424449428915977)),(to_sfixed_a(-0.10650385171175003)),(to_sfixed_a(0.276945024728775)),(to_sfixed_a(0.013648026622831821)),(to_sfixed_a(0.06157433241605759)),(to_sfixed_a(-0.29027488827705383)),(to_sfixed_a(-0.024001045152544975)),(to_sfixed_a(-0.2666182816028595)),(to_sfixed_a(0.018700553104281425)),(to_sfixed_a(-0.20826265215873718)),(to_sfixed_a(-9.070656960830092e-05)),(to_sfixed_a(7.334262045333162e-05)),(to_sfixed_a(0.00010233899229206145)),(to_sfixed_a(-0.0001015513771562837)),(to_sfixed_a(0.00028487257077358663)),(to_sfixed_a(5.9883521316805854e-05)),(to_sfixed_a(-8.902016998035833e-05)),(to_sfixed_a(3.049286169698462e-05)),(to_sfixed_a(0.0142075689509511)),(to_sfixed_a(-0.029760489240288734)),(to_sfixed_a(0.058435726910829544)),(to_sfixed_a(0.07710802555084229)),(to_sfixed_a(0.005365228280425072)),(to_sfixed_a(0.09732210636138916)),(to_sfixed_a(-0.03226049616932869)),(to_sfixed_a(-0.008824504911899567)),(to_sfixed_a(0.4153062701225281)),(to_sfixed_a(0.070221446454525)),(to_sfixed_a(-0.010192930698394775)),(to_sfixed_a(0.09546301513910294)),(to_sfixed_a(-0.00019697847892530262)),(to_sfixed_a(0.15919595956802368)),(to_sfixed_a(0.02213735319674015)),(to_sfixed_a(-0.15011826157569885)),(to_sfixed_a(-0.00037156889447942376)),(to_sfixed_a(-0.22295276820659637)),(to_sfixed_a(-0.10302404314279556)),(to_sfixed_a(0.005628622602671385)),(to_sfixed_a(9.754996426636353e-05)),(to_sfixed_a(0.00011837424244731665)),(to_sfixed_a(-1.9638311641756445e-05)),(to_sfixed_a(-4.1633204091340303e-05)),(to_sfixed_a(-0.00011789338168455288)),(to_sfixed_a(-9.769819007487968e-05)),(to_sfixed_a(-0.0003274580813013017)),(to_sfixed_a(-0.00017465530254412442)),(to_sfixed_a(-0.00026550792972557247)),(to_sfixed_a(-0.010606725700199604)),(to_sfixed_a(0.03564199060201645)),(to_sfixed_a(0.03913162648677826)),(to_sfixed_a(0.211323544383049)),(to_sfixed_a(0.3464414179325104)),(to_sfixed_a(0.037257276475429535)),(to_sfixed_a(-0.04844389855861664)),(to_sfixed_a(0.2565656900405884)),(to_sfixed_a(-0.17305326461791992)),(to_sfixed_a(0.09582558274269104)),(to_sfixed_a(0.12350308895111084)),(to_sfixed_a(-0.11620400846004486)),(to_sfixed_a(0.04571262001991272)),(to_sfixed_a(0.0044852024875581264)),(to_sfixed_a(-0.05714758113026619)),(to_sfixed_a(-0.16532140970230103)),(to_sfixed_a(0.00010208981257164851)),(to_sfixed_a(0.002128991298377514)),(to_sfixed_a(0.0028298450633883476)),(to_sfixed_a(-0.0002179789007641375)),(to_sfixed_a(-2.185610901506152e-05)),(to_sfixed_a(0.0001884523080661893)),(to_sfixed_a(-0.00011825859837699682)),(to_sfixed_a(-0.00011725235526682809)),(to_sfixed_a(-6.012455196469091e-05)),(to_sfixed_a(4.110572626814246e-05)),(to_sfixed_a(-2.484396827640012e-05)),(to_sfixed_a(-0.00014923917478881776)),(to_sfixed_a(-0.001347377896308899)),(to_sfixed_a(-0.0011958335526287556)),(to_sfixed_a(-9.257900092052296e-05)),(to_sfixed_a(0.0002838409272953868)),(to_sfixed_a(-0.00017680363089311868)),(to_sfixed_a(-0.06601423770189285)),(to_sfixed_a(-0.004794837906956673)),(to_sfixed_a(-0.001917428569868207)),(to_sfixed_a(-0.048574019223451614)),(to_sfixed_a(0.0681849792599678)),(to_sfixed_a(-0.0052832867950201035)),(to_sfixed_a(-0.025844009593129158)),(to_sfixed_a(-0.048916690051555634)),(to_sfixed_a(-0.06280507147312164)),(to_sfixed_a(-6.147625390440226e-05)),(to_sfixed_a(-0.0018353356281295419)),(to_sfixed_a(-0.0001264992170035839)),(to_sfixed_a(-0.00014325704250950366)),(to_sfixed_a(-9.586942906025797e-05)),(to_sfixed_a(-0.00013982960081193596)),(to_sfixed_a(3.878126517520286e-05)),(to_sfixed_a(-1.1489966709632427e-05)),(to_sfixed_a(-4.204135620966554e-06)),(to_sfixed_a(-7.790106610627845e-05)),(to_sfixed_a(0.0003822079743258655)),(to_sfixed_a(-3.0453871659119613e-05)),(to_sfixed_a(-2.4977958673844114e-05)),(to_sfixed_a(0.0002562172885518521)),(to_sfixed_a(8.106807217700407e-05)),(to_sfixed_a(-6.414294330170378e-05)),(to_sfixed_a(0.00018922073650173843)),(to_sfixed_a(-0.0003180172643624246)),(to_sfixed_a(0.00010965823457809165)),(to_sfixed_a(0.0001120578235713765)),(to_sfixed_a(0.00012945910566486418)),(to_sfixed_a(3.506078428472392e-05)),(to_sfixed_a(3.7032888940302655e-05)),(to_sfixed_a(-2.0042905816808343e-05)),(to_sfixed_a(-3.619962080847472e-05)),(to_sfixed_a(5.0164471758762375e-05)),(to_sfixed_a(-5.898492599953897e-05)),(to_sfixed_a(-0.00013905971718486398)),(to_sfixed_a(0.00013693551591131836)),(to_sfixed_a(3.1684299756307155e-05)),(to_sfixed_a(-8.017231448320672e-05)),(to_sfixed_a(-7.425401418004185e-05)),(to_sfixed_a(2.28258031711448e-05)),(to_sfixed_a(-0.00018703757086768746)),(to_sfixed_a(-0.00019289780175313354)),(to_sfixed_a(0.00017929892055690289)),(to_sfixed_a(-0.00019969200366176665)));

    constant weight_n0_19 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-0.0002741410571616143)),(to_sfixed_a(9.921361197484657e-05)),(to_sfixed_a(-8.024451381061226e-05)),(to_sfixed_a(-0.00027376547222957015)),(to_sfixed_a(-8.157495176419616e-05)),(to_sfixed_a(0.0003223234380129725)),(to_sfixed_a(0.00012172663991805166)),(to_sfixed_a(-0.00017279107123613358)),(to_sfixed_a(5.385694021242671e-05)),(to_sfixed_a(9.471796511206776e-05)),(to_sfixed_a(-0.00012652957229875028)),(to_sfixed_a(0.0002275631995871663)),(to_sfixed_a(0.00030562514439225197)),(to_sfixed_a(0.00010594905324978754)),(to_sfixed_a(0.0002550584904383868)),(to_sfixed_a(0.00026153726503252983)),(to_sfixed_a(0.0003466022026259452)),(to_sfixed_a(0.00024840724654495716)),(to_sfixed_a(0.00013865575601812452)),(to_sfixed_a(0.00013048724213149399)),(to_sfixed_a(6.625644164159894e-05)),(to_sfixed_a(2.3665417757001705e-05)),(to_sfixed_a(-0.00018739610095508397)),(to_sfixed_a(-4.8283593059750274e-05)),(to_sfixed_a(-9.611475979909301e-05)),(to_sfixed_a(0.00011992752843070775)),(to_sfixed_a(-0.00024178458261303604)),(to_sfixed_a(-0.0002057632664218545)),(to_sfixed_a(-0.00031860239687375724)),(to_sfixed_a(-0.0001816209842218086)),(to_sfixed_a(8.326372335432097e-05)),(to_sfixed_a(0.00011267426452832296)),(to_sfixed_a(0.0002612140087876469)),(to_sfixed_a(8.712882117833942e-05)),(to_sfixed_a(0.0001264891616301611)),(to_sfixed_a(-0.0003948248049709946)),(to_sfixed_a(0.00021363588166423142)),(to_sfixed_a(-0.00013787300849799067)),(to_sfixed_a(0.0002243844064651057)),(to_sfixed_a(-3.1652540201321244e-05)),(to_sfixed_a(-7.3150590651493985e-06)),(to_sfixed_a(1.7539085092721507e-05)),(to_sfixed_a(-0.00012905399489682168)),(to_sfixed_a(-0.00015484585310332477)),(to_sfixed_a(-0.0001191071787616238)),(to_sfixed_a(7.879523036535829e-05)),(to_sfixed_a(-6.681161175947636e-05)),(to_sfixed_a(4.514320971793495e-05)),(to_sfixed_a(0.00018949990044347942)),(to_sfixed_a(-0.00024350045714527369)),(to_sfixed_a(-0.0001751749950926751)),(to_sfixed_a(0.00015878738486208022)),(to_sfixed_a(0.00021679165365640074)),(to_sfixed_a(-3.82642938347999e-05)),(to_sfixed_a(5.235098069533706e-05)),(to_sfixed_a(-6.693279283354059e-05)),(to_sfixed_a(7.680289854761213e-05)),(to_sfixed_a(0.0003837553085759282)),(to_sfixed_a(0.0001369624224025756)),(to_sfixed_a(-5.785754547105171e-05)),(to_sfixed_a(1.2474733921408188e-05)),(to_sfixed_a(4.3654032197082415e-05)),(to_sfixed_a(9.876859257929027e-05)),(to_sfixed_a(-0.0002431790198897943)),(to_sfixed_a(-0.0002581081062089652)),(to_sfixed_a(-2.875838617910631e-06)),(to_sfixed_a(5.033297566114925e-05)),(to_sfixed_a(4.334115510573611e-05)),(to_sfixed_a(7.876747258706018e-05)),(to_sfixed_a(0.00856423657387495)),(to_sfixed_a(-0.00014635520346928388)),(to_sfixed_a(-2.783360287139658e-05)),(to_sfixed_a(-0.0001342909235972911)),(to_sfixed_a(-0.00014637084677815437)),(to_sfixed_a(3.444387766649015e-05)),(to_sfixed_a(8.087839523795992e-05)),(to_sfixed_a(0.00024449144257232547)),(to_sfixed_a(-0.00010349285730626434)),(to_sfixed_a(0.00013372182729654014)),(to_sfixed_a(9.622643847251311e-05)),(to_sfixed_a(-0.00021353985357563943)),(to_sfixed_a(-0.00011764496593968943)),(to_sfixed_a(1.3736846085521393e-05)),(to_sfixed_a(1.9441729818936437e-05)),(to_sfixed_a(0.00016438806778751314)),(to_sfixed_a(7.09295563865453e-05)),(to_sfixed_a(1.4194391951605212e-05)),(to_sfixed_a(-0.0002639994490891695)),(to_sfixed_a(-0.00011565400927793235)),(to_sfixed_a(-0.0001844197540776804)),(to_sfixed_a(0.000166190744494088)),(to_sfixed_a(0.0001429022813681513)),(to_sfixed_a(-0.0798952654004097)),(to_sfixed_a(2.4153136109816842e-05)),(to_sfixed_a(-0.09059152007102966)),(to_sfixed_a(-0.02844223938882351)),(to_sfixed_a(-0.12589497864246368)),(to_sfixed_a(-0.01808454841375351)),(to_sfixed_a(-0.16733941435813904)),(to_sfixed_a(0.07433127611875534)),(to_sfixed_a(-0.0030513606034219265)),(to_sfixed_a(-0.015449819155037403)),(to_sfixed_a(0.07115156948566437)),(to_sfixed_a(-0.0007956466288305819)),(to_sfixed_a(-0.009815641678869724)),(to_sfixed_a(-0.020070476457476616)),(to_sfixed_a(0.0001582843833602965)),(to_sfixed_a(-0.00016150038572959602)),(to_sfixed_a(-7.586408901261166e-05)),(to_sfixed_a(0.00032053980976343155)),(to_sfixed_a(0.0001036305257002823)),(to_sfixed_a(0.00024001175188459456)),(to_sfixed_a(2.9632787118316628e-05)),(to_sfixed_a(-3.6822326364926994e-05)),(to_sfixed_a(0.00032513769110664725)),(to_sfixed_a(-0.00011432357860030606)),(to_sfixed_a(-0.00018029533384833485)),(to_sfixed_a(2.4667147954460233e-05)),(to_sfixed_a(0.000646400498226285)),(to_sfixed_a(-0.06729727983474731)),(to_sfixed_a(0.05596319958567619)),(to_sfixed_a(-0.11405591666698456)),(to_sfixed_a(0.1370743364095688)),(to_sfixed_a(-0.035231009125709534)),(to_sfixed_a(0.10994971543550491)),(to_sfixed_a(0.19182275235652924)),(to_sfixed_a(-0.14172427356243134)),(to_sfixed_a(-0.028496701270341873)),(to_sfixed_a(-0.1426289677619934)),(to_sfixed_a(0.053442154079675674)),(to_sfixed_a(0.07833003997802734)),(to_sfixed_a(-0.050647880882024765)),(to_sfixed_a(-0.005209102761000395)),(to_sfixed_a(-0.03344259411096573)),(to_sfixed_a(-0.03610842302441597)),(to_sfixed_a(-1.0928692972811405e-05)),(to_sfixed_a(0.0013990398729220033)),(to_sfixed_a(-0.00019147062266711146)),(to_sfixed_a(-0.00033853118657134473)),(to_sfixed_a(0.00015641507343389094)),(to_sfixed_a(4.4433931179810315e-05)),(to_sfixed_a(-3.35960321535822e-05)),(to_sfixed_a(-0.00030016389791853726)),(to_sfixed_a(-0.00033244400401599705)),(to_sfixed_a(-4.4708627683576196e-05)),(to_sfixed_a(-0.11753326654434204)),(to_sfixed_a(-0.015012640506029129)),(to_sfixed_a(-0.10097730904817581)),(to_sfixed_a(0.1054028794169426)),(to_sfixed_a(0.07490230351686478)),(to_sfixed_a(-0.09068501740694046)),(to_sfixed_a(-0.05664592236280441)),(to_sfixed_a(-0.06713833659887314)),(to_sfixed_a(-0.3095187842845917)),(to_sfixed_a(-0.13209646940231323)),(to_sfixed_a(-0.2442210167646408)),(to_sfixed_a(-0.2071305215358734)),(to_sfixed_a(-0.05591725930571556)),(to_sfixed_a(-0.017676973715424538)),(to_sfixed_a(0.10831610858440399)),(to_sfixed_a(-0.026481306180357933)),(to_sfixed_a(-0.11136383563280106)),(to_sfixed_a(0.004491083323955536)),(to_sfixed_a(-0.01707392744719982)),(to_sfixed_a(0.002947047585621476)),(to_sfixed_a(-6.0666323406621814e-05)),(to_sfixed_a(-7.02379911672324e-05)),(to_sfixed_a(-1.9585202608141117e-05)),(to_sfixed_a(-0.00013760599540546536)),(to_sfixed_a(-0.00020225900516379625)),(to_sfixed_a(3.5533623304218054e-05)),(to_sfixed_a(-8.324820373672992e-05)),(to_sfixed_a(-0.000230179080972448)),(to_sfixed_a(-0.10909178853034973)),(to_sfixed_a(-0.11068243533372879)),(to_sfixed_a(-0.09392456710338593)),(to_sfixed_a(0.08444876223802567)),(to_sfixed_a(0.2692430019378662)),(to_sfixed_a(0.1726936399936676)),(to_sfixed_a(0.167199969291687)),(to_sfixed_a(0.1403864473104477)),(to_sfixed_a(0.06898113340139389)),(to_sfixed_a(0.21117670834064484)),(to_sfixed_a(0.3440190255641937)),(to_sfixed_a(0.4293091893196106)),(to_sfixed_a(0.39761465787887573)),(to_sfixed_a(0.20783261954784393)),(to_sfixed_a(0.15587136149406433)),(to_sfixed_a(0.11439163237810135)),(to_sfixed_a(-0.058120857924222946)),(to_sfixed_a(-0.15027695894241333)),(to_sfixed_a(-0.13207462430000305)),(to_sfixed_a(-0.0015952049288898706)),(to_sfixed_a(-0.0029945839196443558)),(to_sfixed_a(-0.003580991178750992)),(to_sfixed_a(-0.00017427877173759043)),(to_sfixed_a(-0.0002649606904014945)),(to_sfixed_a(-0.0003883270837832242)),(to_sfixed_a(-7.925659156171605e-05)),(to_sfixed_a(-3.2753781852079555e-05)),(to_sfixed_a(0.00028375835972838104)),(to_sfixed_a(-0.05522590130567551)),(to_sfixed_a(-0.09714993089437485)),(to_sfixed_a(0.12085272371768951)),(to_sfixed_a(0.22330418229103088)),(to_sfixed_a(-0.19005702435970306)),(to_sfixed_a(-0.007019100710749626)),(to_sfixed_a(0.028531895950436592)),(to_sfixed_a(-0.14699801802635193)),(to_sfixed_a(0.15283524990081787)),(to_sfixed_a(0.1364307850599289)),(to_sfixed_a(0.697439968585968)),(to_sfixed_a(0.23037776350975037)),(to_sfixed_a(0.2280334234237671)),(to_sfixed_a(0.2636263072490692)),(to_sfixed_a(0.2711796164512634)),(to_sfixed_a(-0.039485055953264236)),(to_sfixed_a(0.188186377286911)),(to_sfixed_a(-0.006768304854631424)),(to_sfixed_a(0.005829231813549995)),(to_sfixed_a(0.002505436073988676)),(to_sfixed_a(-0.0017856932245194912)),(to_sfixed_a(-0.00014592251682188362)),(to_sfixed_a(-2.8029908207827248e-06)),(to_sfixed_a(1.0639422725944314e-05)),(to_sfixed_a(3.3732474548742175e-05)),(to_sfixed_a(0.00029878117493353784)),(to_sfixed_a(4.893524237559177e-05)),(to_sfixed_a(0.04136353358626366)),(to_sfixed_a(-0.0037649571895599365)),(to_sfixed_a(0.04307657107710838)),(to_sfixed_a(0.00018563777848612517)),(to_sfixed_a(0.4649650752544403)),(to_sfixed_a(0.10238200426101685)),(to_sfixed_a(0.16551218926906586)),(to_sfixed_a(0.12373966723680496)),(to_sfixed_a(-0.09805717319250107)),(to_sfixed_a(0.1506848782300949)),(to_sfixed_a(0.28661900758743286)),(to_sfixed_a(0.3430649936199188)),(to_sfixed_a(0.08823369443416595)),(to_sfixed_a(-0.08464370667934418)),(to_sfixed_a(0.08466022461652756)),(to_sfixed_a(-0.008527787402272224)),(to_sfixed_a(-0.08037252724170685)),(to_sfixed_a(-0.11159085482358932)),(to_sfixed_a(0.0903736874461174)),(to_sfixed_a(-0.09554062783718109)),(to_sfixed_a(-0.10754655301570892)),(to_sfixed_a(-0.002154735615476966)),(to_sfixed_a(-0.0003311455948278308)),(to_sfixed_a(0.00015054087270982563)),(to_sfixed_a(-6.502594624180347e-05)),(to_sfixed_a(0.0003992176498286426)),(to_sfixed_a(-0.00012277578935027122)),(to_sfixed_a(0.00012654505553655326)),(to_sfixed_a(0.0010639243992045522)),(to_sfixed_a(0.11723367124795914)),(to_sfixed_a(-0.03486420959234238)),(to_sfixed_a(0.12294622510671616)),(to_sfixed_a(0.11116334795951843)),(to_sfixed_a(0.0980958640575409)),(to_sfixed_a(0.366086483001709)),(to_sfixed_a(-0.06173108145594597)),(to_sfixed_a(-0.3127533793449402)),(to_sfixed_a(-0.189723938703537)),(to_sfixed_a(0.10572188347578049)),(to_sfixed_a(0.24566136300563812)),(to_sfixed_a(0.0017440502997487783)),(to_sfixed_a(-0.15944337844848633)),(to_sfixed_a(-0.09828659147024155)),(to_sfixed_a(0.3235398530960083)),(to_sfixed_a(0.2849023640155792)),(to_sfixed_a(0.18227297067642212)),(to_sfixed_a(0.03807384520769119)),(to_sfixed_a(0.019581839442253113)),(to_sfixed_a(0.07476798444986343)),(to_sfixed_a(3.871640365105122e-05)),(to_sfixed_a(-0.0001905026292661205)),(to_sfixed_a(3.7549874832620844e-05)),(to_sfixed_a(1.529505243524909e-05)),(to_sfixed_a(-6.600526830879971e-05)),(to_sfixed_a(0.00018008863844443113)),(to_sfixed_a(-0.00031392797245644033)),(to_sfixed_a(0.005895114038139582)),(to_sfixed_a(-0.040427133440971375)),(to_sfixed_a(0.08000235259532928)),(to_sfixed_a(0.1708010733127594)),(to_sfixed_a(0.29088208079338074)),(to_sfixed_a(0.2656892240047455)),(to_sfixed_a(0.18406161665916443)),(to_sfixed_a(-0.45944035053253174)),(to_sfixed_a(-0.2695850431919098)),(to_sfixed_a(-0.13806357979774475)),(to_sfixed_a(0.18247491121292114)),(to_sfixed_a(-0.07405711710453033)),(to_sfixed_a(-0.11223152279853821)),(to_sfixed_a(0.054536204785108566)),(to_sfixed_a(0.06304143369197845)),(to_sfixed_a(0.09483183175325394)),(to_sfixed_a(0.14666688442230225)),(to_sfixed_a(0.17856402695178986)),(to_sfixed_a(0.02895107865333557)),(to_sfixed_a(0.13000796735286713)),(to_sfixed_a(-0.0948496162891388)),(to_sfixed_a(-0.010815724730491638)),(to_sfixed_a(-9.62404374149628e-05)),(to_sfixed_a(-4.663498475565575e-05)),(to_sfixed_a(0.00021875246602576226)),(to_sfixed_a(0.00011587038898142055)),(to_sfixed_a(9.249098366126418e-05)),(to_sfixed_a(-0.048459868878126144)),(to_sfixed_a(0.05771166831254959)),(to_sfixed_a(0.25089508295059204)),(to_sfixed_a(0.11158878356218338)),(to_sfixed_a(0.28827694058418274)),(to_sfixed_a(0.12336590886116028)),(to_sfixed_a(0.2234523892402649)),(to_sfixed_a(0.03611702471971512)),(to_sfixed_a(-0.006173479370772839)),(to_sfixed_a(-0.017484426498413086)),(to_sfixed_a(0.12541070580482483)),(to_sfixed_a(0.36104580760002136)),(to_sfixed_a(-0.050771668553352356)),(to_sfixed_a(-0.0018997330917045474)),(to_sfixed_a(0.026344195008277893)),(to_sfixed_a(0.21108661592006683)),(to_sfixed_a(0.2890656292438507)),(to_sfixed_a(0.3821299970149994)),(to_sfixed_a(0.12240998446941376)),(to_sfixed_a(0.05575832352042198)),(to_sfixed_a(-0.0054121557623147964)),(to_sfixed_a(-0.17973151803016663)),(to_sfixed_a(4.1320989112136886e-05)),(to_sfixed_a(-0.00011609750072238967)),(to_sfixed_a(0.00017232762183994055)),(to_sfixed_a(-2.7150381356477737e-05)),(to_sfixed_a(5.434222111944109e-05)),(to_sfixed_a(-1.6982288798317313e-05)),(to_sfixed_a(0.00021468993509188294)),(to_sfixed_a(0.08279018104076385)),(to_sfixed_a(0.05493045598268509)),(to_sfixed_a(0.11330568790435791)),(to_sfixed_a(-0.030336756259202957)),(to_sfixed_a(-0.13942943513393402)),(to_sfixed_a(0.08515981584787369)),(to_sfixed_a(-0.2786863148212433)),(to_sfixed_a(0.07080908864736557)),(to_sfixed_a(0.3809564411640167)),(to_sfixed_a(0.21568866074085236)),(to_sfixed_a(-0.2632811963558197)),(to_sfixed_a(-0.06078510358929634)),(to_sfixed_a(0.06422178447246552)),(to_sfixed_a(0.013422446325421333)),(to_sfixed_a(-0.004573035053908825)),(to_sfixed_a(0.3427664339542389)),(to_sfixed_a(0.36914268136024475)),(to_sfixed_a(0.13459517061710358)),(to_sfixed_a(0.2913501560688019)),(to_sfixed_a(-0.05560578778386116)),(to_sfixed_a(0.04476276785135269)),(to_sfixed_a(-0.00010153243783861399)),(to_sfixed_a(-1.091195190383587e-05)),(to_sfixed_a(-0.00020184363529551774)),(to_sfixed_a(0.0002902151027228683)),(to_sfixed_a(-0.00016172790492419153)),(to_sfixed_a(0.00014725890650879592)),(to_sfixed_a(0.0002804800751619041)),(to_sfixed_a(-0.0729350820183754)),(to_sfixed_a(-0.0724204033613205)),(to_sfixed_a(-0.07815007865428925)),(to_sfixed_a(0.01715203933417797)),(to_sfixed_a(0.03286800533533096)),(to_sfixed_a(0.19992254674434662)),(to_sfixed_a(0.033821649849414825)),(to_sfixed_a(0.3594505488872528)),(to_sfixed_a(0.14804606139659882)),(to_sfixed_a(-0.17116037011146545)),(to_sfixed_a(0.19534996151924133)),(to_sfixed_a(0.0760875940322876)),(to_sfixed_a(0.08033794909715652)),(to_sfixed_a(0.09701826423406601)),(to_sfixed_a(0.07211912423372269)),(to_sfixed_a(0.14808982610702515)),(to_sfixed_a(0.01276666671037674)),(to_sfixed_a(0.08624260127544403)),(to_sfixed_a(-0.11975906044244766)),(to_sfixed_a(-0.13597150146961212)),(to_sfixed_a(-0.10382897406816483)),(to_sfixed_a(-0.0012605779338628054)),(to_sfixed_a(-0.0023696287535130978)),(to_sfixed_a(0.00011277373414486647)),(to_sfixed_a(6.0771599237341434e-05)),(to_sfixed_a(-0.00021669759007636458)),(to_sfixed_a(-0.00021176804148126394)),(to_sfixed_a(3.146850212942809e-05)),(to_sfixed_a(-0.0010026897070929408)),(to_sfixed_a(0.03438941389322281)),(to_sfixed_a(-0.03297470510005951)),(to_sfixed_a(0.007498402614146471)),(to_sfixed_a(0.10593336075544357)),(to_sfixed_a(0.09490528702735901)),(to_sfixed_a(0.22970308363437653)),(to_sfixed_a(-0.0020324818324297667)),(to_sfixed_a(-0.11407975852489471)),(to_sfixed_a(0.01302525494247675)),(to_sfixed_a(0.2061779499053955)),(to_sfixed_a(0.14682349562644958)),(to_sfixed_a(0.02555428259074688)),(to_sfixed_a(0.16398002207279205)),(to_sfixed_a(0.22184592485427856)),(to_sfixed_a(0.09479987621307373)),(to_sfixed_a(-0.0664738118648529)),(to_sfixed_a(-0.2702715992927551)),(to_sfixed_a(-0.12855790555477142)),(to_sfixed_a(-0.08662377297878265)),(to_sfixed_a(-0.09222530573606491)),(to_sfixed_a(-3.0419738322962075e-05)),(to_sfixed_a(-1.933306884893682e-05)),(to_sfixed_a(-6.413312803488225e-05)),(to_sfixed_a(1.1276399163762107e-05)),(to_sfixed_a(1.2542218428279739e-05)),(to_sfixed_a(7.701135473325849e-05)),(to_sfixed_a(0.00015999445167835802)),(to_sfixed_a(-0.0012792133493348956)),(to_sfixed_a(0.023318324238061905)),(to_sfixed_a(0.06986644864082336)),(to_sfixed_a(-0.09864131361246109)),(to_sfixed_a(0.08078283816576004)),(to_sfixed_a(0.14169473946094513)),(to_sfixed_a(0.08673965185880661)),(to_sfixed_a(-0.0335497222840786)),(to_sfixed_a(-0.12101513892412186)),(to_sfixed_a(0.23099565505981445)),(to_sfixed_a(0.32818928360939026)),(to_sfixed_a(0.1561681628227234)),(to_sfixed_a(0.08592555671930313)),(to_sfixed_a(0.064724862575531)),(to_sfixed_a(-0.08053167164325714)),(to_sfixed_a(-0.247431218624115)),(to_sfixed_a(-0.08261183649301529)),(to_sfixed_a(-0.022062484174966812)),(to_sfixed_a(0.16660673916339874)),(to_sfixed_a(-0.10871514678001404)),(to_sfixed_a(0.006422244478017092)),(to_sfixed_a(-0.00038651813520118594)),(to_sfixed_a(-0.00010111371375387534)),(to_sfixed_a(5.7582186855142936e-05)),(to_sfixed_a(-8.464219718007371e-05)),(to_sfixed_a(-0.0001198009485960938)),(to_sfixed_a(0.00016758155834395438)),(to_sfixed_a(0.0029087322764098644)),(to_sfixed_a(0.18342050909996033)),(to_sfixed_a(0.07307769358158112)),(to_sfixed_a(0.01397128589451313)),(to_sfixed_a(0.18059031665325165)),(to_sfixed_a(0.260612815618515)),(to_sfixed_a(-0.06322582811117172)),(to_sfixed_a(-0.19437232613563538)),(to_sfixed_a(-0.21115441620349884)),(to_sfixed_a(-0.46504124999046326)),(to_sfixed_a(0.03378276526927948)),(to_sfixed_a(0.05512036010622978)),(to_sfixed_a(-0.018831992521882057)),(to_sfixed_a(0.04671928286552429)),(to_sfixed_a(0.11993923038244247)),(to_sfixed_a(-0.23840755224227905)),(to_sfixed_a(-0.3216148912906647)),(to_sfixed_a(-0.3302062153816223)),(to_sfixed_a(-0.2810553014278412)),(to_sfixed_a(-0.15789097547531128)),(to_sfixed_a(0.07946617901325226)),(to_sfixed_a(-0.09440146386623383)),(to_sfixed_a(-0.009812005795538425)),(to_sfixed_a(-0.0002465667494107038)),(to_sfixed_a(-9.480433800490573e-05)),(to_sfixed_a(-9.396744280820712e-05)),(to_sfixed_a(-0.00012462363520171493)),(to_sfixed_a(0.0025916281156241894)),(to_sfixed_a(0.0033592619001865387)),(to_sfixed_a(-0.14157550036907196)),(to_sfixed_a(0.11887854337692261)),(to_sfixed_a(-0.011626964434981346)),(to_sfixed_a(-0.08890563994646072)),(to_sfixed_a(0.27714410424232483)),(to_sfixed_a(0.04280896484851837)),(to_sfixed_a(-0.09654790163040161)),(to_sfixed_a(-0.45721539855003357)),(to_sfixed_a(-0.24041438102722168)),(to_sfixed_a(-0.04851772263646126)),(to_sfixed_a(-0.006899170111864805)),(to_sfixed_a(0.3796718418598175)),(to_sfixed_a(0.12797360122203827)),(to_sfixed_a(-0.10406394302845001)),(to_sfixed_a(-0.20899342000484467)),(to_sfixed_a(-0.4903997480869293)),(to_sfixed_a(-0.23209330439567566)),(to_sfixed_a(0.01285207737237215)),(to_sfixed_a(-0.14504685997962952)),(to_sfixed_a(-0.0152954813092947)),(to_sfixed_a(-0.0002150659856852144)),(to_sfixed_a(1.6001782569219358e-05)),(to_sfixed_a(-0.00012889740173704922)),(to_sfixed_a(9.879013668978587e-05)),(to_sfixed_a(1.2434458767529577e-05)),(to_sfixed_a(0.00010976789781125262)),(to_sfixed_a(-9.757409861776978e-05)),(to_sfixed_a(0.01038326695561409)),(to_sfixed_a(0.019483551383018494)),(to_sfixed_a(0.16680221259593964)),(to_sfixed_a(0.09907418489456177)),(to_sfixed_a(-0.10425978153944016)),(to_sfixed_a(0.11914639919996262)),(to_sfixed_a(-0.09411564469337463)),(to_sfixed_a(-0.12013483047485352)),(to_sfixed_a(0.031581632792949677)),(to_sfixed_a(0.0038119822274893522)),(to_sfixed_a(0.14845839142799377)),(to_sfixed_a(0.16545401513576508)),(to_sfixed_a(-0.11341828852891922)),(to_sfixed_a(0.1002822294831276)),(to_sfixed_a(-0.0026304125785827637)),(to_sfixed_a(-0.12182163447141647)),(to_sfixed_a(-0.33735859394073486)),(to_sfixed_a(-0.03988572582602501)),(to_sfixed_a(0.25928711891174316)),(to_sfixed_a(-0.1532348394393921)),(to_sfixed_a(-0.1257760375738144)),(to_sfixed_a(-0.012375893071293831)),(to_sfixed_a(0.00015286738926079124)),(to_sfixed_a(-4.237256507622078e-05)),(to_sfixed_a(4.6144891712174285e-06)),(to_sfixed_a(3.7003828765591606e-05)),(to_sfixed_a(0.00025483217905275524)),(to_sfixed_a(-5.453435369418003e-05)),(to_sfixed_a(0.06429444253444672)),(to_sfixed_a(0.001807172317057848)),(to_sfixed_a(0.11266036331653595)),(to_sfixed_a(0.06634758412837982)),(to_sfixed_a(0.12436096370220184)),(to_sfixed_a(-0.10848995298147202)),(to_sfixed_a(0.21992522478103638)),(to_sfixed_a(0.44670453667640686)),(to_sfixed_a(0.11103774607181549)),(to_sfixed_a(-0.07920640707015991)),(to_sfixed_a(0.08856220543384552)),(to_sfixed_a(0.11243633180856705)),(to_sfixed_a(0.14948797225952148)),(to_sfixed_a(-0.1474774032831192)),(to_sfixed_a(-0.20039910078048706)),(to_sfixed_a(-0.12321451306343079)),(to_sfixed_a(0.026189785450696945)),(to_sfixed_a(0.0874502956867218)),(to_sfixed_a(0.28561607003211975)),(to_sfixed_a(-0.054535478353500366)),(to_sfixed_a(-0.3155257999897003)),(to_sfixed_a(-3.358598769409582e-05)),(to_sfixed_a(1.8174545402871445e-05)),(to_sfixed_a(1.2095976671844255e-05)),(to_sfixed_a(-3.922842552128714e-06)),(to_sfixed_a(-3.66204149031546e-05)),(to_sfixed_a(-0.00011556276149349287)),(to_sfixed_a(0.00022681395057588816)),(to_sfixed_a(-5.5584536312380806e-05)),(to_sfixed_a(0.005532704293727875)),(to_sfixed_a(-0.027401765808463097)),(to_sfixed_a(0.11260396242141724)),(to_sfixed_a(0.24614201486110687)),(to_sfixed_a(-0.06280829012393951)),(to_sfixed_a(0.0802132859826088)),(to_sfixed_a(-0.1305728554725647)),(to_sfixed_a(-0.040936440229415894)),(to_sfixed_a(0.06777364760637283)),(to_sfixed_a(-0.1189751923084259)),(to_sfixed_a(-0.11376161128282547)),(to_sfixed_a(-0.00328060332685709)),(to_sfixed_a(0.24718280136585236)),(to_sfixed_a(-0.15212880074977875)),(to_sfixed_a(-0.18328729271888733)),(to_sfixed_a(0.2598326802253723)),(to_sfixed_a(0.030988037586212158)),(to_sfixed_a(-0.19225120544433594)),(to_sfixed_a(-0.11765579879283905)),(to_sfixed_a(-0.12891031801700592)),(to_sfixed_a(-0.07924965023994446)),(to_sfixed_a(-4.525809708866291e-05)),(to_sfixed_a(6.079221930122003e-05)),(to_sfixed_a(2.981091893161647e-05)),(to_sfixed_a(-0.00014794705202803016)),(to_sfixed_a(7.79848123784177e-05)),(to_sfixed_a(-5.4306339734466746e-05)),(to_sfixed_a(-0.00016247029998339713)),(to_sfixed_a(-0.01964118890464306)),(to_sfixed_a(0.0006803981377743185)),(to_sfixed_a(0.045023396611213684)),(to_sfixed_a(0.1857362985610962)),(to_sfixed_a(0.18801410496234894)),(to_sfixed_a(0.02674981579184532)),(to_sfixed_a(0.13939303159713745)),(to_sfixed_a(-0.06246937811374664)),(to_sfixed_a(-0.16167370975017548)),(to_sfixed_a(-0.014449615962803364)),(to_sfixed_a(-0.005742230918258429)),(to_sfixed_a(0.060378044843673706)),(to_sfixed_a(-0.039100684225559235)),(to_sfixed_a(0.09001344442367554)),(to_sfixed_a(-0.11805714666843414)),(to_sfixed_a(0.06583777815103531)),(to_sfixed_a(-0.41142383217811584)),(to_sfixed_a(-0.13475999236106873)),(to_sfixed_a(-0.20621728897094727)),(to_sfixed_a(-0.0011608863715082407)),(to_sfixed_a(-0.01065812911838293)),(to_sfixed_a(-0.00011987634206889197)),(to_sfixed_a(0.00015290601004380733)),(to_sfixed_a(-0.00014951106277294457)),(to_sfixed_a(2.604361725389026e-05)),(to_sfixed_a(-6.434341776184738e-05)),(to_sfixed_a(-5.997331390972249e-05)),(to_sfixed_a(3.5147244489053264e-05)),(to_sfixed_a(-0.00024906493490561843)),(to_sfixed_a(0.10462278127670288)),(to_sfixed_a(0.07230917364358902)),(to_sfixed_a(0.17865590751171112)),(to_sfixed_a(0.10313618183135986)),(to_sfixed_a(0.005723987706005573)),(to_sfixed_a(0.052615754306316376)),(to_sfixed_a(-0.08847609162330627)),(to_sfixed_a(-0.0909397229552269)),(to_sfixed_a(0.0015107858926057816)),(to_sfixed_a(-0.006646226160228252)),(to_sfixed_a(-0.0034025334753096104)),(to_sfixed_a(-0.03258560970425606)),(to_sfixed_a(0.28091341257095337)),(to_sfixed_a(0.35967937111854553)),(to_sfixed_a(0.20544150471687317)),(to_sfixed_a(-0.05327916145324707)),(to_sfixed_a(0.0004347253998275846)),(to_sfixed_a(0.004315023776143789)),(to_sfixed_a(-0.007437442895025015)),(to_sfixed_a(-1.78575464815367e-05)),(to_sfixed_a(-0.00023183110170066357)),(to_sfixed_a(-0.00011759916378650814)),(to_sfixed_a(-9.569583926349878e-05)),(to_sfixed_a(0.00017246489005628973)),(to_sfixed_a(-3.212386218365282e-05)),(to_sfixed_a(0.00014249597734306008)),(to_sfixed_a(-3.86338506359607e-05)),(to_sfixed_a(-0.0002852746983990073)),(to_sfixed_a(0.003521847305819392)),(to_sfixed_a(0.058834753930568695)),(to_sfixed_a(0.22591425478458405)),(to_sfixed_a(-0.0996127650141716)),(to_sfixed_a(0.08835846185684204)),(to_sfixed_a(-0.06948301941156387)),(to_sfixed_a(0.01230558194220066)),(to_sfixed_a(0.018007496371865273)),(to_sfixed_a(-0.00894426740705967)),(to_sfixed_a(0.023180721327662468)),(to_sfixed_a(0.1878196895122528)),(to_sfixed_a(0.2087540477514267)),(to_sfixed_a(0.3282504975795746)),(to_sfixed_a(-0.07073628902435303)),(to_sfixed_a(-0.05077078193426132)),(to_sfixed_a(0.09558673948049545)),(to_sfixed_a(-0.05198622867465019)),(to_sfixed_a(-0.006327747832983732)),(to_sfixed_a(-0.034326113760471344)),(to_sfixed_a(0.00011185697076143697)),(to_sfixed_a(-8.345951937371865e-05)),(to_sfixed_a(2.6946595426124986e-06)),(to_sfixed_a(5.516894088941626e-05)),(to_sfixed_a(-1.6348034478141926e-05)),(to_sfixed_a(7.84394251240883e-06)),(to_sfixed_a(-0.00012733660696540028)),(to_sfixed_a(0.00018353214545641094)),(to_sfixed_a(0.012952552177011967)),(to_sfixed_a(0.004910452291369438)),(to_sfixed_a(0.054898325353860855)),(to_sfixed_a(-0.1101529523730278)),(to_sfixed_a(-0.12248607724905014)),(to_sfixed_a(-0.030938059091567993)),(to_sfixed_a(0.08739389479160309)),(to_sfixed_a(0.10078460723161697)),(to_sfixed_a(-0.23040525615215302)),(to_sfixed_a(0.14531175792217255)),(to_sfixed_a(0.06403934955596924)),(to_sfixed_a(0.028272489085793495)),(to_sfixed_a(-0.1781429797410965)),(to_sfixed_a(-0.10478933155536652)),(to_sfixed_a(-0.07666032016277313)),(to_sfixed_a(-0.06155017390847206)),(to_sfixed_a(-0.012008593417704105)),(to_sfixed_a(-0.04046212509274483)),(to_sfixed_a(-0.01799394004046917)),(to_sfixed_a(0.0039717708714306355)),(to_sfixed_a(0.00011360512144165114)),(to_sfixed_a(-0.0002755279710981995)),(to_sfixed_a(-9.408008918398991e-05)),(to_sfixed_a(3.726442810148001e-05)),(to_sfixed_a(1.8319726677873405e-06)),(to_sfixed_a(-0.00017350375128444284)),(to_sfixed_a(-8.554747182643041e-05)),(to_sfixed_a(-2.2609366112646967e-07)),(to_sfixed_a(-0.00015957839787006378)),(to_sfixed_a(-0.020437851548194885)),(to_sfixed_a(0.032681290060281754)),(to_sfixed_a(0.0625031441450119)),(to_sfixed_a(-0.0031644096598029137)),(to_sfixed_a(0.08676464110612869)),(to_sfixed_a(-0.020312899723649025)),(to_sfixed_a(0.05576645955443382)),(to_sfixed_a(0.08766211569309235)),(to_sfixed_a(-0.05914780870079994)),(to_sfixed_a(-0.004544203635305166)),(to_sfixed_a(0.02456613816320896)),(to_sfixed_a(0.06432884931564331)),(to_sfixed_a(-0.02304689958691597)),(to_sfixed_a(0.005342530086636543)),(to_sfixed_a(0.13095848262310028)),(to_sfixed_a(0.03474458307027817)),(to_sfixed_a(-0.001949957455508411)),(to_sfixed_a(-0.0005135233514010906)),(to_sfixed_a(-0.0002933467330876738)),(to_sfixed_a(4.815966167370789e-05)),(to_sfixed_a(0.0002624169865157455)),(to_sfixed_a(7.543472747784108e-05)),(to_sfixed_a(-4.869539770879783e-05)),(to_sfixed_a(0.00019316091493237764)),(to_sfixed_a(-9.962026524590328e-05)),(to_sfixed_a(0.00015132992120925337)),(to_sfixed_a(-2.2909294784767553e-05)),(to_sfixed_a(0.00010775063128676265)),(to_sfixed_a(0.0016512532019987702)),(to_sfixed_a(0.001462645479477942)),(to_sfixed_a(-0.00010678569378796965)),(to_sfixed_a(0.0002299516199855134)),(to_sfixed_a(-0.00027990539092570543)),(to_sfixed_a(0.04216180741786957)),(to_sfixed_a(0.003697935026139021)),(to_sfixed_a(0.00040355612873099744)),(to_sfixed_a(0.0340036004781723)),(to_sfixed_a(0.17329449951648712)),(to_sfixed_a(0.007484195288270712)),(to_sfixed_a(0.09746396541595459)),(to_sfixed_a(0.03248074650764465)),(to_sfixed_a(0.045328155159950256)),(to_sfixed_a(0.0035259302239865065)),(to_sfixed_a(7.439499313477427e-05)),(to_sfixed_a(-4.128000000491738e-05)),(to_sfixed_a(0.00013614268391393125)),(to_sfixed_a(-9.306208812631667e-05)),(to_sfixed_a(2.2666210497845896e-05)),(to_sfixed_a(0.0001810889079933986)),(to_sfixed_a(-8.77081311045913e-06)),(to_sfixed_a(0.00010709856724133715)),(to_sfixed_a(0.0001398407039232552)),(to_sfixed_a(0.00011289623216725886)),(to_sfixed_a(-0.00014762271894142032)),(to_sfixed_a(0.00012581217742990702)),(to_sfixed_a(0.0002349128626519814)),(to_sfixed_a(-0.00011682980402838439)),(to_sfixed_a(0.00036010026815347373)),(to_sfixed_a(7.164295675465837e-05)),(to_sfixed_a(-0.00011087587336078286)),(to_sfixed_a(-5.4479929531225935e-05)),(to_sfixed_a(0.0001383542112307623)),(to_sfixed_a(-0.00012502724712248892)),(to_sfixed_a(-2.9426970286294818e-05)),(to_sfixed_a(-3.277572614024393e-05)),(to_sfixed_a(5.188133582123555e-05)),(to_sfixed_a(1.732945383992046e-05)),(to_sfixed_a(-0.00015572045231238008)),(to_sfixed_a(-2.8717298846459016e-05)),(to_sfixed_a(2.7137935830978677e-05)),(to_sfixed_a(0.00027630478143692017)),(to_sfixed_a(-0.00017945253057405353)),(to_sfixed_a(0.00025136888143606484)),(to_sfixed_a(-5.540979327633977e-05)),(to_sfixed_a(-0.00017450738232582808)),(to_sfixed_a(0.00020804960513487458)),(to_sfixed_a(-0.00010705753084039316)),(to_sfixed_a(-0.00018655238091014326)),(to_sfixed_a(-0.00010714095697039738)));

    constant weight_n0_20 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(0.00012536464782897383)),(to_sfixed_a(-1.2107447219023015e-05)),(to_sfixed_a(3.9239628677023575e-05)),(to_sfixed_a(3.206163091817871e-05)),(to_sfixed_a(-9.514205885352567e-05)),(to_sfixed_a(-0.00011592986265895888)),(to_sfixed_a(7.610081229358912e-05)),(to_sfixed_a(-7.581894897157326e-05)),(to_sfixed_a(0.0001371445250697434)),(to_sfixed_a(-9.128804231295362e-05)),(to_sfixed_a(4.6230499719968066e-05)),(to_sfixed_a(0.000247832213062793)),(to_sfixed_a(-9.40041572903283e-05)),(to_sfixed_a(-3.41367231158074e-05)),(to_sfixed_a(-9.225304529536515e-05)),(to_sfixed_a(0.0002516078529879451)),(to_sfixed_a(0.00018670344434212893)),(to_sfixed_a(6.113809649832547e-05)),(to_sfixed_a(-3.380468115210533e-05)),(to_sfixed_a(9.876306285150349e-05)),(to_sfixed_a(6.512118125101551e-05)),(to_sfixed_a(7.273726077983156e-05)),(to_sfixed_a(0.00012013055675197393)),(to_sfixed_a(5.300616248860024e-05)),(to_sfixed_a(0.00016154356126207858)),(to_sfixed_a(0.00013676715025212616)),(to_sfixed_a(0.0001893384469440207)),(to_sfixed_a(0.00017619428399484605)),(to_sfixed_a(-0.0004688926273956895)),(to_sfixed_a(0.00020430532458703965)),(to_sfixed_a(-8.757108298595995e-05)),(to_sfixed_a(-0.00027747623971663415)),(to_sfixed_a(0.00010257036774419248)),(to_sfixed_a(-1.0518900126044173e-05)),(to_sfixed_a(4.700766294263303e-05)),(to_sfixed_a(-5.570935536525212e-05)),(to_sfixed_a(0.00014560241834260523)),(to_sfixed_a(0.00010028523684013635)),(to_sfixed_a(0.00011968462786171585)),(to_sfixed_a(0.00012375650112517178)),(to_sfixed_a(-0.00013681322161573917)),(to_sfixed_a(-0.000169165781699121)),(to_sfixed_a(-5.735210288548842e-05)),(to_sfixed_a(-0.00016116305778268725)),(to_sfixed_a(0.00018417534010950476)),(to_sfixed_a(2.8185779228806496e-05)),(to_sfixed_a(0.00014487706357613206)),(to_sfixed_a(-0.00016571245214436203)),(to_sfixed_a(-0.00021330731397029012)),(to_sfixed_a(-9.281514212489128e-05)),(to_sfixed_a(-0.0003048184444196522)),(to_sfixed_a(-0.00014826840197201818)),(to_sfixed_a(-6.13498268648982e-05)),(to_sfixed_a(0.0003033755347132683)),(to_sfixed_a(-1.1325792002025992e-05)),(to_sfixed_a(6.059676888980903e-05)),(to_sfixed_a(0.0002015055069932714)),(to_sfixed_a(-0.0002113864029524848)),(to_sfixed_a(0.00013457149907480925)),(to_sfixed_a(2.9330654797377065e-05)),(to_sfixed_a(-0.00039521133294329047)),(to_sfixed_a(-9.804506407817826e-05)),(to_sfixed_a(0.00019965007959399372)),(to_sfixed_a(4.037158578285016e-05)),(to_sfixed_a(5.59331092517823e-05)),(to_sfixed_a(-0.00014669356460217386)),(to_sfixed_a(0.00021677723270840943)),(to_sfixed_a(-0.0001296142872888595)),(to_sfixed_a(7.547475979663432e-05)),(to_sfixed_a(-0.00691543985158205)),(to_sfixed_a(0.00010100812505697832)),(to_sfixed_a(0.00010429327812744305)),(to_sfixed_a(-2.6128431272809394e-05)),(to_sfixed_a(-0.00020652066450566053)),(to_sfixed_a(-7.540943624917418e-05)),(to_sfixed_a(-0.00019798180437646806)),(to_sfixed_a(-3.834102608379908e-05)),(to_sfixed_a(0.00022910944244358689)),(to_sfixed_a(-3.4712582419160753e-05)),(to_sfixed_a(-4.8581758164800704e-05)),(to_sfixed_a(6.948258669581264e-05)),(to_sfixed_a(8.675747085362673e-05)),(to_sfixed_a(-0.00010175833449466154)),(to_sfixed_a(-4.8853991756914183e-05)),(to_sfixed_a(4.582476685754955e-05)),(to_sfixed_a(-0.00021009058400522918)),(to_sfixed_a(1.5630288544343784e-05)),(to_sfixed_a(-8.830478327581659e-05)),(to_sfixed_a(-7.400592585327104e-05)),(to_sfixed_a(1.279203479498392e-05)),(to_sfixed_a(5.412485552369617e-05)),(to_sfixed_a(-8.002274989848956e-05)),(to_sfixed_a(0.0651337206363678)),(to_sfixed_a(8.527484897058457e-05)),(to_sfixed_a(0.07343969494104385)),(to_sfixed_a(-0.022142408415675163)),(to_sfixed_a(0.02419697307050228)),(to_sfixed_a(0.002266489900648594)),(to_sfixed_a(0.0913434624671936)),(to_sfixed_a(0.006467632483690977)),(to_sfixed_a(-0.030042072758078575)),(to_sfixed_a(-0.07970396429300308)),(to_sfixed_a(-0.06364718824625015)),(to_sfixed_a(0.04629051312804222)),(to_sfixed_a(0.03383995220065117)),(to_sfixed_a(0.06853369623422623)),(to_sfixed_a(-1.809988680179231e-05)),(to_sfixed_a(-0.00017715264402795583)),(to_sfixed_a(6.794669752707705e-05)),(to_sfixed_a(9.737468644743785e-05)),(to_sfixed_a(7.030020788079128e-05)),(to_sfixed_a(-0.00029841504874639213)),(to_sfixed_a(2.968158332805615e-05)),(to_sfixed_a(0.00014170700160320848)),(to_sfixed_a(0.0001965090341400355)),(to_sfixed_a(4.420880213729106e-05)),(to_sfixed_a(6.758757081115618e-06)),(to_sfixed_a(-0.00017580624262336642)),(to_sfixed_a(-0.0011334751034155488)),(to_sfixed_a(-0.01666237786412239)),(to_sfixed_a(-0.04906130209565163)),(to_sfixed_a(0.09287887066602707)),(to_sfixed_a(0.11494611948728561)),(to_sfixed_a(-0.023078152909874916)),(to_sfixed_a(-0.11048334836959839)),(to_sfixed_a(-0.13146398961544037)),(to_sfixed_a(-0.21919351816177368)),(to_sfixed_a(0.04458348825573921)),(to_sfixed_a(0.017299972474575043)),(to_sfixed_a(-0.033596768975257874)),(to_sfixed_a(0.061950232833623886)),(to_sfixed_a(-0.03440923988819122)),(to_sfixed_a(0.016139410436153412)),(to_sfixed_a(-0.05210332199931145)),(to_sfixed_a(-0.0026978901587426662)),(to_sfixed_a(7.00197197147645e-05)),(to_sfixed_a(-0.0011341844219714403)),(to_sfixed_a(-0.00011533211363712326)),(to_sfixed_a(-9.647782280808315e-05)),(to_sfixed_a(-0.00010342942550778389)),(to_sfixed_a(-5.0311946324654855e-06)),(to_sfixed_a(0.0003742648405022919)),(to_sfixed_a(0.0002569119387771934)),(to_sfixed_a(0.000110307963041123)),(to_sfixed_a(-0.0015512093668803573)),(to_sfixed_a(-0.04004305973649025)),(to_sfixed_a(-0.018228763714432716)),(to_sfixed_a(-0.07489564269781113)),(to_sfixed_a(-0.029033271595835686)),(to_sfixed_a(0.019814016297459602)),(to_sfixed_a(-0.04449257254600525)),(to_sfixed_a(-0.030768338590860367)),(to_sfixed_a(-0.034930601716041565)),(to_sfixed_a(-0.1874258816242218)),(to_sfixed_a(-0.06846826523542404)),(to_sfixed_a(-0.032838620245456696)),(to_sfixed_a(-0.07975400984287262)),(to_sfixed_a(0.07222291082143784)),(to_sfixed_a(-0.043606534600257874)),(to_sfixed_a(0.03372346609830856)),(to_sfixed_a(-0.07912414520978928)),(to_sfixed_a(0.15797226130962372)),(to_sfixed_a(-0.0014203810133039951)),(to_sfixed_a(0.05712167173624039)),(to_sfixed_a(-0.004327904433012009)),(to_sfixed_a(-0.00021597841987386346)),(to_sfixed_a(0.00012356704974081367)),(to_sfixed_a(0.0001095575062208809)),(to_sfixed_a(-0.00025916300364769995)),(to_sfixed_a(0.00018575810827314854)),(to_sfixed_a(-2.260875362480874e-06)),(to_sfixed_a(9.104425407713279e-05)),(to_sfixed_a(3.458213905105367e-05)),(to_sfixed_a(-0.03413194790482521)),(to_sfixed_a(0.07629909366369247)),(to_sfixed_a(0.015023160725831985)),(to_sfixed_a(0.08434377610683441)),(to_sfixed_a(0.029382064938545227)),(to_sfixed_a(0.06303965300321579)),(to_sfixed_a(-0.031319696456193924)),(to_sfixed_a(0.04098097234964371)),(to_sfixed_a(-0.0688929334282875)),(to_sfixed_a(0.06759103387594223)),(to_sfixed_a(-0.11243125796318054)),(to_sfixed_a(0.11723656952381134)),(to_sfixed_a(0.013923716731369495)),(to_sfixed_a(-0.07756710797548294)),(to_sfixed_a(-0.1480013132095337)),(to_sfixed_a(0.17432266473770142)),(to_sfixed_a(0.005508624482899904)),(to_sfixed_a(-0.045093830674886703)),(to_sfixed_a(-0.1660265177488327)),(to_sfixed_a(7.180206011980772e-05)),(to_sfixed_a(0.00035651595680974424)),(to_sfixed_a(0.001611283514648676)),(to_sfixed_a(2.9662753149750642e-05)),(to_sfixed_a(2.4148295779014006e-05)),(to_sfixed_a(0.0002658739686012268)),(to_sfixed_a(0.00017536283121444285)),(to_sfixed_a(8.292732672998682e-05)),(to_sfixed_a(-7.011520210653543e-05)),(to_sfixed_a(0.030824579298496246)),(to_sfixed_a(0.02772153727710247)),(to_sfixed_a(0.013255741447210312)),(to_sfixed_a(0.0012965328060090542)),(to_sfixed_a(-0.014655087143182755)),(to_sfixed_a(-0.06200461462140083)),(to_sfixed_a(-0.2517933249473572)),(to_sfixed_a(-0.09237191826105118)),(to_sfixed_a(-0.09873495250940323)),(to_sfixed_a(0.04692740738391876)),(to_sfixed_a(0.10975795239210129)),(to_sfixed_a(-0.18821948766708374)),(to_sfixed_a(-0.016058871522545815)),(to_sfixed_a(0.011790123768150806)),(to_sfixed_a(-0.07854815572500229)),(to_sfixed_a(0.12603458762168884)),(to_sfixed_a(-0.27659040689468384)),(to_sfixed_a(0.08562543988227844)),(to_sfixed_a(-0.1431204378604889)),(to_sfixed_a(-0.00527580501511693)),(to_sfixed_a(-0.0018128042574971914)),(to_sfixed_a(-5.421271634986624e-05)),(to_sfixed_a(-2.9235536203486845e-05)),(to_sfixed_a(5.664316631737165e-06)),(to_sfixed_a(-0.00018335357890464365)),(to_sfixed_a(-0.00011021925456589088)),(to_sfixed_a(-0.00011646490747807547)),(to_sfixed_a(-0.058116212487220764)),(to_sfixed_a(0.0010842165211215615)),(to_sfixed_a(0.02444022335112095)),(to_sfixed_a(0.17631952464580536)),(to_sfixed_a(0.038729287683963776)),(to_sfixed_a(-0.15727034211158752)),(to_sfixed_a(-0.10022763907909393)),(to_sfixed_a(-0.010932350531220436)),(to_sfixed_a(-0.1890251189470291)),(to_sfixed_a(-0.18644960224628448)),(to_sfixed_a(0.11161366105079651)),(to_sfixed_a(0.027140047401189804)),(to_sfixed_a(0.15028716623783112)),(to_sfixed_a(-0.12055611610412598)),(to_sfixed_a(0.021445099264383316)),(to_sfixed_a(0.1567540168762207)),(to_sfixed_a(0.16391780972480774)),(to_sfixed_a(-0.07805463671684265)),(to_sfixed_a(-0.16767218708992004)),(to_sfixed_a(0.10721073299646378)),(to_sfixed_a(0.03574333339929581)),(to_sfixed_a(-0.1062270775437355)),(to_sfixed_a(-2.4943969947344158e-06)),(to_sfixed_a(3.9416030631400645e-05)),(to_sfixed_a(-3.9499638660345227e-05)),(to_sfixed_a(0.0004019125481136143)),(to_sfixed_a(0.00018452842778060585)),(to_sfixed_a(8.413856266997755e-05)),(to_sfixed_a(-0.0018946846248582006)),(to_sfixed_a(-0.08684205263853073)),(to_sfixed_a(0.0060214814729988575)),(to_sfixed_a(-0.02354259043931961)),(to_sfixed_a(0.13839568197727203)),(to_sfixed_a(0.004784027114510536)),(to_sfixed_a(0.07043642550706863)),(to_sfixed_a(0.006791336461901665)),(to_sfixed_a(-0.14995403587818146)),(to_sfixed_a(0.21106362342834473)),(to_sfixed_a(0.2825857996940613)),(to_sfixed_a(0.08142221719026566)),(to_sfixed_a(0.4062405526638031)),(to_sfixed_a(-0.0869695171713829)),(to_sfixed_a(0.1316094845533371)),(to_sfixed_a(0.2847481667995453)),(to_sfixed_a(-0.009833608753979206)),(to_sfixed_a(0.012934036552906036)),(to_sfixed_a(0.0022373783867806196)),(to_sfixed_a(-0.3640934228897095)),(to_sfixed_a(-0.26714229583740234)),(to_sfixed_a(-1.4334373190649785e-05)),(to_sfixed_a(-7.629444007761776e-05)),(to_sfixed_a(0.00024479557760059834)),(to_sfixed_a(9.580483606441703e-08)),(to_sfixed_a(0.00021161313634365797)),(to_sfixed_a(-0.00022523061488755047)),(to_sfixed_a(-8.985718159237877e-05)),(to_sfixed_a(-0.007493758574128151)),(to_sfixed_a(0.05072988569736481)),(to_sfixed_a(-0.19433769583702087)),(to_sfixed_a(0.05939451977610588)),(to_sfixed_a(-0.015864264219999313)),(to_sfixed_a(0.002981245517730713)),(to_sfixed_a(-0.05195599049329758)),(to_sfixed_a(0.11481322348117828)),(to_sfixed_a(0.06833179295063019)),(to_sfixed_a(0.17264889180660248)),(to_sfixed_a(0.14145086705684662)),(to_sfixed_a(-0.5975003242492676)),(to_sfixed_a(-0.2497156262397766)),(to_sfixed_a(-0.1845465749502182)),(to_sfixed_a(0.17964161932468414)),(to_sfixed_a(-0.0686245709657669)),(to_sfixed_a(0.03354200720787048)),(to_sfixed_a(-0.006937668193131685)),(to_sfixed_a(-0.11951565742492676)),(to_sfixed_a(-0.4594510793685913)),(to_sfixed_a(-0.10952682048082352)),(to_sfixed_a(0.0014789134729653597)),(to_sfixed_a(-2.565631439210847e-05)),(to_sfixed_a(4.8466547013958916e-05)),(to_sfixed_a(0.00012005594180664048)),(to_sfixed_a(-0.0001318162976531312)),(to_sfixed_a(-0.0003558879834599793)),(to_sfixed_a(-0.029366154223680496)),(to_sfixed_a(-0.0190743375569582)),(to_sfixed_a(0.16407689452171326)),(to_sfixed_a(-0.008780032396316528)),(to_sfixed_a(-0.031812358647584915)),(to_sfixed_a(-0.05203450098633766)),(to_sfixed_a(0.07594229280948639)),(to_sfixed_a(0.07803197205066681)),(to_sfixed_a(0.16177822649478912)),(to_sfixed_a(0.061091575771570206)),(to_sfixed_a(0.2951401472091675)),(to_sfixed_a(-0.09847186505794525)),(to_sfixed_a(-0.09481649845838547)),(to_sfixed_a(-0.15812364220619202)),(to_sfixed_a(0.3457990884780884)),(to_sfixed_a(0.5019026398658752)),(to_sfixed_a(-0.2746347188949585)),(to_sfixed_a(-0.13198481500148773)),(to_sfixed_a(-0.07500281929969788)),(to_sfixed_a(-0.0882895365357399)),(to_sfixed_a(-0.3389888405799866)),(to_sfixed_a(-0.12863054871559143)),(to_sfixed_a(7.056443428155035e-05)),(to_sfixed_a(0.0002468482998665422)),(to_sfixed_a(0.0002270063996547833)),(to_sfixed_a(7.827753142919391e-05)),(to_sfixed_a(5.622874232358299e-05)),(to_sfixed_a(0.00011312533752061427)),(to_sfixed_a(0.00013725385360885412)),(to_sfixed_a(0.18558308482170105)),(to_sfixed_a(0.11796024441719055)),(to_sfixed_a(0.09104876965284348)),(to_sfixed_a(-0.16793403029441833)),(to_sfixed_a(-0.10276991128921509)),(to_sfixed_a(0.06494864821434021)),(to_sfixed_a(0.05729643628001213)),(to_sfixed_a(-0.16969451308250427)),(to_sfixed_a(0.1769874095916748)),(to_sfixed_a(-0.028318505734205246)),(to_sfixed_a(-0.07753996551036835)),(to_sfixed_a(-0.49422964453697205)),(to_sfixed_a(0.12674611806869507)),(to_sfixed_a(0.6473947763442993)),(to_sfixed_a(0.25616031885147095)),(to_sfixed_a(0.21128307282924652)),(to_sfixed_a(-0.22164173424243927)),(to_sfixed_a(-0.14130578935146332)),(to_sfixed_a(-0.14115789532661438)),(to_sfixed_a(-0.02403693087399006)),(to_sfixed_a(-0.06894046068191528)),(to_sfixed_a(-0.00010386545909568667)),(to_sfixed_a(9.078061702894047e-05)),(to_sfixed_a(6.744639540556818e-05)),(to_sfixed_a(0.0003592232533264905)),(to_sfixed_a(8.63347013364546e-05)),(to_sfixed_a(-0.00022965052630752325)),(to_sfixed_a(0.00015866640023887157)),(to_sfixed_a(-0.010998370125889778)),(to_sfixed_a(0.1252477616071701)),(to_sfixed_a(0.11122828722000122)),(to_sfixed_a(-0.01970929093658924)),(to_sfixed_a(0.028061987832188606)),(to_sfixed_a(-0.15913830697536469)),(to_sfixed_a(-0.1693321168422699)),(to_sfixed_a(0.13474206626415253)),(to_sfixed_a(-0.08482702821493149)),(to_sfixed_a(0.03360350430011749)),(to_sfixed_a(-0.19419990479946136)),(to_sfixed_a(0.016926461830735207)),(to_sfixed_a(0.07631279528141022)),(to_sfixed_a(0.4444698989391327)),(to_sfixed_a(0.17307806015014648)),(to_sfixed_a(0.1519119292497635)),(to_sfixed_a(0.037601031363010406)),(to_sfixed_a(0.19984391331672668)),(to_sfixed_a(-0.12840953469276428)),(to_sfixed_a(-0.15497148036956787)),(to_sfixed_a(0.08430768549442291)),(to_sfixed_a(0.0020231378730386496)),(to_sfixed_a(0.0022486294619739056)),(to_sfixed_a(-6.517582369269803e-05)),(to_sfixed_a(1.9684279322973453e-05)),(to_sfixed_a(-0.00019222831178922206)),(to_sfixed_a(-0.00039335727342404425)),(to_sfixed_a(9.726217103889212e-05)),(to_sfixed_a(-0.0010644809808582067)),(to_sfixed_a(-0.16724129021167755)),(to_sfixed_a(-0.15388692915439606)),(to_sfixed_a(-0.39797401428222656)),(to_sfixed_a(-0.11936885118484497)),(to_sfixed_a(-0.18274563550949097)),(to_sfixed_a(0.11712056398391724)),(to_sfixed_a(0.16458848118782043)),(to_sfixed_a(-0.2094154953956604)),(to_sfixed_a(-0.025119761005043983)),(to_sfixed_a(0.15918052196502686)),(to_sfixed_a(-0.1990981101989746)),(to_sfixed_a(0.07050256431102753)),(to_sfixed_a(0.24464379251003265)),(to_sfixed_a(0.10135284811258316)),(to_sfixed_a(-0.01801108941435814)),(to_sfixed_a(0.2422734498977661)),(to_sfixed_a(0.09134563058614731)),(to_sfixed_a(0.08305395394563675)),(to_sfixed_a(-0.1953340470790863)),(to_sfixed_a(0.13768482208251953)),(to_sfixed_a(-0.00027550317463465035)),(to_sfixed_a(-0.0001819590397644788)),(to_sfixed_a(-0.00022818367870058864)),(to_sfixed_a(-0.00018289363652002066)),(to_sfixed_a(-6.530146492877975e-05)),(to_sfixed_a(0.00027786302962340415)),(to_sfixed_a(-9.778505773283541e-05)),(to_sfixed_a(-0.012603502720594406)),(to_sfixed_a(-0.19953791797161102)),(to_sfixed_a(0.01182022225111723)),(to_sfixed_a(0.017346559092402458)),(to_sfixed_a(0.09275370836257935)),(to_sfixed_a(0.12167034298181534)),(to_sfixed_a(-0.0010388153605163097)),(to_sfixed_a(0.027658432722091675)),(to_sfixed_a(-0.15427210927009583)),(to_sfixed_a(0.1621948927640915)),(to_sfixed_a(-0.21556951105594635)),(to_sfixed_a(-0.21465951204299927)),(to_sfixed_a(0.31728288531303406)),(to_sfixed_a(0.03284728154540062)),(to_sfixed_a(0.16751781105995178)),(to_sfixed_a(-0.30083218216896057)),(to_sfixed_a(0.15831713378429413)),(to_sfixed_a(0.16103723645210266)),(to_sfixed_a(-0.05449046194553375)),(to_sfixed_a(-0.13860639929771423)),(to_sfixed_a(-0.23528866469860077)),(to_sfixed_a(-0.00032309783273376524)),(to_sfixed_a(0.00011796656326623634)),(to_sfixed_a(-6.216868314368185e-06)),(to_sfixed_a(-0.00023949475144036114)),(to_sfixed_a(1.1053777598135639e-05)),(to_sfixed_a(4.705226274381857e-06)),(to_sfixed_a(0.001176738180220127)),(to_sfixed_a(0.16897845268249512)),(to_sfixed_a(0.2831612229347229)),(to_sfixed_a(0.3634142279624939)),(to_sfixed_a(0.16178399324417114)),(to_sfixed_a(0.0722392350435257)),(to_sfixed_a(-0.09229356050491333)),(to_sfixed_a(-0.13626517355442047)),(to_sfixed_a(0.1912323236465454)),(to_sfixed_a(-0.13766595721244812)),(to_sfixed_a(-0.023953676223754883)),(to_sfixed_a(0.012040539644658566)),(to_sfixed_a(-0.32034003734588623)),(to_sfixed_a(0.23114310204982758)),(to_sfixed_a(-0.26991453766822815)),(to_sfixed_a(-0.13980668783187866)),(to_sfixed_a(-0.08290374279022217)),(to_sfixed_a(-0.023510858416557312)),(to_sfixed_a(0.18257616460323334)),(to_sfixed_a(-0.15825314819812775)),(to_sfixed_a(-0.06674107909202576)),(to_sfixed_a(0.013705329969525337)),(to_sfixed_a(-0.005888373591005802)),(to_sfixed_a(-7.453514263033867e-05)),(to_sfixed_a(0.00011038490629289299)),(to_sfixed_a(6.540618051076308e-05)),(to_sfixed_a(0.00024951985687948763)),(to_sfixed_a(-7.639092655153945e-05)),(to_sfixed_a(0.0010054714512079954)),(to_sfixed_a(-0.006123484577983618)),(to_sfixed_a(0.1342388242483139)),(to_sfixed_a(0.031825724989175797)),(to_sfixed_a(-0.41580983996391296)),(to_sfixed_a(-0.0015465931501239538)),(to_sfixed_a(-0.06860006600618362)),(to_sfixed_a(0.04082668572664261)),(to_sfixed_a(0.2301381379365921)),(to_sfixed_a(-0.2508836090564728)),(to_sfixed_a(-0.13031229376792908)),(to_sfixed_a(0.02961418218910694)),(to_sfixed_a(-0.13653495907783508)),(to_sfixed_a(0.028277654200792313)),(to_sfixed_a(-0.04034902900457382)),(to_sfixed_a(-0.07457315176725388)),(to_sfixed_a(-0.2987327575683594)),(to_sfixed_a(-0.025815272703766823)),(to_sfixed_a(0.022407805547118187)),(to_sfixed_a(-0.05305134132504463)),(to_sfixed_a(-0.05745478346943855)),(to_sfixed_a(7.436938176397234e-05)),(to_sfixed_a(2.6326790248276666e-05)),(to_sfixed_a(0.00011379843635950238)),(to_sfixed_a(0.00017020621453411877)),(to_sfixed_a(6.492524698842317e-05)),(to_sfixed_a(0.00024129828670993447)),(to_sfixed_a(0.00019893386343028396)),(to_sfixed_a(-0.02631177380681038)),(to_sfixed_a(-0.24346792697906494)),(to_sfixed_a(-0.08156460523605347)),(to_sfixed_a(-0.06960797309875488)),(to_sfixed_a(-0.12894946336746216)),(to_sfixed_a(-0.2587544620037079)),(to_sfixed_a(0.09907878935337067)),(to_sfixed_a(0.2581261992454529)),(to_sfixed_a(-0.0801934078335762)),(to_sfixed_a(-0.1712346225976944)),(to_sfixed_a(-0.005986941047012806)),(to_sfixed_a(-0.13312534987926483)),(to_sfixed_a(-0.16679735481739044)),(to_sfixed_a(0.1400398164987564)),(to_sfixed_a(-0.10244570672512054)),(to_sfixed_a(-0.07433643192052841)),(to_sfixed_a(-0.3151029348373413)),(to_sfixed_a(-0.042139291763305664)),(to_sfixed_a(-0.022784002125263214)),(to_sfixed_a(0.05855691060423851)),(to_sfixed_a(-0.05689307674765587)),(to_sfixed_a(-0.016684263944625854)),(to_sfixed_a(0.00011505718430271372)),(to_sfixed_a(0.0001216107266373001)),(to_sfixed_a(0.0001045255339704454)),(to_sfixed_a(-8.628370551377884e-07)),(to_sfixed_a(0.0003040030424017459)),(to_sfixed_a(0.0001740873558446765)),(to_sfixed_a(0.022373734042048454)),(to_sfixed_a(0.0011715881992131472)),(to_sfixed_a(-0.1746080070734024)),(to_sfixed_a(-0.04271088168025017)),(to_sfixed_a(-0.014683462679386139)),(to_sfixed_a(0.015953030437231064)),(to_sfixed_a(0.04414721950888634)),(to_sfixed_a(0.03222300857305527)),(to_sfixed_a(0.2744600772857666)),(to_sfixed_a(0.34210824966430664)),(to_sfixed_a(-0.04684832692146301)),(to_sfixed_a(-0.019809041172266006)),(to_sfixed_a(-0.20435504615306854)),(to_sfixed_a(0.10514184087514877)),(to_sfixed_a(0.04823381081223488)),(to_sfixed_a(0.03687683120369911)),(to_sfixed_a(-0.011831595562398434)),(to_sfixed_a(-0.02908836118876934)),(to_sfixed_a(0.0047159562818706036)),(to_sfixed_a(0.1558796465396881)),(to_sfixed_a(-0.03353143483400345)),(to_sfixed_a(2.2977057597017847e-05)),(to_sfixed_a(-1.8957567590405233e-05)),(to_sfixed_a(-8.817698108032346e-05)),(to_sfixed_a(0.00011933904170291498)),(to_sfixed_a(-0.0001025977690005675)),(to_sfixed_a(-0.00015443425218109041)),(to_sfixed_a(0.00024127648794092238)),(to_sfixed_a(-0.00011372451263014227)),(to_sfixed_a(-0.05856938287615776)),(to_sfixed_a(0.11632875353097916)),(to_sfixed_a(-0.35023850202560425)),(to_sfixed_a(-0.02140149660408497)),(to_sfixed_a(0.040344756096601486)),(to_sfixed_a(0.09557082504034042)),(to_sfixed_a(0.09648086130619049)),(to_sfixed_a(-0.13270887732505798)),(to_sfixed_a(0.5577953457832336)),(to_sfixed_a(0.03758041933178902)),(to_sfixed_a(0.06727302074432373)),(to_sfixed_a(-0.22287382185459137)),(to_sfixed_a(-0.18106165528297424)),(to_sfixed_a(-0.11391285806894302)),(to_sfixed_a(-0.20369145274162292)),(to_sfixed_a(0.05392296239733696)),(to_sfixed_a(0.07351481169462204)),(to_sfixed_a(0.08028221875429153)),(to_sfixed_a(0.12238864600658417)),(to_sfixed_a(-0.06428699195384979)),(to_sfixed_a(-0.08869951218366623)),(to_sfixed_a(6.453705282183364e-05)),(to_sfixed_a(0.00024240960192400962)),(to_sfixed_a(1.8551983885117806e-05)),(to_sfixed_a(0.00022915621229913086)),(to_sfixed_a(0.0002675370196811855)),(to_sfixed_a(-3.999097771156812e-06)),(to_sfixed_a(0.00026557815726846457)),(to_sfixed_a(0.021810289472341537)),(to_sfixed_a(-0.0006101081962697208)),(to_sfixed_a(-0.021545765921473503)),(to_sfixed_a(0.11709344387054443)),(to_sfixed_a(0.019497158005833626)),(to_sfixed_a(0.16432811319828033)),(to_sfixed_a(0.02047029882669449)),(to_sfixed_a(0.13971185684204102)),(to_sfixed_a(0.3867495656013489)),(to_sfixed_a(0.28315964341163635)),(to_sfixed_a(0.5568668842315674)),(to_sfixed_a(0.04057060927152634)),(to_sfixed_a(-0.13276250660419464)),(to_sfixed_a(-0.4872337281703949)),(to_sfixed_a(-0.08561637997627258)),(to_sfixed_a(-0.1375926434993744)),(to_sfixed_a(0.14889968931674957)),(to_sfixed_a(0.06473004817962646)),(to_sfixed_a(-0.07373230159282684)),(to_sfixed_a(-0.00045451975893229246)),(to_sfixed_a(0.07685015350580215)),(to_sfixed_a(-0.00020464749832171947)),(to_sfixed_a(-6.30038557574153e-05)),(to_sfixed_a(1.0089073839480989e-05)),(to_sfixed_a(-0.00011063212878070772)),(to_sfixed_a(-4.772425654664403e-06)),(to_sfixed_a(9.109059465117753e-05)),(to_sfixed_a(6.948621830815682e-06)),(to_sfixed_a(0.0002807371492963284)),(to_sfixed_a(-0.030469922348856926)),(to_sfixed_a(-0.015446358360350132)),(to_sfixed_a(-0.07775571197271347)),(to_sfixed_a(-0.017325207591056824)),(to_sfixed_a(0.07348459213972092)),(to_sfixed_a(0.2110881805419922)),(to_sfixed_a(0.01268912572413683)),(to_sfixed_a(0.1403743475675583)),(to_sfixed_a(0.1224861890077591)),(to_sfixed_a(0.06487976014614105)),(to_sfixed_a(-0.0928497165441513)),(to_sfixed_a(-0.0038204779848456383)),(to_sfixed_a(-0.09041616320610046)),(to_sfixed_a(-0.41784054040908813)),(to_sfixed_a(-0.08393657952547073)),(to_sfixed_a(0.10607387870550156)),(to_sfixed_a(0.014431439340114594)),(to_sfixed_a(0.08078774809837341)),(to_sfixed_a(0.0001047556652338244)),(to_sfixed_a(-9.094947017729282e-05)),(to_sfixed_a(4.410795008880086e-05)),(to_sfixed_a(0.0001144525595009327)),(to_sfixed_a(-0.00027608650270849466)),(to_sfixed_a(3.6493827792583033e-05)),(to_sfixed_a(-0.00025637002545408905)),(to_sfixed_a(0.00018886695033870637)),(to_sfixed_a(-3.875211041304283e-05)),(to_sfixed_a(0.00034971427521668375)),(to_sfixed_a(-0.00871448777616024)),(to_sfixed_a(0.14147591590881348)),(to_sfixed_a(0.1049787625670433)),(to_sfixed_a(0.16835801303386688)),(to_sfixed_a(-0.0358387790620327)),(to_sfixed_a(0.07225659489631653)),(to_sfixed_a(0.0351504310965538)),(to_sfixed_a(0.019446907564997673)),(to_sfixed_a(0.033386681228876114)),(to_sfixed_a(-0.10750021785497665)),(to_sfixed_a(-0.24935971200466156)),(to_sfixed_a(-0.3181408643722534)),(to_sfixed_a(-0.1885640174150467)),(to_sfixed_a(0.18568067252635956)),(to_sfixed_a(0.11829642206430435)),(to_sfixed_a(-0.04696933552622795)),(to_sfixed_a(-0.04256577044725418)),(to_sfixed_a(-0.0014124090084806085)),(to_sfixed_a(-0.02970566228032112)),(to_sfixed_a(0.0001510953006800264)),(to_sfixed_a(-0.0002526077441871166)),(to_sfixed_a(-0.00019784030155278742)),(to_sfixed_a(-1.0196999937761575e-05)),(to_sfixed_a(1.1509527212183457e-05)),(to_sfixed_a(7.377001020358875e-05)),(to_sfixed_a(0.00010621608089422807)),(to_sfixed_a(0.0003065505006816238)),(to_sfixed_a(0.0409223847091198)),(to_sfixed_a(0.04161253198981285)),(to_sfixed_a(0.1711123287677765)),(to_sfixed_a(0.21899035573005676)),(to_sfixed_a(0.12420684099197388)),(to_sfixed_a(0.0005329055129550397)),(to_sfixed_a(-0.16805097460746765)),(to_sfixed_a(0.026299117133021355)),(to_sfixed_a(0.3600512742996216)),(to_sfixed_a(-0.12018606066703796)),(to_sfixed_a(-0.024363379925489426)),(to_sfixed_a(-0.12177571654319763)),(to_sfixed_a(0.0032665159087628126)),(to_sfixed_a(-0.05657036229968071)),(to_sfixed_a(-0.068828284740448)),(to_sfixed_a(-0.1582849621772766)),(to_sfixed_a(-0.010549749247729778)),(to_sfixed_a(-0.03840145468711853)),(to_sfixed_a(-0.01796114444732666)),(to_sfixed_a(0.00047071289736777544)),(to_sfixed_a(-0.00019264071306679398)),(to_sfixed_a(2.2634552806266584e-05)),(to_sfixed_a(-0.00011245912901358679)),(to_sfixed_a(-0.00022081124188844115)),(to_sfixed_a(-0.0001589888270245865)),(to_sfixed_a(0.0002345326211070642)),(to_sfixed_a(0.00016315326502081007)),(to_sfixed_a(0.00035618102992884815)),(to_sfixed_a(-5.523225263459608e-05)),(to_sfixed_a(0.0979580357670784)),(to_sfixed_a(0.1029713973402977)),(to_sfixed_a(0.11845555901527405)),(to_sfixed_a(0.451373428106308)),(to_sfixed_a(-0.0002407534484518692)),(to_sfixed_a(0.15196895599365234)),(to_sfixed_a(-0.0026596563402563334)),(to_sfixed_a(-0.1952301561832428)),(to_sfixed_a(-0.06454235315322876)),(to_sfixed_a(0.16518744826316833)),(to_sfixed_a(0.18358302116394043)),(to_sfixed_a(-0.08686354011297226)),(to_sfixed_a(-0.03720966726541519)),(to_sfixed_a(-0.010293272323906422)),(to_sfixed_a(-0.1074720174074173)),(to_sfixed_a(-0.08107996731996536)),(to_sfixed_a(-5.094124935567379e-05)),(to_sfixed_a(0.0009765035938471556)),(to_sfixed_a(0.0015186492819339037)),(to_sfixed_a(-1.660968700889498e-05)),(to_sfixed_a(-4.062327207066119e-05)),(to_sfixed_a(4.6648601710330695e-05)),(to_sfixed_a(-0.0001598750241100788)),(to_sfixed_a(-9.925026097334921e-05)),(to_sfixed_a(0.00018257532792631537)),(to_sfixed_a(0.00013794464757665992)),(to_sfixed_a(-0.00022458888997789472)),(to_sfixed_a(3.844469756586477e-05)),(to_sfixed_a(-0.0009055154514499009)),(to_sfixed_a(-0.0010507910046726465)),(to_sfixed_a(-0.00012523698387667537)),(to_sfixed_a(-0.00015071494271978736)),(to_sfixed_a(0.0004053952870890498)),(to_sfixed_a(-0.08338742703199387)),(to_sfixed_a(-0.002980040153488517)),(to_sfixed_a(-0.000255352322710678)),(to_sfixed_a(-0.06575381010770798)),(to_sfixed_a(-0.0021542729809880257)),(to_sfixed_a(0.011150140315294266)),(to_sfixed_a(-0.01566474884748459)),(to_sfixed_a(-0.0642942264676094)),(to_sfixed_a(-0.09082547575235367)),(to_sfixed_a(-0.008083444088697433)),(to_sfixed_a(-0.0038494677282869816)),(to_sfixed_a(-0.0002448185405228287)),(to_sfixed_a(-0.00019444370991550386)),(to_sfixed_a(-1.9159044313710183e-05)),(to_sfixed_a(-2.7246811441727914e-05)),(to_sfixed_a(-9.806089656194672e-05)),(to_sfixed_a(-1.2000129572697915e-05)),(to_sfixed_a(0.00023316867009270936)),(to_sfixed_a(0.00012126742512919009)),(to_sfixed_a(-7.040468335617334e-05)),(to_sfixed_a(3.7907364003331168e-06)),(to_sfixed_a(4.474437082535587e-05)),(to_sfixed_a(4.7167199227260426e-05)),(to_sfixed_a(0.00023184233577921987)),(to_sfixed_a(-1.8100916349794716e-05)),(to_sfixed_a(0.0001397517480654642)),(to_sfixed_a(-1.6830586901050992e-05)),(to_sfixed_a(-0.00014571574865840375)),(to_sfixed_a(-1.7311762348981574e-05)),(to_sfixed_a(-0.00014178818673826754)),(to_sfixed_a(0.0001353387488052249)),(to_sfixed_a(-1.3384054000198375e-05)),(to_sfixed_a(0.00024141668109223247)),(to_sfixed_a(-0.00031681088148616254)),(to_sfixed_a(0.0001822404592530802)),(to_sfixed_a(0.00012662564404308796)),(to_sfixed_a(4.78399197163526e-05)),(to_sfixed_a(-1.3466607924783602e-05)),(to_sfixed_a(-3.921389361494221e-05)),(to_sfixed_a(-7.963907410157844e-05)),(to_sfixed_a(-2.5183857360389084e-05)),(to_sfixed_a(6.783738353988156e-05)),(to_sfixed_a(4.74667212984059e-05)),(to_sfixed_a(3.1194573239190504e-05)),(to_sfixed_a(-0.0003191028372384608)),(to_sfixed_a(0.00015730343875475228)));

    constant weight_n0_21 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(0.00025928555987775326)),(to_sfixed_a(-5.9552068705670536e-05)),(to_sfixed_a(5.475727448356338e-05)),(to_sfixed_a(-0.0002624854096211493)),(to_sfixed_a(-0.0002966233005281538)),(to_sfixed_a(-1.625890399736818e-05)),(to_sfixed_a(-0.0003513609990477562)),(to_sfixed_a(5.8003617596114054e-05)),(to_sfixed_a(-1.232818431162741e-05)),(to_sfixed_a(-0.00025538037880323827)),(to_sfixed_a(4.585003625834361e-05)),(to_sfixed_a(2.0590467102010734e-05)),(to_sfixed_a(-1.167254686151864e-05)),(to_sfixed_a(1.7850908989203162e-05)),(to_sfixed_a(-0.00014482776168733835)),(to_sfixed_a(3.0396279271371895e-06)),(to_sfixed_a(-0.00026891898596659303)),(to_sfixed_a(-7.173296762630343e-05)),(to_sfixed_a(0.00028819876024499536)),(to_sfixed_a(-3.361056587891653e-05)),(to_sfixed_a(-2.6888959837378934e-05)),(to_sfixed_a(-0.00025048726820386946)),(to_sfixed_a(-6.353530625347048e-05)),(to_sfixed_a(2.7856736778630875e-05)),(to_sfixed_a(-0.000114569062134251)),(to_sfixed_a(-0.00029198164702393115)),(to_sfixed_a(-0.00023259797308128327)),(to_sfixed_a(0.00013183290138840675)),(to_sfixed_a(-0.0001265766186406836)),(to_sfixed_a(4.3526553781703115e-05)),(to_sfixed_a(1.4857048881822266e-05)),(to_sfixed_a(-1.1033997907361481e-05)),(to_sfixed_a(4.8640122258802876e-05)),(to_sfixed_a(0.00012800453987438232)),(to_sfixed_a(2.7438491088105366e-05)),(to_sfixed_a(-0.000275070546194911)),(to_sfixed_a(2.115361439791741e-06)),(to_sfixed_a(5.8539753808872774e-05)),(to_sfixed_a(0.00018492339586373419)),(to_sfixed_a(7.736066618235782e-05)),(to_sfixed_a(0.0001230919879162684)),(to_sfixed_a(0.0001313749235123396)),(to_sfixed_a(0.00013220368418842554)),(to_sfixed_a(-0.00014470412861555815)),(to_sfixed_a(-0.00010458287579240277)),(to_sfixed_a(4.4489872379926965e-05)),(to_sfixed_a(-0.00017080656834878027)),(to_sfixed_a(-0.00017172691877931356)),(to_sfixed_a(5.728470569010824e-05)),(to_sfixed_a(9.957594011211768e-05)),(to_sfixed_a(0.00022403769253287464)),(to_sfixed_a(0.0003034053079318255)),(to_sfixed_a(-0.00027392670745030046)),(to_sfixed_a(0.00015548645751550794)),(to_sfixed_a(6.75896808388643e-05)),(to_sfixed_a(-7.012751302681863e-05)),(to_sfixed_a(0.00022279616678133607)),(to_sfixed_a(-7.529290451202542e-05)),(to_sfixed_a(-8.347051334567368e-06)),(to_sfixed_a(4.902047658106312e-05)),(to_sfixed_a(-0.00038903558743186295)),(to_sfixed_a(-0.00013204218703322113)),(to_sfixed_a(-5.439612505142577e-05)),(to_sfixed_a(5.997886546538211e-06)),(to_sfixed_a(-7.189375173766166e-05)),(to_sfixed_a(-0.00021033620578236878)),(to_sfixed_a(9.143250645138323e-05)),(to_sfixed_a(0.00010250125342281535)),(to_sfixed_a(2.854238118743524e-05)),(to_sfixed_a(-0.01625903882086277)),(to_sfixed_a(-6.070026574889198e-05)),(to_sfixed_a(5.0903639930766076e-05)),(to_sfixed_a(-0.0002493398205842823)),(to_sfixed_a(1.1712982995959464e-05)),(to_sfixed_a(4.2551226215437055e-05)),(to_sfixed_a(0.0003005194303113967)),(to_sfixed_a(6.72742971801199e-05)),(to_sfixed_a(0.00026304140919819474)),(to_sfixed_a(7.712216029176489e-05)),(to_sfixed_a(0.00017927275621332228)),(to_sfixed_a(0.0001494802418164909)),(to_sfixed_a(-3.285918865003623e-05)),(to_sfixed_a(4.5621451135957614e-05)),(to_sfixed_a(-5.959076588624157e-05)),(to_sfixed_a(-0.0001868056715466082)),(to_sfixed_a(-6.471871165558696e-05)),(to_sfixed_a(0.00010050038690678775)),(to_sfixed_a(-0.00010981466039083898)),(to_sfixed_a(3.216482946299948e-05)),(to_sfixed_a(-0.00013161961396690458)),(to_sfixed_a(-9.924684127327055e-05)),(to_sfixed_a(-0.00010946505062747747)),(to_sfixed_a(-0.004740920849144459)),(to_sfixed_a(-4.771841486217454e-05)),(to_sfixed_a(-0.005492247175425291)),(to_sfixed_a(0.020746929571032524)),(to_sfixed_a(-0.05264810845255852)),(to_sfixed_a(-0.07333434373140335)),(to_sfixed_a(-0.04802880808711052)),(to_sfixed_a(-0.12109837681055069)),(to_sfixed_a(-0.0384988859295845)),(to_sfixed_a(-0.23649904131889343)),(to_sfixed_a(0.03972470387816429)),(to_sfixed_a(0.05590447783470154)),(to_sfixed_a(0.049318987876176834)),(to_sfixed_a(0.09991946071386337)),(to_sfixed_a(4.6691431634826586e-05)),(to_sfixed_a(3.2159154216060415e-05)),(to_sfixed_a(-0.00017095392104238272)),(to_sfixed_a(8.836082997731864e-05)),(to_sfixed_a(-7.967578881107329e-07)),(to_sfixed_a(8.358016930287704e-05)),(to_sfixed_a(0.0001083448514691554)),(to_sfixed_a(7.636059308424592e-05)),(to_sfixed_a(-6.81239616824314e-05)),(to_sfixed_a(6.902373570483178e-05)),(to_sfixed_a(0.0001107780117308721)),(to_sfixed_a(3.150324846501462e-05)),(to_sfixed_a(-0.0002632064279168844)),(to_sfixed_a(0.014848168939352036)),(to_sfixed_a(0.047400496900081635)),(to_sfixed_a(-0.011213457211852074)),(to_sfixed_a(-0.00459044286981225)),(to_sfixed_a(0.0645870566368103)),(to_sfixed_a(0.12238168716430664)),(to_sfixed_a(0.33813589811325073)),(to_sfixed_a(-0.04110218957066536)),(to_sfixed_a(-0.14745384454727173)),(to_sfixed_a(-0.1967514604330063)),(to_sfixed_a(-0.312728613615036)),(to_sfixed_a(-0.1370757669210434)),(to_sfixed_a(0.02402648702263832)),(to_sfixed_a(0.0012464983155950904)),(to_sfixed_a(0.15355801582336426)),(to_sfixed_a(0.0012744656996801496)),(to_sfixed_a(-0.0003506129141896963)),(to_sfixed_a(0.0024253397714346647)),(to_sfixed_a(1.2298050023673568e-05)),(to_sfixed_a(0.00015778926899656653)),(to_sfixed_a(9.053573739947751e-05)),(to_sfixed_a(-0.00015739047375973314)),(to_sfixed_a(0.00012833750224672258)),(to_sfixed_a(-0.0002506136952433735)),(to_sfixed_a(7.963941607158631e-05)),(to_sfixed_a(-0.0008217424619942904)),(to_sfixed_a(0.04282037541270256)),(to_sfixed_a(0.015379605814814568)),(to_sfixed_a(0.04744705557823181)),(to_sfixed_a(0.017306741327047348)),(to_sfixed_a(0.048294611275196075)),(to_sfixed_a(0.11953724920749664)),(to_sfixed_a(-0.018237201496958733)),(to_sfixed_a(-0.052163124084472656)),(to_sfixed_a(-0.09157314896583557)),(to_sfixed_a(-0.0037398517597466707)),(to_sfixed_a(-0.018201692029833794)),(to_sfixed_a(-0.07537280768156052)),(to_sfixed_a(-0.2648015320301056)),(to_sfixed_a(-0.5679922699928284)),(to_sfixed_a(-0.144174262881279)),(to_sfixed_a(-0.05514451488852501)),(to_sfixed_a(0.03455618396401405)),(to_sfixed_a(0.00019783992320299149)),(to_sfixed_a(0.08609548211097717)),(to_sfixed_a(0.0030602412298321724)),(to_sfixed_a(-0.00020108158059883863)),(to_sfixed_a(-0.0002727456740103662)),(to_sfixed_a(0.0002763878437690437)),(to_sfixed_a(0.0001018689144984819)),(to_sfixed_a(0.00011057090159738436)),(to_sfixed_a(-0.00012245056859683245)),(to_sfixed_a(-1.920039494507364e-06)),(to_sfixed_a(-0.00024278908676933497)),(to_sfixed_a(0.03702200949192047)),(to_sfixed_a(0.03016366995871067)),(to_sfixed_a(0.11837593466043472)),(to_sfixed_a(0.08590561151504517)),(to_sfixed_a(-0.19312940537929535)),(to_sfixed_a(0.10564280301332474)),(to_sfixed_a(0.17102332413196564)),(to_sfixed_a(-0.023444637656211853)),(to_sfixed_a(-0.11544600874185562)),(to_sfixed_a(-0.3791291415691376)),(to_sfixed_a(-0.3545615077018738)),(to_sfixed_a(-0.21426862478256226)),(to_sfixed_a(-0.13164447247982025)),(to_sfixed_a(0.16018731892108917)),(to_sfixed_a(-0.2837485671043396)),(to_sfixed_a(0.010194987989962101)),(to_sfixed_a(0.08601147681474686)),(to_sfixed_a(0.16690096259117126)),(to_sfixed_a(0.09970343112945557)),(to_sfixed_a(-0.002888140268623829)),(to_sfixed_a(-0.0035947442520409822)),(to_sfixed_a(-0.0020992399659007788)),(to_sfixed_a(-0.00014182005543261766)),(to_sfixed_a(8.469433669233695e-05)),(to_sfixed_a(-0.0001640360860619694)),(to_sfixed_a(-0.00027946149930357933)),(to_sfixed_a(-5.2818220865447074e-05)),(to_sfixed_a(-0.00022544067178387195)),(to_sfixed_a(0.013708135113120079)),(to_sfixed_a(0.057330142706632614)),(to_sfixed_a(-0.17497044801712036)),(to_sfixed_a(-0.29492172598838806)),(to_sfixed_a(-0.25119972229003906)),(to_sfixed_a(-0.050311263650655746)),(to_sfixed_a(-0.08919188380241394)),(to_sfixed_a(-0.05673670396208763)),(to_sfixed_a(-0.254330575466156)),(to_sfixed_a(-0.011497417464852333)),(to_sfixed_a(0.08988818526268005)),(to_sfixed_a(-0.20401132106781006)),(to_sfixed_a(0.22996920347213745)),(to_sfixed_a(-0.24420420825481415)),(to_sfixed_a(0.023053186014294624)),(to_sfixed_a(0.03821799159049988)),(to_sfixed_a(-0.22266073524951935)),(to_sfixed_a(0.04830234497785568)),(to_sfixed_a(0.10067880898714066)),(to_sfixed_a(-0.022621655836701393)),(to_sfixed_a(0.00500843208283186)),(to_sfixed_a(1.4717116755491588e-05)),(to_sfixed_a(0.00022148151765577495)),(to_sfixed_a(-1.5695750334998593e-05)),(to_sfixed_a(5.824863819725579e-06)),(to_sfixed_a(6.42477025394328e-05)),(to_sfixed_a(0.0001969681034097448)),(to_sfixed_a(0.05608171969652176)),(to_sfixed_a(0.09889239072799683)),(to_sfixed_a(-0.0006701114471070468)),(to_sfixed_a(0.19932833313941956)),(to_sfixed_a(-0.5035852789878845)),(to_sfixed_a(0.11318990588188171)),(to_sfixed_a(-0.09491558372974396)),(to_sfixed_a(-0.023271556943655014)),(to_sfixed_a(-0.02690996415913105)),(to_sfixed_a(-0.13689777255058289)),(to_sfixed_a(-0.054512858390808105)),(to_sfixed_a(0.05402924492955208)),(to_sfixed_a(-0.03757702186703682)),(to_sfixed_a(0.17064355313777924)),(to_sfixed_a(-0.05031612887978554)),(to_sfixed_a(-0.3706546723842621)),(to_sfixed_a(0.018359586596488953)),(to_sfixed_a(0.03640052303671837)),(to_sfixed_a(-0.06700880825519562)),(to_sfixed_a(-0.021643539890646935)),(to_sfixed_a(0.15285944938659668)),(to_sfixed_a(-0.010365213267505169)),(to_sfixed_a(-8.309072291012853e-05)),(to_sfixed_a(0.00015813398931641132)),(to_sfixed_a(-0.00017734307039063424)),(to_sfixed_a(0.0003033879038412124)),(to_sfixed_a(-8.897289080778137e-05)),(to_sfixed_a(-0.00010486614337423816)),(to_sfixed_a(0.0005869943997822702)),(to_sfixed_a(0.06628266721963882)),(to_sfixed_a(0.024185005575418472)),(to_sfixed_a(-0.42093178629875183)),(to_sfixed_a(0.007216583006083965)),(to_sfixed_a(0.04973834753036499)),(to_sfixed_a(-0.3226125240325928)),(to_sfixed_a(-0.10312707722187042)),(to_sfixed_a(-0.24898287653923035)),(to_sfixed_a(-0.17488929629325867)),(to_sfixed_a(0.34962934255599976)),(to_sfixed_a(0.3649357855319977)),(to_sfixed_a(0.5031697750091553)),(to_sfixed_a(0.4919888973236084)),(to_sfixed_a(-0.012303302995860577)),(to_sfixed_a(-0.33566105365753174)),(to_sfixed_a(-0.4075891077518463)),(to_sfixed_a(-0.19141386449337006)),(to_sfixed_a(-0.0712873786687851)),(to_sfixed_a(-0.16543272137641907)),(to_sfixed_a(0.21259988844394684)),(to_sfixed_a(3.0676910682814196e-06)),(to_sfixed_a(3.246022606617771e-05)),(to_sfixed_a(9.146705451712478e-06)),(to_sfixed_a(-2.5045232177944854e-05)),(to_sfixed_a(-0.0001385981304338202)),(to_sfixed_a(-0.0003371489292476326)),(to_sfixed_a(-0.000142062664963305)),(to_sfixed_a(-0.010757866315543652)),(to_sfixed_a(0.0047709401696920395)),(to_sfixed_a(-0.16160418093204498)),(to_sfixed_a(-0.03537489101290703)),(to_sfixed_a(-0.055710483342409134)),(to_sfixed_a(0.16792574524879456)),(to_sfixed_a(0.06855892390012741)),(to_sfixed_a(0.0936473086476326)),(to_sfixed_a(-0.07665478438138962)),(to_sfixed_a(-0.21958692371845245)),(to_sfixed_a(-0.2796209454536438)),(to_sfixed_a(-0.034203872084617615)),(to_sfixed_a(0.04068446904420853)),(to_sfixed_a(0.3710005581378937)),(to_sfixed_a(-0.07259123772382736)),(to_sfixed_a(-0.05322062969207764)),(to_sfixed_a(-0.21205295622348785)),(to_sfixed_a(-0.2525855004787445)),(to_sfixed_a(-0.23417797684669495)),(to_sfixed_a(-0.2014458030462265)),(to_sfixed_a(0.13862253725528717)),(to_sfixed_a(0.09980859607458115)),(to_sfixed_a(-1.480416722188238e-05)),(to_sfixed_a(-0.00016361012239940464)),(to_sfixed_a(0.000228515564231202)),(to_sfixed_a(-0.00019331061048433185)),(to_sfixed_a(1.6329388017766178e-05)),(to_sfixed_a(-0.02318771928548813)),(to_sfixed_a(0.08932403475046158)),(to_sfixed_a(-0.057342808693647385)),(to_sfixed_a(-0.03242816776037216)),(to_sfixed_a(-0.058130085468292236)),(to_sfixed_a(-0.00399004016071558)),(to_sfixed_a(0.007494933437556028)),(to_sfixed_a(0.02002035267651081)),(to_sfixed_a(-0.14674223959445953)),(to_sfixed_a(-0.061974216252565384)),(to_sfixed_a(0.13391482830047607)),(to_sfixed_a(0.1399969905614853)),(to_sfixed_a(-0.15906326472759247)),(to_sfixed_a(-0.0380549281835556)),(to_sfixed_a(-0.0796322450041771)),(to_sfixed_a(0.14356033504009247)),(to_sfixed_a(0.011743471957743168)),(to_sfixed_a(0.05331237241625786)),(to_sfixed_a(-0.09304972738027573)),(to_sfixed_a(0.025771083310246468)),(to_sfixed_a(-0.23077192902565002)),(to_sfixed_a(-0.09031244367361069)),(to_sfixed_a(6.8264314904809e-05)),(to_sfixed_a(-3.6454959627008066e-05)),(to_sfixed_a(0.00021599698811769485)),(to_sfixed_a(-1.8203963918494992e-05)),(to_sfixed_a(-0.00012145782238803804)),(to_sfixed_a(0.00010545150144025683)),(to_sfixed_a(0.00013911457790527493)),(to_sfixed_a(0.054781295359134674)),(to_sfixed_a(-0.023907221853733063)),(to_sfixed_a(-0.004333888180553913)),(to_sfixed_a(0.08961702883243561)),(to_sfixed_a(0.07422558963298798)),(to_sfixed_a(0.0012181397760286927)),(to_sfixed_a(0.04184086248278618)),(to_sfixed_a(0.04921971261501312)),(to_sfixed_a(0.015322697348892689)),(to_sfixed_a(0.014598746784031391)),(to_sfixed_a(-0.15135090053081512)),(to_sfixed_a(-0.22825512290000916)),(to_sfixed_a(-0.4510616064071655)),(to_sfixed_a(-0.007338681258261204)),(to_sfixed_a(0.1523909568786621)),(to_sfixed_a(0.018882090225815773)),(to_sfixed_a(0.21669520437717438)),(to_sfixed_a(0.06852854043245316)),(to_sfixed_a(0.1376100778579712)),(to_sfixed_a(0.11676635593175888)),(to_sfixed_a(0.27973732352256775)),(to_sfixed_a(0.00014847578131593764)),(to_sfixed_a(0.0001472662843298167)),(to_sfixed_a(4.2511470383033156e-05)),(to_sfixed_a(7.641417323611677e-05)),(to_sfixed_a(0.000403240614105016)),(to_sfixed_a(-0.00010904553346335888)),(to_sfixed_a(6.090052556828596e-05)),(to_sfixed_a(0.015914320945739746)),(to_sfixed_a(-0.021115010604262352)),(to_sfixed_a(-0.002310573821887374)),(to_sfixed_a(0.10512273013591766)),(to_sfixed_a(0.069325752556324)),(to_sfixed_a(0.13206060230731964)),(to_sfixed_a(-0.026432253420352936)),(to_sfixed_a(-0.002352170879021287)),(to_sfixed_a(0.06769653409719467)),(to_sfixed_a(0.046482060104608536)),(to_sfixed_a(-0.04608961194753647)),(to_sfixed_a(-0.15319857001304626)),(to_sfixed_a(-0.10428662598133087)),(to_sfixed_a(0.03097306564450264)),(to_sfixed_a(-0.07670240849256516)),(to_sfixed_a(0.25524330139160156)),(to_sfixed_a(0.07001887261867523)),(to_sfixed_a(0.15133731067180634)),(to_sfixed_a(-0.11343078315258026)),(to_sfixed_a(0.3177182078361511)),(to_sfixed_a(-0.011401359923183918)),(to_sfixed_a(-0.0049027022905647755)),(to_sfixed_a(-0.006464232224971056)),(to_sfixed_a(0.00030511413933709264)),(to_sfixed_a(-0.0002489588223397732)),(to_sfixed_a(-9.374361980007961e-05)),(to_sfixed_a(-3.4210781450383365e-05)),(to_sfixed_a(-4.3199092033319175e-05)),(to_sfixed_a(0.0010573853505775332)),(to_sfixed_a(0.011993122287094593)),(to_sfixed_a(-0.05595504119992256)),(to_sfixed_a(-0.14473144710063934)),(to_sfixed_a(0.07286503911018372)),(to_sfixed_a(0.020053930580615997)),(to_sfixed_a(0.08051274716854095)),(to_sfixed_a(-0.25528407096862793)),(to_sfixed_a(0.03908450901508331)),(to_sfixed_a(-0.09276099503040314)),(to_sfixed_a(0.2726605236530304)),(to_sfixed_a(-0.056530315428972244)),(to_sfixed_a(0.0828884169459343)),(to_sfixed_a(0.16568569839000702)),(to_sfixed_a(-0.07243119180202484)),(to_sfixed_a(-0.04651764780282974)),(to_sfixed_a(0.18979506194591522)),(to_sfixed_a(-0.07458440959453583)),(to_sfixed_a(0.04667448624968529)),(to_sfixed_a(-0.28194037079811096)),(to_sfixed_a(-0.0057602240704)),(to_sfixed_a(-0.0007080165087245405)),(to_sfixed_a(-0.00040961994091048837)),(to_sfixed_a(2.6099149181391113e-05)),(to_sfixed_a(7.183009438449517e-05)),(to_sfixed_a(5.7519344409229234e-05)),(to_sfixed_a(-0.00019936379976570606)),(to_sfixed_a(0.00010701821156544611)),(to_sfixed_a(0.04336414486169815)),(to_sfixed_a(-0.11653456091880798)),(to_sfixed_a(-0.1043611466884613)),(to_sfixed_a(-0.10613272339105606)),(to_sfixed_a(0.008541435934603214)),(to_sfixed_a(-0.10703528672456741)),(to_sfixed_a(0.22175872325897217)),(to_sfixed_a(-0.019579140469431877)),(to_sfixed_a(0.026703177019953728)),(to_sfixed_a(0.5599189400672913)),(to_sfixed_a(0.17482547461986542)),(to_sfixed_a(-0.04910438880324364)),(to_sfixed_a(0.001432823366485536)),(to_sfixed_a(0.0001261216530110687)),(to_sfixed_a(-0.06668388843536377)),(to_sfixed_a(0.07674332708120346)),(to_sfixed_a(-0.5904951691627502)),(to_sfixed_a(-0.041142530739307404)),(to_sfixed_a(-0.045699216425418854)),(to_sfixed_a(-0.042439766228199005)),(to_sfixed_a(-0.16427429020404816)),(to_sfixed_a(-0.0008091286290436983)),(to_sfixed_a(0.00010448820830788463)),(to_sfixed_a(7.715426181675866e-05)),(to_sfixed_a(-7.381082104984671e-05)),(to_sfixed_a(0.00013411804684437811)),(to_sfixed_a(-0.0002476725494489074)),(to_sfixed_a(-8.315374725498259e-05)),(to_sfixed_a(-0.04873171076178551)),(to_sfixed_a(-0.10110625624656677)),(to_sfixed_a(-0.14630462229251862)),(to_sfixed_a(-0.004755463916808367)),(to_sfixed_a(0.05160599574446678)),(to_sfixed_a(0.18158480525016785)),(to_sfixed_a(0.18054215610027313)),(to_sfixed_a(-0.15061607956886292)),(to_sfixed_a(0.08312070369720459)),(to_sfixed_a(-0.11313369870185852)),(to_sfixed_a(-0.13870228826999664)),(to_sfixed_a(-0.08362846821546555)),(to_sfixed_a(0.16934214532375336)),(to_sfixed_a(0.028521688655018806)),(to_sfixed_a(0.035528384149074554)),(to_sfixed_a(-0.12097427994012833)),(to_sfixed_a(-0.344373881816864)),(to_sfixed_a(-0.2750609815120697)),(to_sfixed_a(-0.07201551645994186)),(to_sfixed_a(0.0569738894701004)),(to_sfixed_a(-0.048147182911634445)),(to_sfixed_a(0.015397918410599232)),(to_sfixed_a(3.7682082620449364e-05)),(to_sfixed_a(1.3357497664401308e-05)),(to_sfixed_a(3.695025225169957e-05)),(to_sfixed_a(5.662448165821843e-05)),(to_sfixed_a(-0.0009257636265829206)),(to_sfixed_a(-0.0002699917822610587)),(to_sfixed_a(0.013420617207884789)),(to_sfixed_a(-0.10755418986082077)),(to_sfixed_a(0.028293361887335777)),(to_sfixed_a(0.10730896145105362)),(to_sfixed_a(0.2717908024787903)),(to_sfixed_a(0.0809880942106247)),(to_sfixed_a(0.0861823782324791)),(to_sfixed_a(-0.15908923745155334)),(to_sfixed_a(-0.24880726635456085)),(to_sfixed_a(0.12905386090278625)),(to_sfixed_a(-2.9584558433271013e-05)),(to_sfixed_a(0.021218592301011086)),(to_sfixed_a(0.1208379715681076)),(to_sfixed_a(0.14554822444915771)),(to_sfixed_a(-0.010839846916496754)),(to_sfixed_a(-0.00932400394231081)),(to_sfixed_a(-0.018097491934895515)),(to_sfixed_a(0.05644354224205017)),(to_sfixed_a(-0.2604585289955139)),(to_sfixed_a(-0.04975027218461037)),(to_sfixed_a(-3.82621919925441e-06)),(to_sfixed_a(-0.00015673066081944853)),(to_sfixed_a(-0.0002708645770326257)),(to_sfixed_a(0.0002767164842225611)),(to_sfixed_a(-8.338595216628164e-05)),(to_sfixed_a(0.00018861578428186476)),(to_sfixed_a(1.3751178812526632e-05)),(to_sfixed_a(0.012958605773746967)),(to_sfixed_a(-0.13303618133068085)),(to_sfixed_a(0.04673122987151146)),(to_sfixed_a(0.18980242311954498)),(to_sfixed_a(-0.04289611801505089)),(to_sfixed_a(0.17880207300186157)),(to_sfixed_a(0.056504663079977036)),(to_sfixed_a(0.003132391255348921)),(to_sfixed_a(-0.008388284593820572)),(to_sfixed_a(-0.3260388970375061)),(to_sfixed_a(0.12883919477462769)),(to_sfixed_a(-0.13131728768348694)),(to_sfixed_a(0.10279985517263412)),(to_sfixed_a(0.011951022781431675)),(to_sfixed_a(0.11410005390644073)),(to_sfixed_a(-0.011077096685767174)),(to_sfixed_a(0.04590088129043579)),(to_sfixed_a(-0.03384442254900932)),(to_sfixed_a(-0.1312377154827118)),(to_sfixed_a(-0.027051683515310287)),(to_sfixed_a(-0.003833228722214699)),(to_sfixed_a(0.029569145292043686)),(to_sfixed_a(-1.294423418585211e-05)),(to_sfixed_a(-0.0003330152540002018)),(to_sfixed_a(-2.198950642195996e-05)),(to_sfixed_a(-0.00013313782983459532)),(to_sfixed_a(1.9988972780993208e-05)),(to_sfixed_a(7.762737368466333e-05)),(to_sfixed_a(0.010589977726340294)),(to_sfixed_a(-0.002121192403137684)),(to_sfixed_a(-0.053897809237241745)),(to_sfixed_a(0.06268282234668732)),(to_sfixed_a(0.1936526596546173)),(to_sfixed_a(0.04113848879933357)),(to_sfixed_a(0.2833409011363983)),(to_sfixed_a(0.14103083312511444)),(to_sfixed_a(-0.1158403605222702)),(to_sfixed_a(-0.41905128955841064)),(to_sfixed_a(-0.10548026114702225)),(to_sfixed_a(-0.03406346216797829)),(to_sfixed_a(-0.2152481973171234)),(to_sfixed_a(0.15578851103782654)),(to_sfixed_a(0.3428555727005005)),(to_sfixed_a(0.005046642851084471)),(to_sfixed_a(-0.08015602827072144)),(to_sfixed_a(-0.04581378027796745)),(to_sfixed_a(0.06825253367424011)),(to_sfixed_a(-0.037287648767232895)),(to_sfixed_a(0.03697354346513748)),(to_sfixed_a(-0.00013763979950454086)),(to_sfixed_a(0.00021411065245047212)),(to_sfixed_a(-3.4505519579397514e-05)),(to_sfixed_a(-0.0002182258467655629)),(to_sfixed_a(0.00029095844365656376)),(to_sfixed_a(6.62562160869129e-05)),(to_sfixed_a(0.00011969717888860032)),(to_sfixed_a(-7.900640775915235e-05)),(to_sfixed_a(-0.012929445132613182)),(to_sfixed_a(0.1844288408756256)),(to_sfixed_a(0.04158915579319)),(to_sfixed_a(0.26462647318840027)),(to_sfixed_a(0.21475735306739807)),(to_sfixed_a(0.15146154165267944)),(to_sfixed_a(0.01465977169573307)),(to_sfixed_a(-0.1662999838590622)),(to_sfixed_a(-0.22640961408615112)),(to_sfixed_a(-0.009881172329187393)),(to_sfixed_a(0.001369866426102817)),(to_sfixed_a(0.23769861459732056)),(to_sfixed_a(0.3923771381378174)),(to_sfixed_a(0.074399933218956)),(to_sfixed_a(0.25577419996261597)),(to_sfixed_a(0.18017421662807465)),(to_sfixed_a(0.014910561963915825)),(to_sfixed_a(-0.057492695748806)),(to_sfixed_a(-0.05071872100234032)),(to_sfixed_a(-0.001021790667437017)),(to_sfixed_a(-0.0035059915389865637)),(to_sfixed_a(-0.00010917324834736064)),(to_sfixed_a(-9.473746467847377e-05)),(to_sfixed_a(2.3345230601989897e-06)),(to_sfixed_a(0.00031600825604982674)),(to_sfixed_a(-2.598924947960768e-05)),(to_sfixed_a(2.4229737391578965e-05)),(to_sfixed_a(-2.9791570341330953e-05)),(to_sfixed_a(0.024903057143092155)),(to_sfixed_a(-0.0014262419426813722)),(to_sfixed_a(0.0824519544839859)),(to_sfixed_a(0.07429365813732147)),(to_sfixed_a(0.11435872316360474)),(to_sfixed_a(0.06610406190156937)),(to_sfixed_a(0.019042586907744408)),(to_sfixed_a(-0.038542456924915314)),(to_sfixed_a(-0.03409752622246742)),(to_sfixed_a(0.03857200965285301)),(to_sfixed_a(0.06478151679039001)),(to_sfixed_a(0.04847759008407593)),(to_sfixed_a(0.16870610415935516)),(to_sfixed_a(0.3574647903442383)),(to_sfixed_a(-0.16442552208900452)),(to_sfixed_a(0.004379505291581154)),(to_sfixed_a(0.36839836835861206)),(to_sfixed_a(0.17603203654289246)),(to_sfixed_a(0.20184722542762756)),(to_sfixed_a(-0.0010682088322937489)),(to_sfixed_a(0.15257211029529572)),(to_sfixed_a(-1.9413017071201466e-05)),(to_sfixed_a(-0.0002906890877056867)),(to_sfixed_a(-4.360649472801015e-05)),(to_sfixed_a(-0.0003274849441368133)),(to_sfixed_a(0.00014376711624208838)),(to_sfixed_a(6.92443354637362e-05)),(to_sfixed_a(5.588035855907947e-05)),(to_sfixed_a(-0.00011117883695987985)),(to_sfixed_a(0.24582478404045105)),(to_sfixed_a(0.2545233368873596)),(to_sfixed_a(-0.016419218853116035)),(to_sfixed_a(-0.03867952525615692)),(to_sfixed_a(-0.003756338730454445)),(to_sfixed_a(0.09135179966688156)),(to_sfixed_a(-0.108916275203228)),(to_sfixed_a(-0.012486188672482967)),(to_sfixed_a(-0.0533759668469429)),(to_sfixed_a(1.8348568119108677e-05)),(to_sfixed_a(0.17610050737857819)),(to_sfixed_a(0.12341871857643127)),(to_sfixed_a(0.015469444915652275)),(to_sfixed_a(0.03896002098917961)),(to_sfixed_a(0.07298284769058228)),(to_sfixed_a(0.1330508589744568)),(to_sfixed_a(0.018409578129649162)),(to_sfixed_a(0.16744579374790192)),(to_sfixed_a(0.02097965218126774)),(to_sfixed_a(8.267122757388279e-05)),(to_sfixed_a(-0.00016873983258847147)),(to_sfixed_a(0.0004116252239327878)),(to_sfixed_a(1.639819174670265e-06)),(to_sfixed_a(-1.3906823369325139e-05)),(to_sfixed_a(-0.00011293287388980389)),(to_sfixed_a(3.0266312023741193e-05)),(to_sfixed_a(-0.00024305206898134202)),(to_sfixed_a(-2.7813266569864936e-05)),(to_sfixed_a(0.0072787911631166935)),(to_sfixed_a(0.004451913293451071)),(to_sfixed_a(-0.09515495598316193)),(to_sfixed_a(-0.1469343602657318)),(to_sfixed_a(-0.02488250844180584)),(to_sfixed_a(-0.0025541833601891994)),(to_sfixed_a(0.013134806416928768)),(to_sfixed_a(-0.025420647114515305)),(to_sfixed_a(0.08519402891397476)),(to_sfixed_a(0.13762027025222778)),(to_sfixed_a(0.1272856891155243)),(to_sfixed_a(-0.21199771761894226)),(to_sfixed_a(0.19826360046863556)),(to_sfixed_a(0.2076367884874344)),(to_sfixed_a(0.08008814603090286)),(to_sfixed_a(0.06658018380403519)),(to_sfixed_a(0.13540491461753845)),(to_sfixed_a(0.018467610701918602)),(to_sfixed_a(0.0788128674030304)),(to_sfixed_a(6.230349754332565e-06)),(to_sfixed_a(-0.00020818340999539942)),(to_sfixed_a(-7.46997757232748e-05)),(to_sfixed_a(-2.9966875445097685e-05)),(to_sfixed_a(-0.00019185042765457183)),(to_sfixed_a(3.971230034949258e-05)),(to_sfixed_a(1.581774813530501e-05)),(to_sfixed_a(0.00011169433128088713)),(to_sfixed_a(-0.03285805881023407)),(to_sfixed_a(-0.011156320571899414)),(to_sfixed_a(-0.13406720757484436)),(to_sfixed_a(-0.03809838742017746)),(to_sfixed_a(0.040438421070575714)),(to_sfixed_a(0.1288684904575348)),(to_sfixed_a(0.011701575480401516)),(to_sfixed_a(-0.17189621925354004)),(to_sfixed_a(0.19326800107955933)),(to_sfixed_a(0.22991570830345154)),(to_sfixed_a(0.04115697741508484)),(to_sfixed_a(-0.04184042662382126)),(to_sfixed_a(0.054809365421533585)),(to_sfixed_a(0.18336783349514008)),(to_sfixed_a(0.0046334476210176945)),(to_sfixed_a(0.10413216054439545)),(to_sfixed_a(0.014499549753963947)),(to_sfixed_a(0.07107936590909958)),(to_sfixed_a(0.0326787605881691)),(to_sfixed_a(-0.012134594842791557)),(to_sfixed_a(4.1090112063102424e-05)),(to_sfixed_a(6.905145710334182e-05)),(to_sfixed_a(0.00016650703037157655)),(to_sfixed_a(0.00016284985758829862)),(to_sfixed_a(-0.00010284443851560354)),(to_sfixed_a(6.451935769291595e-05)),(to_sfixed_a(3.5118511732434854e-05)),(to_sfixed_a(9.791915363166481e-05)),(to_sfixed_a(0.00029029863071627915)),(to_sfixed_a(0.0007162429974414408)),(to_sfixed_a(-0.08269381523132324)),(to_sfixed_a(-0.1283893585205078)),(to_sfixed_a(0.08709853142499924)),(to_sfixed_a(0.19760243594646454)),(to_sfixed_a(-0.12301374226808548)),(to_sfixed_a(-0.08077728003263474)),(to_sfixed_a(0.17929641902446747)),(to_sfixed_a(0.09760143607854843)),(to_sfixed_a(0.04973122850060463)),(to_sfixed_a(0.0713476687669754)),(to_sfixed_a(-0.007532177958637476)),(to_sfixed_a(0.006305658724159002)),(to_sfixed_a(-0.021281694993376732)),(to_sfixed_a(-0.0529777929186821)),(to_sfixed_a(-0.19995881617069244)),(to_sfixed_a(-0.001227706321515143)),(to_sfixed_a(-0.005968286655843258)),(to_sfixed_a(-0.0069553907960653305)),(to_sfixed_a(0.00017940852558240294)),(to_sfixed_a(-0.0001115266204578802)),(to_sfixed_a(-2.185073753935285e-05)),(to_sfixed_a(-0.0004044943780172616)),(to_sfixed_a(8.787077240413055e-05)),(to_sfixed_a(-2.55371105595259e-05)),(to_sfixed_a(0.00019228372548241168)),(to_sfixed_a(0.0002811064769048244)),(to_sfixed_a(-0.00010533246677368879)),(to_sfixed_a(0.0008664940251037478)),(to_sfixed_a(0.0006665689288638532)),(to_sfixed_a(0.00021238332556094974)),(to_sfixed_a(-0.00028435763670131564)),(to_sfixed_a(0.0003053171094506979)),(to_sfixed_a(-0.03928607702255249)),(to_sfixed_a(-0.0027934580575674772)),(to_sfixed_a(-0.003792807227000594)),(to_sfixed_a(-0.017543014138936996)),(to_sfixed_a(-0.05902692303061485)),(to_sfixed_a(-1.1996325156360399e-05)),(to_sfixed_a(-0.0008678733720444143)),(to_sfixed_a(-0.026924634352326393)),(to_sfixed_a(-0.045989375561475754)),(to_sfixed_a(-0.014488794840872288)),(to_sfixed_a(-0.004388466943055391)),(to_sfixed_a(9.757166844792664e-05)),(to_sfixed_a(-0.0002559603308327496)),(to_sfixed_a(4.489445927902125e-05)),(to_sfixed_a(-0.00017128467152360827)),(to_sfixed_a(-0.00010715303506003693)),(to_sfixed_a(0.00020964397117495537)),(to_sfixed_a(2.0597961338353343e-05)),(to_sfixed_a(-0.0001602998818270862)),(to_sfixed_a(-5.6795634009176865e-05)),(to_sfixed_a(-9.06780333025381e-05)),(to_sfixed_a(4.413025180838304e-06)),(to_sfixed_a(0.00023918855004012585)),(to_sfixed_a(-0.00012374015932437032)),(to_sfixed_a(-2.791054248518776e-05)),(to_sfixed_a(-7.146277494030073e-05)),(to_sfixed_a(-3.6977486161049455e-05)),(to_sfixed_a(-0.0002057609090115875)),(to_sfixed_a(0.00012002480798400939)),(to_sfixed_a(-5.391574450186454e-05)),(to_sfixed_a(-0.00015932343376334757)),(to_sfixed_a(-7.592958809254924e-06)),(to_sfixed_a(3.667029523057863e-05)),(to_sfixed_a(6.853305239928886e-05)),(to_sfixed_a(-5.262075865175575e-05)),(to_sfixed_a(-1.2206746760057285e-05)),(to_sfixed_a(0.0003245816915296018)),(to_sfixed_a(-0.00010634025966282934)),(to_sfixed_a(0.00016566745762247592)),(to_sfixed_a(-9.268173016607761e-05)),(to_sfixed_a(-8.804537355899811e-05)),(to_sfixed_a(0.00033539452124387026)),(to_sfixed_a(9.398693509865552e-05)),(to_sfixed_a(-3.36627708747983e-05)),(to_sfixed_a(-6.536521686939523e-05)),(to_sfixed_a(-0.00018102675676345825)));

    constant weight_n0_22 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(9.30089590838179e-05)),(to_sfixed_a(-0.0001141368193202652)),(to_sfixed_a(0.0003616096219047904)),(to_sfixed_a(-0.0002460931136738509)),(to_sfixed_a(-9.584222425473854e-05)),(to_sfixed_a(-5.920068360865116e-05)),(to_sfixed_a(-5.081542258267291e-05)),(to_sfixed_a(4.9806512834038585e-05)),(to_sfixed_a(1.0653212484612595e-05)),(to_sfixed_a(0.00012668102863244712)),(to_sfixed_a(-0.00012344142305664718)),(to_sfixed_a(-0.00027464330196380615)),(to_sfixed_a(9.60480156209087e-06)),(to_sfixed_a(0.0002739091287367046)),(to_sfixed_a(-9.226102702086791e-05)),(to_sfixed_a(-0.00023443858663085848)),(to_sfixed_a(0.00019868477829732)),(to_sfixed_a(4.876780076301657e-05)),(to_sfixed_a(-8.344750676769763e-05)),(to_sfixed_a(3.064255361096002e-05)),(to_sfixed_a(-0.0002726087695918977)),(to_sfixed_a(0.00023278694425243884)),(to_sfixed_a(-6.591917190235108e-05)),(to_sfixed_a(1.6013087588362396e-05)),(to_sfixed_a(-0.00020669349760282785)),(to_sfixed_a(-1.0575114174571354e-05)),(to_sfixed_a(-5.2806237363256514e-05)),(to_sfixed_a(-2.844433947757352e-05)),(to_sfixed_a(3.1627958378521726e-05)),(to_sfixed_a(4.329051444074139e-05)),(to_sfixed_a(0.0004324782930780202)),(to_sfixed_a(-8.426508429693058e-05)),(to_sfixed_a(6.435617979150265e-05)),(to_sfixed_a(-3.2672000088496134e-05)),(to_sfixed_a(-7.672806532355025e-05)),(to_sfixed_a(0.00027138899895362556)),(to_sfixed_a(0.00038965896237641573)),(to_sfixed_a(-8.637288556201383e-05)),(to_sfixed_a(-0.00014224578626453876)),(to_sfixed_a(7.581055979244411e-05)),(to_sfixed_a(0.0001539283839520067)),(to_sfixed_a(0.0001160949032055214)),(to_sfixed_a(-0.00022118451306596398)),(to_sfixed_a(-8.712905400898308e-05)),(to_sfixed_a(5.103502553538419e-05)),(to_sfixed_a(0.00037841714220121503)),(to_sfixed_a(-6.457876224885695e-06)),(to_sfixed_a(-2.9607124815811403e-05)),(to_sfixed_a(0.00010711258801165968)),(to_sfixed_a(6.695129559375346e-05)),(to_sfixed_a(-0.00013040051271673292)),(to_sfixed_a(2.3618016712134704e-05)),(to_sfixed_a(-7.839460886316374e-05)),(to_sfixed_a(3.0291243092506193e-05)),(to_sfixed_a(7.670580816920847e-05)),(to_sfixed_a(0.00017926760483533144)),(to_sfixed_a(0.00012316204083617777)),(to_sfixed_a(3.640752038336359e-05)),(to_sfixed_a(-0.00016278575640171766)),(to_sfixed_a(-2.5584960894775577e-05)),(to_sfixed_a(-0.0003280450473539531)),(to_sfixed_a(-0.00020112346101086587)),(to_sfixed_a(-0.00017006430425681174)),(to_sfixed_a(-0.00028515179292298853)),(to_sfixed_a(0.00014757686585653573)),(to_sfixed_a(0.00011358861956978217)),(to_sfixed_a(-8.581051224609837e-05)),(to_sfixed_a(-6.0470443713711575e-05)),(to_sfixed_a(0.00014456808276008815)),(to_sfixed_a(0.024647634476423264)),(to_sfixed_a(-3.598910552682355e-06)),(to_sfixed_a(0.0001395200379192829)),(to_sfixed_a(-0.0002056737575912848)),(to_sfixed_a(-0.00011192197416676208)),(to_sfixed_a(0.0001203059364343062)),(to_sfixed_a(0.00024038211267907172)),(to_sfixed_a(-0.00022981151414569467)),(to_sfixed_a(8.460188109893352e-05)),(to_sfixed_a(4.35897454735823e-05)),(to_sfixed_a(-6.741996912751347e-05)),(to_sfixed_a(-0.0002587520284578204)),(to_sfixed_a(1.022926426230697e-05)),(to_sfixed_a(-3.855336763081141e-05)),(to_sfixed_a(-3.7973928556311876e-05)),(to_sfixed_a(5.348454578779638e-05)),(to_sfixed_a(1.829069333325606e-05)),(to_sfixed_a(-0.00021079614816699177)),(to_sfixed_a(-1.5503412214457057e-05)),(to_sfixed_a(-5.9302070440026e-05)),(to_sfixed_a(0.00022502515639644116)),(to_sfixed_a(-6.854889215901494e-05)),(to_sfixed_a(3.5772040973824915e-06)),(to_sfixed_a(0.01219844352453947)),(to_sfixed_a(5.956326276645996e-05)),(to_sfixed_a(0.013868660666048527)),(to_sfixed_a(0.04881562665104866)),(to_sfixed_a(0.03255581855773926)),(to_sfixed_a(-0.15109601616859436)),(to_sfixed_a(0.008372378535568714)),(to_sfixed_a(-0.13469800353050232)),(to_sfixed_a(0.007312300149351358)),(to_sfixed_a(-0.042442820966243744)),(to_sfixed_a(0.24922730028629303)),(to_sfixed_a(0.06959772109985352)),(to_sfixed_a(0.01087377779185772)),(to_sfixed_a(0.0219663567841053)),(to_sfixed_a(-0.00013774668332189322)),(to_sfixed_a(-0.00016123434761539102)),(to_sfixed_a(-0.00014616953558288515)),(to_sfixed_a(-0.000266707269474864)),(to_sfixed_a(-9.040033546625637e-06)),(to_sfixed_a(-0.00024039859999902546)),(to_sfixed_a(-3.810245470958762e-05)),(to_sfixed_a(0.00018608910613693297)),(to_sfixed_a(-0.00020956950902473181)),(to_sfixed_a(0.00018513508257456124)),(to_sfixed_a(-0.00014415837358683348)),(to_sfixed_a(-9.823724394664168e-05)),(to_sfixed_a(-0.0006705757114104927)),(to_sfixed_a(0.0693129375576973)),(to_sfixed_a(-0.009800187312066555)),(to_sfixed_a(0.015948543325066566)),(to_sfixed_a(-0.284808874130249)),(to_sfixed_a(-0.04907196760177612)),(to_sfixed_a(-0.3358887732028961)),(to_sfixed_a(-0.23260930180549622)),(to_sfixed_a(-0.18779656291007996)),(to_sfixed_a(-0.09184843301773071)),(to_sfixed_a(-0.032038234174251556)),(to_sfixed_a(0.12643326818943024)),(to_sfixed_a(0.11633433401584625)),(to_sfixed_a(-0.09148841351270676)),(to_sfixed_a(0.0072692520916461945)),(to_sfixed_a(0.03868453577160835)),(to_sfixed_a(-0.0019318744307383895)),(to_sfixed_a(-5.010911627323367e-05)),(to_sfixed_a(-0.0009440623689442873)),(to_sfixed_a(-6.264814146561548e-05)),(to_sfixed_a(-6.867179763503373e-05)),(to_sfixed_a(2.6972968043992296e-05)),(to_sfixed_a(2.5875815481413156e-05)),(to_sfixed_a(-1.52188267747988e-05)),(to_sfixed_a(-0.0002588619536254555)),(to_sfixed_a(6.148083775769919e-05)),(to_sfixed_a(0.0005580190918408334)),(to_sfixed_a(0.10233543813228607)),(to_sfixed_a(-0.002452944638207555)),(to_sfixed_a(-0.011778880842030048)),(to_sfixed_a(-0.04320696368813515)),(to_sfixed_a(0.009566732682287693)),(to_sfixed_a(0.07546570897102356)),(to_sfixed_a(-0.22852419316768646)),(to_sfixed_a(-0.202217698097229)),(to_sfixed_a(-0.12138873338699341)),(to_sfixed_a(-0.15398913621902466)),(to_sfixed_a(-0.1415228694677353)),(to_sfixed_a(-0.02880019322037697)),(to_sfixed_a(0.10090041160583496)),(to_sfixed_a(0.2936609387397766)),(to_sfixed_a(0.03799547627568245)),(to_sfixed_a(0.3274300694465637)),(to_sfixed_a(0.18120045959949493)),(to_sfixed_a(-0.0011956209782510996)),(to_sfixed_a(0.011463791131973267)),(to_sfixed_a(0.00475549278780818)),(to_sfixed_a(-0.00042452674824744463)),(to_sfixed_a(-0.00021723605459555984)),(to_sfixed_a(-0.00016119393694680184)),(to_sfixed_a(4.581085704558063e-06)),(to_sfixed_a(-0.00013134600885678083)),(to_sfixed_a(-0.00013666812446899712)),(to_sfixed_a(8.282998351205606e-06)),(to_sfixed_a(5.0344326155027375e-05)),(to_sfixed_a(0.1019153818488121)),(to_sfixed_a(0.06096098944544792)),(to_sfixed_a(0.1660737246274948)),(to_sfixed_a(0.07753074914216995)),(to_sfixed_a(0.13474255800247192)),(to_sfixed_a(0.17049920558929443)),(to_sfixed_a(0.15956106781959534)),(to_sfixed_a(-0.1066005676984787)),(to_sfixed_a(-0.015419556759297848)),(to_sfixed_a(-0.19948305189609528)),(to_sfixed_a(-0.3903319835662842)),(to_sfixed_a(-0.0579228401184082)),(to_sfixed_a(0.013467693701386452)),(to_sfixed_a(-0.014831740409135818)),(to_sfixed_a(0.05069788172841072)),(to_sfixed_a(0.12380588054656982)),(to_sfixed_a(-0.20767566561698914)),(to_sfixed_a(-0.06732066720724106)),(to_sfixed_a(0.06301376968622208)),(to_sfixed_a(0.004549616947770119)),(to_sfixed_a(0.0042016590014100075)),(to_sfixed_a(-0.00025391962844878435)),(to_sfixed_a(-0.000135341368149966)),(to_sfixed_a(3.2182972063310444e-05)),(to_sfixed_a(0.00019629354937933385)),(to_sfixed_a(5.853923357790336e-05)),(to_sfixed_a(4.0102786442730576e-05)),(to_sfixed_a(-0.00016119061911012977)),(to_sfixed_a(0.07222189009189606)),(to_sfixed_a(-0.053924981504678726)),(to_sfixed_a(0.015234889462590218)),(to_sfixed_a(0.08677516877651215)),(to_sfixed_a(0.31067150831222534)),(to_sfixed_a(0.38910195231437683)),(to_sfixed_a(0.4425455927848816)),(to_sfixed_a(0.2526502311229706)),(to_sfixed_a(0.1374613344669342)),(to_sfixed_a(0.10911889374256134)),(to_sfixed_a(0.05767231062054634)),(to_sfixed_a(-0.009793683886528015)),(to_sfixed_a(-0.19798848032951355)),(to_sfixed_a(-0.1653621643781662)),(to_sfixed_a(-0.3402492105960846)),(to_sfixed_a(0.11140618473291397)),(to_sfixed_a(0.24905024468898773)),(to_sfixed_a(-0.06104801595211029)),(to_sfixed_a(-0.1050960049033165)),(to_sfixed_a(0.04181892052292824)),(to_sfixed_a(0.00022472476121038198)),(to_sfixed_a(-0.00019469624385237694)),(to_sfixed_a(-0.00016165773558896035)),(to_sfixed_a(0.00013620297249872237)),(to_sfixed_a(0.0002211633836850524)),(to_sfixed_a(0.0001199150865431875)),(to_sfixed_a(0.00013840051542501897)),(to_sfixed_a(-0.0020851443987339735)),(to_sfixed_a(0.017940428107976913)),(to_sfixed_a(0.030383026227355003)),(to_sfixed_a(0.1078280583024025)),(to_sfixed_a(0.2347945123910904)),(to_sfixed_a(0.3086049556732178)),(to_sfixed_a(0.2762575149536133)),(to_sfixed_a(0.07242079824209213)),(to_sfixed_a(0.057319339364767075)),(to_sfixed_a(0.10011457651853561)),(to_sfixed_a(0.12546014785766602)),(to_sfixed_a(0.13999676704406738)),(to_sfixed_a(0.20865195989608765)),(to_sfixed_a(-0.09118477255105972)),(to_sfixed_a(0.10399597883224487)),(to_sfixed_a(0.29384317994117737)),(to_sfixed_a(0.059465859085321426)),(to_sfixed_a(-0.1672525703907013)),(to_sfixed_a(-0.009799527004361153)),(to_sfixed_a(-0.011580814607441425)),(to_sfixed_a(-0.024389464408159256)),(to_sfixed_a(0.0114658884704113)),(to_sfixed_a(0.00039323465898633003)),(to_sfixed_a(0.0003408946213312447)),(to_sfixed_a(-0.00013240572297945619)),(to_sfixed_a(-0.0001535353803774342)),(to_sfixed_a(0.00012428055924829096)),(to_sfixed_a(-3.16730365739204e-05)),(to_sfixed_a(0.000479463255032897)),(to_sfixed_a(-0.029677335172891617)),(to_sfixed_a(-0.021687237545847893)),(to_sfixed_a(-0.023126570507884026)),(to_sfixed_a(0.22425203025341034)),(to_sfixed_a(0.04892399534583092)),(to_sfixed_a(0.13853365182876587)),(to_sfixed_a(0.18135569989681244)),(to_sfixed_a(-0.08734313398599625)),(to_sfixed_a(-0.052634336054325104)),(to_sfixed_a(0.20437629520893097)),(to_sfixed_a(0.15273497998714447)),(to_sfixed_a(-0.17559491097927094)),(to_sfixed_a(-0.09630335867404938)),(to_sfixed_a(-0.10208581387996674)),(to_sfixed_a(0.31354963779449463)),(to_sfixed_a(0.20364800095558167)),(to_sfixed_a(0.009914143942296505)),(to_sfixed_a(-0.0008956214878708124)),(to_sfixed_a(0.09123403578996658)),(to_sfixed_a(0.16543284058570862)),(to_sfixed_a(-0.00015807533054612577)),(to_sfixed_a(5.1459566748235375e-05)),(to_sfixed_a(-1.600013092684094e-05)),(to_sfixed_a(7.925202226033434e-05)),(to_sfixed_a(-1.8018279661191627e-05)),(to_sfixed_a(-3.9419908716809005e-05)),(to_sfixed_a(2.9353266654652543e-05)),(to_sfixed_a(0.00990515761077404)),(to_sfixed_a(0.016339335590600967)),(to_sfixed_a(-0.29518187046051025)),(to_sfixed_a(-0.16708308458328247)),(to_sfixed_a(-0.18562369048595428)),(to_sfixed_a(-0.23123778402805328)),(to_sfixed_a(-0.18557700514793396)),(to_sfixed_a(-0.4898744225502014)),(to_sfixed_a(-0.35857707262039185)),(to_sfixed_a(0.289049357175827)),(to_sfixed_a(0.5149070024490356)),(to_sfixed_a(0.036285486072301865)),(to_sfixed_a(0.24494603276252747)),(to_sfixed_a(-0.04660782217979431)),(to_sfixed_a(0.08417771011590958)),(to_sfixed_a(-0.08540081232786179)),(to_sfixed_a(-0.14247293770313263)),(to_sfixed_a(-0.10634750127792358)),(to_sfixed_a(0.07998712360858917)),(to_sfixed_a(-0.027180997654795647)),(to_sfixed_a(0.12984615564346313)),(to_sfixed_a(0.03070209175348282)),(to_sfixed_a(-0.00014936845400370657)),(to_sfixed_a(0.00015050491492729634)),(to_sfixed_a(-4.275305400369689e-05)),(to_sfixed_a(-5.9971494920318946e-05)),(to_sfixed_a(5.996104300720617e-05)),(to_sfixed_a(-0.0036045562010258436)),(to_sfixed_a(-0.1259225755929947)),(to_sfixed_a(-0.10199978947639465)),(to_sfixed_a(-0.18387305736541748)),(to_sfixed_a(-0.07883468270301819)),(to_sfixed_a(0.07381106168031693)),(to_sfixed_a(0.10955300182104111)),(to_sfixed_a(-0.008014073595404625)),(to_sfixed_a(-0.04219832271337509)),(to_sfixed_a(0.18440407514572144)),(to_sfixed_a(0.1047896146774292)),(to_sfixed_a(0.201969176530838)),(to_sfixed_a(-0.1064540296792984)),(to_sfixed_a(0.011153279803693295)),(to_sfixed_a(0.12067665904760361)),(to_sfixed_a(-0.10398359596729279)),(to_sfixed_a(-0.042236968874931335)),(to_sfixed_a(-0.13083283603191376)),(to_sfixed_a(-0.03119659051299095)),(to_sfixed_a(0.06641563028097153)),(to_sfixed_a(-0.07865721732378006)),(to_sfixed_a(0.05174940451979637)),(to_sfixed_a(2.983902049891185e-05)),(to_sfixed_a(-4.008918403997086e-05)),(to_sfixed_a(0.00030367515864782035)),(to_sfixed_a(-0.00014135695528239012)),(to_sfixed_a(6.812807987444103e-05)),(to_sfixed_a(3.240280784666538e-05)),(to_sfixed_a(6.376351666403934e-05)),(to_sfixed_a(0.25336483120918274)),(to_sfixed_a(0.14236591756343842)),(to_sfixed_a(-0.054858822375535965)),(to_sfixed_a(0.2647669315338135)),(to_sfixed_a(-0.043457649648189545)),(to_sfixed_a(0.06136898323893547)),(to_sfixed_a(-0.07875190675258636)),(to_sfixed_a(-0.06833666563034058)),(to_sfixed_a(-0.17327271401882172)),(to_sfixed_a(0.1456606388092041)),(to_sfixed_a(-0.011066525243222713)),(to_sfixed_a(0.023867595940828323)),(to_sfixed_a(0.06332461535930634)),(to_sfixed_a(0.3348943591117859)),(to_sfixed_a(-0.0791463553905487)),(to_sfixed_a(-0.036112330853939056)),(to_sfixed_a(-0.3225177526473999)),(to_sfixed_a(0.019781839102506638)),(to_sfixed_a(0.031433649361133575)),(to_sfixed_a(0.1364257037639618)),(to_sfixed_a(-0.018336236476898193)),(to_sfixed_a(2.6824589440366253e-05)),(to_sfixed_a(-0.0006280721863731742)),(to_sfixed_a(0.00012217977200634778)),(to_sfixed_a(0.00010190224566031247)),(to_sfixed_a(-0.00012500771845225245)),(to_sfixed_a(-0.00014162086881697178)),(to_sfixed_a(-0.00015502578753512353)),(to_sfixed_a(-0.039011694490909576)),(to_sfixed_a(-0.13534818589687347)),(to_sfixed_a(-0.01299866009503603)),(to_sfixed_a(0.00027083768509328365)),(to_sfixed_a(0.1594996452331543)),(to_sfixed_a(-0.09887503832578659)),(to_sfixed_a(-0.051882632076740265)),(to_sfixed_a(-0.07644803076982498)),(to_sfixed_a(0.10616295039653778)),(to_sfixed_a(-0.02617020532488823)),(to_sfixed_a(-0.05192749202251434)),(to_sfixed_a(0.03534539043903351)),(to_sfixed_a(0.18725520372390747)),(to_sfixed_a(0.10884958505630493)),(to_sfixed_a(-0.045144062489271164)),(to_sfixed_a(-0.12750382721424103)),(to_sfixed_a(-0.11615470051765442)),(to_sfixed_a(-0.07627655565738678)),(to_sfixed_a(-0.0020068271551281214)),(to_sfixed_a(0.0903836116194725)),(to_sfixed_a(0.01319970190525055)),(to_sfixed_a(-0.002442873315885663)),(to_sfixed_a(-0.0028685869183391333)),(to_sfixed_a(-0.00012159493053331971)),(to_sfixed_a(0.00011728472600225359)),(to_sfixed_a(9.923018660629168e-05)),(to_sfixed_a(6.728143489453942e-05)),(to_sfixed_a(-3.975741856265813e-05)),(to_sfixed_a(0.0001464415981899947)),(to_sfixed_a(-0.12971541285514832)),(to_sfixed_a(-0.0987611711025238)),(to_sfixed_a(-0.20295609533786774)),(to_sfixed_a(-0.1597927063703537)),(to_sfixed_a(-0.08072227984666824)),(to_sfixed_a(0.009667185135185719)),(to_sfixed_a(-0.22151312232017517)),(to_sfixed_a(-0.029969481751322746)),(to_sfixed_a(-0.011381293646991253)),(to_sfixed_a(-0.18449227511882782)),(to_sfixed_a(0.001844066078774631)),(to_sfixed_a(-0.037235163152217865)),(to_sfixed_a(0.0003326204896438867)),(to_sfixed_a(-0.10720272362232208)),(to_sfixed_a(-0.14764952659606934)),(to_sfixed_a(-0.10554982721805573)),(to_sfixed_a(-0.14787599444389343)),(to_sfixed_a(-0.029459061101078987)),(to_sfixed_a(-0.08493094891309738)),(to_sfixed_a(-0.006193102803081274)),(to_sfixed_a(0.0003635472967289388)),(to_sfixed_a(-4.376457945909351e-05)),(to_sfixed_a(8.354719466296956e-05)),(to_sfixed_a(0.00017633575771469623)),(to_sfixed_a(-8.676337893120944e-05)),(to_sfixed_a(-0.0001775638374965638)),(to_sfixed_a(-0.000337195087922737)),(to_sfixed_a(-0.043921276926994324)),(to_sfixed_a(-0.08771338313817978)),(to_sfixed_a(0.023932812735438347)),(to_sfixed_a(-0.03733445331454277)),(to_sfixed_a(0.04597567766904831)),(to_sfixed_a(-0.06841777265071869)),(to_sfixed_a(-0.17752227187156677)),(to_sfixed_a(-0.10267313569784164)),(to_sfixed_a(-0.06081016734242439)),(to_sfixed_a(-0.012332557700574398)),(to_sfixed_a(-0.1299552470445633)),(to_sfixed_a(0.059736158698797226)),(to_sfixed_a(0.006783177610486746)),(to_sfixed_a(0.035864654928445816)),(to_sfixed_a(0.10310980677604675)),(to_sfixed_a(0.15410900115966797)),(to_sfixed_a(0.011485210619866848)),(to_sfixed_a(-0.050853170454502106)),(to_sfixed_a(-0.1701941192150116)),(to_sfixed_a(0.040004897862672806)),(to_sfixed_a(-0.12751927971839905)),(to_sfixed_a(0.0007155571947805583)),(to_sfixed_a(-3.975535946665332e-05)),(to_sfixed_a(-2.8507422030088492e-05)),(to_sfixed_a(-9.06995264813304e-05)),(to_sfixed_a(0.00041759980376809835)),(to_sfixed_a(-6.811112689319998e-05)),(to_sfixed_a(-0.004214882384985685)),(to_sfixed_a(-0.016886405646800995)),(to_sfixed_a(-0.03597017750144005)),(to_sfixed_a(-0.24186839163303375)),(to_sfixed_a(-0.09483370184898376)),(to_sfixed_a(0.0724104568362236)),(to_sfixed_a(0.12134937942028046)),(to_sfixed_a(0.13582412898540497)),(to_sfixed_a(-0.25585848093032837)),(to_sfixed_a(0.2465556263923645)),(to_sfixed_a(-0.023829765617847443)),(to_sfixed_a(0.09745382517576218)),(to_sfixed_a(-0.07642970979213715)),(to_sfixed_a(-0.09719064831733704)),(to_sfixed_a(-0.1913670152425766)),(to_sfixed_a(0.025534948334097862)),(to_sfixed_a(-0.17164002358913422)),(to_sfixed_a(-0.04038539528846741)),(to_sfixed_a(-0.21749863028526306)),(to_sfixed_a(-0.09781448543071747)),(to_sfixed_a(0.010479792021214962)),(to_sfixed_a(-0.02449209801852703)),(to_sfixed_a(-0.0016453786520287395)),(to_sfixed_a(8.451308531221002e-05)),(to_sfixed_a(0.00025947586982510984)),(to_sfixed_a(-9.140724432654679e-05)),(to_sfixed_a(9.909171058097854e-05)),(to_sfixed_a(-0.002785260323435068)),(to_sfixed_a(-0.0038725610356777906)),(to_sfixed_a(0.07093852013349533)),(to_sfixed_a(-0.010039770975708961)),(to_sfixed_a(-0.06875471770763397)),(to_sfixed_a(0.2618189752101898)),(to_sfixed_a(0.06872691214084625)),(to_sfixed_a(0.039233457297086716)),(to_sfixed_a(-0.2860114276409149)),(to_sfixed_a(0.04890996217727661)),(to_sfixed_a(0.4123234152793884)),(to_sfixed_a(-0.11677990108728409)),(to_sfixed_a(0.10991005599498749)),(to_sfixed_a(0.2282555252313614)),(to_sfixed_a(-0.19040457904338837)),(to_sfixed_a(0.10140155255794525)),(to_sfixed_a(0.006865955889225006)),(to_sfixed_a(-0.28527089953422546)),(to_sfixed_a(-0.01876949705183506)),(to_sfixed_a(-0.018077600747346878)),(to_sfixed_a(0.08630067110061646)),(to_sfixed_a(0.040802568197250366)),(to_sfixed_a(0.00020577931718435138)),(to_sfixed_a(0.00019858639279846102)),(to_sfixed_a(9.447361662751064e-05)),(to_sfixed_a(5.64411238883622e-05)),(to_sfixed_a(8.969780174084008e-05)),(to_sfixed_a(5.074505679658614e-05)),(to_sfixed_a(6.9964058639016e-05)),(to_sfixed_a(-0.0022156976629048586)),(to_sfixed_a(-0.11657752096652985)),(to_sfixed_a(-0.13130594789981842)),(to_sfixed_a(0.0029342761263251305)),(to_sfixed_a(-0.24000704288482666)),(to_sfixed_a(-0.18136806786060333)),(to_sfixed_a(-0.07793917506933212)),(to_sfixed_a(0.15212339162826538)),(to_sfixed_a(0.015242000110447407)),(to_sfixed_a(0.0632394477725029)),(to_sfixed_a(-0.007535027805715799)),(to_sfixed_a(0.1587533950805664)),(to_sfixed_a(0.3593682050704956)),(to_sfixed_a(0.20389553904533386)),(to_sfixed_a(-0.15051786601543427)),(to_sfixed_a(0.1163177415728569)),(to_sfixed_a(-0.16424985229969025)),(to_sfixed_a(0.03899144381284714)),(to_sfixed_a(-0.1834273487329483)),(to_sfixed_a(0.06265845149755478)),(to_sfixed_a(-0.039057061076164246)),(to_sfixed_a(-0.009998302906751633)),(to_sfixed_a(-0.000152716034790501)),(to_sfixed_a(0.00015931166126392782)),(to_sfixed_a(-0.0002809191064443439)),(to_sfixed_a(-0.0002419100346742198)),(to_sfixed_a(-8.068332681432366e-05)),(to_sfixed_a(-0.00019582179083954543)),(to_sfixed_a(-0.012869230471551418)),(to_sfixed_a(0.000810684752650559)),(to_sfixed_a(0.1713666170835495)),(to_sfixed_a(-0.026378579437732697)),(to_sfixed_a(0.008246710523962975)),(to_sfixed_a(0.027083251625299454)),(to_sfixed_a(-0.09196589142084122)),(to_sfixed_a(0.027077697217464447)),(to_sfixed_a(0.003070717677474022)),(to_sfixed_a(-0.047260332852602005)),(to_sfixed_a(-0.059698425233364105)),(to_sfixed_a(0.451760470867157)),(to_sfixed_a(0.49041086435317993)),(to_sfixed_a(0.18020519614219666)),(to_sfixed_a(0.272995263338089)),(to_sfixed_a(0.03424898907542229)),(to_sfixed_a(-0.014992950484156609)),(to_sfixed_a(-0.022619370371103287)),(to_sfixed_a(-0.041784726083278656)),(to_sfixed_a(0.014433205127716064)),(to_sfixed_a(0.3421419858932495)),(to_sfixed_a(1.8861849184759194e-06)),(to_sfixed_a(-0.00012888462515547872)),(to_sfixed_a(-4.465928668651031e-06)),(to_sfixed_a(0.00011427941353758797)),(to_sfixed_a(0.0003005823236890137)),(to_sfixed_a(0.0003004103491548449)),(to_sfixed_a(-4.05976788897533e-05)),(to_sfixed_a(6.843812298029661e-05)),(to_sfixed_a(0.005720121320337057)),(to_sfixed_a(0.04441573843359947)),(to_sfixed_a(0.007925482466816902)),(to_sfixed_a(0.5325366854667664)),(to_sfixed_a(0.13389436900615692)),(to_sfixed_a(0.06791534274816513)),(to_sfixed_a(0.09827659279108047)),(to_sfixed_a(-0.005236461292952299)),(to_sfixed_a(-0.34002694487571716)),(to_sfixed_a(0.01907675713300705)),(to_sfixed_a(0.30745929479599)),(to_sfixed_a(0.22491039335727692)),(to_sfixed_a(0.19632881879806519)),(to_sfixed_a(0.33680105209350586)),(to_sfixed_a(-0.09965648502111435)),(to_sfixed_a(0.07538405060768127)),(to_sfixed_a(-0.04990169778466225)),(to_sfixed_a(0.0041393679566681385)),(to_sfixed_a(0.2465861290693283)),(to_sfixed_a(0.01374957524240017)),(to_sfixed_a(-0.16459870338439941)),(to_sfixed_a(-0.0002857812214642763)),(to_sfixed_a(-8.141119178617373e-05)),(to_sfixed_a(0.00020461258827708662)),(to_sfixed_a(0.00012402971333358437)),(to_sfixed_a(0.00033902167342603207)),(to_sfixed_a(4.314333273214288e-05)),(to_sfixed_a(-0.00014591576473321766)),(to_sfixed_a(0.05312472954392433)),(to_sfixed_a(-0.00017215139814652503)),(to_sfixed_a(-0.0075328717939555645)),(to_sfixed_a(0.36026400327682495)),(to_sfixed_a(0.14984360337257385)),(to_sfixed_a(-0.1122153103351593)),(to_sfixed_a(0.08481377363204956)),(to_sfixed_a(0.15986576676368713)),(to_sfixed_a(-0.07246430963277817)),(to_sfixed_a(0.10573526471853256)),(to_sfixed_a(0.04066638648509979)),(to_sfixed_a(0.15422116219997406)),(to_sfixed_a(0.162151500582695)),(to_sfixed_a(0.34137243032455444)),(to_sfixed_a(0.07148241251707077)),(to_sfixed_a(-0.02629895508289337)),(to_sfixed_a(0.34702733159065247)),(to_sfixed_a(0.08303367346525192)),(to_sfixed_a(0.07206571102142334)),(to_sfixed_a(0.00011906329018529505)),(to_sfixed_a(0.04034276306629181)),(to_sfixed_a(5.647635043715127e-05)),(to_sfixed_a(0.0002206940989708528)),(to_sfixed_a(-7.319221185753122e-05)),(to_sfixed_a(-1.7661359379417263e-05)),(to_sfixed_a(-0.00011430075392127037)),(to_sfixed_a(1.2156095181126148e-05)),(to_sfixed_a(0.00012526358477771282)),(to_sfixed_a(3.953795021516271e-05)),(to_sfixed_a(0.01944003626704216)),(to_sfixed_a(-0.02217085473239422)),(to_sfixed_a(0.08800029754638672)),(to_sfixed_a(0.08635621517896652)),(to_sfixed_a(0.04208032786846161)),(to_sfixed_a(-0.030663127079606056)),(to_sfixed_a(0.11631830781698227)),(to_sfixed_a(-0.16444368660449982)),(to_sfixed_a(0.024655209854245186)),(to_sfixed_a(-0.01639540307223797)),(to_sfixed_a(0.25524452328681946)),(to_sfixed_a(0.02111034281551838)),(to_sfixed_a(0.024744121357798576)),(to_sfixed_a(-0.31654781103134155)),(to_sfixed_a(-0.18637578189373016)),(to_sfixed_a(0.08033672720193863)),(to_sfixed_a(0.03681833669543266)),(to_sfixed_a(0.07480016350746155)),(to_sfixed_a(-0.010140952654182911)),(to_sfixed_a(-2.8483185815275647e-05)),(to_sfixed_a(0.00014142520376481116)),(to_sfixed_a(4.497356712818146e-05)),(to_sfixed_a(-2.9819122573826462e-05)),(to_sfixed_a(-5.786433757748455e-05)),(to_sfixed_a(4.535575499176048e-05)),(to_sfixed_a(4.182458724244498e-05)),(to_sfixed_a(0.0002631047391332686)),(to_sfixed_a(0.00019794034596998245)),(to_sfixed_a(-0.010996517725288868)),(to_sfixed_a(-0.04898190125823021)),(to_sfixed_a(-0.1685728132724762)),(to_sfixed_a(-0.15049825608730316)),(to_sfixed_a(0.08196621388196945)),(to_sfixed_a(-0.13741335272789001)),(to_sfixed_a(-0.12182663381099701)),(to_sfixed_a(-0.02285337634384632)),(to_sfixed_a(-0.09101757407188416)),(to_sfixed_a(-0.13146838545799255)),(to_sfixed_a(0.16525737941265106)),(to_sfixed_a(0.0806327760219574)),(to_sfixed_a(0.01986563205718994)),(to_sfixed_a(0.020494142547249794)),(to_sfixed_a(-0.10379742085933685)),(to_sfixed_a(0.02661147154867649)),(to_sfixed_a(0.017256129533052444)),(to_sfixed_a(0.0003218049241695553)),(to_sfixed_a(0.012691043317317963)),(to_sfixed_a(5.5614433222217485e-05)),(to_sfixed_a(3.442436025125062e-08)),(to_sfixed_a(0.00015268393326550722)),(to_sfixed_a(-2.6511543183005415e-06)),(to_sfixed_a(-4.253935912856832e-05)),(to_sfixed_a(5.975679596303962e-05)),(to_sfixed_a(5.8130746765527874e-05)),(to_sfixed_a(7.594323960802285e-06)),(to_sfixed_a(0.03196222335100174)),(to_sfixed_a(-0.0644935816526413)),(to_sfixed_a(0.13445308804512024)),(to_sfixed_a(0.18380679190158844)),(to_sfixed_a(0.09661311656236649)),(to_sfixed_a(-0.019024232402443886)),(to_sfixed_a(-0.11327663064002991)),(to_sfixed_a(-0.0741729810833931)),(to_sfixed_a(0.07448500394821167)),(to_sfixed_a(-0.06704815477132797)),(to_sfixed_a(-0.035570528358221054)),(to_sfixed_a(-0.03609415143728256)),(to_sfixed_a(0.5615269541740417)),(to_sfixed_a(0.23427100479602814)),(to_sfixed_a(0.029768040403723717)),(to_sfixed_a(0.01722334884107113)),(to_sfixed_a(0.004962163511663675)),(to_sfixed_a(0.062352780252695084)),(to_sfixed_a(0.031421903520822525)),(to_sfixed_a(0.02399487979710102)),(to_sfixed_a(0.0001340207818429917)),(to_sfixed_a(0.00013712314830627292)),(to_sfixed_a(0.00016027968376874924)),(to_sfixed_a(-0.0001520127261755988)),(to_sfixed_a(0.00017916678916662931)),(to_sfixed_a(6.18074627709575e-05)),(to_sfixed_a(-8.912969497032464e-05)),(to_sfixed_a(-0.00021478622511494905)),(to_sfixed_a(-2.0418006897671148e-05)),(to_sfixed_a(-0.018460597842931747)),(to_sfixed_a(0.0808362290263176)),(to_sfixed_a(0.10591299831867218)),(to_sfixed_a(0.17116376757621765)),(to_sfixed_a(0.13114400207996368)),(to_sfixed_a(0.06567072123289108)),(to_sfixed_a(0.060223303735256195)),(to_sfixed_a(0.16691535711288452)),(to_sfixed_a(0.01424082275480032)),(to_sfixed_a(-0.06598923355340958)),(to_sfixed_a(0.04041671007871628)),(to_sfixed_a(0.28796327114105225)),(to_sfixed_a(-0.01372299250215292)),(to_sfixed_a(0.008942421525716782)),(to_sfixed_a(0.13517266511917114)),(to_sfixed_a(0.06974231451749802)),(to_sfixed_a(1.0653523531800602e-05)),(to_sfixed_a(0.005689979996532202)),(to_sfixed_a(0.006474176421761513)),(to_sfixed_a(-0.00022573959722649306)),(to_sfixed_a(0.0002573678793851286)),(to_sfixed_a(-5.4159660066943616e-05)),(to_sfixed_a(0.0003728085139300674)),(to_sfixed_a(-8.983469160739332e-05)),(to_sfixed_a(3.915772322216071e-05)),(to_sfixed_a(-5.445233909995295e-05)),(to_sfixed_a(-0.00020146858878433704)),(to_sfixed_a(6.61274534650147e-05)),(to_sfixed_a(0.00015104663907550275)),(to_sfixed_a(0.0004006718227174133)),(to_sfixed_a(-0.00013167363067623228)),(to_sfixed_a(0.0003485057095531374)),(to_sfixed_a(0.00034491921542212367)),(to_sfixed_a(0.0992157906293869)),(to_sfixed_a(0.004609346855431795)),(to_sfixed_a(0.0017368432600051165)),(to_sfixed_a(0.0707319900393486)),(to_sfixed_a(-0.05942154303193092)),(to_sfixed_a(-0.0018701571971178055)),(to_sfixed_a(0.012503692880272865)),(to_sfixed_a(0.07664833962917328)),(to_sfixed_a(0.10976691544055939)),(to_sfixed_a(0.01234468724578619)),(to_sfixed_a(0.006216626614332199)),(to_sfixed_a(-0.00015368218009825796)),(to_sfixed_a(-7.868585817050189e-05)),(to_sfixed_a(-0.000268178409896791)),(to_sfixed_a(-9.657781629357487e-05)),(to_sfixed_a(3.220434518880211e-05)),(to_sfixed_a(-0.000283298606518656)),(to_sfixed_a(0.00019519867782946676)),(to_sfixed_a(0.00016058249457273632)),(to_sfixed_a(-0.0001914928579935804)),(to_sfixed_a(0.0002589652722235769)),(to_sfixed_a(0.00042070134077221155)),(to_sfixed_a(-7.56857989472337e-05)),(to_sfixed_a(-0.00018506578635424376)),(to_sfixed_a(6.664393004029989e-05)),(to_sfixed_a(0.0001622998242964968)),(to_sfixed_a(4.238040492055006e-05)),(to_sfixed_a(1.5222558431560174e-05)),(to_sfixed_a(0.00035738194128498435)),(to_sfixed_a(5.620692536467686e-05)),(to_sfixed_a(4.5077584218233824e-05)),(to_sfixed_a(-1.4850415936962236e-05)),(to_sfixed_a(-8.558118133805692e-05)),(to_sfixed_a(9.110999235417694e-05)),(to_sfixed_a(0.00014767656102776527)),(to_sfixed_a(1.2446611435734667e-05)),(to_sfixed_a(-0.00011618408461799845)),(to_sfixed_a(5.4138894483912736e-05)),(to_sfixed_a(-0.00016198652156163007)),(to_sfixed_a(-0.00017696617578621954)),(to_sfixed_a(-0.00012663409870583564)),(to_sfixed_a(-0.0004233877407386899)),(to_sfixed_a(0.00027915631653741)),(to_sfixed_a(-9.95704103843309e-05)),(to_sfixed_a(-0.00028884317725896835)),(to_sfixed_a(9.900127042783424e-05)));

    constant weight_n0_23 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-0.00011601921141846105)),(to_sfixed_a(-0.0002163233730243519)),(to_sfixed_a(-0.00012752681504935026)),(to_sfixed_a(-4.87226752738934e-05)),(to_sfixed_a(6.708334694849327e-05)),(to_sfixed_a(0.0001311140658799559)),(to_sfixed_a(-0.0002564839960541576)),(to_sfixed_a(0.00011129478662041947)),(to_sfixed_a(4.303840978536755e-05)),(to_sfixed_a(0.0001542688114568591)),(to_sfixed_a(-3.006598308274988e-05)),(to_sfixed_a(4.182184056844562e-05)),(to_sfixed_a(-0.00011403690587030724)),(to_sfixed_a(8.790950960246846e-05)),(to_sfixed_a(2.9327038646442816e-05)),(to_sfixed_a(5.495574441738427e-06)),(to_sfixed_a(6.775656856916612e-06)),(to_sfixed_a(-0.00013872585259377956)),(to_sfixed_a(-0.00016244662401732057)),(to_sfixed_a(-0.00027630318072624505)),(to_sfixed_a(1.0967368325509597e-05)),(to_sfixed_a(0.0001474194141337648)),(to_sfixed_a(-2.7294268875266425e-05)),(to_sfixed_a(-2.9463997634593397e-05)),(to_sfixed_a(4.3294025999784935e-06)),(to_sfixed_a(6.0836056945845485e-05)),(to_sfixed_a(-0.000113005364255514)),(to_sfixed_a(1.3677893548447173e-05)),(to_sfixed_a(-0.00012868795602116734)),(to_sfixed_a(-8.912301564123482e-05)),(to_sfixed_a(7.860986079322174e-05)),(to_sfixed_a(0.00010297221160726622)),(to_sfixed_a(2.7232990760239772e-05)),(to_sfixed_a(0.0001807135558919981)),(to_sfixed_a(-0.00022417303989641368)),(to_sfixed_a(-5.060925832367502e-05)),(to_sfixed_a(-4.866716335527599e-05)),(to_sfixed_a(0.00013534356548916548)),(to_sfixed_a(-9.347897866973653e-05)),(to_sfixed_a(2.4629222025396302e-05)),(to_sfixed_a(-5.552994116442278e-05)),(to_sfixed_a(0.00012612409773282707)),(to_sfixed_a(0.00011500652180984616)),(to_sfixed_a(-0.00012510124361142516)),(to_sfixed_a(-9.741366375237703e-05)),(to_sfixed_a(3.769633258343674e-05)),(to_sfixed_a(8.465709106530994e-05)),(to_sfixed_a(-6.391126225935295e-05)),(to_sfixed_a(-3.700645174831152e-05)),(to_sfixed_a(-0.00016745933680795133)),(to_sfixed_a(-0.0003217133926227689)),(to_sfixed_a(-0.00015504955081269145)),(to_sfixed_a(-9.334718197351322e-05)),(to_sfixed_a(-0.00012371204502414912)),(to_sfixed_a(-5.3261013817973435e-05)),(to_sfixed_a(7.848672976251692e-05)),(to_sfixed_a(-1.2027701814076863e-05)),(to_sfixed_a(0.00017244857735931873)),(to_sfixed_a(-0.00012797700765077025)),(to_sfixed_a(0.0001599173410795629)),(to_sfixed_a(-0.00028786188340745866)),(to_sfixed_a(-2.1495387045433745e-05)),(to_sfixed_a(-3.298375304439105e-05)),(to_sfixed_a(2.5353154342155904e-05)),(to_sfixed_a(-2.3879287255113013e-05)),(to_sfixed_a(-7.683264266233891e-05)),(to_sfixed_a(-5.614882866211701e-06)),(to_sfixed_a(0.00028218983788974583)),(to_sfixed_a(2.5502982680336572e-05)),(to_sfixed_a(0.0023344201035797596)),(to_sfixed_a(5.873913687537424e-05)),(to_sfixed_a(-0.00015017272380646318)),(to_sfixed_a(0.0002884062996599823)),(to_sfixed_a(4.660283593693748e-05)),(to_sfixed_a(2.414970913378056e-05)),(to_sfixed_a(7.48398742871359e-05)),(to_sfixed_a(-0.00028304714942350984)),(to_sfixed_a(0.0001475704339100048)),(to_sfixed_a(0.0001621846604393795)),(to_sfixed_a(-0.00011540317791514099)),(to_sfixed_a(-0.00046544085489585996)),(to_sfixed_a(-0.00011759049812098965)),(to_sfixed_a(4.5799464714946225e-05)),(to_sfixed_a(0.00023995644005481154)),(to_sfixed_a(-2.134525857400149e-05)),(to_sfixed_a(4.72955362056382e-05)),(to_sfixed_a(-4.913688462693244e-05)),(to_sfixed_a(6.411961658159271e-05)),(to_sfixed_a(0.00010554873006185517)),(to_sfixed_a(4.6348734031198546e-05)),(to_sfixed_a(-2.577455416030716e-05)),(to_sfixed_a(0.00022430236276704818)),(to_sfixed_a(0.09724798798561096)),(to_sfixed_a(-0.00010383024346083403)),(to_sfixed_a(0.11037927120923996)),(to_sfixed_a(-0.0017339377664029598)),(to_sfixed_a(0.07778099924325943)),(to_sfixed_a(0.04487765580415726)),(to_sfixed_a(0.19556516408920288)),(to_sfixed_a(0.07863347232341766)),(to_sfixed_a(-0.011776736006140709)),(to_sfixed_a(0.09001533687114716)),(to_sfixed_a(0.07185465842485428)),(to_sfixed_a(-0.0074614412151277065)),(to_sfixed_a(-0.007071387488394976)),(to_sfixed_a(-0.014389114454388618)),(to_sfixed_a(-5.792119191028178e-05)),(to_sfixed_a(3.3963751775445417e-05)),(to_sfixed_a(0.0002373716124566272)),(to_sfixed_a(-0.00013692285574506968)),(to_sfixed_a(-0.0002281720080645755)),(to_sfixed_a(0.00012698165664914995)),(to_sfixed_a(1.9292705474072136e-05)),(to_sfixed_a(8.455578790744767e-05)),(to_sfixed_a(-3.10414943669457e-05)),(to_sfixed_a(-3.4628683351911604e-05)),(to_sfixed_a(-0.0001326552010141313)),(to_sfixed_a(-0.00025002218899317086)),(to_sfixed_a(0.0009521523024886847)),(to_sfixed_a(0.007133613806217909)),(to_sfixed_a(0.01862337626516819)),(to_sfixed_a(0.13913661241531372)),(to_sfixed_a(0.35551348328590393)),(to_sfixed_a(0.08017640560865402)),(to_sfixed_a(0.1338694989681244)),(to_sfixed_a(-0.021575266495347023)),(to_sfixed_a(0.05733545497059822)),(to_sfixed_a(0.30877333879470825)),(to_sfixed_a(0.3116661310195923)),(to_sfixed_a(0.3329114317893982)),(to_sfixed_a(0.18127740919589996)),(to_sfixed_a(0.07056828588247299)),(to_sfixed_a(-0.017788561061024666)),(to_sfixed_a(-0.051846858114004135)),(to_sfixed_a(-0.010598143562674522)),(to_sfixed_a(-7.1943386501516216e-06)),(to_sfixed_a(0.0006011728546582162)),(to_sfixed_a(-4.7612469643354416e-05)),(to_sfixed_a(0.00011684210039675236)),(to_sfixed_a(-0.00034790372592397034)),(to_sfixed_a(1.3451453924062662e-05)),(to_sfixed_a(0.00017660604498814791)),(to_sfixed_a(4.007302050013095e-05)),(to_sfixed_a(9.019357094075531e-05)),(to_sfixed_a(2.8128908979851985e-06)),(to_sfixed_a(0.007474400103092194)),(to_sfixed_a(0.0016783711034804583)),(to_sfixed_a(0.09535510092973709)),(to_sfixed_a(-0.006027034018188715)),(to_sfixed_a(-0.06428267806768417)),(to_sfixed_a(-0.09404739737510681)),(to_sfixed_a(-0.025637052953243256)),(to_sfixed_a(-0.40934282541275024)),(to_sfixed_a(-0.11977355927228928)),(to_sfixed_a(-0.22665180265903473)),(to_sfixed_a(-0.10092094540596008)),(to_sfixed_a(-0.023991946130990982)),(to_sfixed_a(-0.05899008363485336)),(to_sfixed_a(0.16349446773529053)),(to_sfixed_a(-0.026150476187467575)),(to_sfixed_a(0.023615822196006775)),(to_sfixed_a(-0.031746912747621536)),(to_sfixed_a(0.0022216401994228363)),(to_sfixed_a(-0.015612839721143246)),(to_sfixed_a(0.0011204268084838986)),(to_sfixed_a(0.0003087248478550464)),(to_sfixed_a(-0.0002550555218476802)),(to_sfixed_a(-0.00014974779332987964)),(to_sfixed_a(4.681356585933827e-05)),(to_sfixed_a(4.345432898844592e-05)),(to_sfixed_a(-0.00042787037091329694)),(to_sfixed_a(-4.509204518399201e-05)),(to_sfixed_a(-0.00017652774113230407)),(to_sfixed_a(0.007105047348886728)),(to_sfixed_a(0.020482584834098816)),(to_sfixed_a(-0.01585615798830986)),(to_sfixed_a(0.036212846636772156)),(to_sfixed_a(0.16422243416309357)),(to_sfixed_a(0.11397995799779892)),(to_sfixed_a(0.04370703920722008)),(to_sfixed_a(-0.1560208946466446)),(to_sfixed_a(-0.08277454227209091)),(to_sfixed_a(0.1298826038837433)),(to_sfixed_a(0.03880167752504349)),(to_sfixed_a(0.050321538001298904)),(to_sfixed_a(0.11749955266714096)),(to_sfixed_a(-0.01834927499294281)),(to_sfixed_a(-0.12614788115024567)),(to_sfixed_a(-0.15375038981437683)),(to_sfixed_a(-0.00585172651335597)),(to_sfixed_a(-0.11014669388532639)),(to_sfixed_a(-0.136493518948555)),(to_sfixed_a(-0.003442747052758932)),(to_sfixed_a(-0.00322755821980536)),(to_sfixed_a(-0.002900080755352974)),(to_sfixed_a(5.434912600321695e-05)),(to_sfixed_a(4.623647691914812e-05)),(to_sfixed_a(-0.0001207706518471241)),(to_sfixed_a(-2.723216857702937e-05)),(to_sfixed_a(7.420017209369689e-05)),(to_sfixed_a(-0.00015408672334160656)),(to_sfixed_a(-0.01666240394115448)),(to_sfixed_a(-0.031475283205509186)),(to_sfixed_a(0.0290627833455801)),(to_sfixed_a(0.04649614915251732)),(to_sfixed_a(-0.2135995328426361)),(to_sfixed_a(-0.11998997628688812)),(to_sfixed_a(-0.15450315177440643)),(to_sfixed_a(-0.069466233253479)),(to_sfixed_a(0.18135258555412292)),(to_sfixed_a(0.10034951567649841)),(to_sfixed_a(0.12344829738140106)),(to_sfixed_a(0.25294095277786255)),(to_sfixed_a(0.25900763273239136)),(to_sfixed_a(0.24541479349136353)),(to_sfixed_a(0.06676257401704788)),(to_sfixed_a(0.1638692021369934)),(to_sfixed_a(-0.1309695541858673)),(to_sfixed_a(-0.09827020019292831)),(to_sfixed_a(-0.4526226222515106)),(to_sfixed_a(-0.08457279950380325)),(to_sfixed_a(-0.00905109103769064)),(to_sfixed_a(-0.00010270836355630308)),(to_sfixed_a(-5.6308959756279364e-05)),(to_sfixed_a(6.101271992520196e-06)),(to_sfixed_a(-3.256669151596725e-05)),(to_sfixed_a(7.765574991935864e-05)),(to_sfixed_a(3.939937596442178e-05)),(to_sfixed_a(0.0021738759241998196)),(to_sfixed_a(-0.04598848521709442)),(to_sfixed_a(-0.05966496467590332)),(to_sfixed_a(0.1266924887895584)),(to_sfixed_a(-0.3605971038341522)),(to_sfixed_a(-0.020767932757735252)),(to_sfixed_a(-0.28436413407325745)),(to_sfixed_a(0.12629416584968567)),(to_sfixed_a(0.07165443897247314)),(to_sfixed_a(0.12867841124534607)),(to_sfixed_a(0.023109255358576775)),(to_sfixed_a(-0.1632278561592102)),(to_sfixed_a(0.26721951365470886)),(to_sfixed_a(-0.1436379849910736)),(to_sfixed_a(-0.21404509246349335)),(to_sfixed_a(-0.024085083976387978)),(to_sfixed_a(0.024155450984835625)),(to_sfixed_a(-0.003145280759781599)),(to_sfixed_a(-0.014050464145839214)),(to_sfixed_a(-0.1154838427901268)),(to_sfixed_a(-0.08328112959861755)),(to_sfixed_a(-0.02812815085053444)),(to_sfixed_a(4.5139589929021895e-05)),(to_sfixed_a(5.941283961874433e-05)),(to_sfixed_a(-0.0002953179646283388)),(to_sfixed_a(-4.870931661571376e-05)),(to_sfixed_a(2.174086148443166e-05)),(to_sfixed_a(0.00029492389876395464)),(to_sfixed_a(0.003222305793315172)),(to_sfixed_a(0.064301498234272)),(to_sfixed_a(0.00987542886286974)),(to_sfixed_a(0.044937923550605774)),(to_sfixed_a(0.13138286769390106)),(to_sfixed_a(-0.15538367629051208)),(to_sfixed_a(0.11980027705430984)),(to_sfixed_a(-0.10654576122760773)),(to_sfixed_a(0.540919303894043)),(to_sfixed_a(0.2362496703863144)),(to_sfixed_a(0.017116351053118706)),(to_sfixed_a(0.14156346023082733)),(to_sfixed_a(-0.006284942850470543)),(to_sfixed_a(0.09166866540908813)),(to_sfixed_a(-0.1487567275762558)),(to_sfixed_a(-0.02943110466003418)),(to_sfixed_a(0.11292458325624466)),(to_sfixed_a(-0.0760803148150444)),(to_sfixed_a(-0.09694190323352814)),(to_sfixed_a(-0.1197168156504631)),(to_sfixed_a(0.0479922890663147)),(to_sfixed_a(0.000129165273392573)),(to_sfixed_a(0.00016676573432050645)),(to_sfixed_a(-7.765492046019062e-05)),(to_sfixed_a(3.810979251284152e-05)),(to_sfixed_a(-8.105679444270208e-05)),(to_sfixed_a(0.00024134249542839825)),(to_sfixed_a(-0.00027666310779750347)),(to_sfixed_a(0.021141327917575836)),(to_sfixed_a(-0.0027612573467195034)),(to_sfixed_a(0.19776250422000885)),(to_sfixed_a(-0.07470208406448364)),(to_sfixed_a(-0.18024477362632751)),(to_sfixed_a(0.01781069114804268)),(to_sfixed_a(-0.25195634365081787)),(to_sfixed_a(0.0323844738304615)),(to_sfixed_a(0.06336932629346848)),(to_sfixed_a(-0.29717370867729187)),(to_sfixed_a(-0.0796896442770958)),(to_sfixed_a(0.3306393027305603)),(to_sfixed_a(0.21728374063968658)),(to_sfixed_a(0.04508262127637863)),(to_sfixed_a(-0.36314257979393005)),(to_sfixed_a(-0.14627042412757874)),(to_sfixed_a(0.09301115572452545)),(to_sfixed_a(-0.008173919282853603)),(to_sfixed_a(-0.01762854866683483)),(to_sfixed_a(0.16442880034446716)),(to_sfixed_a(-0.0591445229947567)),(to_sfixed_a(0.009983588941395283)),(to_sfixed_a(-1.1103807082690764e-05)),(to_sfixed_a(-3.117439700872637e-05)),(to_sfixed_a(0.0001245005551027134)),(to_sfixed_a(-6.385319466062356e-06)),(to_sfixed_a(1.522953334642807e-05)),(to_sfixed_a(-0.025065360590815544)),(to_sfixed_a(0.07186537981033325)),(to_sfixed_a(-0.1092294454574585)),(to_sfixed_a(0.04714890196919441)),(to_sfixed_a(-0.2727525532245636)),(to_sfixed_a(-0.02978779561817646)),(to_sfixed_a(-0.20519722998142242)),(to_sfixed_a(-0.054832104593515396)),(to_sfixed_a(0.10106442868709564)),(to_sfixed_a(-0.0033054142259061337)),(to_sfixed_a(-0.14707084000110626)),(to_sfixed_a(-0.2284073531627655)),(to_sfixed_a(-0.03678172454237938)),(to_sfixed_a(0.02374310977756977)),(to_sfixed_a(-0.2697789669036865)),(to_sfixed_a(-0.23921124637126923)),(to_sfixed_a(0.0890774205327034)),(to_sfixed_a(0.07654868066310883)),(to_sfixed_a(0.19658884406089783)),(to_sfixed_a(-0.11877981573343277)),(to_sfixed_a(0.014411033131182194)),(to_sfixed_a(-0.07780002802610397)),(to_sfixed_a(6.313443009275943e-05)),(to_sfixed_a(0.0003071219543926418)),(to_sfixed_a(-0.00019503181101754308)),(to_sfixed_a(-5.507751848199405e-05)),(to_sfixed_a(-6.278068030951545e-05)),(to_sfixed_a(-1.885706114990171e-05)),(to_sfixed_a(3.625658428063616e-05)),(to_sfixed_a(0.0048341890797019005)),(to_sfixed_a(-0.15632116794586182)),(to_sfixed_a(-0.11027663946151733)),(to_sfixed_a(-0.13350988924503326)),(to_sfixed_a(-0.027463404461741447)),(to_sfixed_a(-0.02904980629682541)),(to_sfixed_a(0.13208475708961487)),(to_sfixed_a(0.5247769951820374)),(to_sfixed_a(0.2589843273162842)),(to_sfixed_a(-0.22197198867797852)),(to_sfixed_a(0.06534204632043839)),(to_sfixed_a(-0.3740203082561493)),(to_sfixed_a(-0.14865508675575256)),(to_sfixed_a(-0.3211682140827179)),(to_sfixed_a(-0.0951349288225174)),(to_sfixed_a(-0.067538321018219)),(to_sfixed_a(0.11821594089269638)),(to_sfixed_a(0.09645209461450577)),(to_sfixed_a(0.11264907568693161)),(to_sfixed_a(0.29909610748291016)),(to_sfixed_a(-0.17839273810386658)),(to_sfixed_a(0.0001882036740425974)),(to_sfixed_a(-0.00017067328735720366)),(to_sfixed_a(0.00017756386660039425)),(to_sfixed_a(0.00022995664039626718)),(to_sfixed_a(0.00015245524991769344)),(to_sfixed_a(0.0003275912895333022)),(to_sfixed_a(4.294584505259991e-05)),(to_sfixed_a(0.04578031226992607)),(to_sfixed_a(0.028119809925556183)),(to_sfixed_a(-0.0002785100368782878)),(to_sfixed_a(0.009320713579654694)),(to_sfixed_a(-0.0719243511557579)),(to_sfixed_a(0.04676957055926323)),(to_sfixed_a(0.1575828343629837)),(to_sfixed_a(0.08363046497106552)),(to_sfixed_a(-0.048917703330516815)),(to_sfixed_a(0.19911973178386688)),(to_sfixed_a(-0.07820521295070648)),(to_sfixed_a(0.12156661599874496)),(to_sfixed_a(0.1501741111278534)),(to_sfixed_a(0.18206779658794403)),(to_sfixed_a(-0.040876906365156174)),(to_sfixed_a(0.22211915254592896)),(to_sfixed_a(-0.04968880116939545)),(to_sfixed_a(0.17950350046157837)),(to_sfixed_a(-0.004274609498679638)),(to_sfixed_a(-0.18112540245056152)),(to_sfixed_a(0.12441283464431763)),(to_sfixed_a(-6.283233960857615e-05)),(to_sfixed_a(-0.00023971145856194198)),(to_sfixed_a(1.0769477739813738e-05)),(to_sfixed_a(2.0254177798051387e-05)),(to_sfixed_a(0.0002547653566580266)),(to_sfixed_a(-3.904472032445483e-05)),(to_sfixed_a(-6.170341748656938e-06)),(to_sfixed_a(0.001375496038235724)),(to_sfixed_a(-0.03318153694272041)),(to_sfixed_a(-0.23976878821849823)),(to_sfixed_a(0.013940836302936077)),(to_sfixed_a(0.2134055644273758)),(to_sfixed_a(0.13549922406673431)),(to_sfixed_a(0.14060814678668976)),(to_sfixed_a(0.2688603401184082)),(to_sfixed_a(0.0928901880979538)),(to_sfixed_a(0.03987569734454155)),(to_sfixed_a(-0.11675358563661575)),(to_sfixed_a(-0.043978024274110794)),(to_sfixed_a(0.2486521601676941)),(to_sfixed_a(-0.08094165474176407)),(to_sfixed_a(-0.012500150129199028)),(to_sfixed_a(-0.12599892914295197)),(to_sfixed_a(0.04883555322885513)),(to_sfixed_a(-0.06986822187900543)),(to_sfixed_a(0.12234953045845032)),(to_sfixed_a(-0.3062070906162262)),(to_sfixed_a(0.028691867366433144)),(to_sfixed_a(0.0003799468104261905)),(to_sfixed_a(0.00030285221873782575)),(to_sfixed_a(0.00010306971671525389)),(to_sfixed_a(4.4573946070158854e-05)),(to_sfixed_a(-0.00013927639520261437)),(to_sfixed_a(0.0003351557534188032)),(to_sfixed_a(-9.63187703746371e-05)),(to_sfixed_a(-0.024195929989218712)),(to_sfixed_a(0.1361846625804901)),(to_sfixed_a(-0.03364657238125801)),(to_sfixed_a(-0.06716403365135193)),(to_sfixed_a(-0.08464756608009338)),(to_sfixed_a(-0.040024399757385254)),(to_sfixed_a(-0.05254259333014488)),(to_sfixed_a(0.09380540996789932)),(to_sfixed_a(-0.11999965459108353)),(to_sfixed_a(0.2246212661266327)),(to_sfixed_a(0.06263768672943115)),(to_sfixed_a(-0.020357992500066757)),(to_sfixed_a(-0.06435814499855042)),(to_sfixed_a(-0.14753445982933044)),(to_sfixed_a(-0.11249081790447235)),(to_sfixed_a(0.16509594023227692)),(to_sfixed_a(0.12188518792390823)),(to_sfixed_a(-0.010669432580471039)),(to_sfixed_a(-0.051444318145513535)),(to_sfixed_a(-0.14515094459056854)),(to_sfixed_a(-0.2654595375061035)),(to_sfixed_a(0.000568930699955672)),(to_sfixed_a(-0.00015473221719730645)),(to_sfixed_a(-0.00025153570459224284)),(to_sfixed_a(-6.408541230484843e-05)),(to_sfixed_a(5.52812525711488e-05)),(to_sfixed_a(-0.0002559498243499547)),(to_sfixed_a(7.773900870233774e-05)),(to_sfixed_a(0.002293638652190566)),(to_sfixed_a(-0.0047296457923948765)),(to_sfixed_a(0.10449273884296417)),(to_sfixed_a(0.08172936737537384)),(to_sfixed_a(-0.06801783293485641)),(to_sfixed_a(-0.08866186439990997)),(to_sfixed_a(-0.05055296793580055)),(to_sfixed_a(0.043419044464826584)),(to_sfixed_a(0.05004557967185974)),(to_sfixed_a(0.029263556003570557)),(to_sfixed_a(-0.04049352556467056)),(to_sfixed_a(-0.15230156481266022)),(to_sfixed_a(-0.17620833218097687)),(to_sfixed_a(-0.19736255705356598)),(to_sfixed_a(0.02573665976524353)),(to_sfixed_a(-0.17293529212474823)),(to_sfixed_a(-0.2367398589849472)),(to_sfixed_a(-0.2548803389072418)),(to_sfixed_a(-0.16667239367961884)),(to_sfixed_a(0.03176944702863693)),(to_sfixed_a(0.01875246874988079)),(to_sfixed_a(0.0015547010116279125)),(to_sfixed_a(0.00019262747082393616)),(to_sfixed_a(-0.0001592258777236566)),(to_sfixed_a(-1.2384119145281147e-05)),(to_sfixed_a(0.00010471702262293547)),(to_sfixed_a(-0.0005484100547619164)),(to_sfixed_a(0.00028453482082113624)),(to_sfixed_a(-0.04384263977408409)),(to_sfixed_a(-0.10504290461540222)),(to_sfixed_a(0.007551724556833506)),(to_sfixed_a(0.014993194490671158)),(to_sfixed_a(0.016213158145546913)),(to_sfixed_a(-0.03341284021735191)),(to_sfixed_a(0.05058441683650017)),(to_sfixed_a(-0.19785720109939575)),(to_sfixed_a(-0.20971670746803284)),(to_sfixed_a(-0.0446113720536232)),(to_sfixed_a(-0.1404525339603424)),(to_sfixed_a(0.2193039506673813)),(to_sfixed_a(-0.5312446355819702)),(to_sfixed_a(-0.09340813755989075)),(to_sfixed_a(0.0866864025592804)),(to_sfixed_a(-0.09967120736837387)),(to_sfixed_a(-0.18967868387699127)),(to_sfixed_a(-0.06969019025564194)),(to_sfixed_a(-0.17361387610435486)),(to_sfixed_a(0.03386196121573448)),(to_sfixed_a(0.00017273356206715107)),(to_sfixed_a(-7.545004336861894e-05)),(to_sfixed_a(-0.0004321052983868867)),(to_sfixed_a(-8.611316297901794e-05)),(to_sfixed_a(-2.9103790438966826e-05)),(to_sfixed_a(8.712432463653386e-05)),(to_sfixed_a(0.0002809561847243458)),(to_sfixed_a(0.027895933017134666)),(to_sfixed_a(-0.20373588800430298)),(to_sfixed_a(-0.12572549283504486)),(to_sfixed_a(0.08179434388875961)),(to_sfixed_a(0.16003870964050293)),(to_sfixed_a(0.09766307473182678)),(to_sfixed_a(0.054809413850307465)),(to_sfixed_a(0.18634019792079926)),(to_sfixed_a(0.05028150975704193)),(to_sfixed_a(0.2396792620420456)),(to_sfixed_a(-0.003532503731548786)),(to_sfixed_a(0.04622005298733711)),(to_sfixed_a(0.01996760629117489)),(to_sfixed_a(-0.10551534593105316)),(to_sfixed_a(0.003987955395132303)),(to_sfixed_a(-0.18161942064762115)),(to_sfixed_a(-0.1462559700012207)),(to_sfixed_a(-0.05133034661412239)),(to_sfixed_a(-0.22281362116336823)),(to_sfixed_a(-0.04242175444960594)),(to_sfixed_a(0.10067948698997498)),(to_sfixed_a(0.0033903021831065416)),(to_sfixed_a(8.322412031702697e-05)),(to_sfixed_a(0.00027378424420021474)),(to_sfixed_a(0.0003886939666699618)),(to_sfixed_a(0.00011091326450696215)),(to_sfixed_a(-0.00012485503975767642)),(to_sfixed_a(6.930870586074889e-05)),(to_sfixed_a(0.06044141575694084)),(to_sfixed_a(0.00577276898548007)),(to_sfixed_a(0.20191659033298492)),(to_sfixed_a(-0.01812433823943138)),(to_sfixed_a(-0.03665059059858322)),(to_sfixed_a(-0.19172973930835724)),(to_sfixed_a(-0.10427819192409515)),(to_sfixed_a(-0.18930666148662567)),(to_sfixed_a(0.06371723860502243)),(to_sfixed_a(0.15997080504894257)),(to_sfixed_a(0.16649824380874634)),(to_sfixed_a(0.03470630198717117)),(to_sfixed_a(-0.14868757128715515)),(to_sfixed_a(-0.04001929983496666)),(to_sfixed_a(0.2761826813220978)),(to_sfixed_a(-0.02147527225315571)),(to_sfixed_a(0.05278904363512993)),(to_sfixed_a(-0.11494406312704086)),(to_sfixed_a(0.07444581389427185)),(to_sfixed_a(-0.11604141443967819)),(to_sfixed_a(0.14370882511138916)),(to_sfixed_a(-2.476258850947488e-05)),(to_sfixed_a(0.0001439959742128849)),(to_sfixed_a(9.207557013723999e-05)),(to_sfixed_a(-0.000322660431265831)),(to_sfixed_a(-8.58221756061539e-05)),(to_sfixed_a(-6.936545833013952e-05)),(to_sfixed_a(-4.630681360140443e-05)),(to_sfixed_a(-9.96361777652055e-05)),(to_sfixed_a(0.024416567757725716)),(to_sfixed_a(-0.006488199811428785)),(to_sfixed_a(-0.1587899625301361)),(to_sfixed_a(-0.2823111414909363)),(to_sfixed_a(-0.19474917650222778)),(to_sfixed_a(-0.1505151391029358)),(to_sfixed_a(-0.18861250579357147)),(to_sfixed_a(0.07085536420345306)),(to_sfixed_a(-0.17378690838813782)),(to_sfixed_a(-0.08840205520391464)),(to_sfixed_a(0.1507178544998169)),(to_sfixed_a(0.2948244512081146)),(to_sfixed_a(0.07699396461248398)),(to_sfixed_a(0.14523746073246002)),(to_sfixed_a(-0.06078154221177101)),(to_sfixed_a(0.06931374222040176)),(to_sfixed_a(-0.22317489981651306)),(to_sfixed_a(0.056232843548059464)),(to_sfixed_a(-0.05023578554391861)),(to_sfixed_a(0.003093951614573598)),(to_sfixed_a(0.12652167677879333)),(to_sfixed_a(-0.00014227665087673813)),(to_sfixed_a(7.716643449384719e-05)),(to_sfixed_a(-0.00016613923071417958)),(to_sfixed_a(-0.00015291559975594282)),(to_sfixed_a(-0.00014635625120718032)),(to_sfixed_a(0.000253301695920527)),(to_sfixed_a(-0.0001462309155613184)),(to_sfixed_a(-0.0013130205916240811)),(to_sfixed_a(0.0004927863483317196)),(to_sfixed_a(-0.04088428243994713)),(to_sfixed_a(-0.24060171842575073)),(to_sfixed_a(-0.11145742982625961)),(to_sfixed_a(-0.050578318536281586)),(to_sfixed_a(-0.026476368308067322)),(to_sfixed_a(-0.24885597825050354)),(to_sfixed_a(-0.12205137312412262)),(to_sfixed_a(-0.06459462642669678)),(to_sfixed_a(0.22424550354480743)),(to_sfixed_a(0.07213301956653595)),(to_sfixed_a(0.04186665639281273)),(to_sfixed_a(0.11184969544410706)),(to_sfixed_a(-0.11414827406406403)),(to_sfixed_a(-0.13776731491088867)),(to_sfixed_a(-0.06855981796979904)),(to_sfixed_a(0.0735459253191948)),(to_sfixed_a(0.23033495247364044)),(to_sfixed_a(0.0008052511257119477)),(to_sfixed_a(0.019948117434978485)),(to_sfixed_a(0.00023411143047269434)),(to_sfixed_a(-8.668060036143288e-05)),(to_sfixed_a(7.20065800123848e-05)),(to_sfixed_a(0.00014792887668590993)),(to_sfixed_a(4.2422409023856744e-05)),(to_sfixed_a(-2.162333476007916e-05)),(to_sfixed_a(7.744703179923818e-05)),(to_sfixed_a(-0.00021525463671423495)),(to_sfixed_a(0.04275611415505409)),(to_sfixed_a(-0.08499788492918015)),(to_sfixed_a(-0.332073450088501)),(to_sfixed_a(0.11793849617242813)),(to_sfixed_a(-0.014469006098806858)),(to_sfixed_a(-0.14406676590442657)),(to_sfixed_a(-0.12183528393507004)),(to_sfixed_a(-0.14129862189292908)),(to_sfixed_a(-0.01267988421022892)),(to_sfixed_a(0.18200498819351196)),(to_sfixed_a(-0.012927298434078693)),(to_sfixed_a(-0.1731422245502472)),(to_sfixed_a(-0.0830303505063057)),(to_sfixed_a(-0.20966677367687225)),(to_sfixed_a(-0.09839139133691788)),(to_sfixed_a(0.13057667016983032)),(to_sfixed_a(0.026961814612150192)),(to_sfixed_a(0.02507905289530754)),(to_sfixed_a(-0.008603466674685478)),(to_sfixed_a(-3.83886435884051e-05)),(to_sfixed_a(2.095842319249641e-05)),(to_sfixed_a(0.0001468400441808626)),(to_sfixed_a(-3.318824019515887e-05)),(to_sfixed_a(0.00017417008348274976)),(to_sfixed_a(-0.00017328813555650413)),(to_sfixed_a(0.00011143913434352726)),(to_sfixed_a(3.319520146760624e-06)),(to_sfixed_a(-0.00040119889308698475)),(to_sfixed_a(0.006050348747521639)),(to_sfixed_a(-0.007562578655779362)),(to_sfixed_a(-0.09167242050170898)),(to_sfixed_a(0.025191530585289)),(to_sfixed_a(-0.055408820509910583)),(to_sfixed_a(-0.15220750868320465)),(to_sfixed_a(-0.2080700844526291)),(to_sfixed_a(-0.1746555119752884)),(to_sfixed_a(-0.10612078011035919)),(to_sfixed_a(-0.19139954447746277)),(to_sfixed_a(-0.29084184765815735)),(to_sfixed_a(0.19713860750198364)),(to_sfixed_a(-0.2856396436691284)),(to_sfixed_a(0.022240687161684036)),(to_sfixed_a(-0.03802013024687767)),(to_sfixed_a(-0.07709935307502747)),(to_sfixed_a(0.19894233345985413)),(to_sfixed_a(-0.010572620667517185)),(to_sfixed_a(0.15118177235126495)),(to_sfixed_a(-0.00011419851216487586)),(to_sfixed_a(0.0001724110043141991)),(to_sfixed_a(-0.00043885939521715045)),(to_sfixed_a(-0.0001221666025230661)),(to_sfixed_a(5.976892862236127e-05)),(to_sfixed_a(-0.000142143209814094)),(to_sfixed_a(-5.740731648984365e-05)),(to_sfixed_a(-0.00014366464165505022)),(to_sfixed_a(0.0369780957698822)),(to_sfixed_a(-0.04713660478591919)),(to_sfixed_a(0.15238763391971588)),(to_sfixed_a(0.27770617604255676)),(to_sfixed_a(0.04121110215783119)),(to_sfixed_a(-0.04372648522257805)),(to_sfixed_a(0.17254088819026947)),(to_sfixed_a(0.037934884428977966)),(to_sfixed_a(0.215419203042984)),(to_sfixed_a(-0.10034813731908798)),(to_sfixed_a(0.033010032027959824)),(to_sfixed_a(-0.11495441198348999)),(to_sfixed_a(0.0001266993349418044)),(to_sfixed_a(0.018884385004639626)),(to_sfixed_a(-0.05913364142179489)),(to_sfixed_a(0.12340523302555084)),(to_sfixed_a(0.00036003440618515015)),(to_sfixed_a(0.1293567717075348)),(to_sfixed_a(0.08557551354169846)),(to_sfixed_a(0.003974581137299538)),(to_sfixed_a(0.0001789087982615456)),(to_sfixed_a(0.00014741564518772066)),(to_sfixed_a(-4.928619091515429e-06)),(to_sfixed_a(0.0002242533810203895)),(to_sfixed_a(7.500473293475807e-05)),(to_sfixed_a(-5.5709100706735626e-05)),(to_sfixed_a(-0.00010869829566217959)),(to_sfixed_a(7.510944669775199e-06)),(to_sfixed_a(-7.76956367189996e-05)),(to_sfixed_a(0.013072728179395199)),(to_sfixed_a(0.09238643944263458)),(to_sfixed_a(0.14362065494060516)),(to_sfixed_a(0.35455530881881714)),(to_sfixed_a(0.2899055480957031)),(to_sfixed_a(0.11856714636087418)),(to_sfixed_a(0.2829822897911072)),(to_sfixed_a(0.1642153561115265)),(to_sfixed_a(0.06058049947023392)),(to_sfixed_a(0.17154797911643982)),(to_sfixed_a(0.167231947183609)),(to_sfixed_a(0.08500435203313828)),(to_sfixed_a(0.06320499628782272)),(to_sfixed_a(0.02634250558912754)),(to_sfixed_a(0.32217520475387573)),(to_sfixed_a(0.3138526380062103)),(to_sfixed_a(0.0005711580161005259)),(to_sfixed_a(-0.0014139498816803098)),(to_sfixed_a(-0.0026305809151381254)),(to_sfixed_a(0.00037914555286988616)),(to_sfixed_a(-3.4465076168999076e-05)),(to_sfixed_a(9.752236110216472e-06)),(to_sfixed_a(-1.9605135094025172e-05)),(to_sfixed_a(-2.800410584313795e-05)),(to_sfixed_a(0.0002945707819890231)),(to_sfixed_a(6.389418558683246e-05)),(to_sfixed_a(-0.0002689041430130601)),(to_sfixed_a(-0.0002940586127806455)),(to_sfixed_a(0.0003386867174413055)),(to_sfixed_a(0.0006525400676764548)),(to_sfixed_a(-4.564370101434179e-06)),(to_sfixed_a(-0.0003390988567844033)),(to_sfixed_a(0.00011253457341808826)),(to_sfixed_a(0.28319963812828064)),(to_sfixed_a(0.01074819266796112)),(to_sfixed_a(0.0022852562833577394)),(to_sfixed_a(0.20132136344909668)),(to_sfixed_a(-0.019236333668231964)),(to_sfixed_a(-0.013021484017372131)),(to_sfixed_a(0.09436935186386108)),(to_sfixed_a(0.21935486793518066)),(to_sfixed_a(0.30421581864356995)),(to_sfixed_a(0.021387863904237747)),(to_sfixed_a(0.011414609849452972)),(to_sfixed_a(-2.0316336303949356e-05)),(to_sfixed_a(0.00015280912339221686)),(to_sfixed_a(3.2144250781129813e-06)),(to_sfixed_a(-0.00013094881433062255)),(to_sfixed_a(0.00029517317307181656)),(to_sfixed_a(-0.0002000125532504171)),(to_sfixed_a(4.8000249080359936e-05)),(to_sfixed_a(-2.9123921194695868e-05)),(to_sfixed_a(4.421739868121222e-05)),(to_sfixed_a(-1.671405516390223e-05)),(to_sfixed_a(-0.00018897383415605873)),(to_sfixed_a(0.00014258715964388102)),(to_sfixed_a(0.00014068002928979695)),(to_sfixed_a(-0.00014673925761599094)),(to_sfixed_a(0.0002112862712237984)),(to_sfixed_a(7.445838855346665e-05)),(to_sfixed_a(0.00017346649838145822)),(to_sfixed_a(-0.00024936310364864767)),(to_sfixed_a(4.416022784425877e-05)),(to_sfixed_a(-6.736723298672587e-05)),(to_sfixed_a(-7.267492765095085e-05)),(to_sfixed_a(-0.0002769306011032313)),(to_sfixed_a(-0.00017202366143465042)),(to_sfixed_a(0.0001409802644047886)),(to_sfixed_a(0.00028754997765645385)),(to_sfixed_a(-2.8437245418899693e-05)),(to_sfixed_a(0.0001466566027374938)),(to_sfixed_a(-4.336787242209539e-05)),(to_sfixed_a(-0.00017471096361987293)),(to_sfixed_a(0.0001547480933368206)),(to_sfixed_a(-0.00021091375674586743)),(to_sfixed_a(-0.00015429315681103617)),(to_sfixed_a(0.00012892937229480594)),(to_sfixed_a(-0.00014111660129856318)),(to_sfixed_a(-0.0003841456491500139)));

    constant weight_n0_24 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-2.4797576770652086e-05)),(to_sfixed_a(-0.0002493081265129149)),(to_sfixed_a(8.995436655823141e-05)),(to_sfixed_a(6.249808211578056e-05)),(to_sfixed_a(0.00021491697407327592)),(to_sfixed_a(0.00012497718853410333)),(to_sfixed_a(0.00014120261766947806)),(to_sfixed_a(0.00017485729767940938)),(to_sfixed_a(-0.0001418017636751756)),(to_sfixed_a(2.6835389235202456e-06)),(to_sfixed_a(7.325374463107437e-05)),(to_sfixed_a(1.6436519217677414e-05)),(to_sfixed_a(-0.00014632764214184135)),(to_sfixed_a(-3.333255153847858e-05)),(to_sfixed_a(0.0002042984269792214)),(to_sfixed_a(3.0404362405533902e-05)),(to_sfixed_a(-2.2252268536249176e-05)),(to_sfixed_a(-0.00011810610885731876)),(to_sfixed_a(-0.00015164022624958307)),(to_sfixed_a(9.69221509876661e-05)),(to_sfixed_a(3.244213803554885e-05)),(to_sfixed_a(-5.2084993512835354e-05)),(to_sfixed_a(-0.0002485871082171798)),(to_sfixed_a(-6.0787446273025125e-05)),(to_sfixed_a(0.00018098601140081882)),(to_sfixed_a(5.715131192118861e-05)),(to_sfixed_a(-0.00014902447583153844)),(to_sfixed_a(1.8166849258705042e-05)),(to_sfixed_a(0.00016285393212456256)),(to_sfixed_a(1.8082113456330262e-05)),(to_sfixed_a(3.318421295261942e-05)),(to_sfixed_a(6.052446042303927e-05)),(to_sfixed_a(-9.126323129748926e-05)),(to_sfixed_a(-0.00040750083280727267)),(to_sfixed_a(-0.0004376503056846559)),(to_sfixed_a(9.229532588506117e-05)),(to_sfixed_a(0.00011433054169174284)),(to_sfixed_a(-9.67293162830174e-05)),(to_sfixed_a(-0.00028556579491123557)),(to_sfixed_a(0.0001405984367011115)),(to_sfixed_a(-8.630078809801489e-05)),(to_sfixed_a(0.00020413131278473884)),(to_sfixed_a(4.9531990953255445e-05)),(to_sfixed_a(-0.00016757794946897775)),(to_sfixed_a(9.346677688881755e-05)),(to_sfixed_a(0.00018770428141579032)),(to_sfixed_a(0.00019037051242776215)),(to_sfixed_a(-0.0002524971787352115)),(to_sfixed_a(0.0003262092359364033)),(to_sfixed_a(-7.594737689942122e-05)),(to_sfixed_a(0.00010562577517703176)),(to_sfixed_a(-6.942140316823497e-06)),(to_sfixed_a(-0.00033559114672243595)),(to_sfixed_a(8.044520654948428e-05)),(to_sfixed_a(-8.32660443847999e-05)),(to_sfixed_a(0.00016890365805011243)),(to_sfixed_a(-5.841208985657431e-05)),(to_sfixed_a(-8.933699427871034e-05)),(to_sfixed_a(0.00012992933625355363)),(to_sfixed_a(-5.86960231885314e-05)),(to_sfixed_a(0.00014720593753736466)),(to_sfixed_a(0.0001960937661351636)),(to_sfixed_a(0.00019038263417314738)),(to_sfixed_a(-4.3352578359190375e-05)),(to_sfixed_a(1.5695843103458174e-05)),(to_sfixed_a(-5.544501618715003e-05)),(to_sfixed_a(-0.0001544766128063202)),(to_sfixed_a(-0.0001246621395694092)),(to_sfixed_a(-9.169708391709719e-06)),(to_sfixed_a(-0.005344949662685394)),(to_sfixed_a(-1.8206206732429564e-05)),(to_sfixed_a(-0.00010434167052153498)),(to_sfixed_a(0.00018173463467974216)),(to_sfixed_a(0.00025079891202040017)),(to_sfixed_a(-8.313719445141032e-05)),(to_sfixed_a(0.0003294808848295361)),(to_sfixed_a(0.0001848601532401517)),(to_sfixed_a(-0.0002199723239755258)),(to_sfixed_a(8.920502295950428e-05)),(to_sfixed_a(-0.00016431468247901648)),(to_sfixed_a(-3.202934021828696e-05)),(to_sfixed_a(-9.875755495158955e-05)),(to_sfixed_a(1.9476970919640735e-05)),(to_sfixed_a(0.00011716829612851143)),(to_sfixed_a(1.3161150491214357e-05)),(to_sfixed_a(-7.981737326190341e-06)),(to_sfixed_a(-0.00015051172522362322)),(to_sfixed_a(-0.00021371233742684126)),(to_sfixed_a(0.00011643369361991063)),(to_sfixed_a(-0.00016417476581409574)),(to_sfixed_a(-0.00012899108696728945)),(to_sfixed_a(-4.324398105381988e-05)),(to_sfixed_a(0.0013928613625466824)),(to_sfixed_a(-7.213074422907084e-05)),(to_sfixed_a(0.0016037828754633665)),(to_sfixed_a(0.03349584341049194)),(to_sfixed_a(-0.0659794807434082)),(to_sfixed_a(-0.06293649226427078)),(to_sfixed_a(0.004998270887881517)),(to_sfixed_a(-0.0967145711183548)),(to_sfixed_a(0.010498994030058384)),(to_sfixed_a(-0.09361764788627625)),(to_sfixed_a(0.09342022985219955)),(to_sfixed_a(0.03066255711019039)),(to_sfixed_a(0.023169655352830887)),(to_sfixed_a(0.04718201234936714)),(to_sfixed_a(-0.00012491906818468124)),(to_sfixed_a(-2.3022421373752877e-06)),(to_sfixed_a(-3.619811832322739e-05)),(to_sfixed_a(-7.467021350748837e-05)),(to_sfixed_a(0.0001404795330017805)),(to_sfixed_a(-0.00014364391972776502)),(to_sfixed_a(8.922335837269202e-06)),(to_sfixed_a(9.33668197831139e-05)),(to_sfixed_a(-4.487738260650076e-05)),(to_sfixed_a(3.4980410418938845e-05)),(to_sfixed_a(-6.778255919925869e-05)),(to_sfixed_a(-0.00013134136679582298)),(to_sfixed_a(-0.00032655600807629526)),(to_sfixed_a(-0.004407562781125307)),(to_sfixed_a(0.020756447687745094)),(to_sfixed_a(0.0033042454160749912)),(to_sfixed_a(0.07849323749542236)),(to_sfixed_a(0.0263740923255682)),(to_sfixed_a(0.02787814848124981)),(to_sfixed_a(0.01169659849256277)),(to_sfixed_a(-0.06731416285037994)),(to_sfixed_a(-0.21486316621303558)),(to_sfixed_a(-0.28013864159584045)),(to_sfixed_a(0.0567668080329895)),(to_sfixed_a(-0.11090391874313354)),(to_sfixed_a(-0.001192005816847086)),(to_sfixed_a(-0.0075174300000071526)),(to_sfixed_a(0.13851867616176605)),(to_sfixed_a(0.00012550092651508749)),(to_sfixed_a(-0.0004439783515408635)),(to_sfixed_a(0.0005331698921509087)),(to_sfixed_a(-6.811659113736823e-05)),(to_sfixed_a(-0.00016895077715162188)),(to_sfixed_a(-7.897286559455097e-05)),(to_sfixed_a(3.426897819736041e-05)),(to_sfixed_a(1.9636650904431008e-05)),(to_sfixed_a(-0.0002220051974290982)),(to_sfixed_a(9.16870340006426e-05)),(to_sfixed_a(0.00017670441593509167)),(to_sfixed_a(0.017662398517131805)),(to_sfixed_a(0.01939469389617443)),(to_sfixed_a(-0.004115790128707886)),(to_sfixed_a(0.0733385756611824)),(to_sfixed_a(0.05960377678275108)),(to_sfixed_a(0.04375535249710083)),(to_sfixed_a(0.07720848172903061)),(to_sfixed_a(-0.08282936364412308)),(to_sfixed_a(-0.2641759216785431)),(to_sfixed_a(-0.3943995237350464)),(to_sfixed_a(-0.3929738402366638)),(to_sfixed_a(-0.20254004001617432)),(to_sfixed_a(-0.20888686180114746)),(to_sfixed_a(-0.15153884887695312)),(to_sfixed_a(-0.02775956690311432)),(to_sfixed_a(0.025536691769957542)),(to_sfixed_a(-0.005988139193505049)),(to_sfixed_a(-0.003066462930291891)),(to_sfixed_a(-0.004319500178098679)),(to_sfixed_a(-0.0005047988379374146)),(to_sfixed_a(-4.066448673256673e-05)),(to_sfixed_a(-9.155410225503147e-05)),(to_sfixed_a(-0.00032420316711068153)),(to_sfixed_a(1.3638798918691464e-05)),(to_sfixed_a(-5.245587817626074e-05)),(to_sfixed_a(-0.00012409724877215922)),(to_sfixed_a(0.0001861590426415205)),(to_sfixed_a(0.00033474480733275414)),(to_sfixed_a(0.012907445430755615)),(to_sfixed_a(-0.024486754089593887)),(to_sfixed_a(0.016593998298048973)),(to_sfixed_a(0.05337072163820267)),(to_sfixed_a(0.1330258697271347)),(to_sfixed_a(-0.1345328837633133)),(to_sfixed_a(0.06411825120449066)),(to_sfixed_a(0.15761293470859528)),(to_sfixed_a(-0.009603243321180344)),(to_sfixed_a(0.057609546929597855)),(to_sfixed_a(0.2738393247127533)),(to_sfixed_a(-0.061340078711509705)),(to_sfixed_a(0.054608531296253204)),(to_sfixed_a(0.2425065040588379)),(to_sfixed_a(-0.07147728651762009)),(to_sfixed_a(0.17924152314662933)),(to_sfixed_a(0.08652497828006744)),(to_sfixed_a(0.10371094942092896)),(to_sfixed_a(0.07115569710731506)),(to_sfixed_a(0.003659409936517477)),(to_sfixed_a(0.0062128761783242226)),(to_sfixed_a(0.0033439071848988533)),(to_sfixed_a(-0.00013714490341953933)),(to_sfixed_a(2.7284038878860883e-05)),(to_sfixed_a(-4.0886839997256175e-05)),(to_sfixed_a(-9.578492608852684e-05)),(to_sfixed_a(-4.319463187130168e-05)),(to_sfixed_a(-0.00031755055533722043)),(to_sfixed_a(-0.005978827364742756)),(to_sfixed_a(-0.07524312287569046)),(to_sfixed_a(0.09406434744596481)),(to_sfixed_a(-0.0822596624493599)),(to_sfixed_a(-0.024325212463736534)),(to_sfixed_a(-0.280898779630661)),(to_sfixed_a(0.03862221539020538)),(to_sfixed_a(0.08342365175485611)),(to_sfixed_a(0.1265680491924286)),(to_sfixed_a(0.16299042105674744)),(to_sfixed_a(0.48231834173202515)),(to_sfixed_a(0.1964389532804489)),(to_sfixed_a(-0.04255671426653862)),(to_sfixed_a(0.15286865830421448)),(to_sfixed_a(0.07310236990451813)),(to_sfixed_a(0.16219675540924072)),(to_sfixed_a(-0.06376779079437256)),(to_sfixed_a(0.12232102453708649)),(to_sfixed_a(0.014311318285763264)),(to_sfixed_a(0.03219222277402878)),(to_sfixed_a(0.0012386933667585254)),(to_sfixed_a(8.695734868524596e-05)),(to_sfixed_a(0.00015586134395562112)),(to_sfixed_a(-0.0002344949170947075)),(to_sfixed_a(5.3789182857144624e-05)),(to_sfixed_a(-6.362948624882847e-05)),(to_sfixed_a(-5.640040853904793e-06)),(to_sfixed_a(0.011982320807874203)),(to_sfixed_a(0.07753680646419525)),(to_sfixed_a(0.010687116533517838)),(to_sfixed_a(0.001985990907996893)),(to_sfixed_a(-0.05267097428441048)),(to_sfixed_a(0.2969520390033722)),(to_sfixed_a(0.3117060661315918)),(to_sfixed_a(0.019702237099409103)),(to_sfixed_a(0.21609273552894592)),(to_sfixed_a(0.10102876275777817)),(to_sfixed_a(0.08317827433347702)),(to_sfixed_a(-0.16686205565929413)),(to_sfixed_a(0.04845631495118141)),(to_sfixed_a(-0.020948894321918488)),(to_sfixed_a(-0.09509772807359695)),(to_sfixed_a(-0.07674302905797958)),(to_sfixed_a(-0.2333507537841797)),(to_sfixed_a(0.03314809128642082)),(to_sfixed_a(0.00011251925025135279)),(to_sfixed_a(-0.05120662599802017)),(to_sfixed_a(0.08042314648628235)),(to_sfixed_a(0.02388397604227066)),(to_sfixed_a(0.00013362836034502834)),(to_sfixed_a(0.00018633334548212588)),(to_sfixed_a(1.0050349374068901e-05)),(to_sfixed_a(-0.00016576313646510243)),(to_sfixed_a(-0.0001591813052073121)),(to_sfixed_a(1.4376467333931942e-05)),(to_sfixed_a(0.001804362633265555)),(to_sfixed_a(-0.030375778675079346)),(to_sfixed_a(0.03741149231791496)),(to_sfixed_a(0.003721445333212614)),(to_sfixed_a(-0.04975805804133415)),(to_sfixed_a(0.13617673516273499)),(to_sfixed_a(-0.032402362674474716)),(to_sfixed_a(0.08069057017564774)),(to_sfixed_a(0.1626041978597641)),(to_sfixed_a(-0.20856823027133942)),(to_sfixed_a(-0.10682805627584457)),(to_sfixed_a(-0.20352724194526672)),(to_sfixed_a(-0.07968060672283173)),(to_sfixed_a(0.14213135838508606)),(to_sfixed_a(-0.04653923213481903)),(to_sfixed_a(0.205153688788414)),(to_sfixed_a(0.03439170867204666)),(to_sfixed_a(-0.19055460393428802)),(to_sfixed_a(-0.14139050245285034)),(to_sfixed_a(-0.00962564256042242)),(to_sfixed_a(0.20086590945720673)),(to_sfixed_a(-7.928546256152913e-05)),(to_sfixed_a(-0.00010642661800375208)),(to_sfixed_a(-0.00023800857889000326)),(to_sfixed_a(-6.248497811611742e-05)),(to_sfixed_a(-0.00027718182536773384)),(to_sfixed_a(4.516535409493372e-05)),(to_sfixed_a(9.299594967160374e-05)),(to_sfixed_a(-0.00011354334856150672)),(to_sfixed_a(-0.019073782488703728)),(to_sfixed_a(-0.036225900053977966)),(to_sfixed_a(0.029424292966723442)),(to_sfixed_a(-0.10040058195590973)),(to_sfixed_a(-0.022962966933846474)),(to_sfixed_a(-0.014989785850048065)),(to_sfixed_a(0.1834455281496048)),(to_sfixed_a(0.2558709681034088)),(to_sfixed_a(-0.17872114479541779)),(to_sfixed_a(-0.0814608708024025)),(to_sfixed_a(-0.17752417922019958)),(to_sfixed_a(-0.2675938606262207)),(to_sfixed_a(-0.05495240539312363)),(to_sfixed_a(0.06381735950708389)),(to_sfixed_a(-0.015515717677772045)),(to_sfixed_a(0.11321806162595749)),(to_sfixed_a(-0.044670648872852325)),(to_sfixed_a(-0.10547402501106262)),(to_sfixed_a(-0.21648664772510529)),(to_sfixed_a(0.10196700692176819)),(to_sfixed_a(0.03857918456196785)),(to_sfixed_a(0.00012543305638246238)),(to_sfixed_a(0.00010400276369182393)),(to_sfixed_a(8.760791388340294e-05)),(to_sfixed_a(8.030587196117267e-05)),(to_sfixed_a(3.79885364054644e-07)),(to_sfixed_a(0.009912877343595028)),(to_sfixed_a(0.013515355065464973)),(to_sfixed_a(0.0002596850972622633)),(to_sfixed_a(0.04018055647611618)),(to_sfixed_a(0.07460466027259827)),(to_sfixed_a(-0.01938367821276188)),(to_sfixed_a(-0.11632487177848816)),(to_sfixed_a(0.0020224410109221935)),(to_sfixed_a(-0.07222261279821396)),(to_sfixed_a(0.22389481961727142)),(to_sfixed_a(0.405611515045166)),(to_sfixed_a(0.0988885909318924)),(to_sfixed_a(-0.10134318470954895)),(to_sfixed_a(-0.07780659198760986)),(to_sfixed_a(-0.03443615138530731)),(to_sfixed_a(0.33088967204093933)),(to_sfixed_a(0.10752074420452118)),(to_sfixed_a(0.012440711259841919)),(to_sfixed_a(-0.13267460465431213)),(to_sfixed_a(0.018769865855574608)),(to_sfixed_a(-0.060581546276807785)),(to_sfixed_a(-0.04158075898885727)),(to_sfixed_a(-0.00019053134019486606)),(to_sfixed_a(2.2514699594466947e-05)),(to_sfixed_a(-4.968982921127463e-06)),(to_sfixed_a(-2.1349148937588325e-06)),(to_sfixed_a(3.904652658093255e-06)),(to_sfixed_a(0.0001991358440136537)),(to_sfixed_a(1.7020543964463286e-05)),(to_sfixed_a(-0.032177072018384933)),(to_sfixed_a(0.0859169289469719)),(to_sfixed_a(0.03250772878527641)),(to_sfixed_a(0.07491950690746307)),(to_sfixed_a(-0.0036016572266817093)),(to_sfixed_a(-0.12137313187122345)),(to_sfixed_a(0.05930416285991669)),(to_sfixed_a(0.04053959250450134)),(to_sfixed_a(0.14049917459487915)),(to_sfixed_a(0.3948712646961212)),(to_sfixed_a(0.21510058641433716)),(to_sfixed_a(0.04972909763455391)),(to_sfixed_a(-0.058446746319532394)),(to_sfixed_a(-0.3375619947910309)),(to_sfixed_a(-0.06907343864440918)),(to_sfixed_a(0.13256359100341797)),(to_sfixed_a(-0.12458764016628265)),(to_sfixed_a(0.06330033391714096)),(to_sfixed_a(-0.15122149884700775)),(to_sfixed_a(-0.19076097011566162)),(to_sfixed_a(-0.2034531533718109)),(to_sfixed_a(-1.5224436538119335e-05)),(to_sfixed_a(3.651446240837686e-05)),(to_sfixed_a(-0.00023131757916416973)),(to_sfixed_a(0.00019555771723389626)),(to_sfixed_a(-0.0001817032170947641)),(to_sfixed_a(-0.0002208244550274685)),(to_sfixed_a(0.00029776926385238767)),(to_sfixed_a(0.0018435210222378373)),(to_sfixed_a(0.014394269324839115)),(to_sfixed_a(0.04906880110502243)),(to_sfixed_a(-0.09774341434240341)),(to_sfixed_a(-0.035166800022125244)),(to_sfixed_a(-0.1970919668674469)),(to_sfixed_a(-0.013660541735589504)),(to_sfixed_a(-0.16692937910556793)),(to_sfixed_a(-0.1805010885000229)),(to_sfixed_a(0.30953991413116455)),(to_sfixed_a(0.2457977533340454)),(to_sfixed_a(-0.026781408116221428)),(to_sfixed_a(-0.322732150554657)),(to_sfixed_a(-0.42859315872192383)),(to_sfixed_a(-0.16051310300827026)),(to_sfixed_a(-0.0825313925743103)),(to_sfixed_a(0.05895790085196495)),(to_sfixed_a(0.013228096999228)),(to_sfixed_a(-0.07405413687229156)),(to_sfixed_a(-0.18260304629802704)),(to_sfixed_a(0.0019152964232489467)),(to_sfixed_a(0.001048683887347579)),(to_sfixed_a(-0.0002349812421016395)),(to_sfixed_a(5.276147567201406e-05)),(to_sfixed_a(-0.00012699708167929202)),(to_sfixed_a(-0.00019191604224033654)),(to_sfixed_a(0.00017707885126583278)),(to_sfixed_a(0.00017207585915457457)),(to_sfixed_a(-0.0030922971200197935)),(to_sfixed_a(-0.12408258765935898)),(to_sfixed_a(-0.06510711461305618)),(to_sfixed_a(0.08290117233991623)),(to_sfixed_a(-0.12555652856826782)),(to_sfixed_a(-0.050622206181287766)),(to_sfixed_a(-0.4853018820285797)),(to_sfixed_a(-0.3401237726211548)),(to_sfixed_a(-0.0314810611307621)),(to_sfixed_a(0.06643538922071457)),(to_sfixed_a(0.011935851536691189)),(to_sfixed_a(-0.0008742918143980205)),(to_sfixed_a(-0.3534829914569855)),(to_sfixed_a(-0.16630946099758148)),(to_sfixed_a(-0.13814370334148407)),(to_sfixed_a(-0.08894473314285278)),(to_sfixed_a(0.06842830777168274)),(to_sfixed_a(0.17228010296821594)),(to_sfixed_a(0.0420045368373394)),(to_sfixed_a(0.09310712665319443)),(to_sfixed_a(-0.1234218180179596)),(to_sfixed_a(0.00046786508755758405)),(to_sfixed_a(0.0001481943327235058)),(to_sfixed_a(5.7088825997198e-05)),(to_sfixed_a(0.00011827399430330843)),(to_sfixed_a(-2.3632970624021254e-05)),(to_sfixed_a(3.2245505281025544e-05)),(to_sfixed_a(-9.620861237635836e-05)),(to_sfixed_a(0.05939008668065071)),(to_sfixed_a(-0.1283065378665924)),(to_sfixed_a(-0.08408626914024353)),(to_sfixed_a(-0.0977533832192421)),(to_sfixed_a(0.0250424612313509)),(to_sfixed_a(-0.07527493685483932)),(to_sfixed_a(-0.0730229914188385)),(to_sfixed_a(0.11506366729736328)),(to_sfixed_a(0.0748305693268776)),(to_sfixed_a(-0.16521278023719788)),(to_sfixed_a(0.05411918833851814)),(to_sfixed_a(0.003043519100174308)),(to_sfixed_a(-0.31288057565689087)),(to_sfixed_a(-0.06272819638252258)),(to_sfixed_a(0.0025207146536558867)),(to_sfixed_a(0.22112174332141876)),(to_sfixed_a(0.04967566579580307)),(to_sfixed_a(0.04741885885596275)),(to_sfixed_a(-0.0878097340464592)),(to_sfixed_a(0.07096780091524124)),(to_sfixed_a(0.1164681538939476)),(to_sfixed_a(0.00018936116248369217)),(to_sfixed_a(-5.862448233528994e-06)),(to_sfixed_a(0.00012391101336106658)),(to_sfixed_a(-5.363877789932303e-05)),(to_sfixed_a(0.00019344307656865567)),(to_sfixed_a(0.00019171411986462772)),(to_sfixed_a(-8.035587234189734e-05)),(to_sfixed_a(0.020975103601813316)),(to_sfixed_a(0.13531315326690674)),(to_sfixed_a(0.1931043267250061)),(to_sfixed_a(0.0862155631184578)),(to_sfixed_a(0.20879237353801727)),(to_sfixed_a(-0.09093798696994781)),(to_sfixed_a(0.2862173914909363)),(to_sfixed_a(-0.12030435353517532)),(to_sfixed_a(-0.2110752910375595)),(to_sfixed_a(-0.09811457991600037)),(to_sfixed_a(0.1667887419462204)),(to_sfixed_a(-0.048527803272008896)),(to_sfixed_a(-0.2673005759716034)),(to_sfixed_a(0.1584862619638443)),(to_sfixed_a(0.13787159323692322)),(to_sfixed_a(-0.07496879249811172)),(to_sfixed_a(-0.217863991856575)),(to_sfixed_a(-0.25677746534347534)),(to_sfixed_a(-0.059305526316165924)),(to_sfixed_a(-0.015244387090206146)),(to_sfixed_a(0.0567634291946888)),(to_sfixed_a(-0.014884291216731071)),(to_sfixed_a(-5.575894465437159e-05)),(to_sfixed_a(-0.0003190815623383969)),(to_sfixed_a(-0.0002684544015210122)),(to_sfixed_a(-7.77783861849457e-05)),(to_sfixed_a(0.000603934342507273)),(to_sfixed_a(-0.0001699892309261486)),(to_sfixed_a(0.004883157089352608)),(to_sfixed_a(0.1874251663684845)),(to_sfixed_a(0.137647345662117)),(to_sfixed_a(0.3412761390209198)),(to_sfixed_a(0.3628777265548706)),(to_sfixed_a(0.09824802726507187)),(to_sfixed_a(-0.2369992583990097)),(to_sfixed_a(-0.0055710747838020325)),(to_sfixed_a(-0.16104629635810852)),(to_sfixed_a(-0.022751718759536743)),(to_sfixed_a(-0.05149796977639198)),(to_sfixed_a(-0.2595163583755493)),(to_sfixed_a(-0.19144576787948608)),(to_sfixed_a(0.010753404349088669)),(to_sfixed_a(0.11128571629524231)),(to_sfixed_a(0.3612508475780487)),(to_sfixed_a(-0.02333858422935009)),(to_sfixed_a(-0.014504139311611652)),(to_sfixed_a(-0.06295792013406754)),(to_sfixed_a(-0.007004988379776478)),(to_sfixed_a(-0.0001214460062328726)),(to_sfixed_a(2.0391826183185913e-05)),(to_sfixed_a(0.0001373653649352491)),(to_sfixed_a(4.119041113881394e-05)),(to_sfixed_a(0.00014732587442267686)),(to_sfixed_a(-0.0003159437037538737)),(to_sfixed_a(-0.0002198079164372757)),(to_sfixed_a(-0.048383165150880814)),(to_sfixed_a(0.05212986841797829)),(to_sfixed_a(-0.04384736344218254)),(to_sfixed_a(-0.11223267018795013)),(to_sfixed_a(-0.13478009402751923)),(to_sfixed_a(-0.18525545299053192)),(to_sfixed_a(-0.09267912060022354)),(to_sfixed_a(0.028250563889741898)),(to_sfixed_a(-0.11764369159936905)),(to_sfixed_a(0.08749982714653015)),(to_sfixed_a(-0.2689025402069092)),(to_sfixed_a(-0.016977818682789803)),(to_sfixed_a(-0.04843095317482948)),(to_sfixed_a(0.06432313472032547)),(to_sfixed_a(0.2468382567167282)),(to_sfixed_a(0.005686550866812468)),(to_sfixed_a(0.09717771410942078)),(to_sfixed_a(-0.05662389099597931)),(to_sfixed_a(-0.06956221908330917)),(to_sfixed_a(-0.05494842305779457)),(to_sfixed_a(0.009847485460340977)),(to_sfixed_a(-0.013047704473137856)),(to_sfixed_a(0.00011423137766541913)),(to_sfixed_a(-0.00014675865531899035)),(to_sfixed_a(0.00015016285760793835)),(to_sfixed_a(-0.00018824462313205004)),(to_sfixed_a(0.00021947217464912683)),(to_sfixed_a(0.0001287525665247813)),(to_sfixed_a(0.03203349933028221)),(to_sfixed_a(0.006583586800843477)),(to_sfixed_a(0.04492245614528656)),(to_sfixed_a(-0.029953710734844208)),(to_sfixed_a(-0.17954015731811523)),(to_sfixed_a(-0.25489041209220886)),(to_sfixed_a(-0.32664674520492554)),(to_sfixed_a(-0.23547759652137756)),(to_sfixed_a(-0.02464151568710804)),(to_sfixed_a(0.08232280611991882)),(to_sfixed_a(0.1959284394979477)),(to_sfixed_a(0.07906598597764969)),(to_sfixed_a(0.12643422186374664)),(to_sfixed_a(0.32931649684906006)),(to_sfixed_a(0.18864953517913818)),(to_sfixed_a(0.07988390326499939)),(to_sfixed_a(0.005940482951700687)),(to_sfixed_a(-0.07212915271520615)),(to_sfixed_a(-0.07592812180519104)),(to_sfixed_a(-0.12230190634727478)),(to_sfixed_a(0.08373624086380005)),(to_sfixed_a(3.221637598471716e-05)),(to_sfixed_a(2.6849582354770973e-05)),(to_sfixed_a(-5.6799948652042076e-05)),(to_sfixed_a(7.054554589558393e-05)),(to_sfixed_a(-0.00011242698383284733)),(to_sfixed_a(-1.1943508297918015e-06)),(to_sfixed_a(-0.000186465447768569)),(to_sfixed_a(2.5657564037828706e-05)),(to_sfixed_a(-0.005356261041015387)),(to_sfixed_a(0.11344993114471436)),(to_sfixed_a(-0.03225213289260864)),(to_sfixed_a(-0.2563006579875946)),(to_sfixed_a(-0.020692629739642143)),(to_sfixed_a(-0.2717704474925995)),(to_sfixed_a(-0.15523160994052887)),(to_sfixed_a(-0.029683634638786316)),(to_sfixed_a(0.1489003747701645)),(to_sfixed_a(0.2301318347454071)),(to_sfixed_a(-0.011184850707650185)),(to_sfixed_a(-0.020123863592743874)),(to_sfixed_a(0.053162831813097)),(to_sfixed_a(0.09692159295082092)),(to_sfixed_a(0.11233580112457275)),(to_sfixed_a(0.088036447763443)),(to_sfixed_a(0.11711946874856949)),(to_sfixed_a(-0.07105372846126556)),(to_sfixed_a(0.25834783911705017)),(to_sfixed_a(0.10816911607980728)),(to_sfixed_a(-0.018817821517586708)),(to_sfixed_a(9.531163959763944e-05)),(to_sfixed_a(0.00016247309395112097)),(to_sfixed_a(-8.202201570384204e-05)),(to_sfixed_a(7.871176057960838e-05)),(to_sfixed_a(0.00011868305591633543)),(to_sfixed_a(-7.789128721924499e-05)),(to_sfixed_a(-0.00010306111653335392)),(to_sfixed_a(-0.023726286366581917)),(to_sfixed_a(0.0026191161014139652)),(to_sfixed_a(-0.2214023321866989)),(to_sfixed_a(-0.0701904222369194)),(to_sfixed_a(-0.011151178739964962)),(to_sfixed_a(0.12128006666898727)),(to_sfixed_a(-0.12178324162960052)),(to_sfixed_a(-0.0691547766327858)),(to_sfixed_a(0.2538486123085022)),(to_sfixed_a(0.46681979298591614)),(to_sfixed_a(0.20611046254634857)),(to_sfixed_a(-0.03933808580040932)),(to_sfixed_a(-0.06939585506916046)),(to_sfixed_a(0.06579797714948654)),(to_sfixed_a(0.12513498961925507)),(to_sfixed_a(0.009879333898425102)),(to_sfixed_a(0.4267095923423767)),(to_sfixed_a(0.11132638156414032)),(to_sfixed_a(-0.28661006689071655)),(to_sfixed_a(-0.001946194563060999)),(to_sfixed_a(0.1193029135465622)),(to_sfixed_a(0.0001766321947798133)),(to_sfixed_a(0.00013693486107513309)),(to_sfixed_a(-2.597360980871599e-05)),(to_sfixed_a(0.00042342464439570904)),(to_sfixed_a(0.00012689479626715183)),(to_sfixed_a(-0.00011696890578605235)),(to_sfixed_a(-5.156509723747149e-05)),(to_sfixed_a(0.00015177465684246272)),(to_sfixed_a(-0.03593485802412033)),(to_sfixed_a(0.016089674085378647)),(to_sfixed_a(-0.027400780469179153)),(to_sfixed_a(-0.16117389500141144)),(to_sfixed_a(-0.07981877028942108)),(to_sfixed_a(0.3099870979785919)),(to_sfixed_a(0.08140619099140167)),(to_sfixed_a(0.2629060745239258)),(to_sfixed_a(-0.018661368638277054)),(to_sfixed_a(0.01131205353885889)),(to_sfixed_a(0.16291911900043488)),(to_sfixed_a(0.11483561992645264)),(to_sfixed_a(0.005021529272198677)),(to_sfixed_a(0.0961901843547821)),(to_sfixed_a(0.14086377620697021)),(to_sfixed_a(0.05094296857714653)),(to_sfixed_a(0.004815702326595783)),(to_sfixed_a(0.13157334923744202)),(to_sfixed_a(-1.3113699424138758e-05)),(to_sfixed_a(2.6324646569264587e-06)),(to_sfixed_a(-0.0001255456736544147)),(to_sfixed_a(-0.00026007040287368)),(to_sfixed_a(-8.85535919223912e-05)),(to_sfixed_a(0.00020542154379654676)),(to_sfixed_a(-4.6692606701981276e-05)),(to_sfixed_a(-0.00012811129272449762)),(to_sfixed_a(-0.0002053633943432942)),(to_sfixed_a(0.0003208066336810589)),(to_sfixed_a(-0.0062112282030284405)),(to_sfixed_a(0.017497166991233826)),(to_sfixed_a(0.033080220222473145)),(to_sfixed_a(-0.09281608462333679)),(to_sfixed_a(0.002431939821690321)),(to_sfixed_a(0.021234504878520966)),(to_sfixed_a(0.02979404479265213)),(to_sfixed_a(0.12705503404140472)),(to_sfixed_a(0.12678469717502594)),(to_sfixed_a(0.1272905021905899)),(to_sfixed_a(0.018486235290765762)),(to_sfixed_a(-0.28563031554222107)),(to_sfixed_a(-0.15203335881233215)),(to_sfixed_a(-0.2392560988664627)),(to_sfixed_a(-0.1836206018924713)),(to_sfixed_a(-0.005655318032950163)),(to_sfixed_a(-0.2556810677051544)),(to_sfixed_a(0.005415629595518112)),(to_sfixed_a(-0.20125916600227356)),(to_sfixed_a(0.00013184305862523615)),(to_sfixed_a(2.7799631425295956e-05)),(to_sfixed_a(-0.0001588188752066344)),(to_sfixed_a(8.035547216422856e-05)),(to_sfixed_a(0.0002445066347718239)),(to_sfixed_a(7.177567749749869e-05)),(to_sfixed_a(-9.234531171387061e-05)),(to_sfixed_a(1.9152257664245553e-05)),(to_sfixed_a(0.04166688397526741)),(to_sfixed_a(-0.01744893752038479)),(to_sfixed_a(0.1716482937335968)),(to_sfixed_a(0.11600859463214874)),(to_sfixed_a(-0.007794809993356466)),(to_sfixed_a(-0.11422119289636612)),(to_sfixed_a(-0.02601052261888981)),(to_sfixed_a(0.041226595640182495)),(to_sfixed_a(-0.09563585370779037)),(to_sfixed_a(-0.2504865527153015)),(to_sfixed_a(-0.01842259056866169)),(to_sfixed_a(-0.05276557058095932)),(to_sfixed_a(-0.3047628700733185)),(to_sfixed_a(-0.26126307249069214)),(to_sfixed_a(-0.012633849866688251)),(to_sfixed_a(-0.24620072543621063)),(to_sfixed_a(0.014188004657626152)),(to_sfixed_a(-0.1990646868944168)),(to_sfixed_a(-0.10120692849159241)),(to_sfixed_a(-0.0006288793520070612)),(to_sfixed_a(-9.747594049258623e-06)),(to_sfixed_a(0.00013880044571124017)),(to_sfixed_a(-0.00014180003199726343)),(to_sfixed_a(-9.26469947444275e-05)),(to_sfixed_a(0.0003967138472944498)),(to_sfixed_a(-9.653793676989153e-05)),(to_sfixed_a(9.816499368753284e-05)),(to_sfixed_a(-0.0003086084616370499)),(to_sfixed_a(-0.00012564804637804627)),(to_sfixed_a(-0.03344043344259262)),(to_sfixed_a(0.10411006957292557)),(to_sfixed_a(0.09297806769609451)),(to_sfixed_a(-0.06677805632352829)),(to_sfixed_a(-0.08299556374549866)),(to_sfixed_a(0.09043069928884506)),(to_sfixed_a(0.11354232579469681)),(to_sfixed_a(-0.06390798091888428)),(to_sfixed_a(0.052523575723171234)),(to_sfixed_a(-0.00916997343301773)),(to_sfixed_a(-0.09819817543029785)),(to_sfixed_a(0.12798379361629486)),(to_sfixed_a(-0.04482415318489075)),(to_sfixed_a(0.0050591169856488705)),(to_sfixed_a(0.22728034853935242)),(to_sfixed_a(0.03496531769633293)),(to_sfixed_a(-0.0020113911014050245)),(to_sfixed_a(-0.004353562835603952)),(to_sfixed_a(-0.004845377989113331)),(to_sfixed_a(4.92435137857683e-05)),(to_sfixed_a(-2.650970964168664e-05)),(to_sfixed_a(-6.620831845793873e-05)),(to_sfixed_a(7.814901618985459e-05)),(to_sfixed_a(4.369279486127198e-05)),(to_sfixed_a(-0.00010303681483492255)),(to_sfixed_a(-0.0002793007006403059)),(to_sfixed_a(2.3306303774006665e-05)),(to_sfixed_a(-0.00015987013466656208)),(to_sfixed_a(0.00033686039387248456)),(to_sfixed_a(0.0002523345756344497)),(to_sfixed_a(8.056726801441982e-05)),(to_sfixed_a(-0.00014563542208634317)),(to_sfixed_a(-0.0003471329982858151)),(to_sfixed_a(0.16136832535266876)),(to_sfixed_a(-0.002431247616186738)),(to_sfixed_a(-0.0018418673425912857)),(to_sfixed_a(0.13112667202949524)),(to_sfixed_a(0.04132568836212158)),(to_sfixed_a(0.005854368209838867)),(to_sfixed_a(0.12309877574443817)),(to_sfixed_a(0.1308542639017105)),(to_sfixed_a(0.17040765285491943)),(to_sfixed_a(-0.0018053584499284625)),(to_sfixed_a(-0.0017827419796958566)),(to_sfixed_a(-0.00014787024701945484)),(to_sfixed_a(-0.00015325276763178408)),(to_sfixed_a(5.052704727859236e-05)),(to_sfixed_a(-4.935803008265793e-05)),(to_sfixed_a(-3.9758688217261806e-05)),(to_sfixed_a(-8.361334766959772e-05)),(to_sfixed_a(0.0002627871872391552)),(to_sfixed_a(9.07730373000959e-06)),(to_sfixed_a(0.00020342155767139047)),(to_sfixed_a(-7.353885303018615e-05)),(to_sfixed_a(-4.272404476068914e-05)),(to_sfixed_a(1.3904080333304591e-05)),(to_sfixed_a(-0.0001794749405235052)),(to_sfixed_a(0.0002461709373164922)),(to_sfixed_a(-0.0001285876496694982)),(to_sfixed_a(9.657142982177902e-06)),(to_sfixed_a(-3.253648173995316e-05)),(to_sfixed_a(-0.00023865712864790112)),(to_sfixed_a(4.434946458786726e-05)),(to_sfixed_a(0.00015080209414009005)),(to_sfixed_a(-1.8515058400225826e-05)),(to_sfixed_a(-0.00022780215658713132)),(to_sfixed_a(5.762487853644416e-05)),(to_sfixed_a(-2.5983126761275344e-05)),(to_sfixed_a(0.00024510722141712904)),(to_sfixed_a(0.00010587175347609445)),(to_sfixed_a(9.412258805241436e-06)),(to_sfixed_a(0.00022451516997534782)),(to_sfixed_a(-0.00016926367243286222)),(to_sfixed_a(-0.00022565570543520153)),(to_sfixed_a(0.00018235680181533098)),(to_sfixed_a(0.00012283245450817049)),(to_sfixed_a(-0.0002324153610970825)),(to_sfixed_a(-7.236383680719882e-06)),(to_sfixed_a(-2.2534857635037042e-05)));

    constant weight_n0_25 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(6.481730088125914e-05)),(to_sfixed_a(-1.702426561678294e-05)),(to_sfixed_a(0.0001217825774801895)),(to_sfixed_a(6.081046012695879e-05)),(to_sfixed_a(-0.0001071228543878533)),(to_sfixed_a(-0.00010655673395376652)),(to_sfixed_a(0.00034662947291508317)),(to_sfixed_a(-2.355523429287132e-05)),(to_sfixed_a(-0.0001529482105979696)),(to_sfixed_a(-0.0002549820637796074)),(to_sfixed_a(0.00020728471281472594)),(to_sfixed_a(-0.00011659295705612749)),(to_sfixed_a(0.00027737035998143256)),(to_sfixed_a(-0.00020460895029827952)),(to_sfixed_a(1.011350286717061e-05)),(to_sfixed_a(9.351280459668487e-05)),(to_sfixed_a(0.00028158153872936964)),(to_sfixed_a(9.36726646614261e-05)),(to_sfixed_a(-0.00013363589823711663)),(to_sfixed_a(-5.393719402491115e-05)),(to_sfixed_a(-5.7106746680801734e-05)),(to_sfixed_a(-0.00015331247413996607)),(to_sfixed_a(-0.00020342555944807827)),(to_sfixed_a(-0.00025480290059931576)),(to_sfixed_a(6.355164805427194e-05)),(to_sfixed_a(9.263669926440343e-05)),(to_sfixed_a(-0.00019458055612631142)),(to_sfixed_a(0.0002779875067062676)),(to_sfixed_a(-1.8160346371587366e-05)),(to_sfixed_a(9.056212002178654e-05)),(to_sfixed_a(-9.179586777463555e-05)),(to_sfixed_a(0.0002503844734746963)),(to_sfixed_a(0.00010923609079327434)),(to_sfixed_a(-9.660454088589177e-05)),(to_sfixed_a(0.0003584277583286166)),(to_sfixed_a(-0.00022188448929227889)),(to_sfixed_a(-0.0002748407714534551)),(to_sfixed_a(-7.901778008090332e-05)),(to_sfixed_a(-8.20362583908718e-06)),(to_sfixed_a(0.00010832941916305572)),(to_sfixed_a(-9.56634248723276e-05)),(to_sfixed_a(-9.217385377269238e-05)),(to_sfixed_a(0.00012293430336285383)),(to_sfixed_a(4.326838461565785e-05)),(to_sfixed_a(8.064101712079719e-05)),(to_sfixed_a(-1.3738466805079952e-05)),(to_sfixed_a(0.00014012174506206065)),(to_sfixed_a(-0.0002444240089971572)),(to_sfixed_a(-3.381001079105772e-05)),(to_sfixed_a(-4.4913576857652515e-06)),(to_sfixed_a(-0.0003229925350751728)),(to_sfixed_a(-1.8219684534415137e-06)),(to_sfixed_a(6.021195440553129e-05)),(to_sfixed_a(-5.432333182397997e-06)),(to_sfixed_a(-4.205599907436408e-05)),(to_sfixed_a(0.00011396635818528011)),(to_sfixed_a(1.2748840163112618e-05)),(to_sfixed_a(-2.1452307919389568e-05)),(to_sfixed_a(-9.792272612685338e-05)),(to_sfixed_a(8.873143815435469e-05)),(to_sfixed_a(4.221909330226481e-05)),(to_sfixed_a(0.00029017258202657104)),(to_sfixed_a(-0.00010620931425364688)),(to_sfixed_a(-2.153577770513948e-05)),(to_sfixed_a(3.18465317832306e-05)),(to_sfixed_a(-6.761230906704441e-05)),(to_sfixed_a(-0.00011456707579782233)),(to_sfixed_a(-0.00017043479601852596)),(to_sfixed_a(-1.9455506844678894e-05)),(to_sfixed_a(0.01178069319576025)),(to_sfixed_a(-0.00010487232793821022)),(to_sfixed_a(-9.847658657236025e-05)),(to_sfixed_a(-0.00020605666213668883)),(to_sfixed_a(9.13114272407256e-05)),(to_sfixed_a(-3.672864113468677e-05)),(to_sfixed_a(9.30443056859076e-05)),(to_sfixed_a(0.00010408461093902588)),(to_sfixed_a(-0.0001384080678690225)),(to_sfixed_a(-0.00014035002095624804)),(to_sfixed_a(-0.0003305410500615835)),(to_sfixed_a(8.318845357280225e-05)),(to_sfixed_a(1.6477979443152435e-05)),(to_sfixed_a(0.0001884610392153263)),(to_sfixed_a(-0.00016246939776465297)),(to_sfixed_a(0.00012911163503304124)),(to_sfixed_a(0.0001240437850356102)),(to_sfixed_a(4.4154607167001814e-05)),(to_sfixed_a(0.00016226543812081218)),(to_sfixed_a(-7.099750655470416e-05)),(to_sfixed_a(7.529697177233174e-05)),(to_sfixed_a(4.723609163193032e-05)),(to_sfixed_a(0.0001510617003077641)),(to_sfixed_a(-0.04907612502574921)),(to_sfixed_a(-0.00015256561164278537)),(to_sfixed_a(-0.055554408580064774)),(to_sfixed_a(0.0395675003528595)),(to_sfixed_a(0.020706651732325554)),(to_sfixed_a(0.04255449026823044)),(to_sfixed_a(-0.06924137473106384)),(to_sfixed_a(0.10660028457641602)),(to_sfixed_a(0.01238318346440792)),(to_sfixed_a(0.025175150483846664)),(to_sfixed_a(0.187956765294075)),(to_sfixed_a(-0.008066827431321144)),(to_sfixed_a(-0.017428221181035042)),(to_sfixed_a(-0.03512861952185631)),(to_sfixed_a(6.295468665484805e-06)),(to_sfixed_a(0.00014439398364629596)),(to_sfixed_a(0.0001297188427997753)),(to_sfixed_a(2.3050208255881444e-05)),(to_sfixed_a(-4.834179344470613e-05)),(to_sfixed_a(-0.00010512315202504396)),(to_sfixed_a(0.00022161929518915713)),(to_sfixed_a(3.686537456815131e-05)),(to_sfixed_a(-0.00025625480338931084)),(to_sfixed_a(-2.4499688151990995e-05)),(to_sfixed_a(-4.9678597861202434e-05)),(to_sfixed_a(-2.288991709065158e-05)),(to_sfixed_a(-0.0003745179274119437)),(to_sfixed_a(-0.0004349968221504241)),(to_sfixed_a(-0.047041866928339005)),(to_sfixed_a(-0.06890061497688293)),(to_sfixed_a(0.1010165885090828)),(to_sfixed_a(0.09436539560556412)),(to_sfixed_a(-0.06335185468196869)),(to_sfixed_a(-0.0992588922381401)),(to_sfixed_a(-0.11335070431232452)),(to_sfixed_a(0.29094359278678894)),(to_sfixed_a(0.2746698558330536)),(to_sfixed_a(0.044000159949064255)),(to_sfixed_a(0.04281828925013542)),(to_sfixed_a(0.002612969372421503)),(to_sfixed_a(0.005892554763704538)),(to_sfixed_a(0.01701723039150238)),(to_sfixed_a(-0.01983150653541088)),(to_sfixed_a(0.00019029852410312742)),(to_sfixed_a(-0.00011499405809445307)),(to_sfixed_a(0.00017393281450495124)),(to_sfixed_a(0.00012672935554292053)),(to_sfixed_a(1.6103953385027125e-05)),(to_sfixed_a(-2.6994257495971397e-07)),(to_sfixed_a(-6.694498006254435e-05)),(to_sfixed_a(4.2892046622000635e-05)),(to_sfixed_a(-4.156327122473158e-05)),(to_sfixed_a(0.0013212673366069794)),(to_sfixed_a(0.00894943717867136)),(to_sfixed_a(0.008842497132718563)),(to_sfixed_a(-0.1013462245464325)),(to_sfixed_a(0.07885760068893433)),(to_sfixed_a(0.054466575384140015)),(to_sfixed_a(0.09416806697845459)),(to_sfixed_a(-0.027116931974887848)),(to_sfixed_a(0.35222965478897095)),(to_sfixed_a(0.2687046229839325)),(to_sfixed_a(0.11219385266304016)),(to_sfixed_a(0.18542347848415375)),(to_sfixed_a(0.12759414315223694)),(to_sfixed_a(0.03588326647877693)),(to_sfixed_a(-0.33771753311157227)),(to_sfixed_a(-0.07897353917360306)),(to_sfixed_a(-0.09972058236598969)),(to_sfixed_a(0.03434407338500023)),(to_sfixed_a(-0.005286782048642635)),(to_sfixed_a(-0.04486212134361267)),(to_sfixed_a(-0.0007774014957249165)),(to_sfixed_a(0.0005297985626384616)),(to_sfixed_a(1.193736261484446e-05)),(to_sfixed_a(3.878560892189853e-05)),(to_sfixed_a(-6.827046308899298e-05)),(to_sfixed_a(0.0001322698954027146)),(to_sfixed_a(-3.155275771860033e-05)),(to_sfixed_a(0.00020139553816989064)),(to_sfixed_a(7.849370740586892e-05)),(to_sfixed_a(0.00964333675801754)),(to_sfixed_a(0.01738824136555195)),(to_sfixed_a(-0.08320740610361099)),(to_sfixed_a(-0.18554924428462982)),(to_sfixed_a(-0.017788611352443695)),(to_sfixed_a(0.40261873602867126)),(to_sfixed_a(0.0021314267069101334)),(to_sfixed_a(0.09904414415359497)),(to_sfixed_a(0.03700677305459976)),(to_sfixed_a(-0.06694943457841873)),(to_sfixed_a(-0.034974340349435806)),(to_sfixed_a(-0.11275185644626617)),(to_sfixed_a(-0.09768505394458771)),(to_sfixed_a(0.17382726073265076)),(to_sfixed_a(-0.04235992953181267)),(to_sfixed_a(-0.2963544726371765)),(to_sfixed_a(-0.14789479970932007)),(to_sfixed_a(-0.03525065630674362)),(to_sfixed_a(-0.05971597880125046)),(to_sfixed_a(0.0007056818576529622)),(to_sfixed_a(0.0024935004767030478)),(to_sfixed_a(0.0006307289004325867)),(to_sfixed_a(7.499897037632763e-05)),(to_sfixed_a(9.813778888201341e-05)),(to_sfixed_a(0.000278063933365047)),(to_sfixed_a(-6.888705684104934e-05)),(to_sfixed_a(-0.00013320428843144327)),(to_sfixed_a(-0.00016592913016211241)),(to_sfixed_a(-0.03049490600824356)),(to_sfixed_a(0.09100782871246338)),(to_sfixed_a(0.10776612162590027)),(to_sfixed_a(-0.07531342655420303)),(to_sfixed_a(-0.1015135869383812)),(to_sfixed_a(0.41625913977622986)),(to_sfixed_a(-0.025895236060023308)),(to_sfixed_a(0.10584563761949539)),(to_sfixed_a(-0.0009537743753753603)),(to_sfixed_a(0.023711541667580605)),(to_sfixed_a(-0.3162284195423126)),(to_sfixed_a(-0.2519983649253845)),(to_sfixed_a(-0.10552534461021423)),(to_sfixed_a(-0.1327953189611435)),(to_sfixed_a(-0.24691173434257507)),(to_sfixed_a(0.15536394715309143)),(to_sfixed_a(0.14911039173603058)),(to_sfixed_a(-0.14306262135505676)),(to_sfixed_a(0.2066895216703415)),(to_sfixed_a(-0.09213754534721375)),(to_sfixed_a(0.0012609409168362617)),(to_sfixed_a(-0.00014137769176159054)),(to_sfixed_a(-7.683794137847144e-06)),(to_sfixed_a(-0.00020650032092817128)),(to_sfixed_a(-0.000152253734995611)),(to_sfixed_a(-0.00017820931680034846)),(to_sfixed_a(0.00014646722411271185)),(to_sfixed_a(-0.04050035402178764)),(to_sfixed_a(-0.024248188361525536)),(to_sfixed_a(-0.04953707754611969)),(to_sfixed_a(0.2010350078344345)),(to_sfixed_a(0.26718252897262573)),(to_sfixed_a(-0.09727661311626434)),(to_sfixed_a(-0.1539340764284134)),(to_sfixed_a(-0.0892440676689148)),(to_sfixed_a(0.20954498648643494)),(to_sfixed_a(-0.07823588699102402)),(to_sfixed_a(0.15090495347976685)),(to_sfixed_a(-0.10553358495235443)),(to_sfixed_a(-0.19602905213832855)),(to_sfixed_a(0.17749130725860596)),(to_sfixed_a(-0.008589527569711208)),(to_sfixed_a(-0.007669689133763313)),(to_sfixed_a(-0.09789624810218811)),(to_sfixed_a(-0.12806260585784912)),(to_sfixed_a(0.0629841536283493)),(to_sfixed_a(-0.06078086793422699)),(to_sfixed_a(-0.07145026326179504)),(to_sfixed_a(-0.03839767351746559)),(to_sfixed_a(6.164731166791171e-05)),(to_sfixed_a(3.106147050857544e-05)),(to_sfixed_a(8.916595106711611e-05)),(to_sfixed_a(-8.776326285442337e-05)),(to_sfixed_a(-0.00016245349252130836)),(to_sfixed_a(8.79599028849043e-05)),(to_sfixed_a(0.0032743068877607584)),(to_sfixed_a(-0.0899762436747551)),(to_sfixed_a(-0.03580377995967865)),(to_sfixed_a(0.1068623885512352)),(to_sfixed_a(-0.018500206992030144)),(to_sfixed_a(0.059483036398887634)),(to_sfixed_a(-0.03709118813276291)),(to_sfixed_a(-0.5009806752204895)),(to_sfixed_a(0.02975388802587986)),(to_sfixed_a(-0.10527507215738297)),(to_sfixed_a(-0.2526892125606537)),(to_sfixed_a(-0.1641821265220642)),(to_sfixed_a(-0.38472944498062134)),(to_sfixed_a(-0.08919624984264374)),(to_sfixed_a(-0.006938298232853413)),(to_sfixed_a(0.057141322642564774)),(to_sfixed_a(0.1825791299343109)),(to_sfixed_a(-0.09064099937677383)),(to_sfixed_a(-0.2123435139656067)),(to_sfixed_a(-0.009446046315133572)),(to_sfixed_a(0.10584690421819687)),(to_sfixed_a(0.00012999045429751277)),(to_sfixed_a(6.716161442454904e-05)),(to_sfixed_a(3.192045141986455e-06)),(to_sfixed_a(-0.00010936854960164055)),(to_sfixed_a(-1.4885520613461267e-05)),(to_sfixed_a(-7.074631139403209e-05)),(to_sfixed_a(-0.0002618605794850737)),(to_sfixed_a(0.01770995371043682)),(to_sfixed_a(-0.020213458687067032)),(to_sfixed_a(0.1804145872592926)),(to_sfixed_a(0.07152252644300461)),(to_sfixed_a(0.12501420080661774)),(to_sfixed_a(0.2035377472639084)),(to_sfixed_a(0.10258619487285614)),(to_sfixed_a(0.06486961990594864)),(to_sfixed_a(0.004259680863469839)),(to_sfixed_a(0.16005957126617432)),(to_sfixed_a(0.22987061738967896)),(to_sfixed_a(-0.13076242804527283)),(to_sfixed_a(0.2592185139656067)),(to_sfixed_a(0.26686352491378784)),(to_sfixed_a(0.08533769845962524)),(to_sfixed_a(0.10640467703342438)),(to_sfixed_a(-0.10511854290962219)),(to_sfixed_a(-0.4157279133796692)),(to_sfixed_a(0.08883801102638245)),(to_sfixed_a(0.11679858714342117)),(to_sfixed_a(-0.07868749648332596)),(to_sfixed_a(0.014575762674212456)),(to_sfixed_a(0.00015258751227520406)),(to_sfixed_a(5.6351302191615105e-05)),(to_sfixed_a(0.0001625817531021312)),(to_sfixed_a(-2.4004519218578935e-05)),(to_sfixed_a(-3.735328937182203e-05)),(to_sfixed_a(0.009430735372006893)),(to_sfixed_a(-0.05017773061990738)),(to_sfixed_a(0.04326552897691727)),(to_sfixed_a(0.14421691000461578)),(to_sfixed_a(0.06846217811107635)),(to_sfixed_a(0.03677031397819519)),(to_sfixed_a(0.05826922133564949)),(to_sfixed_a(-0.04035560414195061)),(to_sfixed_a(-0.2454427182674408)),(to_sfixed_a(-0.3021167516708374)),(to_sfixed_a(0.2665664255619049)),(to_sfixed_a(0.3354712724685669)),(to_sfixed_a(-0.12699510157108307)),(to_sfixed_a(0.17921052873134613)),(to_sfixed_a(0.09354673326015472)),(to_sfixed_a(0.1004042774438858)),(to_sfixed_a(0.08044104278087616)),(to_sfixed_a(-0.07814282178878784)),(to_sfixed_a(0.08936727792024612)),(to_sfixed_a(-0.10038235783576965)),(to_sfixed_a(-0.063966765999794)),(to_sfixed_a(-0.03444501757621765)),(to_sfixed_a(-8.396083285333589e-05)),(to_sfixed_a(0.00013165133714210242)),(to_sfixed_a(0.0003263397957198322)),(to_sfixed_a(5.9123583923792467e-05)),(to_sfixed_a(0.000131231194245629)),(to_sfixed_a(0.0002556419640313834)),(to_sfixed_a(0.00012194879673188552)),(to_sfixed_a(0.046945635229349136)),(to_sfixed_a(0.01384552102535963)),(to_sfixed_a(-0.03369785100221634)),(to_sfixed_a(0.05377597361803055)),(to_sfixed_a(-0.13440071046352386)),(to_sfixed_a(-0.07867632061243057)),(to_sfixed_a(-0.36144930124282837)),(to_sfixed_a(-0.043395839631557465)),(to_sfixed_a(0.0728105902671814)),(to_sfixed_a(0.07799159735441208)),(to_sfixed_a(-0.01188606582581997)),(to_sfixed_a(-0.3914262056350708)),(to_sfixed_a(-0.21939001977443695)),(to_sfixed_a(0.1565730720758438)),(to_sfixed_a(0.026773856952786446)),(to_sfixed_a(-0.6497020721435547)),(to_sfixed_a(0.27744776010513306)),(to_sfixed_a(0.06923356652259827)),(to_sfixed_a(0.028325680643320084)),(to_sfixed_a(0.1110430657863617)),(to_sfixed_a(-0.07000677287578583)),(to_sfixed_a(8.673647971590981e-05)),(to_sfixed_a(-4.722916128230281e-05)),(to_sfixed_a(0.00015211047139018774)),(to_sfixed_a(-0.00023254513507708907)),(to_sfixed_a(-0.0002676461881492287)),(to_sfixed_a(0.00017791705613490194)),(to_sfixed_a(0.00014581199502572417)),(to_sfixed_a(-0.019934864714741707)),(to_sfixed_a(-0.23372885584831238)),(to_sfixed_a(-0.07560135424137115)),(to_sfixed_a(-0.11262017488479614)),(to_sfixed_a(0.05578869581222534)),(to_sfixed_a(0.12083417922258377)),(to_sfixed_a(-0.06756934523582458)),(to_sfixed_a(-0.2482217699289322)),(to_sfixed_a(-0.20973829925060272)),(to_sfixed_a(0.11933156847953796)),(to_sfixed_a(0.0038833252619951963)),(to_sfixed_a(-0.21221622824668884)),(to_sfixed_a(-0.17341011762619019)),(to_sfixed_a(-0.03687603771686554)),(to_sfixed_a(-0.13854719698429108)),(to_sfixed_a(-0.12637455761432648)),(to_sfixed_a(-0.10798342525959015)),(to_sfixed_a(0.3276788592338562)),(to_sfixed_a(-0.06971687078475952)),(to_sfixed_a(0.06565851718187332)),(to_sfixed_a(-0.058332644402980804)),(to_sfixed_a(0.0032776237931102514)),(to_sfixed_a(0.003670050296932459)),(to_sfixed_a(-4.945736691297498e-06)),(to_sfixed_a(9.948847582563758e-05)),(to_sfixed_a(-6.83802500134334e-05)),(to_sfixed_a(0.00033936946419999003)),(to_sfixed_a(7.924932288005948e-05)),(to_sfixed_a(0.0013447353849187493)),(to_sfixed_a(-0.004484530072659254)),(to_sfixed_a(-0.07964642345905304)),(to_sfixed_a(0.04224571958184242)),(to_sfixed_a(0.23702387511730194)),(to_sfixed_a(0.05395108088850975)),(to_sfixed_a(-0.10792452841997147)),(to_sfixed_a(0.016339214518666267)),(to_sfixed_a(0.05519535765051842)),(to_sfixed_a(-0.08731895685195923)),(to_sfixed_a(-0.13837741315364838)),(to_sfixed_a(-0.14365574717521667)),(to_sfixed_a(-0.22484368085861206)),(to_sfixed_a(0.052326492965221405)),(to_sfixed_a(0.05877260863780975)),(to_sfixed_a(0.022376764565706253)),(to_sfixed_a(0.12441986054182053)),(to_sfixed_a(0.033470138907432556)),(to_sfixed_a(-0.003713584505021572)),(to_sfixed_a(-0.05392961949110031)),(to_sfixed_a(0.060307055711746216)),(to_sfixed_a(9.677043999545276e-05)),(to_sfixed_a(0.00021325988927856088)),(to_sfixed_a(-0.00018762375111691654)),(to_sfixed_a(0.000153237851918675)),(to_sfixed_a(-3.196392208337784e-05)),(to_sfixed_a(-3.693102189572528e-05)),(to_sfixed_a(0.00011365484533598647)),(to_sfixed_a(0.09085220843553543)),(to_sfixed_a(-0.1009427011013031)),(to_sfixed_a(-0.1124543845653534)),(to_sfixed_a(-0.15669704973697662)),(to_sfixed_a(-0.017179150134325027)),(to_sfixed_a(-0.14169947803020477)),(to_sfixed_a(-0.13301725685596466)),(to_sfixed_a(0.13505809009075165)),(to_sfixed_a(0.08737882226705551)),(to_sfixed_a(-0.12606240808963776)),(to_sfixed_a(-0.03507613763213158)),(to_sfixed_a(0.0449606329202652)),(to_sfixed_a(-0.013765491545200348)),(to_sfixed_a(0.2513318955898285)),(to_sfixed_a(0.14139987528324127)),(to_sfixed_a(-0.16484686732292175)),(to_sfixed_a(-0.17095299065113068)),(to_sfixed_a(-0.01850154623389244)),(to_sfixed_a(-0.0023494940251111984)),(to_sfixed_a(-0.03883954510092735)),(to_sfixed_a(-0.1424645632505417)),(to_sfixed_a(-0.0002171318483306095)),(to_sfixed_a(0.00010275854583596811)),(to_sfixed_a(-6.713514449074864e-05)),(to_sfixed_a(-8.463399717584252e-05)),(to_sfixed_a(6.345628935378045e-05)),(to_sfixed_a(-9.96026792563498e-05)),(to_sfixed_a(-0.00014624829054810107)),(to_sfixed_a(-0.0722527876496315)),(to_sfixed_a(-0.03058692440390587)),(to_sfixed_a(0.0071885716170072556)),(to_sfixed_a(-0.06291595846414566)),(to_sfixed_a(-0.13626912236213684)),(to_sfixed_a(-0.20204785466194153)),(to_sfixed_a(-0.008662316016852856)),(to_sfixed_a(0.06769534200429916)),(to_sfixed_a(-0.03699927777051926)),(to_sfixed_a(-0.10160506516695023)),(to_sfixed_a(-0.02320645935833454)),(to_sfixed_a(0.1094498485326767)),(to_sfixed_a(-0.020137839019298553)),(to_sfixed_a(0.038854558020830154)),(to_sfixed_a(0.2774175703525543)),(to_sfixed_a(-0.09813079982995987)),(to_sfixed_a(-0.3569122552871704)),(to_sfixed_a(-0.28380125761032104)),(to_sfixed_a(-0.1497260481119156)),(to_sfixed_a(0.04509107396006584)),(to_sfixed_a(-0.10422723740339279)),(to_sfixed_a(0.0227203369140625)),(to_sfixed_a(-0.0002729912812355906)),(to_sfixed_a(-7.471340359188616e-05)),(to_sfixed_a(0.0002026393631240353)),(to_sfixed_a(6.786367885069922e-05)),(to_sfixed_a(-0.00016238028183579445)),(to_sfixed_a(-4.140000601182692e-05)),(to_sfixed_a(-0.06054847687482834)),(to_sfixed_a(-0.14637520909309387)),(to_sfixed_a(-0.03704570606350899)),(to_sfixed_a(-0.16939309239387512)),(to_sfixed_a(-0.050240982323884964)),(to_sfixed_a(0.03669861704111099)),(to_sfixed_a(-0.02264513447880745)),(to_sfixed_a(0.1018364429473877)),(to_sfixed_a(-0.19778920710086823)),(to_sfixed_a(-0.05523020029067993)),(to_sfixed_a(0.07742750644683838)),(to_sfixed_a(0.2905615568161011)),(to_sfixed_a(0.17379949986934662)),(to_sfixed_a(-0.0707581415772438)),(to_sfixed_a(0.023967161774635315)),(to_sfixed_a(0.030592331662774086)),(to_sfixed_a(-0.08421114832162857)),(to_sfixed_a(0.04978439584374428)),(to_sfixed_a(0.1771095246076584)),(to_sfixed_a(-0.036143675446510315)),(to_sfixed_a(0.00010636361548677087)),(to_sfixed_a(0.0001773252006387338)),(to_sfixed_a(7.65257136663422e-05)),(to_sfixed_a(-4.173427078058012e-05)),(to_sfixed_a(-0.00012709178554359823)),(to_sfixed_a(-0.0002723211655393243)),(to_sfixed_a(-3.539460522006266e-05)),(to_sfixed_a(0.016373496502637863)),(to_sfixed_a(-0.10810171067714691)),(to_sfixed_a(-0.1290992647409439)),(to_sfixed_a(-0.13162177801132202)),(to_sfixed_a(-0.04488399624824524)),(to_sfixed_a(-0.05431928113102913)),(to_sfixed_a(0.18971489369869232)),(to_sfixed_a(0.20876820385456085)),(to_sfixed_a(0.2505447566509247)),(to_sfixed_a(-0.001750312396325171)),(to_sfixed_a(-0.02120097726583481)),(to_sfixed_a(0.28544414043426514)),(to_sfixed_a(0.10937691479921341)),(to_sfixed_a(0.11888058483600616)),(to_sfixed_a(0.013105219230055809)),(to_sfixed_a(-0.16096222400665283)),(to_sfixed_a(-0.20659612119197845)),(to_sfixed_a(0.09865277260541916)),(to_sfixed_a(0.06801176816225052)),(to_sfixed_a(-0.053593385964632034)),(to_sfixed_a(-0.03781156614422798)),(to_sfixed_a(0.04003123939037323)),(to_sfixed_a(3.748894414457027e-06)),(to_sfixed_a(-0.0003862811718136072)),(to_sfixed_a(-0.00022765174799133092)),(to_sfixed_a(1.0194358765147626e-05)),(to_sfixed_a(-6.890415534144267e-05)),(to_sfixed_a(-5.19026507390663e-05)),(to_sfixed_a(0.05491182580590248)),(to_sfixed_a(0.002478851703926921)),(to_sfixed_a(0.0376843586564064)),(to_sfixed_a(-0.07154236733913422)),(to_sfixed_a(-0.09682805091142654)),(to_sfixed_a(0.1771346926689148)),(to_sfixed_a(-0.10147280246019363)),(to_sfixed_a(-0.10716277360916138)),(to_sfixed_a(-0.21762162446975708)),(to_sfixed_a(0.28223657608032227)),(to_sfixed_a(0.26457977294921875)),(to_sfixed_a(0.12070006877183914)),(to_sfixed_a(-0.1236153095960617)),(to_sfixed_a(0.06997868418693542)),(to_sfixed_a(0.024630574509501457)),(to_sfixed_a(-0.023227903991937637)),(to_sfixed_a(0.09786926954984665)),(to_sfixed_a(0.03264608234167099)),(to_sfixed_a(0.10124678164720535)),(to_sfixed_a(-0.0336284264922142)),(to_sfixed_a(-0.01837889477610588)),(to_sfixed_a(0.00010274702799506485)),(to_sfixed_a(-0.00013023102656006813)),(to_sfixed_a(-0.00011605180043261498)),(to_sfixed_a(8.363526285393164e-05)),(to_sfixed_a(4.9834747187560424e-05)),(to_sfixed_a(-0.00018919847207143903)),(to_sfixed_a(-0.00012481529847718775)),(to_sfixed_a(-5.7659693993628025e-05)),(to_sfixed_a(0.011843654327094555)),(to_sfixed_a(-0.013022266328334808)),(to_sfixed_a(0.17814910411834717)),(to_sfixed_a(-0.24794544279575348)),(to_sfixed_a(0.014093880541622639)),(to_sfixed_a(-0.25482237339019775)),(to_sfixed_a(-0.07880144566297531)),(to_sfixed_a(-0.029736673459410667)),(to_sfixed_a(0.133488267660141)),(to_sfixed_a(0.15857210755348206)),(to_sfixed_a(-0.02033485844731331)),(to_sfixed_a(-0.05061968043446541)),(to_sfixed_a(-0.17203927040100098)),(to_sfixed_a(-0.15354855358600616)),(to_sfixed_a(-0.14738573133945465)),(to_sfixed_a(0.29363295435905457)),(to_sfixed_a(0.2951367497444153)),(to_sfixed_a(-0.10024823248386383)),(to_sfixed_a(0.09357736259698868)),(to_sfixed_a(0.08449570089578629)),(to_sfixed_a(0.02205587364733219)),(to_sfixed_a(1.99086862266995e-05)),(to_sfixed_a(0.00012218549090903252)),(to_sfixed_a(-0.00013043786748312414)),(to_sfixed_a(-0.00010652787022991106)),(to_sfixed_a(0.00019621977116912603)),(to_sfixed_a(-0.00017059878155123442)),(to_sfixed_a(0.00012069379590684548)),(to_sfixed_a(-0.039379049092531204)),(to_sfixed_a(-0.00023377168690785766)),(to_sfixed_a(0.028409864753484726)),(to_sfixed_a(0.043952591717243195)),(to_sfixed_a(-0.22257673740386963)),(to_sfixed_a(-0.13066235184669495)),(to_sfixed_a(0.05781811475753784)),(to_sfixed_a(-0.12574510276317596)),(to_sfixed_a(-0.2242635041475296)),(to_sfixed_a(-0.10505618155002594)),(to_sfixed_a(0.05345749855041504)),(to_sfixed_a(0.01969820447266102)),(to_sfixed_a(-0.2550663352012634)),(to_sfixed_a(-0.26028332114219666)),(to_sfixed_a(-0.006713464390486479)),(to_sfixed_a(0.05438005551695824)),(to_sfixed_a(0.3569495677947998)),(to_sfixed_a(0.0872032567858696)),(to_sfixed_a(-0.01837342418730259)),(to_sfixed_a(0.0019573590252548456)),(to_sfixed_a(0.06898436695337296)),(to_sfixed_a(0.00014691893011331558)),(to_sfixed_a(5.32966478203889e-05)),(to_sfixed_a(-0.0002353949676034972)),(to_sfixed_a(-6.579815089935437e-05)),(to_sfixed_a(0.00048300213529728353)),(to_sfixed_a(-1.613403219380416e-05)),(to_sfixed_a(-4.7362689656438306e-05)),(to_sfixed_a(-0.0004896041937172413)),(to_sfixed_a(-0.20858760178089142)),(to_sfixed_a(-0.027991842478513718)),(to_sfixed_a(0.18294011056423187)),(to_sfixed_a(0.051506444811820984)),(to_sfixed_a(0.08022239804267883)),(to_sfixed_a(-0.2506335377693176)),(to_sfixed_a(0.037116486579179764)),(to_sfixed_a(-0.12007570266723633)),(to_sfixed_a(-0.028415633365511894)),(to_sfixed_a(0.1450517326593399)),(to_sfixed_a(0.14430108666419983)),(to_sfixed_a(0.007624495308846235)),(to_sfixed_a(0.2284950166940689)),(to_sfixed_a(-0.02426319196820259)),(to_sfixed_a(-0.12989947199821472)),(to_sfixed_a(0.1408388614654541)),(to_sfixed_a(0.03926623985171318)),(to_sfixed_a(0.10744170844554901)),(to_sfixed_a(-0.003284808248281479)),(to_sfixed_a(-0.00030749544384889305)),(to_sfixed_a(5.390749720390886e-06)),(to_sfixed_a(-3.541487603797577e-05)),(to_sfixed_a(-0.00024186729569919407)),(to_sfixed_a(3.712538455147296e-05)),(to_sfixed_a(-4.7974222979974e-05)),(to_sfixed_a(0.00019778904970735312)),(to_sfixed_a(-9.367180609842762e-05)),(to_sfixed_a(-0.0006346168229356408)),(to_sfixed_a(0.025417376309633255)),(to_sfixed_a(0.03811609372496605)),(to_sfixed_a(-0.11729917675256729)),(to_sfixed_a(0.20401063561439514)),(to_sfixed_a(0.009660017676651478)),(to_sfixed_a(0.002365912776440382)),(to_sfixed_a(0.10873643308877945)),(to_sfixed_a(-0.003168728668242693)),(to_sfixed_a(-0.14879584312438965)),(to_sfixed_a(-0.027363933622837067)),(to_sfixed_a(0.008354364894330502)),(to_sfixed_a(0.010013371706008911)),(to_sfixed_a(0.055015679448843)),(to_sfixed_a(-0.3077789843082428)),(to_sfixed_a(-0.1693570911884308)),(to_sfixed_a(0.10588094592094421)),(to_sfixed_a(-0.05274258926510811)),(to_sfixed_a(-0.010522674769163132)),(to_sfixed_a(-0.03781374171376228)),(to_sfixed_a(0.00037927814992144704)),(to_sfixed_a(-0.0001554020564071834)),(to_sfixed_a(-8.790374704403803e-05)),(to_sfixed_a(-0.00013453686551656574)),(to_sfixed_a(-2.152923661924433e-05)),(to_sfixed_a(8.129629350150935e-06)),(to_sfixed_a(-7.852757335058413e-06)),(to_sfixed_a(0.00015863921726122499)),(to_sfixed_a(-0.014852991327643394)),(to_sfixed_a(-0.036959901452064514)),(to_sfixed_a(-0.0637679472565651)),(to_sfixed_a(0.025220666080713272)),(to_sfixed_a(0.12628580629825592)),(to_sfixed_a(0.057026952505111694)),(to_sfixed_a(0.07702764868736267)),(to_sfixed_a(-0.08791375905275345)),(to_sfixed_a(0.1341012716293335)),(to_sfixed_a(0.1862115114927292)),(to_sfixed_a(0.19629140198230743)),(to_sfixed_a(0.20823590457439423)),(to_sfixed_a(-0.3278440535068512)),(to_sfixed_a(-0.4411047697067261)),(to_sfixed_a(-0.07957098633050919)),(to_sfixed_a(-0.09921662509441376)),(to_sfixed_a(0.010912693105638027)),(to_sfixed_a(-0.0034392857924103737)),(to_sfixed_a(-0.02029467560350895)),(to_sfixed_a(-0.005462808534502983)),(to_sfixed_a(-0.00017589567869435996)),(to_sfixed_a(-9.294271876569837e-05)),(to_sfixed_a(-6.949327507754788e-05)),(to_sfixed_a(-1.340791550319409e-05)),(to_sfixed_a(0.0001481941289966926)),(to_sfixed_a(-0.00021555136481765658)),(to_sfixed_a(-0.00018066058692056686)),(to_sfixed_a(-6.049407966202125e-05)),(to_sfixed_a(1.828516360546928e-05)),(to_sfixed_a(0.008593459613621235)),(to_sfixed_a(-0.036951128393411636)),(to_sfixed_a(-0.07570833712816238)),(to_sfixed_a(0.11468472331762314)),(to_sfixed_a(0.1937633901834488)),(to_sfixed_a(-0.16396929323673248)),(to_sfixed_a(-0.13571207225322723)),(to_sfixed_a(-0.03875313699245453)),(to_sfixed_a(-0.0042390841990709305)),(to_sfixed_a(0.20074260234832764)),(to_sfixed_a(0.0663466826081276)),(to_sfixed_a(0.22806331515312195)),(to_sfixed_a(0.054731957614421844)),(to_sfixed_a(0.01519792526960373)),(to_sfixed_a(-0.020305516198277473)),(to_sfixed_a(0.023116355761885643)),(to_sfixed_a(0.001754764816723764)),(to_sfixed_a(0.001166248694062233)),(to_sfixed_a(0.0009448391501791775)),(to_sfixed_a(-0.00019382305617909878)),(to_sfixed_a(-6.717376891174354e-06)),(to_sfixed_a(-0.00013764148752670735)),(to_sfixed_a(-1.3739946552959736e-05)),(to_sfixed_a(0.00019449419050943106)),(to_sfixed_a(0.00017499932437203825)),(to_sfixed_a(9.025770850712433e-06)),(to_sfixed_a(-0.00014051988546270877)),(to_sfixed_a(6.603146903216839e-05)),(to_sfixed_a(0.00015970636741258204)),(to_sfixed_a(0.00010230785846943036)),(to_sfixed_a(0.0003664195246528834)),(to_sfixed_a(0.0003608177066780627)),(to_sfixed_a(6.468498759204522e-05)),(to_sfixed_a(-0.03321106731891632)),(to_sfixed_a(0.0012837446993216872)),(to_sfixed_a(-0.00013506441609933972)),(to_sfixed_a(-0.022982725873589516)),(to_sfixed_a(-0.024330416694283485)),(to_sfixed_a(0.005543678533285856)),(to_sfixed_a(-0.025327341631054878)),(to_sfixed_a(-0.02755497395992279)),(to_sfixed_a(-0.021415522322058678)),(to_sfixed_a(0.016112925484776497)),(to_sfixed_a(0.006288770120590925)),(to_sfixed_a(2.0250581656000577e-05)),(to_sfixed_a(0.00012193135626148432)),(to_sfixed_a(-9.485867849434726e-06)),(to_sfixed_a(0.00014542228018399328)),(to_sfixed_a(-0.0002577135164756328)),(to_sfixed_a(3.860386277665384e-05)),(to_sfixed_a(-0.00046671798918396235)),(to_sfixed_a(4.7165412979666144e-05)),(to_sfixed_a(-6.123810453573242e-05)),(to_sfixed_a(-0.00014686601934954524)),(to_sfixed_a(-8.741358033148572e-05)),(to_sfixed_a(8.419894584221765e-05)),(to_sfixed_a(-0.0002685383951757103)),(to_sfixed_a(-1.796712604118511e-05)),(to_sfixed_a(0.00023607916955370456)),(to_sfixed_a(-8.900179636839312e-06)),(to_sfixed_a(0.00019571537268348038)),(to_sfixed_a(-0.00036632217234000564)),(to_sfixed_a(9.644345118431374e-05)),(to_sfixed_a(-6.994277646299452e-05)),(to_sfixed_a(-9.087020589504391e-05)),(to_sfixed_a(-7.932359585538507e-05)),(to_sfixed_a(4.932797673973255e-05)),(to_sfixed_a(0.00012528113438747823)),(to_sfixed_a(-3.9689737604931e-05)),(to_sfixed_a(-8.21022258605808e-05)),(to_sfixed_a(6.70798763167113e-05)),(to_sfixed_a(7.133685721782967e-05)),(to_sfixed_a(-9.245295223081484e-05)),(to_sfixed_a(-6.96421557222493e-05)),(to_sfixed_a(0.0002675170253496617)),(to_sfixed_a(7.020575867500156e-05)),(to_sfixed_a(6.796455272706226e-05)),(to_sfixed_a(6.48690402158536e-05)),(to_sfixed_a(-6.078995284042321e-05)));

    constant weight_n0_26 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(0.0001999454980250448)),(to_sfixed_a(-0.00022229670139495283)),(to_sfixed_a(-0.00013215177750680596)),(to_sfixed_a(-0.00010179099626839161)),(to_sfixed_a(-0.00010373707482358441)),(to_sfixed_a(-1.1174664905411191e-05)),(to_sfixed_a(6.836800457676873e-05)),(to_sfixed_a(-0.00020279437012504786)),(to_sfixed_a(0.00020548007159959525)),(to_sfixed_a(9.954452252713963e-05)),(to_sfixed_a(-0.00016073035658337176)),(to_sfixed_a(2.0402144400577527e-06)),(to_sfixed_a(0.00011049209570046514)),(to_sfixed_a(0.0001374871499137953)),(to_sfixed_a(-8.207632345147431e-05)),(to_sfixed_a(-0.00016864795179571956)),(to_sfixed_a(7.876416202634573e-05)),(to_sfixed_a(-0.00016836712893564254)),(to_sfixed_a(-2.077632598229684e-05)),(to_sfixed_a(-0.00011123427975689992)),(to_sfixed_a(0.00013156096974853426)),(to_sfixed_a(1.737101047183387e-05)),(to_sfixed_a(0.00012330693425610662)),(to_sfixed_a(1.582661298016319e-06)),(to_sfixed_a(-0.00030112903914414346)),(to_sfixed_a(0.0001519058714620769)),(to_sfixed_a(0.00019692226487677544)),(to_sfixed_a(0.00019663335115183145)),(to_sfixed_a(0.00016310364298988134)),(to_sfixed_a(-0.00013008575479034334)),(to_sfixed_a(0.0003465345362201333)),(to_sfixed_a(0.0001618098613107577)),(to_sfixed_a(-5.080207483842969e-05)),(to_sfixed_a(-0.00013096992915961891)),(to_sfixed_a(0.00012337979569565505)),(to_sfixed_a(-1.8518264823796926e-06)),(to_sfixed_a(0.00017332899733446538)),(to_sfixed_a(-2.2174863261170685e-05)),(to_sfixed_a(0.00011681269097607583)),(to_sfixed_a(-3.232111339457333e-05)),(to_sfixed_a(5.155791586730629e-05)),(to_sfixed_a(0.00019171787425875664)),(to_sfixed_a(0.00013142169336788356)),(to_sfixed_a(-6.633358134422451e-05)),(to_sfixed_a(-0.00018395049846731126)),(to_sfixed_a(-5.880348544451408e-05)),(to_sfixed_a(-3.3371114113833755e-05)),(to_sfixed_a(0.00019801418238785118)),(to_sfixed_a(-0.00020955209038220346)),(to_sfixed_a(-5.907118247705512e-05)),(to_sfixed_a(-0.00019589542353060097)),(to_sfixed_a(4.172475655650487e-06)),(to_sfixed_a(4.007343886769377e-05)),(to_sfixed_a(-0.00031244545243680477)),(to_sfixed_a(3.5941702662967145e-05)),(to_sfixed_a(-0.00028629080043174326)),(to_sfixed_a(-0.00010005972580984235)),(to_sfixed_a(-2.7470491659187246e-06)),(to_sfixed_a(5.8649155107559636e-05)),(to_sfixed_a(-1.41437021738966e-05)),(to_sfixed_a(-5.517981480807066e-05)),(to_sfixed_a(-0.00014928610471542925)),(to_sfixed_a(5.4112915677251294e-05)),(to_sfixed_a(-7.949866994749755e-05)),(to_sfixed_a(-0.00015233297017402947)),(to_sfixed_a(-6.461972225224599e-05)),(to_sfixed_a(0.00014814709720667452)),(to_sfixed_a(-0.0001079876528820023)),(to_sfixed_a(-0.0001843591162469238)),(to_sfixed_a(0.014828840270638466)),(to_sfixed_a(7.233544693008298e-06)),(to_sfixed_a(-0.00015121047908905894)),(to_sfixed_a(-0.00022302720753941685)),(to_sfixed_a(-0.0001398497261106968)),(to_sfixed_a(-6.86088387737982e-05)),(to_sfixed_a(-3.959799505537376e-05)),(to_sfixed_a(0.0003883911413140595)),(to_sfixed_a(-0.00017433414177503437)),(to_sfixed_a(9.777447121450678e-05)),(to_sfixed_a(4.070900831720792e-05)),(to_sfixed_a(-2.147096165572293e-05)),(to_sfixed_a(0.000344800588209182)),(to_sfixed_a(-2.4841150661814027e-05)),(to_sfixed_a(-0.00014550561900250614)),(to_sfixed_a(-0.00024114020925480872)),(to_sfixed_a(0.00021300952357705683)),(to_sfixed_a(-0.00015308837464544922)),(to_sfixed_a(4.347134381532669e-05)),(to_sfixed_a(0.00021433812798932195)),(to_sfixed_a(-1.255398728972068e-05)),(to_sfixed_a(-6.25109751126729e-05)),(to_sfixed_a(-0.0001710178330540657)),(to_sfixed_a(-0.09491025656461716)),(to_sfixed_a(-8.484803402097896e-05)),(to_sfixed_a(-0.10774505883455276)),(to_sfixed_a(-0.13004082441329956)),(to_sfixed_a(-0.10264207422733307)),(to_sfixed_a(0.05362618714570999)),(to_sfixed_a(-0.2295643538236618)),(to_sfixed_a(0.08067347854375839)),(to_sfixed_a(0.013684295117855072)),(to_sfixed_a(-0.018918510526418686)),(to_sfixed_a(-0.055290915071964264)),(to_sfixed_a(0.0005898966337554157)),(to_sfixed_a(-0.016031423583626747)),(to_sfixed_a(-0.032504040747880936)),(to_sfixed_a(-2.4359836970688775e-05)),(to_sfixed_a(-2.8143058443674818e-05)),(to_sfixed_a(-0.00016438961029052734)),(to_sfixed_a(-3.724830094142817e-05)),(to_sfixed_a(6.885408220114186e-05)),(to_sfixed_a(-9.128427336690947e-05)),(to_sfixed_a(-0.00010958842176478356)),(to_sfixed_a(-2.3774218789185397e-05)),(to_sfixed_a(3.0033883376745507e-05)),(to_sfixed_a(-8.10993296909146e-05)),(to_sfixed_a(6.786191079299897e-05)),(to_sfixed_a(-0.0001882726646726951)),(to_sfixed_a(1.2970163879799657e-05)),(to_sfixed_a(-0.081144317984581)),(to_sfixed_a(-0.06712384521961212)),(to_sfixed_a(-0.13972309231758118)),(to_sfixed_a(0.22017359733581543)),(to_sfixed_a(0.12751509249210358)),(to_sfixed_a(0.1600525975227356)),(to_sfixed_a(-0.021186262369155884)),(to_sfixed_a(-0.24167400598526)),(to_sfixed_a(-0.04442495480179787)),(to_sfixed_a(-0.03963949531316757)),(to_sfixed_a(0.03316574916243553)),(to_sfixed_a(0.08284135907888412)),(to_sfixed_a(0.05918530747294426)),(to_sfixed_a(-0.022655760869383812)),(to_sfixed_a(0.010903392918407917)),(to_sfixed_a(0.005441619083285332)),(to_sfixed_a(0.00023928094014991075)),(to_sfixed_a(-0.0011318885954096913)),(to_sfixed_a(0.00016673262871336192)),(to_sfixed_a(-0.00016743056767154485)),(to_sfixed_a(-2.622133251861669e-05)),(to_sfixed_a(-5.076098386780359e-05)),(to_sfixed_a(-8.485040598316118e-05)),(to_sfixed_a(7.286885374924168e-05)),(to_sfixed_a(0.00022433768026530743)),(to_sfixed_a(0.0004177675291430205)),(to_sfixed_a(-0.1089891865849495)),(to_sfixed_a(0.010399390943348408)),(to_sfixed_a(-0.13777552545070648)),(to_sfixed_a(-0.08414456993341446)),(to_sfixed_a(-0.012530442327260971)),(to_sfixed_a(-0.009706809185445309)),(to_sfixed_a(0.14430804550647736)),(to_sfixed_a(-0.25839847326278687)),(to_sfixed_a(-0.2818606197834015)),(to_sfixed_a(-0.04701683670282364)),(to_sfixed_a(0.1169019490480423)),(to_sfixed_a(0.2821023166179657)),(to_sfixed_a(0.047362469136714935)),(to_sfixed_a(-0.21454748511314392)),(to_sfixed_a(0.02371879294514656)),(to_sfixed_a(0.08786734938621521)),(to_sfixed_a(0.04097748175263405)),(to_sfixed_a(-0.0023618671111762524)),(to_sfixed_a(-0.0027912301011383533)),(to_sfixed_a(0.0017283294582739472)),(to_sfixed_a(-0.00018182216444984078)),(to_sfixed_a(-0.0003865792241413146)),(to_sfixed_a(0.0001775143318809569)),(to_sfixed_a(-2.9769631510134786e-05)),(to_sfixed_a(-0.00012777761730831116)),(to_sfixed_a(0.00014970476331654936)),(to_sfixed_a(0.00015069812070578337)),(to_sfixed_a(0.00012598661123774946)),(to_sfixed_a(-0.1060982197523117)),(to_sfixed_a(-0.021391484886407852)),(to_sfixed_a(-0.08476465195417404)),(to_sfixed_a(0.028864145278930664)),(to_sfixed_a(-0.08673494309186935)),(to_sfixed_a(-0.1764543503522873)),(to_sfixed_a(-0.14206181466579437)),(to_sfixed_a(-0.30997714400291443)),(to_sfixed_a(-0.07719191908836365)),(to_sfixed_a(-0.1112106591463089)),(to_sfixed_a(0.03415016457438469)),(to_sfixed_a(0.07656126469373703)),(to_sfixed_a(0.1547996997833252)),(to_sfixed_a(-0.06475851684808731)),(to_sfixed_a(-0.13331788778305054)),(to_sfixed_a(-0.14349424839019775)),(to_sfixed_a(-0.1347503811120987)),(to_sfixed_a(-0.038061290979385376)),(to_sfixed_a(-0.0011356966570019722)),(to_sfixed_a(0.008045501075685024)),(to_sfixed_a(0.008819442242383957)),(to_sfixed_a(0.004222115967422724)),(to_sfixed_a(-6.519390444736928e-05)),(to_sfixed_a(8.893606718629599e-05)),(to_sfixed_a(0.00013053149450570345)),(to_sfixed_a(2.9156597520341165e-05)),(to_sfixed_a(-0.00012436206452548504)),(to_sfixed_a(-2.7465270250104368e-05)),(to_sfixed_a(-0.127059668302536)),(to_sfixed_a(-0.07548502087593079)),(to_sfixed_a(0.005051517393440008)),(to_sfixed_a(-0.15177373588085175)),(to_sfixed_a(-0.2583131194114685)),(to_sfixed_a(-0.243482306599617)),(to_sfixed_a(-0.15256266295909882)),(to_sfixed_a(-0.15183711051940918)),(to_sfixed_a(-0.21688692271709442)),(to_sfixed_a(0.299199640750885)),(to_sfixed_a(0.22090604901313782)),(to_sfixed_a(0.19721436500549316)),(to_sfixed_a(-0.07058901339769363)),(to_sfixed_a(-0.19293776154518127)),(to_sfixed_a(-0.436632364988327)),(to_sfixed_a(0.11746641248464584)),(to_sfixed_a(0.10544264316558838)),(to_sfixed_a(0.09908223897218704)),(to_sfixed_a(0.14890863001346588)),(to_sfixed_a(0.06190814822912216)),(to_sfixed_a(0.004104952793568373)),(to_sfixed_a(0.00010149420268135145)),(to_sfixed_a(0.0003456884587649256)),(to_sfixed_a(-0.0003050978702958673)),(to_sfixed_a(0.00010043518705060706)),(to_sfixed_a(0.0002719504409469664)),(to_sfixed_a(8.952890493674204e-05)),(to_sfixed_a(-0.09413285553455353)),(to_sfixed_a(0.00433392496779561)),(to_sfixed_a(-0.21756069362163544)),(to_sfixed_a(-0.041430357843637466)),(to_sfixed_a(-0.16043652594089508)),(to_sfixed_a(-0.08817259967327118)),(to_sfixed_a(-0.09095655381679535)),(to_sfixed_a(-0.030561259016394615)),(to_sfixed_a(0.06829829514026642)),(to_sfixed_a(-0.005660122260451317)),(to_sfixed_a(0.4324294328689575)),(to_sfixed_a(0.2225203961133957)),(to_sfixed_a(0.4836733639240265)),(to_sfixed_a(0.12348436564207077)),(to_sfixed_a(0.022200562059879303)),(to_sfixed_a(0.0018446464091539383)),(to_sfixed_a(0.08198428899049759)),(to_sfixed_a(-0.1074950322508812)),(to_sfixed_a(-0.03167077898979187)),(to_sfixed_a(0.019231654703617096)),(to_sfixed_a(0.10116279870271683)),(to_sfixed_a(-0.012937294319272041)),(to_sfixed_a(-0.0001597085501998663)),(to_sfixed_a(-6.984721403568983e-05)),(to_sfixed_a(0.00018856636597774923)),(to_sfixed_a(0.00018640393682289869)),(to_sfixed_a(0.00011870837624883279)),(to_sfixed_a(0.00014414088218472898)),(to_sfixed_a(-0.00018002567230723798)),(to_sfixed_a(-0.07064497470855713)),(to_sfixed_a(-0.03159654885530472)),(to_sfixed_a(0.029300281777977943)),(to_sfixed_a(0.0774272158741951)),(to_sfixed_a(0.08454201370477676)),(to_sfixed_a(0.3515510559082031)),(to_sfixed_a(-0.10849560052156448)),(to_sfixed_a(-0.44712480902671814)),(to_sfixed_a(-0.08969613164663315)),(to_sfixed_a(0.04563292860984802)),(to_sfixed_a(0.023533668369054794)),(to_sfixed_a(-0.24402502179145813)),(to_sfixed_a(-0.13237939774990082)),(to_sfixed_a(0.022148428484797478)),(to_sfixed_a(0.03982856869697571)),(to_sfixed_a(-0.006428517866879702)),(to_sfixed_a(-0.0531497560441494)),(to_sfixed_a(-0.15976162254810333)),(to_sfixed_a(-0.09972239285707474)),(to_sfixed_a(-0.03576182574033737)),(to_sfixed_a(0.0002102471044054255)),(to_sfixed_a(0.00014060491230338812)),(to_sfixed_a(-4.1058036003960297e-05)),(to_sfixed_a(0.00012249231804162264)),(to_sfixed_a(-0.00017839013889897615)),(to_sfixed_a(3.259583536419086e-05)),(to_sfixed_a(9.571486771164928e-06)),(to_sfixed_a(-0.009751550853252411)),(to_sfixed_a(-0.11191723495721817)),(to_sfixed_a(0.21774832904338837)),(to_sfixed_a(0.19880273938179016)),(to_sfixed_a(0.11507372558116913)),(to_sfixed_a(0.1370915174484253)),(to_sfixed_a(0.19127145409584045)),(to_sfixed_a(-0.20800051093101501)),(to_sfixed_a(-0.15379726886749268)),(to_sfixed_a(0.07506772875785828)),(to_sfixed_a(-0.22242875397205353)),(to_sfixed_a(-0.0618339478969574)),(to_sfixed_a(-0.07674510776996613)),(to_sfixed_a(-0.17576690018177032)),(to_sfixed_a(0.014970654621720314)),(to_sfixed_a(-0.07455116510391235)),(to_sfixed_a(0.19552327692508698)),(to_sfixed_a(0.05485858768224716)),(to_sfixed_a(0.0748780146241188)),(to_sfixed_a(0.011719482019543648)),(to_sfixed_a(0.04708652198314667)),(to_sfixed_a(0.02699323184788227)),(to_sfixed_a(-1.6123489331221208e-05)),(to_sfixed_a(-7.333028861467028e-06)),(to_sfixed_a(0.0001630302722332999)),(to_sfixed_a(-4.17538067267742e-05)),(to_sfixed_a(-5.485772271640599e-05)),(to_sfixed_a(0.02596184052526951)),(to_sfixed_a(-0.09469860047101974)),(to_sfixed_a(0.07813311368227005)),(to_sfixed_a(0.11615375429391861)),(to_sfixed_a(-0.16578461229801178)),(to_sfixed_a(0.1008119136095047)),(to_sfixed_a(0.03874359652400017)),(to_sfixed_a(-0.07166512310504913)),(to_sfixed_a(0.08075111359357834)),(to_sfixed_a(-0.1655990034341812)),(to_sfixed_a(-0.2927384376525879)),(to_sfixed_a(-0.35161110758781433)),(to_sfixed_a(0.0931018516421318)),(to_sfixed_a(-0.03433145210146904)),(to_sfixed_a(0.15742763876914978)),(to_sfixed_a(0.22878144681453705)),(to_sfixed_a(0.22286787629127502)),(to_sfixed_a(0.20959211885929108)),(to_sfixed_a(-0.1430758833885193)),(to_sfixed_a(-0.046147461980581284)),(to_sfixed_a(-0.02049660123884678)),(to_sfixed_a(0.14350265264511108)),(to_sfixed_a(-5.5011638323776424e-05)),(to_sfixed_a(-1.5061940757732373e-05)),(to_sfixed_a(1.0421015758765861e-05)),(to_sfixed_a(0.00018098125292453915)),(to_sfixed_a(6.276479689404368e-05)),(to_sfixed_a(0.0003172942961100489)),(to_sfixed_a(-9.862964361673221e-05)),(to_sfixed_a(-0.12488076090812683)),(to_sfixed_a(-0.13206195831298828)),(to_sfixed_a(0.02680642530322075)),(to_sfixed_a(-0.09509023278951645)),(to_sfixed_a(0.012929975986480713)),(to_sfixed_a(0.07862875610589981)),(to_sfixed_a(-0.09897401928901672)),(to_sfixed_a(0.1588859260082245)),(to_sfixed_a(-0.049235470592975616)),(to_sfixed_a(0.023081479594111443)),(to_sfixed_a(-0.02913537248969078)),(to_sfixed_a(0.14598466455936432)),(to_sfixed_a(0.22517772018909454)),(to_sfixed_a(0.1880965381860733)),(to_sfixed_a(0.04173428937792778)),(to_sfixed_a(0.2801964581012726)),(to_sfixed_a(0.01611163094639778)),(to_sfixed_a(-0.05682048201560974)),(to_sfixed_a(-0.16136808693408966)),(to_sfixed_a(-0.09491368383169174)),(to_sfixed_a(-0.1572270393371582)),(to_sfixed_a(0.00011563376028789207)),(to_sfixed_a(5.388794306782074e-05)),(to_sfixed_a(-0.00014652828394901007)),(to_sfixed_a(-1.9881414118572138e-05)),(to_sfixed_a(8.259442984126508e-05)),(to_sfixed_a(-0.00015554149285890162)),(to_sfixed_a(-7.497600017813966e-05)),(to_sfixed_a(0.022317299619317055)),(to_sfixed_a(0.3273969888687134)),(to_sfixed_a(0.18056699633598328)),(to_sfixed_a(0.08318305760622025)),(to_sfixed_a(0.04522594064474106)),(to_sfixed_a(0.16121692955493927)),(to_sfixed_a(0.19208040833473206)),(to_sfixed_a(-0.035345617681741714)),(to_sfixed_a(-0.0017892895266413689)),(to_sfixed_a(0.006969154812395573)),(to_sfixed_a(0.001511596841737628)),(to_sfixed_a(-0.06535538285970688)),(to_sfixed_a(-0.03536643832921982)),(to_sfixed_a(0.2233155220746994)),(to_sfixed_a(0.08032961189746857)),(to_sfixed_a(0.0010339041473343968)),(to_sfixed_a(-0.10350719094276428)),(to_sfixed_a(-0.060153406113386154)),(to_sfixed_a(0.0065080029889941216)),(to_sfixed_a(-0.46872052550315857)),(to_sfixed_a(-0.12186112999916077)),(to_sfixed_a(-0.0018966678762808442)),(to_sfixed_a(-0.001408719806931913)),(to_sfixed_a(-0.00028292322531342506)),(to_sfixed_a(5.815719487145543e-05)),(to_sfixed_a(-0.00012417447578627616)),(to_sfixed_a(1.2277068890398368e-05)),(to_sfixed_a(5.946641522314167e-06)),(to_sfixed_a(-0.0009665390243753791)),(to_sfixed_a(0.18330830335617065)),(to_sfixed_a(0.10723206400871277)),(to_sfixed_a(0.3661469519138336)),(to_sfixed_a(0.23326586186885834)),(to_sfixed_a(0.32618391513824463)),(to_sfixed_a(-0.014298946596682072)),(to_sfixed_a(-0.22919495403766632)),(to_sfixed_a(-0.06699240207672119)),(to_sfixed_a(-0.07517488300800323)),(to_sfixed_a(0.09862668812274933)),(to_sfixed_a(-0.001480286824516952)),(to_sfixed_a(-0.136441171169281)),(to_sfixed_a(0.008653988130390644)),(to_sfixed_a(0.12136372923851013)),(to_sfixed_a(-0.367199569940567)),(to_sfixed_a(0.035550251603126526)),(to_sfixed_a(0.003629544284194708)),(to_sfixed_a(-0.10365710407495499)),(to_sfixed_a(-0.11677806079387665)),(to_sfixed_a(0.1285969614982605)),(to_sfixed_a(0.0003454801335465163)),(to_sfixed_a(-0.00013796590792480856)),(to_sfixed_a(-0.0002634157135616988)),(to_sfixed_a(1.2419231097737793e-05)),(to_sfixed_a(8.589446952100843e-05)),(to_sfixed_a(0.00015944741608109325)),(to_sfixed_a(0.00036449506296776235)),(to_sfixed_a(0.004586640279740095)),(to_sfixed_a(0.23573686182498932)),(to_sfixed_a(-0.08663021773099899)),(to_sfixed_a(-0.21798811852931976)),(to_sfixed_a(-0.26024505496025085)),(to_sfixed_a(-0.2847888767719269)),(to_sfixed_a(-0.2360571324825287)),(to_sfixed_a(-0.15101192891597748)),(to_sfixed_a(0.06849990785121918)),(to_sfixed_a(-0.09320139139890671)),(to_sfixed_a(-0.02524043805897236)),(to_sfixed_a(-0.009946668520569801)),(to_sfixed_a(0.18786263465881348)),(to_sfixed_a(0.18740692734718323)),(to_sfixed_a(-0.110118567943573)),(to_sfixed_a(-0.02587198279798031)),(to_sfixed_a(-0.031144632026553154)),(to_sfixed_a(-0.03176211565732956)),(to_sfixed_a(-0.12824350595474243)),(to_sfixed_a(-0.16886137425899506)),(to_sfixed_a(0.0035140197724103928)),(to_sfixed_a(-3.984183058491908e-05)),(to_sfixed_a(0.00020019944349769503)),(to_sfixed_a(5.535277887247503e-05)),(to_sfixed_a(0.0002162413438782096)),(to_sfixed_a(0.00024855972151272)),(to_sfixed_a(0.0004859589971601963)),(to_sfixed_a(0.004337793681770563)),(to_sfixed_a(-0.15075768530368805)),(to_sfixed_a(0.025719739496707916)),(to_sfixed_a(0.24250653386116028)),(to_sfixed_a(-0.16338174045085907)),(to_sfixed_a(-0.2611228823661804)),(to_sfixed_a(-0.24881665408611298)),(to_sfixed_a(-0.18850970268249512)),(to_sfixed_a(-0.17512862384319305)),(to_sfixed_a(0.10726180672645569)),(to_sfixed_a(-0.13475720584392548)),(to_sfixed_a(-0.004690317902714014)),(to_sfixed_a(0.023758476600050926)),(to_sfixed_a(-0.013089686632156372)),(to_sfixed_a(-0.10661100596189499)),(to_sfixed_a(0.17122972011566162)),(to_sfixed_a(-0.07016851007938385)),(to_sfixed_a(0.024406256154179573)),(to_sfixed_a(0.07313776016235352)),(to_sfixed_a(0.02705228701233864)),(to_sfixed_a(-0.013220248743891716)),(to_sfixed_a(-0.10006646066904068)),(to_sfixed_a(-0.00622875802218914)),(to_sfixed_a(9.995286382036284e-05)),(to_sfixed_a(0.00012417492689564824)),(to_sfixed_a(0.00020517231314443052)),(to_sfixed_a(-0.0001980488741537556)),(to_sfixed_a(0.003997665364295244)),(to_sfixed_a(0.00442122295498848)),(to_sfixed_a(0.09915030002593994)),(to_sfixed_a(-0.0889812633395195)),(to_sfixed_a(0.021309882402420044)),(to_sfixed_a(0.008161702193319798)),(to_sfixed_a(-0.1066085696220398)),(to_sfixed_a(-0.04604809358716011)),(to_sfixed_a(0.11790348589420319)),(to_sfixed_a(0.3559632897377014)),(to_sfixed_a(0.08465833961963654)),(to_sfixed_a(-0.13685502111911774)),(to_sfixed_a(-0.20382077991962433)),(to_sfixed_a(-0.001902321120724082)),(to_sfixed_a(-0.10709312558174133)),(to_sfixed_a(0.21431076526641846)),(to_sfixed_a(0.07693078368902206)),(to_sfixed_a(0.0629265084862709)),(to_sfixed_a(-0.05001169815659523)),(to_sfixed_a(0.008727619424462318)),(to_sfixed_a(-0.34683164954185486)),(to_sfixed_a(-0.008199821226298809)),(to_sfixed_a(7.769311923766509e-05)),(to_sfixed_a(-0.000177694033482112)),(to_sfixed_a(-4.7368281229864806e-05)),(to_sfixed_a(-3.8664449675707147e-05)),(to_sfixed_a(2.8952128559467383e-05)),(to_sfixed_a(-6.856438994873315e-05)),(to_sfixed_a(-0.0001252519286936149)),(to_sfixed_a(0.02069118060171604)),(to_sfixed_a(0.025588952004909515)),(to_sfixed_a(-0.057729922235012054)),(to_sfixed_a(-0.02237658016383648)),(to_sfixed_a(-0.0563451312482357)),(to_sfixed_a(0.012174446135759354)),(to_sfixed_a(0.06248760595917702)),(to_sfixed_a(0.0894070565700531)),(to_sfixed_a(0.1557747721672058)),(to_sfixed_a(0.022427869960665703)),(to_sfixed_a(-0.22817988693714142)),(to_sfixed_a(-0.05026736855506897)),(to_sfixed_a(0.1517612189054489)),(to_sfixed_a(0.15557441115379333)),(to_sfixed_a(0.09047327190637589)),(to_sfixed_a(0.09829280525445938)),(to_sfixed_a(0.18705107271671295)),(to_sfixed_a(-0.018230628222227097)),(to_sfixed_a(-0.14103642106056213)),(to_sfixed_a(-0.027890916913747787)),(to_sfixed_a(-0.15873242914676666)),(to_sfixed_a(-0.011685424484312534)),(to_sfixed_a(-0.00019105467072222382)),(to_sfixed_a(0.0003367984900251031)),(to_sfixed_a(-3.4411626984365284e-05)),(to_sfixed_a(-2.6583962608128786e-05)),(to_sfixed_a(0.00010392827243776992)),(to_sfixed_a(-4.2994095565518364e-05)),(to_sfixed_a(0.05822322517633438)),(to_sfixed_a(0.0018559382297098637)),(to_sfixed_a(0.03430197015404701)),(to_sfixed_a(-0.056634772568941116)),(to_sfixed_a(-0.2194392830133438)),(to_sfixed_a(-0.15706689655780792)),(to_sfixed_a(0.015141154639422894)),(to_sfixed_a(-0.16785350441932678)),(to_sfixed_a(-0.07448103278875351)),(to_sfixed_a(-0.023410916328430176)),(to_sfixed_a(0.048859670758247375)),(to_sfixed_a(-0.18598729372024536)),(to_sfixed_a(0.08806023001670837)),(to_sfixed_a(0.04766853526234627)),(to_sfixed_a(-0.10470198094844818)),(to_sfixed_a(0.0697711706161499)),(to_sfixed_a(0.026413489133119583)),(to_sfixed_a(-0.03594690561294556)),(to_sfixed_a(-0.21807153522968292)),(to_sfixed_a(0.11309892684221268)),(to_sfixed_a(0.14971014857292175)),(to_sfixed_a(-0.00018134419224224985)),(to_sfixed_a(-5.861179670318961e-05)),(to_sfixed_a(2.6295436327927746e-05)),(to_sfixed_a(-2.706883788050618e-05)),(to_sfixed_a(0.0003131599514745176)),(to_sfixed_a(-0.00018737409845925868)),(to_sfixed_a(-0.00011137279216200113)),(to_sfixed_a(0.0002632860851008445)),(to_sfixed_a(-0.02638028748333454)),(to_sfixed_a(-0.0388227216899395)),(to_sfixed_a(0.21920406818389893)),(to_sfixed_a(-0.14710019528865814)),(to_sfixed_a(0.05451153218746185)),(to_sfixed_a(-0.007509184535592794)),(to_sfixed_a(0.09937028586864471)),(to_sfixed_a(-0.3084775507450104)),(to_sfixed_a(-0.35399824380874634)),(to_sfixed_a(-0.007542680017650127)),(to_sfixed_a(-0.04163505509495735)),(to_sfixed_a(-0.21708889305591583)),(to_sfixed_a(0.06908073276281357)),(to_sfixed_a(0.3252154290676117)),(to_sfixed_a(0.3989408016204834)),(to_sfixed_a(-0.03704652562737465)),(to_sfixed_a(-0.016225257888436317)),(to_sfixed_a(0.2179899960756302)),(to_sfixed_a(-0.00876513309776783)),(to_sfixed_a(0.11214128136634827)),(to_sfixed_a(0.1173517182469368)),(to_sfixed_a(2.1315993308235193e-06)),(to_sfixed_a(0.00027311115991324186)),(to_sfixed_a(-0.00010206768638454378)),(to_sfixed_a(0.0004034604935441166)),(to_sfixed_a(0.0002631203969940543)),(to_sfixed_a(3.765002838918008e-05)),(to_sfixed_a(-0.00013540519285015762)),(to_sfixed_a(-0.09943125396966934)),(to_sfixed_a(0.0005460316897369921)),(to_sfixed_a(-0.06473939120769501)),(to_sfixed_a(0.13079188764095306)),(to_sfixed_a(0.005652955267578363)),(to_sfixed_a(-0.17242611944675446)),(to_sfixed_a(-0.11498362571001053)),(to_sfixed_a(0.11820201575756073)),(to_sfixed_a(-0.2526434659957886)),(to_sfixed_a(-0.10675276815891266)),(to_sfixed_a(-0.2311362475156784)),(to_sfixed_a(-0.08350574970245361)),(to_sfixed_a(0.009085959754884243)),(to_sfixed_a(-0.10855727642774582)),(to_sfixed_a(0.0382068045437336)),(to_sfixed_a(-0.04521070048213005)),(to_sfixed_a(0.11113139986991882)),(to_sfixed_a(0.05572567880153656)),(to_sfixed_a(0.08039742708206177)),(to_sfixed_a(0.0005765630048699677)),(to_sfixed_a(-0.0007014391594566405)),(to_sfixed_a(-0.00016553871682845056)),(to_sfixed_a(0.00021932840172667056)),(to_sfixed_a(0.0001869366387836635)),(to_sfixed_a(-7.037483737803996e-05)),(to_sfixed_a(0.0001922864030348137)),(to_sfixed_a(0.00017152576765511185)),(to_sfixed_a(0.00012606610835064203)),(to_sfixed_a(0.00026410570717416704)),(to_sfixed_a(0.13620778918266296)),(to_sfixed_a(-0.021158864721655846)),(to_sfixed_a(0.1739482581615448)),(to_sfixed_a(-0.02129165641963482)),(to_sfixed_a(-0.04998987168073654)),(to_sfixed_a(-0.11395248770713806)),(to_sfixed_a(-0.007806016597896814)),(to_sfixed_a(-0.14788614213466644)),(to_sfixed_a(0.02271977625787258)),(to_sfixed_a(0.12265745550394058)),(to_sfixed_a(-0.014196816831827164)),(to_sfixed_a(0.16250191628932953)),(to_sfixed_a(-0.014088338240981102)),(to_sfixed_a(-0.14979737997055054)),(to_sfixed_a(-0.08677711337804794)),(to_sfixed_a(-0.04616611823439598)),(to_sfixed_a(0.006764041725546122)),(to_sfixed_a(0.014962282031774521)),(to_sfixed_a(0.0018713034223765135)),(to_sfixed_a(4.208102109259926e-05)),(to_sfixed_a(0.00012817252718377858)),(to_sfixed_a(-0.00017022107203956693)),(to_sfixed_a(1.7206199117936194e-05)),(to_sfixed_a(-0.00022653907944913954)),(to_sfixed_a(0.00016061463975347579)),(to_sfixed_a(-6.641966319875792e-05)),(to_sfixed_a(-3.691560050356202e-05)),(to_sfixed_a(0.00032484170515090227)),(to_sfixed_a(-0.023594999685883522)),(to_sfixed_a(-0.006709227804094553)),(to_sfixed_a(-0.13363224267959595)),(to_sfixed_a(0.2966100871562958)),(to_sfixed_a(-0.12922155857086182)),(to_sfixed_a(-0.0293686855584383)),(to_sfixed_a(0.2090330421924591)),(to_sfixed_a(0.35407257080078125)),(to_sfixed_a(-0.05880540981888771)),(to_sfixed_a(0.31284549832344055)),(to_sfixed_a(0.3594013750553131)),(to_sfixed_a(-0.16700367629528046)),(to_sfixed_a(0.18269118666648865)),(to_sfixed_a(0.03609749674797058)),(to_sfixed_a(0.047747451812028885)),(to_sfixed_a(0.11408773809671402)),(to_sfixed_a(-0.014487173408269882)),(to_sfixed_a(0.005433632060885429)),(to_sfixed_a(-0.01640094630420208)),(to_sfixed_a(-0.0001077769193216227)),(to_sfixed_a(0.00022005525534041226)),(to_sfixed_a(-0.00046567796380259097)),(to_sfixed_a(-7.592904148623347e-05)),(to_sfixed_a(-0.00020543465507216752)),(to_sfixed_a(-2.7062515073339455e-05)),(to_sfixed_a(0.00018200979684479535)),(to_sfixed_a(9.114266140386462e-05)),(to_sfixed_a(0.004192369524389505)),(to_sfixed_a(0.014970765449106693)),(to_sfixed_a(0.01811199076473713)),(to_sfixed_a(0.10957560688257217)),(to_sfixed_a(0.07551544904708862)),(to_sfixed_a(0.09012763947248459)),(to_sfixed_a(-0.12701237201690674)),(to_sfixed_a(-0.16989187896251678)),(to_sfixed_a(0.07948721200227737)),(to_sfixed_a(0.10976031422615051)),(to_sfixed_a(-0.24972479045391083)),(to_sfixed_a(-0.07077895104885101)),(to_sfixed_a(0.0645999014377594)),(to_sfixed_a(0.09305418282747269)),(to_sfixed_a(0.05452831834554672)),(to_sfixed_a(0.005476146936416626)),(to_sfixed_a(0.009820366278290749)),(to_sfixed_a(0.009291119873523712)),(to_sfixed_a(0.0038732262328267097)),(to_sfixed_a(0.010354064404964447)),(to_sfixed_a(-0.0003087009536102414)),(to_sfixed_a(-3.7365192838478833e-05)),(to_sfixed_a(0.00011584463936742395)),(to_sfixed_a(4.876095408690162e-05)),(to_sfixed_a(0.00028808918432332575)),(to_sfixed_a(9.462352318223566e-05)),(to_sfixed_a(0.0001684449816821143)),(to_sfixed_a(-9.308612789027393e-05)),(to_sfixed_a(0.00020047256839461625)),(to_sfixed_a(0.056452978402376175)),(to_sfixed_a(0.010185039602220058)),(to_sfixed_a(0.05485956370830536)),(to_sfixed_a(0.08025768399238586)),(to_sfixed_a(-0.06553229689598083)),(to_sfixed_a(0.02360093966126442)),(to_sfixed_a(-0.001728271134197712)),(to_sfixed_a(-0.08403819054365158)),(to_sfixed_a(0.10911604762077332)),(to_sfixed_a(-0.03307730704545975)),(to_sfixed_a(0.01857222244143486)),(to_sfixed_a(-0.03382857143878937)),(to_sfixed_a(0.018479425460100174)),(to_sfixed_a(-0.010939007624983788)),(to_sfixed_a(0.07519850134849548)),(to_sfixed_a(0.0020163985900580883)),(to_sfixed_a(0.0009888972854241729)),(to_sfixed_a(0.004612988326698542)),(to_sfixed_a(0.005000225733965635)),(to_sfixed_a(2.049620889010839e-05)),(to_sfixed_a(0.0003105289360973984)),(to_sfixed_a(-0.0001727947237668559)),(to_sfixed_a(0.0001277576229767874)),(to_sfixed_a(-0.000574655132368207)),(to_sfixed_a(8.355608588317409e-05)),(to_sfixed_a(1.0324325558030978e-05)),(to_sfixed_a(0.0002977111143991351)),(to_sfixed_a(-0.00015168609388638288)),(to_sfixed_a(-0.0003322686825413257)),(to_sfixed_a(-8.168126078089699e-05)),(to_sfixed_a(5.9647423768183216e-05)),(to_sfixed_a(-0.0003068180230911821)),(to_sfixed_a(0.0003446244227234274)),(to_sfixed_a(-0.0005154649843461812)),(to_sfixed_a(0.014523802325129509)),(to_sfixed_a(0.0025804005563259125)),(to_sfixed_a(-0.009048416279256344)),(to_sfixed_a(-0.0680728405714035)),(to_sfixed_a(-0.018282683566212654)),(to_sfixed_a(0.05901346355676651)),(to_sfixed_a(-0.0068506523966789246)),(to_sfixed_a(-0.018937241286039352)),(to_sfixed_a(-0.008053101599216461)),(to_sfixed_a(-0.002284456044435501)),(to_sfixed_a(0.00011988640471827239)),(to_sfixed_a(-0.00018027921032626182)),(to_sfixed_a(7.153162005124614e-05)),(to_sfixed_a(0.0001505390537204221)),(to_sfixed_a(0.00015290976443793625)),(to_sfixed_a(-9.221512300428003e-05)),(to_sfixed_a(0.00011705682845786214)),(to_sfixed_a(8.151534530043136e-06)),(to_sfixed_a(-1.097480549105967e-06)),(to_sfixed_a(0.00015659125347156078)),(to_sfixed_a(-0.00014249637024477124)),(to_sfixed_a(2.005080932576675e-05)),(to_sfixed_a(-0.0004621956904884428)),(to_sfixed_a(3.3586631616344675e-05)),(to_sfixed_a(-9.351514017907903e-05)),(to_sfixed_a(0.00012233138841111213)),(to_sfixed_a(2.5297458705608733e-05)),(to_sfixed_a(0.0001782434992492199)),(to_sfixed_a(-8.272493869299069e-05)),(to_sfixed_a(-0.00014487230509985238)),(to_sfixed_a(-1.3695876077690627e-05)),(to_sfixed_a(-0.0001964818948181346)),(to_sfixed_a(4.801939576282166e-05)),(to_sfixed_a(0.0001205906446557492)),(to_sfixed_a(0.0002803892130032182)),(to_sfixed_a(0.00030314011382870376)),(to_sfixed_a(-9.322068945039064e-05)),(to_sfixed_a(2.5620422093197703e-05)),(to_sfixed_a(0.0002384654653724283)),(to_sfixed_a(0.00016558088827878237)),(to_sfixed_a(0.00016145705012604594)),(to_sfixed_a(-0.00015051322407089174)),(to_sfixed_a(2.7352163556315645e-07)),(to_sfixed_a(0.0002147688064724207)),(to_sfixed_a(8.943155080487486e-06)));

    constant weight_n0_27 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-0.0003715312632266432)),(to_sfixed_a(-3.229812500649132e-05)),(to_sfixed_a(-5.068421160103753e-05)),(to_sfixed_a(-0.0001566256396472454)),(to_sfixed_a(9.37236545723863e-05)),(to_sfixed_a(-5.5161483032861724e-05)),(to_sfixed_a(0.0002627712383400649)),(to_sfixed_a(0.00016081801732070744)),(to_sfixed_a(0.0002716754679568112)),(to_sfixed_a(3.615001332946122e-05)),(to_sfixed_a(-1.3659878277394455e-05)),(to_sfixed_a(-9.394837252330035e-05)),(to_sfixed_a(0.0001287570339627564)),(to_sfixed_a(-5.795116521767341e-06)),(to_sfixed_a(0.00012452028749976307)),(to_sfixed_a(5.262588820187375e-05)),(to_sfixed_a(-0.0001390130491927266)),(to_sfixed_a(-2.3851123842177913e-05)),(to_sfixed_a(-6.554967694683e-05)),(to_sfixed_a(-0.00015835986414458603)),(to_sfixed_a(8.36312465253286e-05)),(to_sfixed_a(-0.00036505243042483926)),(to_sfixed_a(-0.0003443902241997421)),(to_sfixed_a(-1.0132072020496707e-05)),(to_sfixed_a(-0.0001351832615910098)),(to_sfixed_a(0.00016827996296342462)),(to_sfixed_a(0.0001443272631149739)),(to_sfixed_a(-7.069305138429627e-05)),(to_sfixed_a(-0.00015600648475810885)),(to_sfixed_a(-0.00013201212277635932)),(to_sfixed_a(-0.000304327200865373)),(to_sfixed_a(-7.762706809444353e-05)),(to_sfixed_a(7.344350160565227e-05)),(to_sfixed_a(-2.197273715864867e-05)),(to_sfixed_a(0.00011930002801818773)),(to_sfixed_a(-0.00021468086924869567)),(to_sfixed_a(-4.4003947550663725e-05)),(to_sfixed_a(-1.2363722817099188e-05)),(to_sfixed_a(-0.0001035499808494933)),(to_sfixed_a(-6.710286834277213e-05)),(to_sfixed_a(4.210203769616783e-05)),(to_sfixed_a(9.516556019661948e-06)),(to_sfixed_a(-2.379886427661404e-05)),(to_sfixed_a(-0.00027832816704176366)),(to_sfixed_a(0.00033483904553577304)),(to_sfixed_a(-0.00015356106450781226)),(to_sfixed_a(8.20917630335316e-05)),(to_sfixed_a(0.00010964293323922902)),(to_sfixed_a(-3.820060010184534e-05)),(to_sfixed_a(2.5587198251741938e-05)),(to_sfixed_a(0.00010670450137695298)),(to_sfixed_a(-3.826840111287311e-05)),(to_sfixed_a(0.00014526555605698377)),(to_sfixed_a(-7.811879186192527e-05)),(to_sfixed_a(0.0001453006116207689)),(to_sfixed_a(5.33874481334351e-05)),(to_sfixed_a(0.000318297155899927)),(to_sfixed_a(1.232567592523992e-05)),(to_sfixed_a(-2.1392809230746934e-06)),(to_sfixed_a(-0.00028411211678758264)),(to_sfixed_a(9.267422683478799e-06)),(to_sfixed_a(-0.0002589701907709241)),(to_sfixed_a(-0.00021607373491860926)),(to_sfixed_a(3.586894308682531e-05)),(to_sfixed_a(-5.7950179325416684e-05)),(to_sfixed_a(-0.00018038311100099236)),(to_sfixed_a(-6.272788141359342e-06)),(to_sfixed_a(3.467746137175709e-05)),(to_sfixed_a(-3.043129800062161e-05)),(to_sfixed_a(-0.00519759813323617)),(to_sfixed_a(0.00019732363580260426)),(to_sfixed_a(-0.00022674018691759557)),(to_sfixed_a(3.093959094258025e-05)),(to_sfixed_a(-0.00020040132221765816)),(to_sfixed_a(-8.085336594376713e-05)),(to_sfixed_a(-5.9464480727910995e-05)),(to_sfixed_a(-1.50073020677155e-07)),(to_sfixed_a(-0.00011537947284523398)),(to_sfixed_a(-1.1905569408554584e-05)),(to_sfixed_a(9.957339352695271e-05)),(to_sfixed_a(-0.0003051319799851626)),(to_sfixed_a(8.537266694474965e-05)),(to_sfixed_a(1.3228361240180675e-05)),(to_sfixed_a(-9.992207196773961e-05)),(to_sfixed_a(-0.00010312467202311382)),(to_sfixed_a(-0.00015393183275591582)),(to_sfixed_a(-4.617136437445879e-05)),(to_sfixed_a(3.813610237557441e-05)),(to_sfixed_a(7.646351878065616e-05)),(to_sfixed_a(-0.00012452754890546203)),(to_sfixed_a(0.00018556129361968488)),(to_sfixed_a(0.00020304664212744683)),(to_sfixed_a(-0.02483232505619526)),(to_sfixed_a(1.016051828628406e-05)),(to_sfixed_a(-0.028354551643133163)),(to_sfixed_a(0.11724592000246048)),(to_sfixed_a(0.03695289418101311)),(to_sfixed_a(0.21596026420593262)),(to_sfixed_a(-0.03699073940515518)),(to_sfixed_a(-0.014515974558889866)),(to_sfixed_a(0.0043806042522192)),(to_sfixed_a(-0.1362762302160263)),(to_sfixed_a(-0.2545757293701172)),(to_sfixed_a(-0.14629799127578735)),(to_sfixed_a(-0.07517294585704803)),(to_sfixed_a(-0.15229982137680054)),(to_sfixed_a(3.0057854019105434e-06)),(to_sfixed_a(2.9512822948163375e-05)),(to_sfixed_a(-0.00012528212391771376)),(to_sfixed_a(-0.00012176825111964718)),(to_sfixed_a(-8.31338456919184e-06)),(to_sfixed_a(-0.00016597429930698127)),(to_sfixed_a(-0.0001667077449383214)),(to_sfixed_a(0.0002898239763453603)),(to_sfixed_a(9.693069296190515e-05)),(to_sfixed_a(5.4752737923990935e-05)),(to_sfixed_a(3.392100188648328e-05)),(to_sfixed_a(-6.554119318025187e-05)),(to_sfixed_a(0.0012103457702323794)),(to_sfixed_a(0.00946476124227047)),(to_sfixed_a(-0.05399880185723305)),(to_sfixed_a(-0.04257579520344734)),(to_sfixed_a(0.041535403579473495)),(to_sfixed_a(0.07335568219423294)),(to_sfixed_a(0.1789671778678894)),(to_sfixed_a(0.1568053960800171)),(to_sfixed_a(-0.017944658175110817)),(to_sfixed_a(-0.1596512347459793)),(to_sfixed_a(-0.08301202952861786)),(to_sfixed_a(-0.23459836840629578)),(to_sfixed_a(-0.07655995339155197)),(to_sfixed_a(-0.05622391030192375)),(to_sfixed_a(0.019421536475419998)),(to_sfixed_a(0.09326197952032089)),(to_sfixed_a(0.020189234986901283)),(to_sfixed_a(0.0005567301996052265)),(to_sfixed_a(0.0010185625869780779)),(to_sfixed_a(0.00010055821621790528)),(to_sfixed_a(4.577859363052994e-05)),(to_sfixed_a(-2.4336785031664476e-07)),(to_sfixed_a(4.5448661694535986e-05)),(to_sfixed_a(0.00025637634098529816)),(to_sfixed_a(4.677986362366937e-05)),(to_sfixed_a(-4.322168751969002e-05)),(to_sfixed_a(0.0003851673100143671)),(to_sfixed_a(0.017296066507697105)),(to_sfixed_a(0.00861979927867651)),(to_sfixed_a(0.05177207291126251)),(to_sfixed_a(0.21126991510391235)),(to_sfixed_a(0.036718692630529404)),(to_sfixed_a(0.004400052595883608)),(to_sfixed_a(0.1130969226360321)),(to_sfixed_a(0.42104822397232056)),(to_sfixed_a(-0.17363251745700836)),(to_sfixed_a(-0.22827701270580292)),(to_sfixed_a(-0.392882376909256)),(to_sfixed_a(-0.16099227964878082)),(to_sfixed_a(-0.11683578789234161)),(to_sfixed_a(-0.15860433876514435)),(to_sfixed_a(0.19339169561862946)),(to_sfixed_a(0.07258350402116776)),(to_sfixed_a(-0.07785731554031372)),(to_sfixed_a(0.0034463920164853334)),(to_sfixed_a(-0.11029475182294846)),(to_sfixed_a(0.003134608268737793)),(to_sfixed_a(0.0006565131479874253)),(to_sfixed_a(0.00011424160038586706)),(to_sfixed_a(9.083569239010103e-06)),(to_sfixed_a(-0.00012662950030062348)),(to_sfixed_a(2.98063168884255e-05)),(to_sfixed_a(3.7062662158859894e-05)),(to_sfixed_a(5.36905208718963e-05)),(to_sfixed_a(-7.399891183013096e-05)),(to_sfixed_a(0.014936254359781742)),(to_sfixed_a(-0.00010247601312585175)),(to_sfixed_a(-0.04309656471014023)),(to_sfixed_a(-0.03616369143128395)),(to_sfixed_a(-0.009654190391302109)),(to_sfixed_a(0.37321141362190247)),(to_sfixed_a(0.1783078908920288)),(to_sfixed_a(0.21339815855026245)),(to_sfixed_a(0.012014547362923622)),(to_sfixed_a(0.04009551927447319)),(to_sfixed_a(0.3404722511768341)),(to_sfixed_a(0.025578157976269722)),(to_sfixed_a(-0.1574067771434784)),(to_sfixed_a(-0.14384476840496063)),(to_sfixed_a(-0.07454836368560791)),(to_sfixed_a(-0.22058042883872986)),(to_sfixed_a(-0.01252590212970972)),(to_sfixed_a(-0.023754460737109184)),(to_sfixed_a(0.0021679287310689688)),(to_sfixed_a(-0.0033757651690393686)),(to_sfixed_a(-0.007034515030682087)),(to_sfixed_a(-0.003073285333812237)),(to_sfixed_a(2.3673726900597103e-05)),(to_sfixed_a(4.9949267122428864e-05)),(to_sfixed_a(-0.0003478078870102763)),(to_sfixed_a(0.00011588061170186847)),(to_sfixed_a(1.683695700194221e-05)),(to_sfixed_a(-8.760942000662908e-05)),(to_sfixed_a(-0.03645534813404083)),(to_sfixed_a(-0.1951514631509781)),(to_sfixed_a(-0.04956609010696411)),(to_sfixed_a(0.040935032069683075)),(to_sfixed_a(0.05583738163113594)),(to_sfixed_a(-0.09353751689195633)),(to_sfixed_a(-0.07906737923622131)),(to_sfixed_a(0.01169128343462944)),(to_sfixed_a(0.1744200885295868)),(to_sfixed_a(0.06756298243999481)),(to_sfixed_a(0.15347608923912048)),(to_sfixed_a(0.014237552881240845)),(to_sfixed_a(-0.2380598783493042)),(to_sfixed_a(0.1048530787229538)),(to_sfixed_a(0.04781375080347061)),(to_sfixed_a(-0.2520885765552521)),(to_sfixed_a(-0.10575734078884125)),(to_sfixed_a(-0.16371408104896545)),(to_sfixed_a(0.07637479901313782)),(to_sfixed_a(-0.0702815130352974)),(to_sfixed_a(-0.004504816606640816)),(to_sfixed_a(0.0002469312457833439)),(to_sfixed_a(0.00032675464171916246)),(to_sfixed_a(2.1104862753418274e-05)),(to_sfixed_a(-4.120559970033355e-05)),(to_sfixed_a(0.00021310789452400059)),(to_sfixed_a(4.401279511512257e-05)),(to_sfixed_a(-0.04126005619764328)),(to_sfixed_a(0.04186633601784706)),(to_sfixed_a(-0.06939026713371277)),(to_sfixed_a(0.04969261214137077)),(to_sfixed_a(-0.176022469997406)),(to_sfixed_a(0.2044084519147873)),(to_sfixed_a(-0.06473451852798462)),(to_sfixed_a(0.30341529846191406)),(to_sfixed_a(0.3927290141582489)),(to_sfixed_a(0.0675075501203537)),(to_sfixed_a(-0.06285962462425232)),(to_sfixed_a(0.14072328805923462)),(to_sfixed_a(-0.19770236313343048)),(to_sfixed_a(0.07960910350084305)),(to_sfixed_a(-0.039760034531354904)),(to_sfixed_a(-0.16067035496234894)),(to_sfixed_a(0.11034879088401794)),(to_sfixed_a(-0.1436391919851303)),(to_sfixed_a(-0.015124850906431675)),(to_sfixed_a(-0.12128896266222)),(to_sfixed_a(-0.2425392121076584)),(to_sfixed_a(0.02191823162138462)),(to_sfixed_a(-9.669276187196374e-05)),(to_sfixed_a(8.27152980491519e-05)),(to_sfixed_a(3.6727054975926876e-05)),(to_sfixed_a(0.0002090998023049906)),(to_sfixed_a(-3.488629954517819e-05)),(to_sfixed_a(-0.0003716387436725199)),(to_sfixed_a(0.0004408147360663861)),(to_sfixed_a(-0.1758815348148346)),(to_sfixed_a(-0.08521164208650589)),(to_sfixed_a(-0.13786816596984863)),(to_sfixed_a(-0.05902669206261635)),(to_sfixed_a(0.038113147020339966)),(to_sfixed_a(0.09445738792419434)),(to_sfixed_a(-0.14847052097320557)),(to_sfixed_a(0.11012321710586548)),(to_sfixed_a(-0.22472162544727325)),(to_sfixed_a(-0.4298388957977295)),(to_sfixed_a(-0.056520555168390274)),(to_sfixed_a(-0.0761164203286171)),(to_sfixed_a(0.3964460492134094)),(to_sfixed_a(0.1472586691379547)),(to_sfixed_a(-0.11174550652503967)),(to_sfixed_a(0.12865124642848969)),(to_sfixed_a(0.23617368936538696)),(to_sfixed_a(0.05416790395975113)),(to_sfixed_a(0.09597564488649368)),(to_sfixed_a(-0.23580391705036163)),(to_sfixed_a(3.57016506313812e-05)),(to_sfixed_a(-7.116964843589813e-05)),(to_sfixed_a(-1.0514725545363035e-05)),(to_sfixed_a(-0.0001503731618868187)),(to_sfixed_a(-1.3167565157345962e-05)),(to_sfixed_a(-7.450700650224462e-05)),(to_sfixed_a(0.0002986482286360115)),(to_sfixed_a(-0.0043726214207708836)),(to_sfixed_a(-0.028375187888741493)),(to_sfixed_a(0.3346134424209595)),(to_sfixed_a(0.031390585005283356)),(to_sfixed_a(-0.02892826870083809)),(to_sfixed_a(0.05652472376823425)),(to_sfixed_a(0.03550659865140915)),(to_sfixed_a(0.2665156424045563)),(to_sfixed_a(0.021546822041273117)),(to_sfixed_a(0.029633106663823128)),(to_sfixed_a(-0.4229170083999634)),(to_sfixed_a(-0.22807416319847107)),(to_sfixed_a(0.22931644320487976)),(to_sfixed_a(0.2011261284351349)),(to_sfixed_a(-0.1075923964381218)),(to_sfixed_a(0.189261332154274)),(to_sfixed_a(0.1293249875307083)),(to_sfixed_a(-0.07826840132474899)),(to_sfixed_a(0.10892773419618607)),(to_sfixed_a(0.11466307193040848)),(to_sfixed_a(-0.12776429951190948)),(to_sfixed_a(-0.06904581189155579)),(to_sfixed_a(-3.197156183887273e-05)),(to_sfixed_a(-4.463069490157068e-05)),(to_sfixed_a(0.0002870875468943268)),(to_sfixed_a(-7.422660564770922e-05)),(to_sfixed_a(-8.536655514035374e-05)),(to_sfixed_a(0.0033534064423292875)),(to_sfixed_a(-0.02503337524831295)),(to_sfixed_a(0.03306398540735245)),(to_sfixed_a(0.12677474319934845)),(to_sfixed_a(0.07632333040237427)),(to_sfixed_a(-0.026870466768741608)),(to_sfixed_a(-0.08408217132091522)),(to_sfixed_a(0.0535733737051487)),(to_sfixed_a(0.22647228837013245)),(to_sfixed_a(0.2315826714038849)),(to_sfixed_a(-0.04569973051548004)),(to_sfixed_a(-0.13463638722896576)),(to_sfixed_a(0.00040401535807177424)),(to_sfixed_a(0.27214792370796204)),(to_sfixed_a(0.0070692868903279305)),(to_sfixed_a(-0.09871247410774231)),(to_sfixed_a(-0.07768667489290237)),(to_sfixed_a(-0.2696380913257599)),(to_sfixed_a(-0.1261039674282074)),(to_sfixed_a(-0.05965534970164299)),(to_sfixed_a(0.02982393279671669)),(to_sfixed_a(-0.008330662734806538)),(to_sfixed_a(8.417768549406901e-05)),(to_sfixed_a(7.582468970213085e-05)),(to_sfixed_a(-0.00017569790361449122)),(to_sfixed_a(-0.0002954126102849841)),(to_sfixed_a(-4.2721826503111515e-06)),(to_sfixed_a(4.0584804082755e-05)),(to_sfixed_a(-0.0001237882097484544)),(to_sfixed_a(0.021275321021676064)),(to_sfixed_a(0.021339602768421173)),(to_sfixed_a(-0.07388332486152649)),(to_sfixed_a(0.13130323588848114)),(to_sfixed_a(0.0036733639426529408)),(to_sfixed_a(-0.06568686664104462)),(to_sfixed_a(-0.0036171735264360905)),(to_sfixed_a(0.2979426980018616)),(to_sfixed_a(0.2771085798740387)),(to_sfixed_a(0.0740019902586937)),(to_sfixed_a(-0.20060376822948456)),(to_sfixed_a(-0.011748969554901123)),(to_sfixed_a(-0.05484785512089729)),(to_sfixed_a(0.06477303802967072)),(to_sfixed_a(0.1685740351676941)),(to_sfixed_a(-0.05640004575252533)),(to_sfixed_a(-0.10197586566209793)),(to_sfixed_a(0.021399805322289467)),(to_sfixed_a(-0.05346447974443436)),(to_sfixed_a(0.10730761289596558)),(to_sfixed_a(0.10862520337104797)),(to_sfixed_a(-0.00015866140893194824)),(to_sfixed_a(0.0003978683380410075)),(to_sfixed_a(-2.342289917578455e-05)),(to_sfixed_a(0.0004149322339799255)),(to_sfixed_a(9.637139737606049e-05)),(to_sfixed_a(0.00013645041326526552)),(to_sfixed_a(-0.00023826188407838345)),(to_sfixed_a(-0.048165060579776764)),(to_sfixed_a(-0.2554265856742859)),(to_sfixed_a(-0.00880427472293377)),(to_sfixed_a(-0.11439240723848343)),(to_sfixed_a(0.02852410078048706)),(to_sfixed_a(-0.023533856496214867)),(to_sfixed_a(0.03756289929151535)),(to_sfixed_a(0.07558088004589081)),(to_sfixed_a(0.05579029396176338)),(to_sfixed_a(-0.21848513185977936)),(to_sfixed_a(-0.3767874836921692)),(to_sfixed_a(-0.10355217009782791)),(to_sfixed_a(-0.025626735761761665)),(to_sfixed_a(0.045225705951452255)),(to_sfixed_a(0.07890085875988007)),(to_sfixed_a(-0.03482525795698166)),(to_sfixed_a(0.10650691390037537)),(to_sfixed_a(-0.040231578052043915)),(to_sfixed_a(-0.11603306233882904)),(to_sfixed_a(0.020578483119606972)),(to_sfixed_a(-0.03319305181503296)),(to_sfixed_a(-0.002254420891404152)),(to_sfixed_a(-0.00192346575204283)),(to_sfixed_a(-4.620613617589697e-05)),(to_sfixed_a(-2.8727041353704408e-05)),(to_sfixed_a(0.00026041228557005525)),(to_sfixed_a(0.00013365925406105816)),(to_sfixed_a(-0.00017079275858122855)),(to_sfixed_a(-0.00042933336226269603)),(to_sfixed_a(0.1085655689239502)),(to_sfixed_a(0.07206621021032333)),(to_sfixed_a(0.04509399086236954)),(to_sfixed_a(0.11605090647935867)),(to_sfixed_a(-0.0350128710269928)),(to_sfixed_a(0.07114572077989578)),(to_sfixed_a(-0.07684914767742157)),(to_sfixed_a(0.13604101538658142)),(to_sfixed_a(-0.16281968355178833)),(to_sfixed_a(-0.21864035725593567)),(to_sfixed_a(-0.04722738638520241)),(to_sfixed_a(-0.04328997805714607)),(to_sfixed_a(0.06899438053369522)),(to_sfixed_a(0.09226100891828537)),(to_sfixed_a(-0.09354854375123978)),(to_sfixed_a(-0.09486372023820877)),(to_sfixed_a(0.07791649550199509)),(to_sfixed_a(-0.052977390587329865)),(to_sfixed_a(0.004645559936761856)),(to_sfixed_a(-0.025904707610607147)),(to_sfixed_a(-0.00015994880232028663)),(to_sfixed_a(0.0003163487708661705)),(to_sfixed_a(0.00021122259204275906)),(to_sfixed_a(-4.506632831180468e-05)),(to_sfixed_a(-0.0001423972862539813)),(to_sfixed_a(-8.91413219505921e-05)),(to_sfixed_a(-0.00017419428331777453)),(to_sfixed_a(0.04004860296845436)),(to_sfixed_a(0.12898345291614532)),(to_sfixed_a(0.05470946058630943)),(to_sfixed_a(0.10838139802217484)),(to_sfixed_a(0.20803984999656677)),(to_sfixed_a(-0.0557120181620121)),(to_sfixed_a(0.2530227303504944)),(to_sfixed_a(0.0972718670964241)),(to_sfixed_a(-0.001424842164851725)),(to_sfixed_a(-0.055153582245111465)),(to_sfixed_a(-0.14638358354568481)),(to_sfixed_a(0.10091271251440048)),(to_sfixed_a(0.029280945658683777)),(to_sfixed_a(0.19721312820911407)),(to_sfixed_a(0.044272102415561676)),(to_sfixed_a(-0.17333407700061798)),(to_sfixed_a(0.5874295830726624)),(to_sfixed_a(0.31783419847488403)),(to_sfixed_a(-0.05296645313501358)),(to_sfixed_a(-0.029295045882463455)),(to_sfixed_a(-0.0075354790315032005)),(to_sfixed_a(9.762057743500918e-05)),(to_sfixed_a(0.00017029505397658795)),(to_sfixed_a(-9.927639621309936e-05)),(to_sfixed_a(-0.0001387698284815997)),(to_sfixed_a(7.683602598262951e-05)),(to_sfixed_a(-0.0001060248541762121)),(to_sfixed_a(-0.0002314277517143637)),(to_sfixed_a(-0.051957543939352036)),(to_sfixed_a(-0.12213905900716782)),(to_sfixed_a(-0.13351298868656158)),(to_sfixed_a(-0.16084034740924835)),(to_sfixed_a(0.012764752842485905)),(to_sfixed_a(0.08864009380340576)),(to_sfixed_a(0.0234213937073946)),(to_sfixed_a(0.29075542092323303)),(to_sfixed_a(0.3454875349998474)),(to_sfixed_a(-0.06430104374885559)),(to_sfixed_a(0.08520655333995819)),(to_sfixed_a(0.0671209841966629)),(to_sfixed_a(-0.16076132655143738)),(to_sfixed_a(-0.07444463670253754)),(to_sfixed_a(-0.131795734167099)),(to_sfixed_a(-0.06536266952753067)),(to_sfixed_a(0.14544054865837097)),(to_sfixed_a(0.20718416571617126)),(to_sfixed_a(-0.09402325749397278)),(to_sfixed_a(0.0023002547677606344)),(to_sfixed_a(-0.018112264573574066)),(to_sfixed_a(-0.00613879319280386)),(to_sfixed_a(4.0697454096516594e-05)),(to_sfixed_a(3.1852068786974996e-05)),(to_sfixed_a(3.288468360551633e-05)),(to_sfixed_a(-0.00020835470058955252)),(to_sfixed_a(-0.0005097283283248544)),(to_sfixed_a(-0.0004956654738634825)),(to_sfixed_a(-0.05300925299525261)),(to_sfixed_a(-0.14509707689285278)),(to_sfixed_a(-0.07001335173845291)),(to_sfixed_a(0.008691282011568546)),(to_sfixed_a(-0.011518350802361965)),(to_sfixed_a(0.008549930527806282)),(to_sfixed_a(0.06850048899650574)),(to_sfixed_a(0.29025694727897644)),(to_sfixed_a(0.16580428183078766)),(to_sfixed_a(0.18597225844860077)),(to_sfixed_a(0.12715567648410797)),(to_sfixed_a(0.1624186635017395)),(to_sfixed_a(-0.10928361117839813)),(to_sfixed_a(-0.012575488537549973)),(to_sfixed_a(-0.09860735386610031)),(to_sfixed_a(0.07040004432201385)),(to_sfixed_a(0.017311498522758484)),(to_sfixed_a(0.11582720279693604)),(to_sfixed_a(-0.028176873922348022)),(to_sfixed_a(-0.031515028327703476)),(to_sfixed_a(-1.0404081876913551e-05)),(to_sfixed_a(0.00011912017362192273)),(to_sfixed_a(-1.752689939849006e-07)),(to_sfixed_a(6.319351814454421e-05)),(to_sfixed_a(0.00010752777598099783)),(to_sfixed_a(0.00027607494848780334)),(to_sfixed_a(-3.728240335476585e-05)),(to_sfixed_a(-0.00921448040753603)),(to_sfixed_a(-0.01721462979912758)),(to_sfixed_a(-0.05425285920500755)),(to_sfixed_a(0.02450341172516346)),(to_sfixed_a(-0.00805254839360714)),(to_sfixed_a(0.0711209699511528)),(to_sfixed_a(0.023496145382523537)),(to_sfixed_a(-0.052337177097797394)),(to_sfixed_a(-0.012800872325897217)),(to_sfixed_a(-0.1961144357919693)),(to_sfixed_a(-0.030181439593434334)),(to_sfixed_a(-0.03912857174873352)),(to_sfixed_a(0.22069062292575836)),(to_sfixed_a(0.1206907108426094)),(to_sfixed_a(0.12544865906238556)),(to_sfixed_a(0.05368172749876976)),(to_sfixed_a(-0.20422956347465515)),(to_sfixed_a(-0.09109564125537872)),(to_sfixed_a(0.02896387130022049)),(to_sfixed_a(0.135060116648674)),(to_sfixed_a(-0.15619942545890808)),(to_sfixed_a(-0.010164008475840092)),(to_sfixed_a(-0.00012329411401879042)),(to_sfixed_a(0.0002443426928948611)),(to_sfixed_a(4.92258150188718e-05)),(to_sfixed_a(-9.147100172413047e-06)),(to_sfixed_a(0.00022214995988178998)),(to_sfixed_a(2.0413604943314567e-05)),(to_sfixed_a(-0.09492386877536774)),(to_sfixed_a(-6.300238601397723e-05)),(to_sfixed_a(-0.10914205014705658)),(to_sfixed_a(0.09054147452116013)),(to_sfixed_a(0.0628025233745575)),(to_sfixed_a(0.2242349088191986)),(to_sfixed_a(0.17420703172683716)),(to_sfixed_a(0.4445320963859558)),(to_sfixed_a(-0.07068406790494919)),(to_sfixed_a(-0.1760336458683014)),(to_sfixed_a(-0.13191209733486176)),(to_sfixed_a(0.2496001273393631)),(to_sfixed_a(0.29048001766204834)),(to_sfixed_a(0.16110652685165405)),(to_sfixed_a(0.017636330798268318)),(to_sfixed_a(-0.015784770250320435)),(to_sfixed_a(0.007204282563179731)),(to_sfixed_a(-0.06244392320513725)),(to_sfixed_a(0.03287937864661217)),(to_sfixed_a(0.22042256593704224)),(to_sfixed_a(-0.0025095846503973007)),(to_sfixed_a(0.00021924851171206683)),(to_sfixed_a(4.068477574037388e-05)),(to_sfixed_a(9.17296638363041e-05)),(to_sfixed_a(3.535665018716827e-05)),(to_sfixed_a(-8.648478979011998e-05)),(to_sfixed_a(0.000145662110298872)),(to_sfixed_a(-7.605400605825707e-05)),(to_sfixed_a(7.12667460902594e-05)),(to_sfixed_a(-0.00010877076420001686)),(to_sfixed_a(-0.1714327037334442)),(to_sfixed_a(-0.10493158549070358)),(to_sfixed_a(0.0254364050924778)),(to_sfixed_a(0.1245187520980835)),(to_sfixed_a(0.2838234305381775)),(to_sfixed_a(0.025792934000492096)),(to_sfixed_a(0.09407814592123032)),(to_sfixed_a(0.07821574062108994)),(to_sfixed_a(-0.07317401468753815)),(to_sfixed_a(0.057913973927497864)),(to_sfixed_a(0.10533850640058517)),(to_sfixed_a(0.0881577581167221)),(to_sfixed_a(0.0995575562119484)),(to_sfixed_a(-0.31209245324134827)),(to_sfixed_a(0.047983285039663315)),(to_sfixed_a(0.17268435657024384)),(to_sfixed_a(0.17914658784866333)),(to_sfixed_a(0.022803159430623055)),(to_sfixed_a(-0.05471311882138252)),(to_sfixed_a(-0.020337583497166634)),(to_sfixed_a(0.0001508975401520729)),(to_sfixed_a(-0.00032245495822280645)),(to_sfixed_a(-4.1907311242539436e-05)),(to_sfixed_a(5.035879439674318e-05)),(to_sfixed_a(0.00019473647989798337)),(to_sfixed_a(-6.277887587202713e-05)),(to_sfixed_a(-4.057897604070604e-05)),(to_sfixed_a(-0.01233641430735588)),(to_sfixed_a(-0.00010176717478316277)),(to_sfixed_a(0.06970594823360443)),(to_sfixed_a(-0.09717825055122375)),(to_sfixed_a(0.2825303077697754)),(to_sfixed_a(0.07052403688430786)),(to_sfixed_a(-0.06490176171064377)),(to_sfixed_a(-0.0774666965007782)),(to_sfixed_a(-0.2550557255744934)),(to_sfixed_a(0.10843772441148758)),(to_sfixed_a(-0.11483261734247208)),(to_sfixed_a(-0.035386163741350174)),(to_sfixed_a(0.17897413671016693)),(to_sfixed_a(-0.03398149833083153)),(to_sfixed_a(-0.12472789734601974)),(to_sfixed_a(-0.08178924024105072)),(to_sfixed_a(0.16460062563419342)),(to_sfixed_a(0.034605056047439575)),(to_sfixed_a(-0.05377667397260666)),(to_sfixed_a(-0.0002081015845760703)),(to_sfixed_a(0.03432993218302727)),(to_sfixed_a(-8.859846275299788e-05)),(to_sfixed_a(-0.0002373824390815571)),(to_sfixed_a(2.1515666958293878e-05)),(to_sfixed_a(5.4514141083927825e-05)),(to_sfixed_a(6.040556854713941e-07)),(to_sfixed_a(2.201757342845667e-05)),(to_sfixed_a(0.00020308820239733905)),(to_sfixed_a(-0.00027248330297879875)),(to_sfixed_a(0.02184692583978176)),(to_sfixed_a(0.0165551770478487)),(to_sfixed_a(0.15831111371517181)),(to_sfixed_a(0.09823784232139587)),(to_sfixed_a(-0.11048243939876556)),(to_sfixed_a(-0.01624358631670475)),(to_sfixed_a(0.034757792949676514)),(to_sfixed_a(0.01964326575398445)),(to_sfixed_a(-0.12851688265800476)),(to_sfixed_a(-0.007429850287735462)),(to_sfixed_a(0.0604063905775547)),(to_sfixed_a(-0.053831350058317184)),(to_sfixed_a(-0.2121724784374237)),(to_sfixed_a(-0.2679692804813385)),(to_sfixed_a(0.12413857132196426)),(to_sfixed_a(-0.003996941726654768)),(to_sfixed_a(0.011818818747997284)),(to_sfixed_a(0.028017688542604446)),(to_sfixed_a(0.0008370340801775455)),(to_sfixed_a(-1.8046092009171844e-05)),(to_sfixed_a(-0.00020703284826595336)),(to_sfixed_a(-0.0001875873567769304)),(to_sfixed_a(4.8735040763858706e-05)),(to_sfixed_a(8.815726323518902e-05)),(to_sfixed_a(-0.00012738621444441378)),(to_sfixed_a(3.8646787288598716e-05)),(to_sfixed_a(-0.00016808668442536145)),(to_sfixed_a(-0.0004341749590821564)),(to_sfixed_a(0.005668429657816887)),(to_sfixed_a(-0.0024552391842007637)),(to_sfixed_a(0.16450318694114685)),(to_sfixed_a(0.21570391952991486)),(to_sfixed_a(0.11518966406583786)),(to_sfixed_a(-0.06959978491067886)),(to_sfixed_a(0.07689774036407471)),(to_sfixed_a(0.010368473827838898)),(to_sfixed_a(-0.05441694334149361)),(to_sfixed_a(0.15464290976524353)),(to_sfixed_a(0.19552092254161835)),(to_sfixed_a(-0.15017098188400269)),(to_sfixed_a(-0.1297905594110489)),(to_sfixed_a(0.1456204056739807)),(to_sfixed_a(0.14735697209835052)),(to_sfixed_a(0.045178819447755814)),(to_sfixed_a(0.014239327982068062)),(to_sfixed_a(0.0026166026946157217)),(to_sfixed_a(0.004594358615577221)),(to_sfixed_a(0.00017717793525662273)),(to_sfixed_a(7.767011993564665e-05)),(to_sfixed_a(-4.620000981958583e-05)),(to_sfixed_a(-6.296155333984643e-05)),(to_sfixed_a(-9.08057190827094e-05)),(to_sfixed_a(-1.8134856873075478e-05)),(to_sfixed_a(-1.3514600141206756e-05)),(to_sfixed_a(0.00015377072850242257)),(to_sfixed_a(0.06074340268969536)),(to_sfixed_a(-0.040539517998695374)),(to_sfixed_a(0.25341761112213135)),(to_sfixed_a(0.01962975226342678)),(to_sfixed_a(0.05300761014223099)),(to_sfixed_a(-0.052535802125930786)),(to_sfixed_a(-0.11010687053203583)),(to_sfixed_a(0.0906866043806076)),(to_sfixed_a(0.09005498141050339)),(to_sfixed_a(0.14643943309783936)),(to_sfixed_a(-0.06522737443447113)),(to_sfixed_a(-0.06858963519334793)),(to_sfixed_a(-0.016897419467568398)),(to_sfixed_a(0.2691550552845001)),(to_sfixed_a(-0.040950316935777664)),(to_sfixed_a(-0.11130780726671219)),(to_sfixed_a(0.006042467895895243)),(to_sfixed_a(-0.026087578386068344)),(to_sfixed_a(0.009851701557636261)),(to_sfixed_a(0.004175115376710892)),(to_sfixed_a(-0.00016237862291745842)),(to_sfixed_a(-0.0001602247211849317)),(to_sfixed_a(-0.0005010216846130788)),(to_sfixed_a(1.987705400097184e-05)),(to_sfixed_a(0.00022160151274874806)),(to_sfixed_a(0.00028426380595192313)),(to_sfixed_a(-9.749182208906859e-05)),(to_sfixed_a(0.00015977172006387264)),(to_sfixed_a(0.0001518687349744141)),(to_sfixed_a(-0.011408327147364616)),(to_sfixed_a(0.1522732675075531)),(to_sfixed_a(0.12535744905471802)),(to_sfixed_a(0.12268055230379105)),(to_sfixed_a(-0.21604251861572266)),(to_sfixed_a(0.1989886611700058)),(to_sfixed_a(0.16534435749053955)),(to_sfixed_a(-0.39359477162361145)),(to_sfixed_a(-0.19158881902694702)),(to_sfixed_a(-0.037498556077480316)),(to_sfixed_a(-0.07846421003341675)),(to_sfixed_a(0.0647687241435051)),(to_sfixed_a(-0.06712375581264496)),(to_sfixed_a(-0.0016963592497631907)),(to_sfixed_a(0.1943986564874649)),(to_sfixed_a(0.10487143695354462)),(to_sfixed_a(-0.00021021097199991345)),(to_sfixed_a(-0.002971076173707843)),(to_sfixed_a(-0.0038874272722750902)),(to_sfixed_a(0.0001445620582671836)),(to_sfixed_a(5.324900848791003e-05)),(to_sfixed_a(2.3491809770348482e-05)),(to_sfixed_a(-4.953062216372928e-06)),(to_sfixed_a(0.00012899284774903208)),(to_sfixed_a(-1.108548076445004e-05)),(to_sfixed_a(-2.2890495529281907e-05)),(to_sfixed_a(0.00018704355170484632)),(to_sfixed_a(1.6485482774442062e-05)),(to_sfixed_a(0.00023971201153472066)),(to_sfixed_a(0.00018987777002621442)),(to_sfixed_a(0.00013987720012664795)),(to_sfixed_a(0.00017810010467655957)),(to_sfixed_a(-0.00029545321012847126)),(to_sfixed_a(0.19563238322734833)),(to_sfixed_a(-0.00044980592792853713)),(to_sfixed_a(-0.0005421306123025715)),(to_sfixed_a(0.15078580379486084)),(to_sfixed_a(0.03231361135840416)),(to_sfixed_a(0.01826798915863037)),(to_sfixed_a(0.09863188862800598)),(to_sfixed_a(0.15576672554016113)),(to_sfixed_a(0.1991361528635025)),(to_sfixed_a(-0.002005958463996649)),(to_sfixed_a(-0.00021756466594524682)),(to_sfixed_a(-9.696850611362606e-05)),(to_sfixed_a(0.00036798897781409323)),(to_sfixed_a(-1.2605837582668755e-05)),(to_sfixed_a(-7.740721775917336e-05)),(to_sfixed_a(-2.6910427550319582e-05)),(to_sfixed_a(-8.864022674970329e-05)),(to_sfixed_a(4.810390237253159e-05)),(to_sfixed_a(-0.0001906339020933956)),(to_sfixed_a(8.928435272537172e-05)),(to_sfixed_a(0.00018352046026848257)),(to_sfixed_a(-2.9461312806233764e-05)),(to_sfixed_a(-0.00011708407691912726)),(to_sfixed_a(0.00011366623948561028)),(to_sfixed_a(0.00019131832232233137)),(to_sfixed_a(8.729174624022562e-06)),(to_sfixed_a(-7.00773261996801e-06)),(to_sfixed_a(6.27889166935347e-05)),(to_sfixed_a(-0.00023747525119688362)),(to_sfixed_a(-8.247324876720086e-05)),(to_sfixed_a(0.00010653806384652853)),(to_sfixed_a(0.0003707311989273876)),(to_sfixed_a(0.00040812158840708435)),(to_sfixed_a(-7.270849891938269e-05)),(to_sfixed_a(3.7592967601085547e-06)),(to_sfixed_a(-0.00026430096477270126)),(to_sfixed_a(6.384179869201034e-05)),(to_sfixed_a(7.241286220960319e-05)),(to_sfixed_a(9.680385119281709e-05)),(to_sfixed_a(-0.0002202988980570808)),(to_sfixed_a(0.000109563407022506)),(to_sfixed_a(-8.70456569828093e-05)),(to_sfixed_a(-0.00010042203211924061)),(to_sfixed_a(-1.988697022170527e-06)),(to_sfixed_a(1.9019711544387974e-05)),(to_sfixed_a(0.00033277407055720687)));

    constant weight_n0_28 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-0.00011219259613426402)),(to_sfixed_a(-1.0710748483688803e-06)),(to_sfixed_a(-6.647493137279525e-05)),(to_sfixed_a(-0.00013603625120595098)),(to_sfixed_a(-0.0001587823498994112)),(to_sfixed_a(-7.904718950157985e-05)),(to_sfixed_a(-5.375383989303373e-05)),(to_sfixed_a(-5.937476544204401e-06)),(to_sfixed_a(6.775544170523062e-05)),(to_sfixed_a(0.00011685425124596804)),(to_sfixed_a(-0.00038641528226435184)),(to_sfixed_a(-0.0001508343848399818)),(to_sfixed_a(4.9927861255127937e-05)),(to_sfixed_a(0.0002687934902496636)),(to_sfixed_a(-0.00013018667232245207)),(to_sfixed_a(0.0001513713359599933)),(to_sfixed_a(-4.178784365649335e-05)),(to_sfixed_a(6.222605588845909e-05)),(to_sfixed_a(0.00017002287495415658)),(to_sfixed_a(-3.997868770966306e-05)),(to_sfixed_a(-0.00025099326740019023)),(to_sfixed_a(-9.448706259718165e-05)),(to_sfixed_a(0.0001322180760325864)),(to_sfixed_a(0.00014810479478910565)),(to_sfixed_a(-0.00020570633932948112)),(to_sfixed_a(-0.00019201052782591432)),(to_sfixed_a(-0.00022201672254595906)),(to_sfixed_a(-0.00010296475375071168)),(to_sfixed_a(0.00013796929852105677)),(to_sfixed_a(0.00024368244339711964)),(to_sfixed_a(-9.149641846306622e-05)),(to_sfixed_a(-0.00022855299175716937)),(to_sfixed_a(5.113784936838783e-05)),(to_sfixed_a(8.532070205546916e-05)),(to_sfixed_a(-1.2386410162434913e-05)),(to_sfixed_a(0.00011315091251162812)),(to_sfixed_a(-0.00025631097378209233)),(to_sfixed_a(-0.00019513373263180256)),(to_sfixed_a(-2.9897364584030584e-05)),(to_sfixed_a(-0.00014230862143449485)),(to_sfixed_a(8.966301538748667e-05)),(to_sfixed_a(-0.00018622385687194765)),(to_sfixed_a(-0.0002083528379444033)),(to_sfixed_a(-0.0002936155360657722)),(to_sfixed_a(0.00022276390518527478)),(to_sfixed_a(7.762242603348568e-05)),(to_sfixed_a(4.1902334487531334e-05)),(to_sfixed_a(-2.0516843051154865e-06)),(to_sfixed_a(-0.0001891988213174045)),(to_sfixed_a(2.247461634397041e-05)),(to_sfixed_a(-3.8362635677913204e-05)),(to_sfixed_a(-0.0003441623121034354)),(to_sfixed_a(0.00011818052735179663)),(to_sfixed_a(2.6526018700678833e-05)),(to_sfixed_a(-6.906977796461433e-05)),(to_sfixed_a(2.8890564863104373e-05)),(to_sfixed_a(-1.5132173757592682e-05)),(to_sfixed_a(-0.00016723696899134666)),(to_sfixed_a(-2.6858780984184705e-05)),(to_sfixed_a(-2.032218617387116e-05)),(to_sfixed_a(-0.00021141592878848314)),(to_sfixed_a(-2.3997543394216336e-05)),(to_sfixed_a(-5.850122761330567e-05)),(to_sfixed_a(7.175975042628124e-05)),(to_sfixed_a(0.00021852429199498147)),(to_sfixed_a(6.253376341192052e-05)),(to_sfixed_a(6.912785465829074e-05)),(to_sfixed_a(3.597471004468389e-05)),(to_sfixed_a(-5.2820771088590845e-05)),(to_sfixed_a(0.0002567082701716572)),(to_sfixed_a(0.00012384235742501915)),(to_sfixed_a(-3.41589875461068e-05)),(to_sfixed_a(-0.00011872452887473628)),(to_sfixed_a(-7.3888772931240965e-06)),(to_sfixed_a(4.036106929561356e-06)),(to_sfixed_a(-0.0002063213032670319)),(to_sfixed_a(-1.5972269466146827e-05)),(to_sfixed_a(0.00013571458111982793)),(to_sfixed_a(5.569694621954113e-05)),(to_sfixed_a(9.047573985299096e-05)),(to_sfixed_a(-0.00027961385785602033)),(to_sfixed_a(0.00021863140864297748)),(to_sfixed_a(3.688210927066393e-05)),(to_sfixed_a(-2.1697880583815277e-05)),(to_sfixed_a(8.116762910503894e-05)),(to_sfixed_a(7.299599383259192e-05)),(to_sfixed_a(-8.909321331884712e-05)),(to_sfixed_a(-9.87536259344779e-05)),(to_sfixed_a(0.00010109526192536578)),(to_sfixed_a(-0.0001391091791447252)),(to_sfixed_a(0.00011154262028867379)),(to_sfixed_a(-0.00013103029050398618)),(to_sfixed_a(0.021161744371056557)),(to_sfixed_a(5.7000870583578944e-05)),(to_sfixed_a(0.02391100861132145)),(to_sfixed_a(0.004910513758659363)),(to_sfixed_a(0.021285492926836014)),(to_sfixed_a(0.04408125951886177)),(to_sfixed_a(0.08859771490097046)),(to_sfixed_a(0.03449273481965065)),(to_sfixed_a(-0.008058645762503147)),(to_sfixed_a(-0.01164939533919096)),(to_sfixed_a(0.14197500050067902)),(to_sfixed_a(-0.020028045400977135)),(to_sfixed_a(-0.01119392178952694)),(to_sfixed_a(-0.02236921340227127)),(to_sfixed_a(-2.4339045921806246e-05)),(to_sfixed_a(-2.9735918360529467e-05)),(to_sfixed_a(0.00010180650861002505)),(to_sfixed_a(8.649737719679251e-05)),(to_sfixed_a(0.0002680823381524533)),(to_sfixed_a(4.033161894767545e-05)),(to_sfixed_a(4.061574873048812e-05)),(to_sfixed_a(5.077537571196444e-05)),(to_sfixed_a(-7.11351094651036e-06)),(to_sfixed_a(-1.997787330765277e-05)),(to_sfixed_a(-0.0001753088436089456)),(to_sfixed_a(-0.00010702929284889251)),(to_sfixed_a(0.00034244207199662924)),(to_sfixed_a(-0.00806700624525547)),(to_sfixed_a(0.032977648079395294)),(to_sfixed_a(0.01791364885866642)),(to_sfixed_a(0.026176564395427704)),(to_sfixed_a(-0.015907548367977142)),(to_sfixed_a(0.0011144678574055433)),(to_sfixed_a(-0.237979456782341)),(to_sfixed_a(-0.31651920080184937)),(to_sfixed_a(-0.14272207021713257)),(to_sfixed_a(0.13384279608726501)),(to_sfixed_a(0.1462896168231964)),(to_sfixed_a(0.04711971804499626)),(to_sfixed_a(-0.03436577692627907)),(to_sfixed_a(-0.0001934575557243079)),(to_sfixed_a(0.0771043449640274)),(to_sfixed_a(0.043429598212242126)),(to_sfixed_a(5.6285967730218545e-05)),(to_sfixed_a(0.0006502109463326633)),(to_sfixed_a(8.08163094916381e-05)),(to_sfixed_a(-8.552511280868202e-05)),(to_sfixed_a(8.718007302377373e-05)),(to_sfixed_a(-7.501501386286691e-05)),(to_sfixed_a(-2.1736384951509535e-05)),(to_sfixed_a(0.00013740187569055706)),(to_sfixed_a(0.00015431649808306247)),(to_sfixed_a(0.0019928012043237686)),(to_sfixed_a(-0.009480195119976997)),(to_sfixed_a(0.0019905949011445045)),(to_sfixed_a(-0.05998396500945091)),(to_sfixed_a(0.03982880711555481)),(to_sfixed_a(-0.023568376898765564)),(to_sfixed_a(0.03532673791050911)),(to_sfixed_a(-0.13069725036621094)),(to_sfixed_a(0.10321901738643646)),(to_sfixed_a(-0.0385671928524971)),(to_sfixed_a(-0.07203811407089233)),(to_sfixed_a(-0.02493952214717865)),(to_sfixed_a(-0.028768135234713554)),(to_sfixed_a(0.188007190823555)),(to_sfixed_a(0.20674888789653778)),(to_sfixed_a(0.2062523365020752)),(to_sfixed_a(-0.08251121640205383)),(to_sfixed_a(-0.03724805638194084)),(to_sfixed_a(0.0021398202516138554)),(to_sfixed_a(-0.05405106022953987)),(to_sfixed_a(0.0001751529925968498)),(to_sfixed_a(0.00010963539534714073)),(to_sfixed_a(-4.239542977302335e-05)),(to_sfixed_a(-0.00015571167750749737)),(to_sfixed_a(-8.860446541802958e-05)),(to_sfixed_a(-0.0002157406706828624)),(to_sfixed_a(2.5455510694882832e-05)),(to_sfixed_a(8.1152371421922e-05)),(to_sfixed_a(8.735973096918315e-05)),(to_sfixed_a(-0.009172563441097736)),(to_sfixed_a(-0.025290146470069885)),(to_sfixed_a(-0.007821865379810333)),(to_sfixed_a(0.03356810286641121)),(to_sfixed_a(0.024588681757450104)),(to_sfixed_a(0.08992139995098114)),(to_sfixed_a(-0.04731125012040138)),(to_sfixed_a(-0.013708023354411125)),(to_sfixed_a(0.128766268491745)),(to_sfixed_a(-0.11946578323841095)),(to_sfixed_a(0.15472598373889923)),(to_sfixed_a(0.11238960921764374)),(to_sfixed_a(-0.0755874365568161)),(to_sfixed_a(-0.09721438586711884)),(to_sfixed_a(-0.016597731038928032)),(to_sfixed_a(-0.1702081710100174)),(to_sfixed_a(-0.08181845396757126)),(to_sfixed_a(-0.05755998566746712)),(to_sfixed_a(-0.09503672271966934)),(to_sfixed_a(0.0011915875365957618)),(to_sfixed_a(0.000977474614046514)),(to_sfixed_a(0.001135513884946704)),(to_sfixed_a(-0.00032655912218615413)),(to_sfixed_a(0.00030059050186537206)),(to_sfixed_a(0.00016713133663870394)),(to_sfixed_a(-6.092546391300857e-05)),(to_sfixed_a(0.00016238940588664263)),(to_sfixed_a(-6.599785410799086e-05)),(to_sfixed_a(0.04932224005460739)),(to_sfixed_a(0.02178770676255226)),(to_sfixed_a(0.11463051289319992)),(to_sfixed_a(0.15319490432739258)),(to_sfixed_a(-0.026054659858345985)),(to_sfixed_a(0.053296975791454315)),(to_sfixed_a(-0.12294474989175797)),(to_sfixed_a(-0.024932237342000008)),(to_sfixed_a(0.20126046240329742)),(to_sfixed_a(0.047632914036512375)),(to_sfixed_a(-0.060031384229660034)),(to_sfixed_a(0.10964758694171906)),(to_sfixed_a(0.10366448760032654)),(to_sfixed_a(-0.17809034883975983)),(to_sfixed_a(-0.3916774094104767)),(to_sfixed_a(-0.169958233833313)),(to_sfixed_a(-0.13024397194385529)),(to_sfixed_a(0.0542297437787056)),(to_sfixed_a(-0.20241695642471313)),(to_sfixed_a(-0.03576777130365372)),(to_sfixed_a(-0.003455034689977765)),(to_sfixed_a(4.265043025952764e-05)),(to_sfixed_a(-7.001386256888509e-05)),(to_sfixed_a(0.00012430292554199696)),(to_sfixed_a(4.5088389015290886e-05)),(to_sfixed_a(-0.0003451732627581805)),(to_sfixed_a(-6.659447535639629e-05)),(to_sfixed_a(0.04117690026760101)),(to_sfixed_a(0.0035335589200258255)),(to_sfixed_a(0.10529173165559769)),(to_sfixed_a(-0.17859193682670593)),(to_sfixed_a(0.028870999813079834)),(to_sfixed_a(-0.039754871279001236)),(to_sfixed_a(-0.22496116161346436)),(to_sfixed_a(0.22940610349178314)),(to_sfixed_a(0.014057371765375137)),(to_sfixed_a(-0.14472541213035583)),(to_sfixed_a(0.07198368012905121)),(to_sfixed_a(0.03650582581758499)),(to_sfixed_a(-0.22435808181762695)),(to_sfixed_a(-0.13669437170028687)),(to_sfixed_a(0.057191669940948486)),(to_sfixed_a(-0.07912538945674896)),(to_sfixed_a(0.13463561236858368)),(to_sfixed_a(-0.21561019122600555)),(to_sfixed_a(-0.12878771126270294)),(to_sfixed_a(0.14008302986621857)),(to_sfixed_a(-0.15549281239509583)),(to_sfixed_a(-0.0239242110401392)),(to_sfixed_a(7.916560571175069e-05)),(to_sfixed_a(0.00030208000680431724)),(to_sfixed_a(-3.8300964661175385e-05)),(to_sfixed_a(0.00028603587998077273)),(to_sfixed_a(-0.0001083279203157872)),(to_sfixed_a(0.0001173044292954728)),(to_sfixed_a(0.0013677324168384075)),(to_sfixed_a(0.13926130533218384)),(to_sfixed_a(0.17645207047462463)),(to_sfixed_a(-0.0031183494720607996)),(to_sfixed_a(0.07387630641460419)),(to_sfixed_a(0.051759637892246246)),(to_sfixed_a(0.37022560834884644)),(to_sfixed_a(0.14600838720798492)),(to_sfixed_a(0.35363954305648804)),(to_sfixed_a(-0.001244796090759337)),(to_sfixed_a(-0.1509246975183487)),(to_sfixed_a(-0.19515246152877808)),(to_sfixed_a(0.06801824271678925)),(to_sfixed_a(0.2811303436756134)),(to_sfixed_a(0.05694486200809479)),(to_sfixed_a(-0.12032291293144226)),(to_sfixed_a(0.13472343981266022)),(to_sfixed_a(-0.08339313417673111)),(to_sfixed_a(-0.23543088138103485)),(to_sfixed_a(0.13564623892307281)),(to_sfixed_a(0.06898637861013412)),(to_sfixed_a(-0.00014942357665859163)),(to_sfixed_a(8.271380465885159e-06)),(to_sfixed_a(-0.00011896937940036878)),(to_sfixed_a(1.3387390254138154e-06)),(to_sfixed_a(0.00023710272216703743)),(to_sfixed_a(5.6499859056202695e-05)),(to_sfixed_a(-0.00016656309890095145)),(to_sfixed_a(0.015705272555351257)),(to_sfixed_a(0.07224202901124954)),(to_sfixed_a(-0.07223115116357803)),(to_sfixed_a(0.03711544722318649)),(to_sfixed_a(-0.08017787337303162)),(to_sfixed_a(-0.022207120433449745)),(to_sfixed_a(-0.04957488551735878)),(to_sfixed_a(-0.014222613535821438)),(to_sfixed_a(0.09521081298589706)),(to_sfixed_a(-0.20647849142551422)),(to_sfixed_a(-0.25432339310646057)),(to_sfixed_a(0.018074534833431244)),(to_sfixed_a(0.28258630633354187)),(to_sfixed_a(0.1641162782907486)),(to_sfixed_a(-0.004116381518542767)),(to_sfixed_a(-0.08139218389987946)),(to_sfixed_a(-0.17519988119602203)),(to_sfixed_a(-0.2080390304327011)),(to_sfixed_a(0.09181611239910126)),(to_sfixed_a(0.11026490479707718)),(to_sfixed_a(-0.06210875138640404)),(to_sfixed_a(-0.039773162454366684)),(to_sfixed_a(5.412788232206367e-05)),(to_sfixed_a(-4.405266008689068e-05)),(to_sfixed_a(6.303811096586287e-05)),(to_sfixed_a(4.104967229068279e-05)),(to_sfixed_a(0.0001265788305317983)),(to_sfixed_a(0.019702021032571793)),(to_sfixed_a(0.10189444571733475)),(to_sfixed_a(0.07705690711736679)),(to_sfixed_a(-0.050772957503795624)),(to_sfixed_a(0.03887425363063812)),(to_sfixed_a(-0.01969306357204914)),(to_sfixed_a(-0.12215588241815567)),(to_sfixed_a(-0.016987143084406853)),(to_sfixed_a(0.045409757643938065)),(to_sfixed_a(0.2626795470714569)),(to_sfixed_a(0.09749516099691391)),(to_sfixed_a(0.15263786911964417)),(to_sfixed_a(-0.15588828921318054)),(to_sfixed_a(0.08971536159515381)),(to_sfixed_a(-0.10890400409698486)),(to_sfixed_a(0.17762252688407898)),(to_sfixed_a(0.026593979448080063)),(to_sfixed_a(0.04858774319291115)),(to_sfixed_a(0.00016393253463320434)),(to_sfixed_a(0.03427701070904732)),(to_sfixed_a(-0.06582305580377579)),(to_sfixed_a(0.04631996527314186)),(to_sfixed_a(-0.00012121935287723318)),(to_sfixed_a(0.0001698378036962822)),(to_sfixed_a(-5.2230683650122955e-05)),(to_sfixed_a(-0.00013886213127989322)),(to_sfixed_a(-1.2798961506632622e-05)),(to_sfixed_a(-0.00012632727157324553)),(to_sfixed_a(-7.401173934340477e-05)),(to_sfixed_a(-0.008293762803077698)),(to_sfixed_a(0.15493996441364288)),(to_sfixed_a(0.07838767766952515)),(to_sfixed_a(-0.05452815815806389)),(to_sfixed_a(0.06424622237682343)),(to_sfixed_a(-0.09762127697467804)),(to_sfixed_a(0.08311427384614944)),(to_sfixed_a(0.06080068647861481)),(to_sfixed_a(0.25247645378112793)),(to_sfixed_a(0.045154865831136703)),(to_sfixed_a(0.0874706283211708)),(to_sfixed_a(-0.2551818788051605)),(to_sfixed_a(-0.18358337879180908)),(to_sfixed_a(-0.1456701010465622)),(to_sfixed_a(-0.040558669716119766)),(to_sfixed_a(-0.05251552537083626)),(to_sfixed_a(0.12170573323965073)),(to_sfixed_a(0.11757203191518784)),(to_sfixed_a(0.02375897392630577)),(to_sfixed_a(-0.18582728505134583)),(to_sfixed_a(-0.06568489223718643)),(to_sfixed_a(-8.116111712297425e-05)),(to_sfixed_a(-0.00021495450346264988)),(to_sfixed_a(-0.00017257336003240198)),(to_sfixed_a(1.655427331570536e-05)),(to_sfixed_a(0.00010652842320268974)),(to_sfixed_a(1.063257241185056e-05)),(to_sfixed_a(-3.1056876537149947e-07)),(to_sfixed_a(0.12239763140678406)),(to_sfixed_a(0.2094360589981079)),(to_sfixed_a(0.1039338931441307)),(to_sfixed_a(-0.12039700895547867)),(to_sfixed_a(-0.015774061903357506)),(to_sfixed_a(-0.03639842942357063)),(to_sfixed_a(-0.15505994856357574)),(to_sfixed_a(0.295168936252594)),(to_sfixed_a(0.23608148097991943)),(to_sfixed_a(-0.0066789621487259865)),(to_sfixed_a(0.14914347231388092)),(to_sfixed_a(-0.2252197414636612)),(to_sfixed_a(-0.2875562310218811)),(to_sfixed_a(-0.10403226315975189)),(to_sfixed_a(-0.1186390221118927)),(to_sfixed_a(-0.1697855144739151)),(to_sfixed_a(-0.10587270557880402)),(to_sfixed_a(-0.10114704817533493)),(to_sfixed_a(0.017816592007875443)),(to_sfixed_a(-0.03404468297958374)),(to_sfixed_a(0.02757377363741398)),(to_sfixed_a(0.0007214086363092065)),(to_sfixed_a(0.001325466320849955)),(to_sfixed_a(0.0003822515136562288)),(to_sfixed_a(-7.308972999453545e-05)),(to_sfixed_a(0.00017118651885539293)),(to_sfixed_a(-0.0006186705431900918)),(to_sfixed_a(-3.316647052997723e-05)),(to_sfixed_a(0.0005119115812703967)),(to_sfixed_a(-0.3497597277164459)),(to_sfixed_a(-0.018833909183740616)),(to_sfixed_a(-0.2260565161705017)),(to_sfixed_a(-0.24318741261959076)),(to_sfixed_a(-0.047668810933828354)),(to_sfixed_a(0.01599312014877796)),(to_sfixed_a(-0.014919052831828594)),(to_sfixed_a(-0.5030843615531921)),(to_sfixed_a(-0.3561365008354187)),(to_sfixed_a(0.1409849375486374)),(to_sfixed_a(-0.14757481217384338)),(to_sfixed_a(-0.19172027707099915)),(to_sfixed_a(0.0008390876464545727)),(to_sfixed_a(0.05802981182932854)),(to_sfixed_a(0.00919664278626442)),(to_sfixed_a(-0.008617214858531952)),(to_sfixed_a(-0.13406462967395782)),(to_sfixed_a(-0.01717517152428627)),(to_sfixed_a(0.0899631530046463)),(to_sfixed_a(0.03123917616903782)),(to_sfixed_a(0.0008847241988405585)),(to_sfixed_a(-9.299354132963344e-05)),(to_sfixed_a(-6.5669919422362e-05)),(to_sfixed_a(0.00015595901641063392)),(to_sfixed_a(-4.769655424752273e-05)),(to_sfixed_a(0.00017796210886444896)),(to_sfixed_a(-4.482404619920999e-06)),(to_sfixed_a(0.0012523324694484472)),(to_sfixed_a(-0.19647032022476196)),(to_sfixed_a(0.07335346937179565)),(to_sfixed_a(-0.15140964090824127)),(to_sfixed_a(0.18465331196784973)),(to_sfixed_a(0.12245024740695953)),(to_sfixed_a(0.10996879637241364)),(to_sfixed_a(-0.13069050014019012)),(to_sfixed_a(-0.2664380967617035)),(to_sfixed_a(-0.12603218853473663)),(to_sfixed_a(0.06222568079829216)),(to_sfixed_a(-0.17043396830558777)),(to_sfixed_a(-0.12322843074798584)),(to_sfixed_a(0.04593046382069588)),(to_sfixed_a(-0.055018700659275055)),(to_sfixed_a(-0.027206875383853912)),(to_sfixed_a(-0.13939662277698517)),(to_sfixed_a(-0.14133089780807495)),(to_sfixed_a(-0.02898513898253441)),(to_sfixed_a(0.013678285293281078)),(to_sfixed_a(0.17401741445064545)),(to_sfixed_a(0.0005255380528979003)),(to_sfixed_a(-0.00012381686246953905)),(to_sfixed_a(0.00021082768216729164)),(to_sfixed_a(-0.0004002971691079438)),(to_sfixed_a(-9.602423961041495e-05)),(to_sfixed_a(-6.367157766362652e-05)),(to_sfixed_a(0.0013217757223173976)),(to_sfixed_a(0.19557899236679077)),(to_sfixed_a(0.1728820502758026)),(to_sfixed_a(0.01150953397154808)),(to_sfixed_a(0.28734079003334045)),(to_sfixed_a(0.10360363870859146)),(to_sfixed_a(0.06537726521492004)),(to_sfixed_a(-0.2816019058227539)),(to_sfixed_a(-0.19094306230545044)),(to_sfixed_a(0.20218482613563538)),(to_sfixed_a(0.2719271183013916)),(to_sfixed_a(0.052640315145254135)),(to_sfixed_a(0.013888491317629814)),(to_sfixed_a(-0.02323331870138645)),(to_sfixed_a(0.2872627377510071)),(to_sfixed_a(0.1795283555984497)),(to_sfixed_a(0.08467366546392441)),(to_sfixed_a(-0.06830362230539322)),(to_sfixed_a(-0.09482534229755402)),(to_sfixed_a(-0.021535934880375862)),(to_sfixed_a(0.01857919804751873)),(to_sfixed_a(0.07764506340026855)),(to_sfixed_a(-0.022389346733689308)),(to_sfixed_a(3.626446414273232e-05)),(to_sfixed_a(-0.0003845408500637859)),(to_sfixed_a(0.0001985810522455722)),(to_sfixed_a(-5.813141251564957e-05)),(to_sfixed_a(0.0010584571864455938)),(to_sfixed_a(0.001618517329916358)),(to_sfixed_a(0.0017366205574944615)),(to_sfixed_a(0.25760188698768616)),(to_sfixed_a(0.0005921438569203019)),(to_sfixed_a(-0.3914545476436615)),(to_sfixed_a(-0.1969822347164154)),(to_sfixed_a(-0.3367108404636383)),(to_sfixed_a(-0.007679938338696957)),(to_sfixed_a(0.16701196134090424)),(to_sfixed_a(0.4726778566837311)),(to_sfixed_a(0.26821181178092957)),(to_sfixed_a(-0.030508875846862793)),(to_sfixed_a(-0.0014314750442281365)),(to_sfixed_a(0.3307654857635498)),(to_sfixed_a(0.07679431885480881)),(to_sfixed_a(0.16112597286701202)),(to_sfixed_a(-0.42614203691482544)),(to_sfixed_a(0.002325674518942833)),(to_sfixed_a(-0.13430288434028625)),(to_sfixed_a(-0.1542471945285797)),(to_sfixed_a(0.006436957977712154)),(to_sfixed_a(0.00023463176330551505)),(to_sfixed_a(0.00019183382391929626)),(to_sfixed_a(-0.00013955720351077616)),(to_sfixed_a(0.00034537503961473703)),(to_sfixed_a(-4.4780106691177934e-05)),(to_sfixed_a(0.00013704836601391435)),(to_sfixed_a(-0.0001305223413510248)),(to_sfixed_a(-0.00701395096257329)),(to_sfixed_a(0.1433660089969635)),(to_sfixed_a(0.07136858254671097)),(to_sfixed_a(0.050509680062532425)),(to_sfixed_a(-0.01653781719505787)),(to_sfixed_a(-0.31182199716567993)),(to_sfixed_a(-0.16240431368350983)),(to_sfixed_a(0.012111268937587738)),(to_sfixed_a(-0.04750802367925644)),(to_sfixed_a(-0.10381150990724564)),(to_sfixed_a(-0.39655542373657227)),(to_sfixed_a(-0.2977997362613678)),(to_sfixed_a(0.11970686912536621)),(to_sfixed_a(0.19707100093364716)),(to_sfixed_a(0.23659104108810425)),(to_sfixed_a(0.034142568707466125)),(to_sfixed_a(0.10286834836006165)),(to_sfixed_a(0.017713874578475952)),(to_sfixed_a(-0.10822948813438416)),(to_sfixed_a(-0.08768510073423386)),(to_sfixed_a(0.01323873270303011)),(to_sfixed_a(-0.020638544112443924)),(to_sfixed_a(5.267697633826174e-05)),(to_sfixed_a(9.792107448447496e-06)),(to_sfixed_a(4.1543000406818464e-05)),(to_sfixed_a(0.00020928250160068274)),(to_sfixed_a(2.5163468308164738e-05)),(to_sfixed_a(6.896749255247414e-05)),(to_sfixed_a(-0.005733346566557884)),(to_sfixed_a(-0.00509326858446002)),(to_sfixed_a(0.03645303472876549)),(to_sfixed_a(-0.017772939056158066)),(to_sfixed_a(-0.012974786572158337)),(to_sfixed_a(-0.17515935003757477)),(to_sfixed_a(0.16806355118751526)),(to_sfixed_a(0.1855297088623047)),(to_sfixed_a(0.15526774525642395)),(to_sfixed_a(-0.04548611864447594)),(to_sfixed_a(-0.2626492977142334)),(to_sfixed_a(-0.29621201753616333)),(to_sfixed_a(-0.15006019175052643)),(to_sfixed_a(-0.10237781703472137)),(to_sfixed_a(0.2718367278575897)),(to_sfixed_a(0.15873847901821136)),(to_sfixed_a(-0.01863882876932621)),(to_sfixed_a(-0.011973556131124496)),(to_sfixed_a(-0.21955284476280212)),(to_sfixed_a(0.13321611285209656)),(to_sfixed_a(0.025327958166599274)),(to_sfixed_a(-0.0001562737743370235)),(to_sfixed_a(2.96285143122077e-05)),(to_sfixed_a(0.0001446146343369037)),(to_sfixed_a(-0.00011318210454192013)),(to_sfixed_a(0.00019882824562955648)),(to_sfixed_a(-6.156504969112575e-05)),(to_sfixed_a(-0.0001456040481571108)),(to_sfixed_a(0.00011370570427970961)),(to_sfixed_a(-0.022833088412880898)),(to_sfixed_a(-0.028798017650842667)),(to_sfixed_a(0.050296884030103683)),(to_sfixed_a(0.029749298468232155)),(to_sfixed_a(0.1603870540857315)),(to_sfixed_a(0.07728276401758194)),(to_sfixed_a(0.005611879751086235)),(to_sfixed_a(-0.0011956039816141129)),(to_sfixed_a(0.08874614536762238)),(to_sfixed_a(-0.061638783663511276)),(to_sfixed_a(-0.36554405093193054)),(to_sfixed_a(-0.08888375014066696)),(to_sfixed_a(-0.10289794206619263)),(to_sfixed_a(0.20952090620994568)),(to_sfixed_a(0.1343274861574173)),(to_sfixed_a(-0.0029525465797632933)),(to_sfixed_a(-0.13294552266597748)),(to_sfixed_a(-0.028214046731591225)),(to_sfixed_a(0.015591409988701344)),(to_sfixed_a(0.03541883826255798)),(to_sfixed_a(-0.04651978984475136)),(to_sfixed_a(4.60416322312085e-06)),(to_sfixed_a(-0.00017695188580546528)),(to_sfixed_a(-0.0002632525283843279)),(to_sfixed_a(-5.444553244160488e-05)),(to_sfixed_a(-0.00014172600640449673)),(to_sfixed_a(7.016966992523521e-05)),(to_sfixed_a(-5.219196100370027e-05)),(to_sfixed_a(0.009716030210256577)),(to_sfixed_a(-0.0015108699444681406)),(to_sfixed_a(-0.10422660410404205)),(to_sfixed_a(-0.07344979792833328)),(to_sfixed_a(-0.211146742105484)),(to_sfixed_a(-0.12964299321174622)),(to_sfixed_a(0.14248508214950562)),(to_sfixed_a(0.014664733782410622)),(to_sfixed_a(-0.010222646407783031)),(to_sfixed_a(-0.18757201731204987)),(to_sfixed_a(-0.20517441630363464)),(to_sfixed_a(0.12829093635082245)),(to_sfixed_a(-0.10284440219402313)),(to_sfixed_a(0.12342140078544617)),(to_sfixed_a(0.0005166250630281866)),(to_sfixed_a(-0.022046416997909546)),(to_sfixed_a(-0.039500411599874496)),(to_sfixed_a(-0.04325852915644646)),(to_sfixed_a(0.15582741796970367)),(to_sfixed_a(0.0013783450704067945)),(to_sfixed_a(0.005535063799470663)),(to_sfixed_a(4.441718556336127e-05)),(to_sfixed_a(9.434983803657815e-05)),(to_sfixed_a(-5.029155727243051e-05)),(to_sfixed_a(-0.0001014042500173673)),(to_sfixed_a(3.080724854953587e-05)),(to_sfixed_a(-0.00018495209224056453)),(to_sfixed_a(-0.00017411820590496063)),(to_sfixed_a(6.545033556903945e-06)),(to_sfixed_a(0.0656638890504837)),(to_sfixed_a(0.05395599827170372)),(to_sfixed_a(-0.16683219373226166)),(to_sfixed_a(0.11007986217737198)),(to_sfixed_a(-0.0772109404206276)),(to_sfixed_a(0.00552563788369298)),(to_sfixed_a(0.002209128811955452)),(to_sfixed_a(0.1411404013633728)),(to_sfixed_a(0.2802782356739044)),(to_sfixed_a(-0.018861893564462662)),(to_sfixed_a(0.0383651964366436)),(to_sfixed_a(-0.0007211787160485983)),(to_sfixed_a(0.039942581206560135)),(to_sfixed_a(-0.02784908190369606)),(to_sfixed_a(-0.2317049354314804)),(to_sfixed_a(0.05774703994393349)),(to_sfixed_a(0.022681239992380142)),(to_sfixed_a(0.04285405948758125)),(to_sfixed_a(-0.006391448900103569)),(to_sfixed_a(1.403631267749006e-05)),(to_sfixed_a(-0.00021928637579549104)),(to_sfixed_a(0.0001371280668536201)),(to_sfixed_a(5.331053034751676e-05)),(to_sfixed_a(2.4579359887866303e-05)),(to_sfixed_a(0.0002763337397482246)),(to_sfixed_a(2.2287909814622253e-05)),(to_sfixed_a(0.00018881898722611368)),(to_sfixed_a(2.4625413061585277e-05)),(to_sfixed_a(-0.006188318599015474)),(to_sfixed_a(0.0021312804892659187)),(to_sfixed_a(-0.15899786353111267)),(to_sfixed_a(0.15993964672088623)),(to_sfixed_a(-0.09775649756193161)),(to_sfixed_a(0.1482178121805191)),(to_sfixed_a(0.12153592705726624)),(to_sfixed_a(0.19023466110229492)),(to_sfixed_a(0.22723275423049927)),(to_sfixed_a(0.0706222727894783)),(to_sfixed_a(-0.07393626868724823)),(to_sfixed_a(-0.045813847333192825)),(to_sfixed_a(0.07412543892860413)),(to_sfixed_a(-0.12526676058769226)),(to_sfixed_a(-0.035600341856479645)),(to_sfixed_a(-0.07308799028396606)),(to_sfixed_a(0.1476975977420807)),(to_sfixed_a(-0.00449042534455657)),(to_sfixed_a(0.1119806244969368)),(to_sfixed_a(-0.00015874688688199967)),(to_sfixed_a(-0.00014534607180394232)),(to_sfixed_a(8.198522846214473e-05)),(to_sfixed_a(0.00038199906703084707)),(to_sfixed_a(6.632547865592642e-06)),(to_sfixed_a(-0.0001226250606123358)),(to_sfixed_a(-2.2914353394298814e-05)),(to_sfixed_a(-3.8522262912010774e-05)),(to_sfixed_a(-0.02809486724436283)),(to_sfixed_a(0.023064875975251198)),(to_sfixed_a(-0.11536544561386108)),(to_sfixed_a(-0.17917640507221222)),(to_sfixed_a(0.1326785534620285)),(to_sfixed_a(0.1479307860136032)),(to_sfixed_a(-0.06882661581039429)),(to_sfixed_a(-0.01355838030576706)),(to_sfixed_a(-0.09890058636665344)),(to_sfixed_a(0.014797184616327286)),(to_sfixed_a(0.24568572640419006)),(to_sfixed_a(0.14233851432800293)),(to_sfixed_a(0.032866135239601135)),(to_sfixed_a(0.012659186497330666)),(to_sfixed_a(0.07842768728733063)),(to_sfixed_a(0.2559314966201782)),(to_sfixed_a(0.006679476238787174)),(to_sfixed_a(0.16105453670024872)),(to_sfixed_a(0.06838031858205795)),(to_sfixed_a(0.007074775639921427)),(to_sfixed_a(-2.7151692847837694e-05)),(to_sfixed_a(2.453219349263236e-05)),(to_sfixed_a(0.0001271013607038185)),(to_sfixed_a(7.334995461860672e-05)),(to_sfixed_a(-7.777728751534596e-05)),(to_sfixed_a(2.648015106387902e-05)),(to_sfixed_a(-0.00012391549535095692)),(to_sfixed_a(0.00016365297778975219)),(to_sfixed_a(0.00012994938879273832)),(to_sfixed_a(-0.017020149156451225)),(to_sfixed_a(-0.06983418017625809)),(to_sfixed_a(-0.037653543055057526)),(to_sfixed_a(-0.25086647272109985)),(to_sfixed_a(0.04983493313193321)),(to_sfixed_a(-0.05492143705487251)),(to_sfixed_a(-0.04560493305325508)),(to_sfixed_a(0.04961289465427399)),(to_sfixed_a(0.023480849340558052)),(to_sfixed_a(-0.11810418963432312)),(to_sfixed_a(-0.06025439873337746)),(to_sfixed_a(0.016096124425530434)),(to_sfixed_a(0.06603699177503586)),(to_sfixed_a(0.013860584236681461)),(to_sfixed_a(0.15255986154079437)),(to_sfixed_a(0.05731939151883125)),(to_sfixed_a(0.0013697708491235971)),(to_sfixed_a(0.0033969939686357975)),(to_sfixed_a(0.003295603906735778)),(to_sfixed_a(0.00011951386841246858)),(to_sfixed_a(-0.00012048431381117553)),(to_sfixed_a(-5.194992627366446e-05)),(to_sfixed_a(4.790213642991148e-05)),(to_sfixed_a(5.1510603952920064e-05)),(to_sfixed_a(0.00011919344979105517)),(to_sfixed_a(-0.00016477241297252476)),(to_sfixed_a(5.8236520999344066e-05)),(to_sfixed_a(3.0144427000777796e-05)),(to_sfixed_a(0.0009426379110664129)),(to_sfixed_a(0.0007687056786380708)),(to_sfixed_a(-0.0001774979755282402)),(to_sfixed_a(-0.00020148695330135524)),(to_sfixed_a(-0.0004578721127472818)),(to_sfixed_a(0.0559612400829792)),(to_sfixed_a(0.005312848836183548)),(to_sfixed_a(0.0032419280614703894)),(to_sfixed_a(0.03737592324614525)),(to_sfixed_a(0.014629202894866467)),(to_sfixed_a(-0.00146026024594903)),(to_sfixed_a(0.02707945927977562)),(to_sfixed_a(0.041285548359155655)),(to_sfixed_a(0.06886980682611465)),(to_sfixed_a(0.016589587554335594)),(to_sfixed_a(0.011282253079116344)),(to_sfixed_a(4.1790102841332555e-05)),(to_sfixed_a(0.0002570381620898843)),(to_sfixed_a(-5.9459212025103625e-06)),(to_sfixed_a(-3.175190067850053e-05)),(to_sfixed_a(0.0001395759463775903)),(to_sfixed_a(-0.000176624656887725)),(to_sfixed_a(-0.00010789986117742956)),(to_sfixed_a(0.00012473580136429518)),(to_sfixed_a(-0.00020085289725102484)),(to_sfixed_a(1.4946879673516378e-05)),(to_sfixed_a(0.0001319673756370321)),(to_sfixed_a(0.00010073991870740429)),(to_sfixed_a(-0.00013500168279279023)),(to_sfixed_a(-9.792405762709677e-05)),(to_sfixed_a(0.00016193484771065414)),(to_sfixed_a(0.0002710564876906574)),(to_sfixed_a(-1.9593353499658406e-05)),(to_sfixed_a(3.6180837923893705e-05)),(to_sfixed_a(-0.00014701664622407407)),(to_sfixed_a(-0.00011168574565090239)),(to_sfixed_a(-0.00014402477245312184)),(to_sfixed_a(0.0001852344867074862)),(to_sfixed_a(7.372565596597269e-05)),(to_sfixed_a(8.935562800616026e-05)),(to_sfixed_a(4.5224114728625864e-05)),(to_sfixed_a(-0.0001552031608298421)),(to_sfixed_a(-1.482316838519182e-05)),(to_sfixed_a(0.0001609531173016876)),(to_sfixed_a(-9.885572944767773e-05)),(to_sfixed_a(-0.00022324682504404336)),(to_sfixed_a(-1.4145090062811505e-05)),(to_sfixed_a(-5.916260488447733e-05)),(to_sfixed_a(-4.306475602788851e-05)),(to_sfixed_a(-0.00031203325488604605)),(to_sfixed_a(-0.0001398600434185937)));

    constant weight_n0_29 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(3.156435923301615e-05)),(to_sfixed_a(6.314710481092334e-05)),(to_sfixed_a(-0.00013043551007285714)),(to_sfixed_a(-7.056555477902293e-05)),(to_sfixed_a(0.0002538799890317023)),(to_sfixed_a(0.0002971882640849799)),(to_sfixed_a(0.00011336996249156073)),(to_sfixed_a(0.00015691232692915946)),(to_sfixed_a(-7.403649942716584e-05)),(to_sfixed_a(2.33526452575461e-06)),(to_sfixed_a(4.2752657464006916e-05)),(to_sfixed_a(-0.00016393691475968808)),(to_sfixed_a(-0.00017975505033973604)),(to_sfixed_a(-0.00013147119898349047)),(to_sfixed_a(0.00027792557375505567)),(to_sfixed_a(8.774646266829222e-05)),(to_sfixed_a(-6.48073764750734e-05)),(to_sfixed_a(6.020612272550352e-05)),(to_sfixed_a(-6.393328931153519e-06)),(to_sfixed_a(8.571326907258481e-05)),(to_sfixed_a(0.0001605322031537071)),(to_sfixed_a(-8.282552153104916e-05)),(to_sfixed_a(1.057392728398554e-05)),(to_sfixed_a(2.307295835635159e-05)),(to_sfixed_a(-0.0002598022110760212)),(to_sfixed_a(5.431778117781505e-05)),(to_sfixed_a(-0.0001038451082422398)),(to_sfixed_a(-6.995613512117416e-05)),(to_sfixed_a(0.0001441876229364425)),(to_sfixed_a(3.406971518415958e-05)),(to_sfixed_a(-0.00012186440289951861)),(to_sfixed_a(-0.00023493717890232801)),(to_sfixed_a(-7.617669325554743e-05)),(to_sfixed_a(-0.00016063950897660106)),(to_sfixed_a(0.00012481104931794107)),(to_sfixed_a(5.0583686970639974e-05)),(to_sfixed_a(0.00019982288358733058)),(to_sfixed_a(-0.00028763682348653674)),(to_sfixed_a(-1.1121906936750747e-05)),(to_sfixed_a(-3.596211172407493e-05)),(to_sfixed_a(8.670632814755663e-05)),(to_sfixed_a(-0.00022946708486415446)),(to_sfixed_a(0.00012355820217635483)),(to_sfixed_a(-5.6377157306997105e-05)),(to_sfixed_a(3.2883897802094e-05)),(to_sfixed_a(-9.002425213111565e-05)),(to_sfixed_a(-4.239404734107666e-05)),(to_sfixed_a(3.299291347502731e-05)),(to_sfixed_a(0.00010221677803201601)),(to_sfixed_a(0.00014741785707883537)),(to_sfixed_a(0.00018328221631236374)),(to_sfixed_a(-0.00011446033022366464)),(to_sfixed_a(-0.00017900973034556955)),(to_sfixed_a(0.0002258971508126706)),(to_sfixed_a(1.67841135407798e-05)),(to_sfixed_a(-0.0001722374581731856)),(to_sfixed_a(-0.0002333763986825943)),(to_sfixed_a(-1.7169137208838947e-05)),(to_sfixed_a(0.00012748751032631844)),(to_sfixed_a(-0.00010332415695302188)),(to_sfixed_a(-8.512428757967427e-05)),(to_sfixed_a(-0.00012371654156595469)),(to_sfixed_a(4.647714376915246e-05)),(to_sfixed_a(-0.00012133464770158753)),(to_sfixed_a(-0.00019600271480157971)),(to_sfixed_a(-2.1518924768315628e-05)),(to_sfixed_a(6.569896504515782e-05)),(to_sfixed_a(4.192402775515802e-05)),(to_sfixed_a(4.6976889279903844e-05)),(to_sfixed_a(0.005666322540491819)),(to_sfixed_a(0.00012445778702385724)),(to_sfixed_a(2.0377170585561544e-05)),(to_sfixed_a(-6.644405857514357e-06)),(to_sfixed_a(-0.00020083079289179295)),(to_sfixed_a(-1.9317507394589484e-05)),(to_sfixed_a(0.0001500039652455598)),(to_sfixed_a(-0.00015364159480668604)),(to_sfixed_a(0.0001593700872035697)),(to_sfixed_a(5.674416752299294e-05)),(to_sfixed_a(0.0002061837731162086)),(to_sfixed_a(-0.00014648932847194374)),(to_sfixed_a(-0.00024510303046554327)),(to_sfixed_a(8.273295293292904e-07)),(to_sfixed_a(6.361439591273665e-05)),(to_sfixed_a(0.00021384950377978384)),(to_sfixed_a(-0.0002929832844529301)),(to_sfixed_a(-5.557864369620802e-06)),(to_sfixed_a(-7.332443146879086e-06)),(to_sfixed_a(-0.00031148517155088484)),(to_sfixed_a(-5.1214839913882315e-05)),(to_sfixed_a(5.7888944866135716e-05)),(to_sfixed_a(-0.00018291074957232922)),(to_sfixed_a(-0.010187949985265732)),(to_sfixed_a(5.284100552671589e-05)),(to_sfixed_a(-0.011557608842849731)),(to_sfixed_a(-0.08067233115434647)),(to_sfixed_a(0.02633138746023178)),(to_sfixed_a(0.05535319820046425)),(to_sfixed_a(-0.06070278212428093)),(to_sfixed_a(0.04472927749156952)),(to_sfixed_a(0.00984770804643631)),(to_sfixed_a(0.04793308302760124)),(to_sfixed_a(0.0533936433494091)),(to_sfixed_a(-0.000457349990028888)),(to_sfixed_a(-0.006276921834796667)),(to_sfixed_a(-0.012887374497950077)),(to_sfixed_a(1.6049581972765736e-05)),(to_sfixed_a(0.00010294056119164452)),(to_sfixed_a(7.407878729281947e-05)),(to_sfixed_a(-9.378825052408502e-05)),(to_sfixed_a(0.00023931314353831112)),(to_sfixed_a(-3.708697477122769e-05)),(to_sfixed_a(-0.00023592177603859454)),(to_sfixed_a(-0.00044049075222574174)),(to_sfixed_a(6.372507777996361e-05)),(to_sfixed_a(-0.00023454203619621694)),(to_sfixed_a(-3.165358793921769e-05)),(to_sfixed_a(0.00015813681238796562)),(to_sfixed_a(-9.439772111363709e-05)),(to_sfixed_a(-0.01580914855003357)),(to_sfixed_a(0.08742450177669525)),(to_sfixed_a(-0.01577894203364849)),(to_sfixed_a(-0.22247079014778137)),(to_sfixed_a(-0.09193170815706253)),(to_sfixed_a(0.08438681811094284)),(to_sfixed_a(0.08721417188644409)),(to_sfixed_a(-0.10510136187076569)),(to_sfixed_a(-0.03637247160077095)),(to_sfixed_a(0.06114813685417175)),(to_sfixed_a(-0.05283329635858536)),(to_sfixed_a(-0.13053542375564575)),(to_sfixed_a(0.08329127728939056)),(to_sfixed_a(0.008199539966881275)),(to_sfixed_a(-0.03178548067808151)),(to_sfixed_a(0.06618008762598038)),(to_sfixed_a(-8.013653132366017e-05)),(to_sfixed_a(0.0015940011944621801)),(to_sfixed_a(1.6640078683849424e-05)),(to_sfixed_a(-4.596007420332171e-05)),(to_sfixed_a(-0.00010123787069460377)),(to_sfixed_a(-3.4677930671023205e-05)),(to_sfixed_a(-8.775894821155816e-05)),(to_sfixed_a(-3.1227989438775694e-06)),(to_sfixed_a(-0.00011380094656487927)),(to_sfixed_a(0.0006562462658621371)),(to_sfixed_a(-0.03970389813184738)),(to_sfixed_a(-0.014367313124239445)),(to_sfixed_a(0.05699021369218826)),(to_sfixed_a(-0.11619768291711807)),(to_sfixed_a(-0.05516131594777107)),(to_sfixed_a(0.021572768688201904)),(to_sfixed_a(-0.07661721855401993)),(to_sfixed_a(0.07119082659482956)),(to_sfixed_a(-0.1921265572309494)),(to_sfixed_a(0.021309828385710716)),(to_sfixed_a(-0.047634538263082504)),(to_sfixed_a(0.25758758187294006)),(to_sfixed_a(-0.0982288345694542)),(to_sfixed_a(0.2546771466732025)),(to_sfixed_a(0.1517488956451416)),(to_sfixed_a(-0.18060192465782166)),(to_sfixed_a(-0.0009215610916726291)),(to_sfixed_a(0.004584541544318199)),(to_sfixed_a(-0.02764323726296425)),(to_sfixed_a(0.00529339537024498)),(to_sfixed_a(-6.494456101791002e-06)),(to_sfixed_a(0.000170347819221206)),(to_sfixed_a(0.00010287566692568362)),(to_sfixed_a(5.6541724916314706e-05)),(to_sfixed_a(-0.00044517958303913474)),(to_sfixed_a(-2.609364855743479e-05)),(to_sfixed_a(0.0002251797850476578)),(to_sfixed_a(0.0002824387629516423)),(to_sfixed_a(-0.03444429859519005)),(to_sfixed_a(0.007438788656145334)),(to_sfixed_a(-0.15464921295642853)),(to_sfixed_a(-0.12023711949586868)),(to_sfixed_a(0.019091088324785233)),(to_sfixed_a(-0.3594309687614441)),(to_sfixed_a(-0.22542302310466766)),(to_sfixed_a(-0.08205114305019379)),(to_sfixed_a(-0.004798075649887323)),(to_sfixed_a(-0.049493178725242615)),(to_sfixed_a(-0.08639176189899445)),(to_sfixed_a(-0.1604354977607727)),(to_sfixed_a(0.07316214591264725)),(to_sfixed_a(0.019018445163965225)),(to_sfixed_a(0.14756056666374207)),(to_sfixed_a(-0.09323146939277649)),(to_sfixed_a(-0.036016013473272324)),(to_sfixed_a(0.10784746706485748)),(to_sfixed_a(0.0562007911503315)),(to_sfixed_a(0.0034402005840092897)),(to_sfixed_a(0.002617781050503254)),(to_sfixed_a(-2.3152679204940796e-05)),(to_sfixed_a(-1.9876984879374504e-05)),(to_sfixed_a(6.814183052483713e-06)),(to_sfixed_a(-6.168241816340014e-05)),(to_sfixed_a(0.00016712893557269126)),(to_sfixed_a(-5.3808795200893655e-05)),(to_sfixed_a(7.710009413131047e-06)),(to_sfixed_a(0.02726261503994465)),(to_sfixed_a(0.0085692023858428)),(to_sfixed_a(-0.07259085774421692)),(to_sfixed_a(0.26660335063934326)),(to_sfixed_a(-0.0006642520893365145)),(to_sfixed_a(-0.4258037507534027)),(to_sfixed_a(-0.13496187329292297)),(to_sfixed_a(-0.2060931921005249)),(to_sfixed_a(0.030770713463425636)),(to_sfixed_a(-0.07532794773578644)),(to_sfixed_a(-0.16356228291988373)),(to_sfixed_a(0.06946789473295212)),(to_sfixed_a(-0.10010635107755661)),(to_sfixed_a(-0.01015841867774725)),(to_sfixed_a(0.01684771291911602)),(to_sfixed_a(-0.1560220569372177)),(to_sfixed_a(0.024036793038249016)),(to_sfixed_a(-0.018634527921676636)),(to_sfixed_a(0.06512220948934555)),(to_sfixed_a(0.018752777948975563)),(to_sfixed_a(0.0005595005350187421)),(to_sfixed_a(-0.0003904833283741027)),(to_sfixed_a(-0.00013538580969907343)),(to_sfixed_a(-0.00012370712647680193)),(to_sfixed_a(0.00012450468784663826)),(to_sfixed_a(0.00021701439982280135)),(to_sfixed_a(0.00012253952445462346)),(to_sfixed_a(0.11598850041627884)),(to_sfixed_a(-0.020909911021590233)),(to_sfixed_a(0.05739913135766983)),(to_sfixed_a(0.07240770757198334)),(to_sfixed_a(-0.06870610266923904)),(to_sfixed_a(-0.2525152266025543)),(to_sfixed_a(0.030685806646943092)),(to_sfixed_a(0.0006196548929437995)),(to_sfixed_a(-0.18054978549480438)),(to_sfixed_a(-0.0091312937438488)),(to_sfixed_a(-0.2473258227109909)),(to_sfixed_a(0.20725665986537933)),(to_sfixed_a(-0.1764872521162033)),(to_sfixed_a(0.02126338705420494)),(to_sfixed_a(0.0470692403614521)),(to_sfixed_a(0.015561697073280811)),(to_sfixed_a(-0.0560673289000988)),(to_sfixed_a(0.021762799471616745)),(to_sfixed_a(-0.14913302659988403)),(to_sfixed_a(0.04770006611943245)),(to_sfixed_a(-0.044709425419569016)),(to_sfixed_a(-0.030745776370167732)),(to_sfixed_a(7.681834540562704e-05)),(to_sfixed_a(-0.00016221652913372964)),(to_sfixed_a(0.00027426762972027063)),(to_sfixed_a(-2.0802861399715766e-05)),(to_sfixed_a(0.00010975446639349684)),(to_sfixed_a(0.0002304131630808115)),(to_sfixed_a(-0.0033903908915817738)),(to_sfixed_a(0.15762671828269958)),(to_sfixed_a(0.11844495683908463)),(to_sfixed_a(-0.03651195764541626)),(to_sfixed_a(0.02904103882610798)),(to_sfixed_a(-0.07100037485361099)),(to_sfixed_a(0.005244469735771418)),(to_sfixed_a(0.09080135822296143)),(to_sfixed_a(-0.34058427810668945)),(to_sfixed_a(0.006511251907795668)),(to_sfixed_a(-0.16090945899486542)),(to_sfixed_a(0.04962240532040596)),(to_sfixed_a(-0.12642303109169006)),(to_sfixed_a(-0.08721126616001129)),(to_sfixed_a(-0.22041961550712585)),(to_sfixed_a(0.10857818275690079)),(to_sfixed_a(0.030932899564504623)),(to_sfixed_a(-0.11666633933782578)),(to_sfixed_a(-0.07485195994377136)),(to_sfixed_a(-0.036311399191617966)),(to_sfixed_a(-0.10578804463148117)),(to_sfixed_a(-0.00017105057486332953)),(to_sfixed_a(0.0002800889778882265)),(to_sfixed_a(-6.661169027211145e-05)),(to_sfixed_a(3.278064468759112e-05)),(to_sfixed_a(7.25032077752985e-05)),(to_sfixed_a(5.7702010963112116e-05)),(to_sfixed_a(-0.00027592838159762323)),(to_sfixed_a(-0.008174271322786808)),(to_sfixed_a(0.04789947345852852)),(to_sfixed_a(0.13140438497066498)),(to_sfixed_a(-0.02965395525097847)),(to_sfixed_a(0.01919218711555004)),(to_sfixed_a(0.1424449235200882)),(to_sfixed_a(-0.28323256969451904)),(to_sfixed_a(-0.23400761187076569)),(to_sfixed_a(-0.12567633390426636)),(to_sfixed_a(-0.15568988025188446)),(to_sfixed_a(0.1665995717048645)),(to_sfixed_a(0.21776072680950165)),(to_sfixed_a(0.07223228365182877)),(to_sfixed_a(-0.15446960926055908)),(to_sfixed_a(0.04584461823105812)),(to_sfixed_a(0.025591403245925903)),(to_sfixed_a(0.1924332231283188)),(to_sfixed_a(0.12577587366104126)),(to_sfixed_a(-0.11776454001665115)),(to_sfixed_a(-0.08425664156675339)),(to_sfixed_a(-0.19117675721645355)),(to_sfixed_a(-0.028675345703959465)),(to_sfixed_a(-5.001391036785208e-05)),(to_sfixed_a(6.474826659541577e-05)),(to_sfixed_a(0.00012081852037226781)),(to_sfixed_a(0.000245071278186515)),(to_sfixed_a(9.00764498510398e-05)),(to_sfixed_a(0.00863696914166212)),(to_sfixed_a(0.15695251524448395)),(to_sfixed_a(-0.06911136955022812)),(to_sfixed_a(-0.1182747483253479)),(to_sfixed_a(-0.32224205136299133)),(to_sfixed_a(-0.1203211322426796)),(to_sfixed_a(-0.0149606391787529)),(to_sfixed_a(-0.028295814990997314)),(to_sfixed_a(-0.25613993406295776)),(to_sfixed_a(-0.29702720046043396)),(to_sfixed_a(0.06451807916164398)),(to_sfixed_a(0.05239500105381012)),(to_sfixed_a(0.26065340638160706)),(to_sfixed_a(0.04389648139476776)),(to_sfixed_a(0.06858538836240768)),(to_sfixed_a(-0.06496483832597733)),(to_sfixed_a(-0.01888723112642765)),(to_sfixed_a(0.06833220273256302)),(to_sfixed_a(-0.11219225078821182)),(to_sfixed_a(0.06522410362958908)),(to_sfixed_a(-0.021529069170355797)),(to_sfixed_a(-0.18369999527931213)),(to_sfixed_a(0.0001043963129632175)),(to_sfixed_a(-0.00020161693100817502)),(to_sfixed_a(0.00020628640777431428)),(to_sfixed_a(-5.5140168115030974e-05)),(to_sfixed_a(0.00030523582245223224)),(to_sfixed_a(-3.7436540878843516e-05)),(to_sfixed_a(-2.9438184355967678e-05)),(to_sfixed_a(-0.11155444383621216)),(to_sfixed_a(-0.06218530982732773)),(to_sfixed_a(0.022560128942131996)),(to_sfixed_a(-0.23378176987171173)),(to_sfixed_a(-0.052237361669540405)),(to_sfixed_a(0.0821155533194542)),(to_sfixed_a(0.06102835386991501)),(to_sfixed_a(-0.1548730432987213)),(to_sfixed_a(0.1401333063840866)),(to_sfixed_a(-0.017198750749230385)),(to_sfixed_a(-0.08726760745048523)),(to_sfixed_a(-0.06647126376628876)),(to_sfixed_a(0.2280881255865097)),(to_sfixed_a(-0.04049720987677574)),(to_sfixed_a(-0.0037701199762523174)),(to_sfixed_a(-0.34485697746276855)),(to_sfixed_a(-0.005585567560046911)),(to_sfixed_a(-0.016383826732635498)),(to_sfixed_a(-0.09539927542209625)),(to_sfixed_a(0.0915367379784584)),(to_sfixed_a(0.19067855179309845)),(to_sfixed_a(-3.3354939660057425e-05)),(to_sfixed_a(8.603602327639237e-05)),(to_sfixed_a(-0.0001579667441546917)),(to_sfixed_a(-0.0001683542359387502)),(to_sfixed_a(2.3124450308387168e-05)),(to_sfixed_a(0.00013730608043260872)),(to_sfixed_a(-0.00011032123438781127)),(to_sfixed_a(0.017577864229679108)),(to_sfixed_a(0.3094046413898468)),(to_sfixed_a(0.17768211662769318)),(to_sfixed_a(0.11017709970474243)),(to_sfixed_a(-0.12100809067487717)),(to_sfixed_a(0.08582709729671478)),(to_sfixed_a(0.005527353845536709)),(to_sfixed_a(-0.04673777520656586)),(to_sfixed_a(-0.14414085447788239)),(to_sfixed_a(-0.2197561413049698)),(to_sfixed_a(0.1081867665052414)),(to_sfixed_a(0.0661223903298378)),(to_sfixed_a(-0.022612901404500008)),(to_sfixed_a(0.03134362772107124)),(to_sfixed_a(0.0049207089468836784)),(to_sfixed_a(0.0205130223184824)),(to_sfixed_a(-0.1334802210330963)),(to_sfixed_a(-0.059249114245176315)),(to_sfixed_a(0.06741289794445038)),(to_sfixed_a(0.29080161452293396)),(to_sfixed_a(-0.01054106093943119)),(to_sfixed_a(0.0033123421017080545)),(to_sfixed_a(0.003984073176980019)),(to_sfixed_a(0.0002189108490711078)),(to_sfixed_a(-8.345827154698782e-06)),(to_sfixed_a(9.431238140678033e-05)),(to_sfixed_a(-0.00025969199487008154)),(to_sfixed_a(-0.00022887876548338681)),(to_sfixed_a(-0.0022556516341865063)),(to_sfixed_a(-0.18278154730796814)),(to_sfixed_a(-0.0564558170735836)),(to_sfixed_a(-0.07637440413236618)),(to_sfixed_a(-0.3353980481624603)),(to_sfixed_a(0.12789827585220337)),(to_sfixed_a(-0.15575620532035828)),(to_sfixed_a(-0.03465179726481438)),(to_sfixed_a(-0.308187335729599)),(to_sfixed_a(-0.09543883800506592)),(to_sfixed_a(-0.1667911857366562)),(to_sfixed_a(-0.01876380294561386)),(to_sfixed_a(-0.10709226131439209)),(to_sfixed_a(-0.0865432396531105)),(to_sfixed_a(0.09542150050401688)),(to_sfixed_a(-0.2970161437988281)),(to_sfixed_a(0.03310111165046692)),(to_sfixed_a(-0.04085146263241768)),(to_sfixed_a(-0.0720210000872612)),(to_sfixed_a(-0.05390245467424393)),(to_sfixed_a(0.07059715688228607)),(to_sfixed_a(-0.00039090175414457917)),(to_sfixed_a(-8.924851135816425e-05)),(to_sfixed_a(2.58678355748998e-05)),(to_sfixed_a(0.0001834233698900789)),(to_sfixed_a(-0.00021397232194431126)),(to_sfixed_a(-3.143620415357873e-05)),(to_sfixed_a(0.00020693353144451976)),(to_sfixed_a(-0.03311583027243614)),(to_sfixed_a(-0.19275832176208496)),(to_sfixed_a(-0.09165656566619873)),(to_sfixed_a(-0.058953311294317245)),(to_sfixed_a(-0.07636290043592453)),(to_sfixed_a(-0.18447627127170563)),(to_sfixed_a(0.03973674774169922)),(to_sfixed_a(0.18257655203342438)),(to_sfixed_a(-0.1629517823457718)),(to_sfixed_a(-0.15255314111709595)),(to_sfixed_a(0.1866319328546524)),(to_sfixed_a(-0.0076370760798454285)),(to_sfixed_a(-0.04173152148723602)),(to_sfixed_a(0.08077305555343628)),(to_sfixed_a(-0.05757131054997444)),(to_sfixed_a(0.3821927607059479)),(to_sfixed_a(0.041385501623153687)),(to_sfixed_a(0.036383938044309616)),(to_sfixed_a(-0.030469704419374466)),(to_sfixed_a(-0.05225098878145218)),(to_sfixed_a(-0.09420386701822281)),(to_sfixed_a(-0.0002399160439381376)),(to_sfixed_a(-0.00024540466256439686)),(to_sfixed_a(-4.476879985304549e-05)),(to_sfixed_a(4.393606286612339e-05)),(to_sfixed_a(-0.00013664213474839926)),(to_sfixed_a(-9.525342647975776e-06)),(to_sfixed_a(0.0011543172877281904)),(to_sfixed_a(-0.04190153256058693)),(to_sfixed_a(-0.06983841955661774)),(to_sfixed_a(0.2594474256038666)),(to_sfixed_a(-0.1412207931280136)),(to_sfixed_a(-0.033738769590854645)),(to_sfixed_a(0.10816653817892075)),(to_sfixed_a(-0.13088954985141754)),(to_sfixed_a(-0.0820608139038086)),(to_sfixed_a(-0.0787457525730133)),(to_sfixed_a(0.06411077827215195)),(to_sfixed_a(0.13910514116287231)),(to_sfixed_a(0.03666769713163376)),(to_sfixed_a(0.17032556235790253)),(to_sfixed_a(0.05042000859975815)),(to_sfixed_a(-0.14040036499500275)),(to_sfixed_a(0.036800023168325424)),(to_sfixed_a(-0.4437674582004547)),(to_sfixed_a(-0.1400931179523468)),(to_sfixed_a(-0.15631839632987976)),(to_sfixed_a(0.013073193840682507)),(to_sfixed_a(-0.02711801789700985)),(to_sfixed_a(-0.0020382441580295563)),(to_sfixed_a(4.235217784298584e-05)),(to_sfixed_a(6.559232133440673e-05)),(to_sfixed_a(5.806893022963777e-05)),(to_sfixed_a(2.906977715610992e-05)),(to_sfixed_a(0.000786357675679028)),(to_sfixed_a(0.001326213008724153)),(to_sfixed_a(-0.14897353947162628)),(to_sfixed_a(-0.1521713137626648)),(to_sfixed_a(0.13936837017536163)),(to_sfixed_a(0.41415587067604065)),(to_sfixed_a(-0.12786930799484253)),(to_sfixed_a(-0.08744335174560547)),(to_sfixed_a(0.342824250459671)),(to_sfixed_a(0.048812150955200195)),(to_sfixed_a(0.2669486105442047)),(to_sfixed_a(0.19590184092521667)),(to_sfixed_a(0.22279690206050873)),(to_sfixed_a(0.032540012151002884)),(to_sfixed_a(-0.10769931226968765)),(to_sfixed_a(0.16633039712905884)),(to_sfixed_a(0.19612126052379608)),(to_sfixed_a(0.22141744196414948)),(to_sfixed_a(0.022091301158070564)),(to_sfixed_a(-0.12418970465660095)),(to_sfixed_a(0.010462949983775616)),(to_sfixed_a(0.023333372548222542)),(to_sfixed_a(6.545090582221746e-05)),(to_sfixed_a(-0.0002819414949044585)),(to_sfixed_a(9.263665560865775e-05)),(to_sfixed_a(9.025659892358817e-06)),(to_sfixed_a(-0.0001810553076211363)),(to_sfixed_a(-0.00021057864069007337)),(to_sfixed_a(1.970538323803339e-05)),(to_sfixed_a(-0.04782478138804436)),(to_sfixed_a(-0.14142990112304688)),(to_sfixed_a(-0.18657678365707397)),(to_sfixed_a(-0.08727846294641495)),(to_sfixed_a(0.06711170077323914)),(to_sfixed_a(0.24298420548439026)),(to_sfixed_a(0.004922022577375174)),(to_sfixed_a(-0.21945390105247498)),(to_sfixed_a(-0.4004337787628174)),(to_sfixed_a(-0.08469138294458389)),(to_sfixed_a(0.27370598912239075)),(to_sfixed_a(-0.12234128266572952)),(to_sfixed_a(0.04368283227086067)),(to_sfixed_a(0.004351820796728134)),(to_sfixed_a(0.24555133283138275)),(to_sfixed_a(0.007982033304870129)),(to_sfixed_a(-0.11497195065021515)),(to_sfixed_a(-0.1235538199543953)),(to_sfixed_a(0.019253848120570183)),(to_sfixed_a(-0.07193409651517868)),(to_sfixed_a(-0.0684918463230133)),(to_sfixed_a(-0.03671446442604065)),(to_sfixed_a(-4.673115836340003e-05)),(to_sfixed_a(-2.0994410078856163e-05)),(to_sfixed_a(0.0001449619303457439)),(to_sfixed_a(-0.00019733470981009305)),(to_sfixed_a(4.5131459046388045e-05)),(to_sfixed_a(0.00015218491898849607)),(to_sfixed_a(-0.01114098634570837)),(to_sfixed_a(0.0016326219774782658)),(to_sfixed_a(-0.021379681304097176)),(to_sfixed_a(0.03800645470619202)),(to_sfixed_a(0.07300923019647598)),(to_sfixed_a(0.1741705983877182)),(to_sfixed_a(0.18886537849903107)),(to_sfixed_a(0.1038249284029007)),(to_sfixed_a(-0.10404026508331299)),(to_sfixed_a(-0.20402543246746063)),(to_sfixed_a(-0.014520996250212193)),(to_sfixed_a(0.14517618715763092)),(to_sfixed_a(0.08686797320842743)),(to_sfixed_a(0.03949863463640213)),(to_sfixed_a(-0.09968294948339462)),(to_sfixed_a(-0.1273888200521469)),(to_sfixed_a(0.030486779287457466)),(to_sfixed_a(-0.011281708255410194)),(to_sfixed_a(0.07134205847978592)),(to_sfixed_a(-0.014466200955212116)),(to_sfixed_a(0.025697194039821625)),(to_sfixed_a(0.00016095487808343023)),(to_sfixed_a(-4.7446825192309916e-05)),(to_sfixed_a(-0.0001160983374575153)),(to_sfixed_a(0.00019416341092437506)),(to_sfixed_a(-7.94316019891994e-06)),(to_sfixed_a(-6.378314719768241e-05)),(to_sfixed_a(0.0001449708070140332)),(to_sfixed_a(3.8101497921161354e-05)),(to_sfixed_a(0.012105504050850868)),(to_sfixed_a(-0.03499707579612732)),(to_sfixed_a(-0.12092127650976181)),(to_sfixed_a(0.37116944789886475)),(to_sfixed_a(0.10225903242826462)),(to_sfixed_a(-0.08742546290159225)),(to_sfixed_a(0.015953708440065384)),(to_sfixed_a(0.047426700592041016)),(to_sfixed_a(-0.07681483030319214)),(to_sfixed_a(0.031775735318660736)),(to_sfixed_a(-0.28731516003608704)),(to_sfixed_a(0.046941958367824554)),(to_sfixed_a(-0.017615843564271927)),(to_sfixed_a(-0.05426885560154915)),(to_sfixed_a(-0.44740551710128784)),(to_sfixed_a(0.013892842456698418)),(to_sfixed_a(0.20386214554309845)),(to_sfixed_a(-0.03999069333076477)),(to_sfixed_a(0.007239798083901405)),(to_sfixed_a(0.10595967620611191)),(to_sfixed_a(0.14633473753929138)),(to_sfixed_a(-3.6657755117630586e-05)),(to_sfixed_a(4.618826278601773e-05)),(to_sfixed_a(0.00012397152022458613)),(to_sfixed_a(9.40298632485792e-05)),(to_sfixed_a(0.0002119302371283993)),(to_sfixed_a(-4.4783231714973226e-05)),(to_sfixed_a(0.00026838938356377184)),(to_sfixed_a(0.011922073550522327)),(to_sfixed_a(0.00018134246056433767)),(to_sfixed_a(-0.09315373748540878)),(to_sfixed_a(0.07981285452842712)),(to_sfixed_a(-0.23293565213680267)),(to_sfixed_a(-0.12184949964284897)),(to_sfixed_a(-0.023156223818659782)),(to_sfixed_a(-0.09583106637001038)),(to_sfixed_a(0.03779471293091774)),(to_sfixed_a(0.0777057632803917)),(to_sfixed_a(0.0002998335985466838)),(to_sfixed_a(-0.20177911221981049)),(to_sfixed_a(0.05090966075658798)),(to_sfixed_a(-0.08745915442705154)),(to_sfixed_a(-0.2855875492095947)),(to_sfixed_a(-0.0941564217209816)),(to_sfixed_a(0.26621493697166443)),(to_sfixed_a(0.025186149403452873)),(to_sfixed_a(-0.058039937168359756)),(to_sfixed_a(0.0007146333809942007)),(to_sfixed_a(-0.04825032129883766)),(to_sfixed_a(-2.8529178962344304e-05)),(to_sfixed_a(7.849769463064149e-05)),(to_sfixed_a(0.0003566565574146807)),(to_sfixed_a(-0.00016829425294417888)),(to_sfixed_a(-0.00020631799998227507)),(to_sfixed_a(-0.0001545010891277343)),(to_sfixed_a(0.0002815229818224907)),(to_sfixed_a(-1.7857979401014745e-05)),(to_sfixed_a(-0.04236586019396782)),(to_sfixed_a(0.12418334186077118)),(to_sfixed_a(-0.10923215001821518)),(to_sfixed_a(0.013381551019847393)),(to_sfixed_a(-0.061787981539964676)),(to_sfixed_a(0.005843574646860361)),(to_sfixed_a(0.14958326518535614)),(to_sfixed_a(0.212044820189476)),(to_sfixed_a(0.05396995693445206)),(to_sfixed_a(0.015982307493686676)),(to_sfixed_a(0.19949062168598175)),(to_sfixed_a(-0.07330404222011566)),(to_sfixed_a(0.017358554527163506)),(to_sfixed_a(-0.10978661477565765)),(to_sfixed_a(-0.03366231545805931)),(to_sfixed_a(-0.0671946257352829)),(to_sfixed_a(-0.0012905538314953446)),(to_sfixed_a(-0.03562704473733902)),(to_sfixed_a(-0.002311933785676956)),(to_sfixed_a(-0.00013223894347902387)),(to_sfixed_a(0.0002483432472217828)),(to_sfixed_a(-0.0001900609495351091)),(to_sfixed_a(4.660641207010485e-05)),(to_sfixed_a(-8.017272921279073e-05)),(to_sfixed_a(-0.00010703552834456787)),(to_sfixed_a(-0.0001147395305451937)),(to_sfixed_a(0.00011223852925468236)),(to_sfixed_a(-1.554623509036901e-06)),(to_sfixed_a(0.006677032448351383)),(to_sfixed_a(0.21903498470783234)),(to_sfixed_a(0.26666736602783203)),(to_sfixed_a(-0.15839883685112)),(to_sfixed_a(-0.13284973800182343)),(to_sfixed_a(0.12794749438762665)),(to_sfixed_a(0.20122100412845612)),(to_sfixed_a(0.18338139355182648)),(to_sfixed_a(0.14996422827243805)),(to_sfixed_a(0.029751725494861603)),(to_sfixed_a(0.0938263013958931)),(to_sfixed_a(0.2379962056875229)),(to_sfixed_a(-0.21603061258792877)),(to_sfixed_a(-0.06832371652126312)),(to_sfixed_a(-0.11950844526290894)),(to_sfixed_a(0.03038899600505829)),(to_sfixed_a(-0.08905816078186035)),(to_sfixed_a(-0.0031855779234319925)),(to_sfixed_a(-0.06098377704620361)),(to_sfixed_a(4.9047077482100576e-05)),(to_sfixed_a(-0.00010994987678714097)),(to_sfixed_a(7.071314757922664e-05)),(to_sfixed_a(3.502497565932572e-05)),(to_sfixed_a(-6.199502240633592e-05)),(to_sfixed_a(6.234296597540379e-05)),(to_sfixed_a(1.1351207831467036e-05)),(to_sfixed_a(1.1409729268052615e-06)),(to_sfixed_a(0.031172674149274826)),(to_sfixed_a(0.06413954496383667)),(to_sfixed_a(0.13111111521720886)),(to_sfixed_a(0.19067928194999695)),(to_sfixed_a(0.17287009954452515)),(to_sfixed_a(0.09635550528764725)),(to_sfixed_a(0.1097196564078331)),(to_sfixed_a(0.39895138144493103)),(to_sfixed_a(0.17183972895145416)),(to_sfixed_a(0.23944172263145447)),(to_sfixed_a(0.24973970651626587)),(to_sfixed_a(-0.05708009749650955)),(to_sfixed_a(-0.08109764009714127)),(to_sfixed_a(-0.211222305893898)),(to_sfixed_a(-0.15521618723869324)),(to_sfixed_a(-0.13716939091682434)),(to_sfixed_a(-0.004528935067355633)),(to_sfixed_a(-0.05164425075054169)),(to_sfixed_a(-0.035029370337724686)),(to_sfixed_a(0.0004155414062552154)),(to_sfixed_a(-0.00010237949027214199)),(to_sfixed_a(-0.00016354175750166178)),(to_sfixed_a(4.588594674714841e-05)),(to_sfixed_a(-0.00011241959873586893)),(to_sfixed_a(-0.0002715769223868847)),(to_sfixed_a(0.00010929053678410128)),(to_sfixed_a(-0.00020315490837674588)),(to_sfixed_a(6.168138497741893e-05)),(to_sfixed_a(-0.0001557948417030275)),(to_sfixed_a(0.033010367304086685)),(to_sfixed_a(0.0782206803560257)),(to_sfixed_a(0.05633290857076645)),(to_sfixed_a(0.20459268987178802)),(to_sfixed_a(0.13490793108940125)),(to_sfixed_a(0.2720469534397125)),(to_sfixed_a(0.07838620990514755)),(to_sfixed_a(-0.05367041751742363)),(to_sfixed_a(-0.036483801901340485)),(to_sfixed_a(0.09927093982696533)),(to_sfixed_a(0.09194100648164749)),(to_sfixed_a(-0.27973097562789917)),(to_sfixed_a(0.02792162261903286)),(to_sfixed_a(-0.0019342608284205198)),(to_sfixed_a(0.018860170617699623)),(to_sfixed_a(0.0517691969871521)),(to_sfixed_a(0.0006933800177648664)),(to_sfixed_a(0.0035607723984867334)),(to_sfixed_a(0.003626491641625762)),(to_sfixed_a(6.176168244564906e-05)),(to_sfixed_a(0.00012923240137752146)),(to_sfixed_a(4.358097066869959e-05)),(to_sfixed_a(-5.966818571323529e-05)),(to_sfixed_a(8.771420652919915e-06)),(to_sfixed_a(-0.00020995309751015157)),(to_sfixed_a(7.018560427241027e-05)),(to_sfixed_a(0.0001618043752387166)),(to_sfixed_a(-0.0001398866588715464)),(to_sfixed_a(0.00019803130999207497)),(to_sfixed_a(8.101030834950507e-05)),(to_sfixed_a(-0.00010472087888047099)),(to_sfixed_a(0.00020749376562889665)),(to_sfixed_a(0.0001838015450630337)),(to_sfixed_a(0.005903182085603476)),(to_sfixed_a(2.0744266294059344e-05)),(to_sfixed_a(-0.00022421810717787594)),(to_sfixed_a(0.015527268871665001)),(to_sfixed_a(-0.04703077673912048)),(to_sfixed_a(0.00428682891651988)),(to_sfixed_a(-0.01460761297494173)),(to_sfixed_a(0.0036272930447012186)),(to_sfixed_a(0.001393587444908917)),(to_sfixed_a(-0.00022806735069025308)),(to_sfixed_a(0.0014858768554404378)),(to_sfixed_a(-8.71011616254691e-06)),(to_sfixed_a(-8.864609117154032e-05)),(to_sfixed_a(-0.0001621125848032534)),(to_sfixed_a(-0.00011307349632261321)),(to_sfixed_a(-2.7320242224959657e-05)),(to_sfixed_a(9.70721521298401e-05)),(to_sfixed_a(0.0002879289095290005)),(to_sfixed_a(7.575712515972555e-05)),(to_sfixed_a(-3.35640215780586e-05)),(to_sfixed_a(-0.0002161585580324754)),(to_sfixed_a(7.821864710422233e-05)),(to_sfixed_a(0.00029139002435840666)),(to_sfixed_a(-7.062646909616888e-05)),(to_sfixed_a(-3.936321445507929e-05)),(to_sfixed_a(-0.00010459913755767047)),(to_sfixed_a(0.0001273179950658232)),(to_sfixed_a(-7.989656296558678e-05)),(to_sfixed_a(8.486200385959819e-06)),(to_sfixed_a(0.0004111240559723228)),(to_sfixed_a(-0.0001818994351197034)),(to_sfixed_a(-0.0001414269208908081)),(to_sfixed_a(-6.625885725952685e-05)),(to_sfixed_a(-5.829032670590095e-05)),(to_sfixed_a(-0.0001516850752523169)),(to_sfixed_a(-0.0001690880162641406)),(to_sfixed_a(-9.330510511063039e-05)),(to_sfixed_a(0.00011002090468537062)),(to_sfixed_a(4.978364449925721e-05)),(to_sfixed_a(-1.140183667303063e-05)),(to_sfixed_a(7.022186036920175e-05)),(to_sfixed_a(0.0001527986314613372)),(to_sfixed_a(-0.00017032015603035688)),(to_sfixed_a(-0.0001063186427927576)),(to_sfixed_a(0.00012932418030686677)),(to_sfixed_a(-6.275979103520513e-05)));

    constant weight_n0_30 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(5.995195169816725e-05)),(to_sfixed_a(9.513008990325034e-05)),(to_sfixed_a(-0.0002548981865402311)),(to_sfixed_a(1.9914516087737866e-05)),(to_sfixed_a(-0.0001865003869170323)),(to_sfixed_a(-6.267474236665294e-05)),(to_sfixed_a(-3.947301229345612e-05)),(to_sfixed_a(-0.0002887072041630745)),(to_sfixed_a(-2.18551758734975e-05)),(to_sfixed_a(-0.00022211538453120738)),(to_sfixed_a(3.561260018614121e-05)),(to_sfixed_a(-0.0001325562479905784)),(to_sfixed_a(-0.000249084725510329)),(to_sfixed_a(3.1190844310913235e-05)),(to_sfixed_a(-0.0003786127199418843)),(to_sfixed_a(2.253138882224448e-05)),(to_sfixed_a(0.00022543713566847146)),(to_sfixed_a(-0.00013850290270056576)),(to_sfixed_a(9.185940871248022e-05)),(to_sfixed_a(-6.429538188967854e-06)),(to_sfixed_a(2.1243129594950005e-05)),(to_sfixed_a(-8.613317186245695e-05)),(to_sfixed_a(-7.077434929669835e-06)),(to_sfixed_a(-0.00010300211579306051)),(to_sfixed_a(6.390109047060832e-05)),(to_sfixed_a(-0.00018231815192848444)),(to_sfixed_a(-4.042478394694626e-05)),(to_sfixed_a(1.4869458027533256e-05)),(to_sfixed_a(0.00014997863036114722)),(to_sfixed_a(-9.399009286426008e-05)),(to_sfixed_a(9.051612869370729e-05)),(to_sfixed_a(0.00015451900253538042)),(to_sfixed_a(-0.00021070432558190078)),(to_sfixed_a(-4.6124823711579666e-05)),(to_sfixed_a(7.972442836035043e-05)),(to_sfixed_a(-3.372139690327458e-05)),(to_sfixed_a(-0.00010452159040141851)),(to_sfixed_a(-0.00013382422912400216)),(to_sfixed_a(-7.073186679917853e-06)),(to_sfixed_a(-0.00030229255207814276)),(to_sfixed_a(-0.0002078348770737648)),(to_sfixed_a(-0.00023521548428107053)),(to_sfixed_a(-0.00022545717365574092)),(to_sfixed_a(3.015992660948541e-05)),(to_sfixed_a(0.0001762126194080338)),(to_sfixed_a(-1.155496920546284e-05)),(to_sfixed_a(4.927023474010639e-05)),(to_sfixed_a(-3.8521349779330194e-05)),(to_sfixed_a(0.00011409250873839483)),(to_sfixed_a(-0.00034378498094156384)),(to_sfixed_a(0.00013399311865214258)),(to_sfixed_a(-0.00031682534608989954)),(to_sfixed_a(8.028178126551211e-05)),(to_sfixed_a(-0.00012592034181579947)),(to_sfixed_a(0.00017025764100253582)),(to_sfixed_a(-2.5517445465084165e-05)),(to_sfixed_a(0.00020392442820593715)),(to_sfixed_a(0.00019922404317185283)),(to_sfixed_a(4.116200943826698e-05)),(to_sfixed_a(-8.940422412706539e-05)),(to_sfixed_a(0.00015560179599560797)),(to_sfixed_a(-0.0001944918476510793)),(to_sfixed_a(0.0001506399712525308)),(to_sfixed_a(0.0002593646931927651)),(to_sfixed_a(0.00015645610983483493)),(to_sfixed_a(0.00011983102012891322)),(to_sfixed_a(-2.065564103759243e-06)),(to_sfixed_a(-6.564677460119128e-05)),(to_sfixed_a(-0.00022905704099684954)),(to_sfixed_a(0.009311962872743607)),(to_sfixed_a(-4.9256930651608855e-05)),(to_sfixed_a(0.00020704031339846551)),(to_sfixed_a(-0.00016378566215280443)),(to_sfixed_a(-1.4527107850881293e-05)),(to_sfixed_a(-0.00020434973703231663)),(to_sfixed_a(8.989017078420147e-05)),(to_sfixed_a(-2.9026650736341253e-05)),(to_sfixed_a(-0.00013591091556008905)),(to_sfixed_a(-0.000129003994516097)),(to_sfixed_a(0.000329373317072168)),(to_sfixed_a(-0.00015018768317531794)),(to_sfixed_a(-1.871945642051287e-05)),(to_sfixed_a(9.744057024363428e-05)),(to_sfixed_a(5.543747101910412e-05)),(to_sfixed_a(1.357981363980798e-05)),(to_sfixed_a(0.0002529807388782501)),(to_sfixed_a(-8.549758786102757e-05)),(to_sfixed_a(-0.0002396100026089698)),(to_sfixed_a(-7.352290595008526e-06)),(to_sfixed_a(-1.2248963685124181e-05)),(to_sfixed_a(-8.604955655755475e-05)),(to_sfixed_a(-0.0002577301347628236)),(to_sfixed_a(-0.00596463680267334)),(to_sfixed_a(4.088547939318232e-05)),(to_sfixed_a(-0.006679490674287081)),(to_sfixed_a(0.09514734894037247)),(to_sfixed_a(-0.01636999286711216)),(to_sfixed_a(0.17874841392040253)),(to_sfixed_a(-0.06767395883798599)),(to_sfixed_a(-0.11587409675121307)),(to_sfixed_a(0.017160266637802124)),(to_sfixed_a(-0.024303752928972244)),(to_sfixed_a(-0.009919706732034683)),(to_sfixed_a(0.02328597567975521)),(to_sfixed_a(0.0023728609085083008)),(to_sfixed_a(0.004861206281930208)),(to_sfixed_a(3.08641538140364e-05)),(to_sfixed_a(0.00018222643120680004)),(to_sfixed_a(-0.00013522992958314717)),(to_sfixed_a(3.6075951356906444e-05)),(to_sfixed_a(-0.0001954878680408001)),(to_sfixed_a(0.0001463063235860318)),(to_sfixed_a(-0.00019089320267084986)),(to_sfixed_a(-1.2909996257803869e-05)),(to_sfixed_a(-3.0989322112873197e-05)),(to_sfixed_a(-0.00010872832353925332)),(to_sfixed_a(-0.00020848003623541445)),(to_sfixed_a(-0.00010339564323658124)),(to_sfixed_a(0.0004931568400934339)),(to_sfixed_a(0.04531596973538399)),(to_sfixed_a(0.020373070612549782)),(to_sfixed_a(-0.014934767037630081)),(to_sfixed_a(0.3333325684070587)),(to_sfixed_a(0.04823649674654007)),(to_sfixed_a(0.18554647266864777)),(to_sfixed_a(0.026990480720996857)),(to_sfixed_a(0.12272577732801437)),(to_sfixed_a(0.12634283304214478)),(to_sfixed_a(0.11443400382995605)),(to_sfixed_a(0.0044938912615180016)),(to_sfixed_a(0.004540227819234133)),(to_sfixed_a(0.03521546348929405)),(to_sfixed_a(-0.01825595274567604)),(to_sfixed_a(0.03291332721710205)),(to_sfixed_a(-0.007502967957407236)),(to_sfixed_a(6.976328677410493e-06)),(to_sfixed_a(-0.0006734690396115184)),(to_sfixed_a(-0.0001404242211719975)),(to_sfixed_a(-0.00021562153415288776)),(to_sfixed_a(-5.488780152518302e-05)),(to_sfixed_a(0.0001580760581418872)),(to_sfixed_a(0.000274190359050408)),(to_sfixed_a(-2.104752820741851e-05)),(to_sfixed_a(-0.00011753961734939367)),(to_sfixed_a(0.0002963792940136045)),(to_sfixed_a(0.06357400864362717)),(to_sfixed_a(0.0005828283028677106)),(to_sfixed_a(0.02118712104856968)),(to_sfixed_a(0.08265134692192078)),(to_sfixed_a(0.07745412737131119)),(to_sfixed_a(0.012026500888168812)),(to_sfixed_a(0.10977014899253845)),(to_sfixed_a(-0.15571968257427216)),(to_sfixed_a(-0.33917325735092163)),(to_sfixed_a(-0.1211489662528038)),(to_sfixed_a(-0.25130870938301086)),(to_sfixed_a(-0.060493409633636475)),(to_sfixed_a(-0.3407427668571472)),(to_sfixed_a(-0.03791217505931854)),(to_sfixed_a(-0.18570944666862488)),(to_sfixed_a(-0.10849427431821823)),(to_sfixed_a(0.05757622420787811)),(to_sfixed_a(-0.0019349176436662674)),(to_sfixed_a(-0.011922555975615978)),(to_sfixed_a(0.0014809968415647745)),(to_sfixed_a(0.00029872756567783654)),(to_sfixed_a(0.00026642956072464585)),(to_sfixed_a(-5.368422353058122e-05)),(to_sfixed_a(5.4871059546712786e-05)),(to_sfixed_a(-9.472934152654489e-07)),(to_sfixed_a(-6.62568854750134e-05)),(to_sfixed_a(4.7220190026564524e-05)),(to_sfixed_a(0.00019192528270650655)),(to_sfixed_a(0.0618518590927124)),(to_sfixed_a(0.01696493849158287)),(to_sfixed_a(-0.008125507272779942)),(to_sfixed_a(-0.06008242070674896)),(to_sfixed_a(-0.12288959324359894)),(to_sfixed_a(0.006590061355382204)),(to_sfixed_a(0.011995482258498669)),(to_sfixed_a(0.33636540174484253)),(to_sfixed_a(-0.0640493854880333)),(to_sfixed_a(-0.1201271116733551)),(to_sfixed_a(-0.018010888248682022)),(to_sfixed_a(-0.1604992300271988)),(to_sfixed_a(0.038989901542663574)),(to_sfixed_a(0.18125393986701965)),(to_sfixed_a(-0.06887784600257874)),(to_sfixed_a(0.18216171860694885)),(to_sfixed_a(-0.08778386563062668)),(to_sfixed_a(0.012488791719079018)),(to_sfixed_a(0.11938051134347916)),(to_sfixed_a(0.006416977848857641)),(to_sfixed_a(0.007386524695903063)),(to_sfixed_a(0.0045639099553227425)),(to_sfixed_a(-0.00011573931988095865)),(to_sfixed_a(1.2630238416022621e-05)),(to_sfixed_a(8.17891996121034e-05)),(to_sfixed_a(-0.0001193235075334087)),(to_sfixed_a(7.983366231201217e-05)),(to_sfixed_a(-1.4035775166121311e-05)),(to_sfixed_a(0.04211767762899399)),(to_sfixed_a(0.06496969610452652)),(to_sfixed_a(-0.07201654464006424)),(to_sfixed_a(-0.29676687717437744)),(to_sfixed_a(-0.12173476815223694)),(to_sfixed_a(-0.29078638553619385)),(to_sfixed_a(-0.14355672895908356)),(to_sfixed_a(-0.3426940143108368)),(to_sfixed_a(-0.17815391719341278)),(to_sfixed_a(-0.1031656265258789)),(to_sfixed_a(0.009085150435566902)),(to_sfixed_a(0.06049596518278122)),(to_sfixed_a(-0.05705372244119644)),(to_sfixed_a(0.2550045847892761)),(to_sfixed_a(-0.33221590518951416)),(to_sfixed_a(-0.19579219818115234)),(to_sfixed_a(-0.03931012004613876)),(to_sfixed_a(0.10227926075458527)),(to_sfixed_a(0.16465021669864655)),(to_sfixed_a(0.07484395056962967)),(to_sfixed_a(0.007561410777270794)),(to_sfixed_a(-1.0310269317415077e-05)),(to_sfixed_a(-8.366362453671172e-05)),(to_sfixed_a(3.060084054595791e-05)),(to_sfixed_a(0.00019286497263237834)),(to_sfixed_a(4.315282785682939e-05)),(to_sfixed_a(-0.00018445128807798028)),(to_sfixed_a(0.051146309822797775)),(to_sfixed_a(0.023060791194438934)),(to_sfixed_a(0.03850318118929863)),(to_sfixed_a(0.04161949083209038)),(to_sfixed_a(0.20990628004074097)),(to_sfixed_a(0.05146069824695587)),(to_sfixed_a(-0.07119085639715195)),(to_sfixed_a(0.0679146870970726)),(to_sfixed_a(0.06209219619631767)),(to_sfixed_a(0.33233046531677246)),(to_sfixed_a(-0.25946685671806335)),(to_sfixed_a(-0.11403334140777588)),(to_sfixed_a(0.05071668326854706)),(to_sfixed_a(0.031214505434036255)),(to_sfixed_a(0.18460145592689514)),(to_sfixed_a(0.08774584531784058)),(to_sfixed_a(0.07623022049665451)),(to_sfixed_a(0.25675278902053833)),(to_sfixed_a(-0.08360791951417923)),(to_sfixed_a(0.032518673688173294)),(to_sfixed_a(0.26617133617401123)),(to_sfixed_a(-0.03369995206594467)),(to_sfixed_a(0.0002310312702320516)),(to_sfixed_a(0.0001240493729710579)),(to_sfixed_a(-0.000229534663958475)),(to_sfixed_a(1.4038056178833358e-05)),(to_sfixed_a(-2.18776949623134e-05)),(to_sfixed_a(-0.00039441618719138205)),(to_sfixed_a(0.0004820761096198112)),(to_sfixed_a(0.051472533494234085)),(to_sfixed_a(-0.07265615463256836)),(to_sfixed_a(-0.004182924050837755)),(to_sfixed_a(-0.0411420501768589)),(to_sfixed_a(-0.1028120294213295)),(to_sfixed_a(-0.3354724645614624)),(to_sfixed_a(-0.20652812719345093)),(to_sfixed_a(-0.05644773319363594)),(to_sfixed_a(-0.22924110293388367)),(to_sfixed_a(0.04510029777884483)),(to_sfixed_a(0.07472486793994904)),(to_sfixed_a(-0.2683236002922058)),(to_sfixed_a(-0.0378701314330101)),(to_sfixed_a(0.07965248823165894)),(to_sfixed_a(0.20289133489131927)),(to_sfixed_a(-0.19270552694797516)),(to_sfixed_a(-0.08974165469408035)),(to_sfixed_a(-0.019444165751338005)),(to_sfixed_a(0.016055211424827576)),(to_sfixed_a(0.10007775574922562)),(to_sfixed_a(-9.189242700813338e-05)),(to_sfixed_a(-8.178073039744049e-05)),(to_sfixed_a(-1.4657888414149056e-06)),(to_sfixed_a(5.704072827938944e-05)),(to_sfixed_a(-0.0002193273394368589)),(to_sfixed_a(-9.293823677580804e-05)),(to_sfixed_a(-0.00017270375974476337)),(to_sfixed_a(0.003645971417427063)),(to_sfixed_a(0.07316093146800995)),(to_sfixed_a(0.1748632788658142)),(to_sfixed_a(-0.15922562777996063)),(to_sfixed_a(-0.12687726318836212)),(to_sfixed_a(0.005059765186160803)),(to_sfixed_a(-0.1496773213148117)),(to_sfixed_a(-0.004718979354947805)),(to_sfixed_a(-0.21364304423332214)),(to_sfixed_a(0.2656905949115753)),(to_sfixed_a(-0.2392091602087021)),(to_sfixed_a(-0.04556189849972725)),(to_sfixed_a(-0.019370131194591522)),(to_sfixed_a(-0.05893542617559433)),(to_sfixed_a(0.3193657100200653)),(to_sfixed_a(0.07170826941728592)),(to_sfixed_a(0.12315332889556885)),(to_sfixed_a(0.08175406605005264)),(to_sfixed_a(0.01821023039519787)),(to_sfixed_a(-0.25764036178588867)),(to_sfixed_a(0.1771373599767685)),(to_sfixed_a(0.07194047421216965)),(to_sfixed_a(-7.714382263657171e-06)),(to_sfixed_a(0.00013496687461156398)),(to_sfixed_a(0.0001491490111220628)),(to_sfixed_a(-0.00010020592890214175)),(to_sfixed_a(6.112435221439227e-05)),(to_sfixed_a(0.03858788311481476)),(to_sfixed_a(0.1826266199350357)),(to_sfixed_a(-0.004289939533919096)),(to_sfixed_a(-0.04486587271094322)),(to_sfixed_a(-0.15660937130451202)),(to_sfixed_a(-0.14381051063537598)),(to_sfixed_a(-0.13304917514324188)),(to_sfixed_a(0.048218730837106705)),(to_sfixed_a(0.028519073501229286)),(to_sfixed_a(-0.04672722890973091)),(to_sfixed_a(0.24856144189834595)),(to_sfixed_a(0.029716236516833305)),(to_sfixed_a(0.12912768125534058)),(to_sfixed_a(-0.030497968196868896)),(to_sfixed_a(0.14827165007591248)),(to_sfixed_a(-0.02596915140748024)),(to_sfixed_a(-0.14383564889431)),(to_sfixed_a(0.13622133433818817)),(to_sfixed_a(-0.009638849645853043)),(to_sfixed_a(0.25456926226615906)),(to_sfixed_a(-0.0456230603158474)),(to_sfixed_a(0.026505082845687866)),(to_sfixed_a(-5.865407729288563e-05)),(to_sfixed_a(7.117739005479962e-05)),(to_sfixed_a(-1.784848063834943e-05)),(to_sfixed_a(0.0005678804009221494)),(to_sfixed_a(-0.00015249809075612575)),(to_sfixed_a(1.2294599400775041e-05)),(to_sfixed_a(-0.00013471329293679446)),(to_sfixed_a(-0.036534037441015244)),(to_sfixed_a(-0.1634678989648819)),(to_sfixed_a(-0.18094202876091003)),(to_sfixed_a(-0.21359999477863312)),(to_sfixed_a(0.04179469123482704)),(to_sfixed_a(-0.043141692876815796)),(to_sfixed_a(0.021629462018609047)),(to_sfixed_a(-0.13075754046440125)),(to_sfixed_a(0.21093305945396423)),(to_sfixed_a(-0.02947418764233589)),(to_sfixed_a(-0.06561283767223358)),(to_sfixed_a(0.1537475436925888)),(to_sfixed_a(0.17164935171604156)),(to_sfixed_a(-0.01823590137064457)),(to_sfixed_a(0.06181211397051811)),(to_sfixed_a(0.027446454390883446)),(to_sfixed_a(0.050151411443948746)),(to_sfixed_a(0.047230515629053116)),(to_sfixed_a(0.013716581277549267)),(to_sfixed_a(0.06372468918561935)),(to_sfixed_a(0.11444141715765)),(to_sfixed_a(1.2150598195148632e-05)),(to_sfixed_a(0.0006914034602232277)),(to_sfixed_a(-1.0702214240154717e-05)),(to_sfixed_a(-0.0001415376173099503)),(to_sfixed_a(-5.878560114069842e-05)),(to_sfixed_a(8.83332613739185e-05)),(to_sfixed_a(-2.473989297868684e-05)),(to_sfixed_a(-0.07221734523773193)),(to_sfixed_a(-0.24913141131401062)),(to_sfixed_a(0.024321602657437325)),(to_sfixed_a(0.10333902388811111)),(to_sfixed_a(0.11564669758081436)),(to_sfixed_a(-0.08585769683122635)),(to_sfixed_a(-0.14780767261981964)),(to_sfixed_a(0.17535698413848877)),(to_sfixed_a(0.06847172230482101)),(to_sfixed_a(-0.023319728672504425)),(to_sfixed_a(0.3649630546569824)),(to_sfixed_a(0.1070961281657219)),(to_sfixed_a(0.03455033153295517)),(to_sfixed_a(-0.05565008521080017)),(to_sfixed_a(0.06064480170607567)),(to_sfixed_a(0.273858904838562)),(to_sfixed_a(-0.0738007128238678)),(to_sfixed_a(0.017259327694773674)),(to_sfixed_a(0.027980925515294075)),(to_sfixed_a(0.057770222425460815)),(to_sfixed_a(-0.006086588371545076)),(to_sfixed_a(0.00014455945347435772)),(to_sfixed_a(0.001220356090925634)),(to_sfixed_a(-8.122896542772651e-05)),(to_sfixed_a(4.1343755583511665e-05)),(to_sfixed_a(-1.8930519217974506e-05)),(to_sfixed_a(-0.0005035165813751519)),(to_sfixed_a(0.0001274371170438826)),(to_sfixed_a(0.0010967188281938434)),(to_sfixed_a(0.07680420577526093)),(to_sfixed_a(-0.12500768899917603)),(to_sfixed_a(-0.403109610080719)),(to_sfixed_a(-0.19578781723976135)),(to_sfixed_a(-0.29446497559547424)),(to_sfixed_a(0.21589818596839905)),(to_sfixed_a(0.3244796097278595)),(to_sfixed_a(-0.31009039282798767)),(to_sfixed_a(-0.22562295198440552)),(to_sfixed_a(-0.015107940882444382)),(to_sfixed_a(0.06767220050096512)),(to_sfixed_a(0.15664109587669373)),(to_sfixed_a(-0.07350456714630127)),(to_sfixed_a(0.017718195915222168)),(to_sfixed_a(-0.11561340093612671)),(to_sfixed_a(0.0821373239159584)),(to_sfixed_a(-0.060233525931835175)),(to_sfixed_a(0.007744429633021355)),(to_sfixed_a(0.009495080448687077)),(to_sfixed_a(-0.07661917805671692)),(to_sfixed_a(0.00044158779201097786)),(to_sfixed_a(0.0002722414501477033)),(to_sfixed_a(-0.00015246414113789797)),(to_sfixed_a(0.0001584031415404752)),(to_sfixed_a(-0.00010059096530312672)),(to_sfixed_a(-0.00016356620471924543)),(to_sfixed_a(-8.76548801898025e-05)),(to_sfixed_a(-0.06813779473304749)),(to_sfixed_a(-0.05211099609732628)),(to_sfixed_a(-0.04258546233177185)),(to_sfixed_a(0.07436986267566681)),(to_sfixed_a(0.005391546059399843)),(to_sfixed_a(0.14162211120128632)),(to_sfixed_a(0.02872348204255104)),(to_sfixed_a(-0.2131376713514328)),(to_sfixed_a(-0.1204444169998169)),(to_sfixed_a(-0.24555493891239166)),(to_sfixed_a(0.073274165391922)),(to_sfixed_a(0.07069030404090881)),(to_sfixed_a(-0.1433010697364807)),(to_sfixed_a(0.088135726749897)),(to_sfixed_a(0.23091493546962738)),(to_sfixed_a(0.18385683000087738)),(to_sfixed_a(-0.04386857524514198)),(to_sfixed_a(0.09623110294342041)),(to_sfixed_a(-0.024380162358283997)),(to_sfixed_a(0.055349647998809814)),(to_sfixed_a(-0.03773941099643707)),(to_sfixed_a(0.0004241941496729851)),(to_sfixed_a(8.363732922589406e-05)),(to_sfixed_a(-4.032189099234529e-05)),(to_sfixed_a(0.0001202977800858207)),(to_sfixed_a(-9.162690548691899e-05)),(to_sfixed_a(-9.220178617397323e-05)),(to_sfixed_a(-0.0024425783194601536)),(to_sfixed_a(0.0850520208477974)),(to_sfixed_a(0.030605677515268326)),(to_sfixed_a(-0.22500371932983398)),(to_sfixed_a(0.01150232832878828)),(to_sfixed_a(-0.15288566052913666)),(to_sfixed_a(-0.009174119681119919)),(to_sfixed_a(0.1721038818359375)),(to_sfixed_a(-0.02103608474135399)),(to_sfixed_a(0.06253215670585632)),(to_sfixed_a(0.028230562806129456)),(to_sfixed_a(-0.0033998535946011543)),(to_sfixed_a(0.06151773780584335)),(to_sfixed_a(-0.20424127578735352)),(to_sfixed_a(0.0515841580927372)),(to_sfixed_a(-0.0021753376349806786)),(to_sfixed_a(0.04420031979680061)),(to_sfixed_a(0.09120268374681473)),(to_sfixed_a(-0.2439413219690323)),(to_sfixed_a(0.13617902994155884)),(to_sfixed_a(-0.05526156350970268)),(to_sfixed_a(0.022108646109700203)),(to_sfixed_a(-0.01326209306716919)),(to_sfixed_a(1.2769985914928839e-05)),(to_sfixed_a(-0.00028181663947179914)),(to_sfixed_a(0.0001283213496208191)),(to_sfixed_a(7.587347681692336e-06)),(to_sfixed_a(-0.0015923298196867108)),(to_sfixed_a(-0.0025866699870675802)),(to_sfixed_a(0.07272370904684067)),(to_sfixed_a(0.027653325349092484)),(to_sfixed_a(-0.12729397416114807)),(to_sfixed_a(-0.41935181617736816)),(to_sfixed_a(-0.3843044936656952)),(to_sfixed_a(-0.14439821243286133)),(to_sfixed_a(-0.011474202387034893)),(to_sfixed_a(0.038590144366025925)),(to_sfixed_a(0.09770379960536957)),(to_sfixed_a(-0.05205145850777626)),(to_sfixed_a(-0.16701288521289825)),(to_sfixed_a(0.02010349929332733)),(to_sfixed_a(-0.030232710763812065)),(to_sfixed_a(-0.04076157137751579)),(to_sfixed_a(-0.02689874731004238)),(to_sfixed_a(-0.08784065395593643)),(to_sfixed_a(-0.07083629071712494)),(to_sfixed_a(0.10243366658687592)),(to_sfixed_a(0.22905780375003815)),(to_sfixed_a(0.0021444465965032578)),(to_sfixed_a(3.9472030266551883e-07)),(to_sfixed_a(0.00010152862523682415)),(to_sfixed_a(-2.56830044236267e-05)),(to_sfixed_a(5.354125096346252e-05)),(to_sfixed_a(-3.52995175489923e-06)),(to_sfixed_a(-2.5637609724071808e-05)),(to_sfixed_a(3.484457192826085e-05)),(to_sfixed_a(0.03395986557006836)),(to_sfixed_a(0.005403503775596619)),(to_sfixed_a(-0.03712531179189682)),(to_sfixed_a(-0.1037578210234642)),(to_sfixed_a(0.03063492849469185)),(to_sfixed_a(-0.03361712768673897)),(to_sfixed_a(0.0749870017170906)),(to_sfixed_a(0.2550322711467743)),(to_sfixed_a(0.1299639642238617)),(to_sfixed_a(0.005376286339014769)),(to_sfixed_a(0.1756570190191269)),(to_sfixed_a(0.29952213168144226)),(to_sfixed_a(0.11648906767368317)),(to_sfixed_a(0.06473768502473831)),(to_sfixed_a(-0.044118888676166534)),(to_sfixed_a(-0.06628396362066269)),(to_sfixed_a(0.3705504238605499)),(to_sfixed_a(0.21854150295257568)),(to_sfixed_a(0.12000924348831177)),(to_sfixed_a(0.1419893205165863)),(to_sfixed_a(-0.03690635412931442)),(to_sfixed_a(-0.0395759716629982)),(to_sfixed_a(-0.00013307596964295954)),(to_sfixed_a(-0.0001370764512103051)),(to_sfixed_a(-0.0001924301468534395)),(to_sfixed_a(-0.000285892077954486)),(to_sfixed_a(-2.9540053219534457e-05)),(to_sfixed_a(2.3163174773799255e-05)),(to_sfixed_a(-0.029934624210000038)),(to_sfixed_a(0.00209266459569335)),(to_sfixed_a(-0.11999061703681946)),(to_sfixed_a(-0.07901546359062195)),(to_sfixed_a(-0.021337686106562614)),(to_sfixed_a(0.038393355906009674)),(to_sfixed_a(-0.06919688731431961)),(to_sfixed_a(-0.06279977411031723)),(to_sfixed_a(-0.0011659328592941165)),(to_sfixed_a(0.07265640795230865)),(to_sfixed_a(0.14375105500221252)),(to_sfixed_a(-0.132818341255188)),(to_sfixed_a(0.029103873297572136)),(to_sfixed_a(-0.05138666555285454)),(to_sfixed_a(-0.1502888947725296)),(to_sfixed_a(0.03445471078157425)),(to_sfixed_a(-0.05708318203687668)),(to_sfixed_a(0.16743719577789307)),(to_sfixed_a(-0.051066525280475616)),(to_sfixed_a(0.09726685285568237)),(to_sfixed_a(0.10976973176002502)),(to_sfixed_a(-1.88430003618123e-05)),(to_sfixed_a(0.00014667438517790288)),(to_sfixed_a(0.0002903361455537379)),(to_sfixed_a(0.0001419051841367036)),(to_sfixed_a(0.0004413595306687057)),(to_sfixed_a(-0.00014575125533156097)),(to_sfixed_a(-1.7631287846597843e-05)),(to_sfixed_a(-1.3733952982875053e-05)),(to_sfixed_a(-0.005875247996300459)),(to_sfixed_a(-0.023822562769055367)),(to_sfixed_a(-0.19084575772285461)),(to_sfixed_a(0.18679653108119965)),(to_sfixed_a(0.17899073660373688)),(to_sfixed_a(0.04037634655833244)),(to_sfixed_a(-0.07464815676212311)),(to_sfixed_a(0.12976409494876862)),(to_sfixed_a(-0.03370009362697601)),(to_sfixed_a(0.0025697879027575254)),(to_sfixed_a(-0.24855536222457886)),(to_sfixed_a(-0.2223893105983734)),(to_sfixed_a(-0.22955499589443207)),(to_sfixed_a(-0.32884618639945984)),(to_sfixed_a(0.21874946355819702)),(to_sfixed_a(-0.07471497356891632)),(to_sfixed_a(0.06940804421901703)),(to_sfixed_a(0.03960607573390007)),(to_sfixed_a(0.061112526804208755)),(to_sfixed_a(0.03800328075885773)),(to_sfixed_a(0.06748023629188538)),(to_sfixed_a(0.0002482305862940848)),(to_sfixed_a(-0.00010728371853474528)),(to_sfixed_a(6.172922894620569e-06)),(to_sfixed_a(-4.8306657845387235e-05)),(to_sfixed_a(-7.910142448963597e-05)),(to_sfixed_a(-1.6840140233398415e-05)),(to_sfixed_a(0.00019793721730820835)),(to_sfixed_a(0.015141179785132408)),(to_sfixed_a(-0.0002554735983721912)),(to_sfixed_a(0.13701343536376953)),(to_sfixed_a(0.11570291966199875)),(to_sfixed_a(0.09330694377422333)),(to_sfixed_a(-0.0577617883682251)),(to_sfixed_a(0.18255022168159485)),(to_sfixed_a(-0.04035503417253494)),(to_sfixed_a(-0.16560165584087372)),(to_sfixed_a(-0.10290580987930298)),(to_sfixed_a(-0.01995495893061161)),(to_sfixed_a(-0.4013480544090271)),(to_sfixed_a(-0.06507942825555801)),(to_sfixed_a(0.13085323572158813)),(to_sfixed_a(0.21516795456409454)),(to_sfixed_a(0.2520298659801483)),(to_sfixed_a(-0.06194833293557167)),(to_sfixed_a(-0.045871540904045105)),(to_sfixed_a(0.07965445518493652)),(to_sfixed_a(-0.0010005440562963486)),(to_sfixed_a(-0.07223626226186752)),(to_sfixed_a(-2.771182516880799e-05)),(to_sfixed_a(-5.401948874350637e-05)),(to_sfixed_a(-0.0003607632825151086)),(to_sfixed_a(3.766479130717926e-05)),(to_sfixed_a(0.00023549352772533894)),(to_sfixed_a(-7.846082735341042e-05)),(to_sfixed_a(-0.00022546514810528606)),(to_sfixed_a(-0.00014077707601245493)),(to_sfixed_a(-0.05702289938926697)),(to_sfixed_a(0.03099755384027958)),(to_sfixed_a(0.09852530807256699)),(to_sfixed_a(0.008181600831449032)),(to_sfixed_a(-0.07377147674560547)),(to_sfixed_a(0.03967529162764549)),(to_sfixed_a(-0.013603756204247475)),(to_sfixed_a(-0.21030190587043762)),(to_sfixed_a(-0.11348940432071686)),(to_sfixed_a(-0.0724344253540039)),(to_sfixed_a(-0.08739209175109863)),(to_sfixed_a(0.056030455976724625)),(to_sfixed_a(0.0890517309308052)),(to_sfixed_a(0.2616061866283417)),(to_sfixed_a(0.13484947383403778)),(to_sfixed_a(0.022504445165395737)),(to_sfixed_a(-0.006621550768613815)),(to_sfixed_a(-0.08658242225646973)),(to_sfixed_a(-0.007656922098249197)),(to_sfixed_a(2.296620368724689e-05)),(to_sfixed_a(0.00020979912369512022)),(to_sfixed_a(-0.00014442384417634457)),(to_sfixed_a(9.191697608912364e-05)),(to_sfixed_a(-0.0001385301147820428)),(to_sfixed_a(0.00010382881737314165)),(to_sfixed_a(-7.67658420954831e-05)),(to_sfixed_a(-0.00021510370424948633)),(to_sfixed_a(-0.0001239480043295771)),(to_sfixed_a(-0.007041467819362879)),(to_sfixed_a(-0.021929852664470673)),(to_sfixed_a(-0.2842399775981903)),(to_sfixed_a(-0.0030202423222362995)),(to_sfixed_a(0.01840362325310707)),(to_sfixed_a(-0.09985557198524475)),(to_sfixed_a(-0.11116241663694382)),(to_sfixed_a(0.00044446534593589604)),(to_sfixed_a(-0.059480227530002594)),(to_sfixed_a(0.020558224990963936)),(to_sfixed_a(-0.017285361886024475)),(to_sfixed_a(-0.05662418156862259)),(to_sfixed_a(-0.0630202516913414)),(to_sfixed_a(0.02367706224322319)),(to_sfixed_a(0.07844600826501846)),(to_sfixed_a(0.01871039718389511)),(to_sfixed_a(0.09431704878807068)),(to_sfixed_a(0.0010280886199325323)),(to_sfixed_a(0.06957370042800903)),(to_sfixed_a(0.00029113859636709094)),(to_sfixed_a(0.00018433183140587062)),(to_sfixed_a(-7.295070645341184e-07)),(to_sfixed_a(-0.00016658428648952395)),(to_sfixed_a(-7.380187889793888e-05)),(to_sfixed_a(-0.00018069565703626722)),(to_sfixed_a(0.0002279109467053786)),(to_sfixed_a(4.116927448194474e-05)),(to_sfixed_a(0.023161068558692932)),(to_sfixed_a(0.03740272670984268)),(to_sfixed_a(0.0955473780632019)),(to_sfixed_a(0.11086209118366241)),(to_sfixed_a(0.06844388693571091)),(to_sfixed_a(0.13436701893806458)),(to_sfixed_a(-0.02626716159284115)),(to_sfixed_a(-0.1543971747159958)),(to_sfixed_a(0.03250999003648758)),(to_sfixed_a(-0.010986017994582653)),(to_sfixed_a(0.0887916311621666)),(to_sfixed_a(0.12392356991767883)),(to_sfixed_a(0.1181836798787117)),(to_sfixed_a(0.01846439577639103)),(to_sfixed_a(0.09093455970287323)),(to_sfixed_a(0.15565325319766998)),(to_sfixed_a(-0.000467782374471426)),(to_sfixed_a(0.14450187981128693)),(to_sfixed_a(0.05333111062645912)),(to_sfixed_a(0.018261078745126724)),(to_sfixed_a(-1.6184158084797673e-05)),(to_sfixed_a(-6.092572948546149e-05)),(to_sfixed_a(7.929916318971664e-05)),(to_sfixed_a(0.0001642329734750092)),(to_sfixed_a(0.00036016356898471713)),(to_sfixed_a(0.00013127631973475218)),(to_sfixed_a(-0.0001527466083643958)),(to_sfixed_a(-0.00022519720369018614)),(to_sfixed_a(-7.718388951616362e-05)),(to_sfixed_a(-0.031215468421578407)),(to_sfixed_a(0.057934924960136414)),(to_sfixed_a(0.02901594713330269)),(to_sfixed_a(0.049771059304475784)),(to_sfixed_a(-0.03156093880534172)),(to_sfixed_a(0.04861724004149437)),(to_sfixed_a(0.16415870189666748)),(to_sfixed_a(-0.066916324198246)),(to_sfixed_a(0.019974414259195328)),(to_sfixed_a(0.11296647787094116)),(to_sfixed_a(0.07471900433301926)),(to_sfixed_a(0.31688371300697327)),(to_sfixed_a(-0.05338042229413986)),(to_sfixed_a(0.0055212462320923805)),(to_sfixed_a(0.33100223541259766)),(to_sfixed_a(0.13531000912189484)),(to_sfixed_a(-0.0006184601224958897)),(to_sfixed_a(-0.0010254087392240763)),(to_sfixed_a(-0.0009008576162159443)),(to_sfixed_a(-0.0001269956264877692)),(to_sfixed_a(-6.135176226962358e-05)),(to_sfixed_a(-0.00028276685043238103)),(to_sfixed_a(-0.00022773556702304631)),(to_sfixed_a(0.00014154832751955837)),(to_sfixed_a(-0.00034426175989210606)),(to_sfixed_a(-8.962858555605635e-05)),(to_sfixed_a(-8.810379949864e-05)),(to_sfixed_a(-0.00019720352429430932)),(to_sfixed_a(-0.0006706432905048132)),(to_sfixed_a(-0.0007597960066050291)),(to_sfixed_a(0.00019881386833731085)),(to_sfixed_a(-6.240334187168628e-05)),(to_sfixed_a(5.7901856052922085e-05)),(to_sfixed_a(0.19090315699577332)),(to_sfixed_a(-0.009502032771706581)),(to_sfixed_a(-0.0016892249695956707)),(to_sfixed_a(0.14847080409526825)),(to_sfixed_a(0.02155783213675022)),(to_sfixed_a(0.013479688204824924)),(to_sfixed_a(0.08599981665611267)),(to_sfixed_a(0.15477395057678223)),(to_sfixed_a(0.20406727492809296)),(to_sfixed_a(0.006858388893306255)),(to_sfixed_a(0.004693267866969109)),(to_sfixed_a(0.00011198454012628645)),(to_sfixed_a(-4.4427528337109834e-05)),(to_sfixed_a(-5.1870312745450065e-05)),(to_sfixed_a(-9.946286445483565e-05)),(to_sfixed_a(6.172609573695809e-05)),(to_sfixed_a(-5.2381717978278175e-05)),(to_sfixed_a(0.0002720073389355093)),(to_sfixed_a(-0.00024472735822200775)),(to_sfixed_a(9.063223842531443e-05)),(to_sfixed_a(2.6806579626281746e-05)),(to_sfixed_a(-6.107433728175238e-05)),(to_sfixed_a(-0.00023719963792245835)),(to_sfixed_a(0.00020877935457974672)),(to_sfixed_a(7.928962077130564e-06)),(to_sfixed_a(-1.8664582967176102e-05)),(to_sfixed_a(-0.00023001596855465323)),(to_sfixed_a(7.52976193325594e-05)),(to_sfixed_a(-0.00018024069140665233)),(to_sfixed_a(-0.0003467547066975385)),(to_sfixed_a(-1.0335126717109233e-05)),(to_sfixed_a(6.076959834899753e-05)),(to_sfixed_a(0.00010288512567058206)),(to_sfixed_a(8.669702219776809e-05)),(to_sfixed_a(9.543958003632724e-05)),(to_sfixed_a(-0.00010379749437561259)),(to_sfixed_a(4.447656465345062e-06)),(to_sfixed_a(0.00012564955977723002)),(to_sfixed_a(0.00010884186485782266)),(to_sfixed_a(0.0001319009461440146)),(to_sfixed_a(0.00011900687968591228)),(to_sfixed_a(0.00014157130499370396)),(to_sfixed_a(-3.863774691126309e-05)),(to_sfixed_a(-3.248716893722303e-05)),(to_sfixed_a(-1.4671356439066585e-05)),(to_sfixed_a(0.0001512609451310709)));

    constant weight_n0_31 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(0.0001789199304766953)),(to_sfixed_a(-4.864115544478409e-05)),(to_sfixed_a(0.00010102221858687699)),(to_sfixed_a(-1.4368129086506087e-05)),(to_sfixed_a(0.00015171848644968122)),(to_sfixed_a(-1.4215748706192244e-05)),(to_sfixed_a(2.6239955332130194e-05)),(to_sfixed_a(-0.0001703430461930111)),(to_sfixed_a(0.00014088806346990168)),(to_sfixed_a(-0.00010098538768943399)),(to_sfixed_a(2.6254949261783622e-05)),(to_sfixed_a(-5.947496902081184e-05)),(to_sfixed_a(-6.577106250915676e-05)),(to_sfixed_a(7.861085759941489e-05)),(to_sfixed_a(-8.37774932733737e-05)),(to_sfixed_a(4.733470632345416e-06)),(to_sfixed_a(-7.42764605092816e-05)),(to_sfixed_a(0.0001548565342091024)),(to_sfixed_a(-3.996202940470539e-05)),(to_sfixed_a(0.00011428291327320039)),(to_sfixed_a(0.00012494025577325374)),(to_sfixed_a(0.00032776963780634105)),(to_sfixed_a(-2.3505088392994367e-05)),(to_sfixed_a(-3.5171986382920295e-05)),(to_sfixed_a(-0.0002085081796394661)),(to_sfixed_a(0.0001467079418944195)),(to_sfixed_a(-7.970822480274364e-05)),(to_sfixed_a(-0.00013305139145813882)),(to_sfixed_a(0.0003873302775900811)),(to_sfixed_a(-0.00012172860442660749)),(to_sfixed_a(2.789003701764159e-05)),(to_sfixed_a(-2.2008309315424412e-05)),(to_sfixed_a(-0.00027507171034812927)),(to_sfixed_a(7.253674993989989e-05)),(to_sfixed_a(-0.00018935654952656478)),(to_sfixed_a(5.164929825696163e-05)),(to_sfixed_a(-9.506460628472269e-05)),(to_sfixed_a(-6.025868060532957e-05)),(to_sfixed_a(-0.00018476517288945615)),(to_sfixed_a(2.2810518203186803e-05)),(to_sfixed_a(0.0002643547486513853)),(to_sfixed_a(-0.0001847021485446021)),(to_sfixed_a(-0.0001938142959261313)),(to_sfixed_a(0.00024753392790444195)),(to_sfixed_a(-0.00034835634869523346)),(to_sfixed_a(-0.00018386193551123142)),(to_sfixed_a(-8.754297596169636e-05)),(to_sfixed_a(-0.00011012232425855473)),(to_sfixed_a(0.0001666979951551184)),(to_sfixed_a(0.00021341476531233639)),(to_sfixed_a(5.2839597628917545e-05)),(to_sfixed_a(-0.00010074403689941391)),(to_sfixed_a(0.00019476847955957055)),(to_sfixed_a(-8.187667117454112e-05)),(to_sfixed_a(-0.0001598170056240633)),(to_sfixed_a(-5.387240162235685e-05)),(to_sfixed_a(-0.00011994690430583432)),(to_sfixed_a(5.705763032892719e-05)),(to_sfixed_a(-0.0001509688445366919)),(to_sfixed_a(-0.00018001471471507102)),(to_sfixed_a(3.0334991606650874e-05)),(to_sfixed_a(-0.00013625442807096988)),(to_sfixed_a(0.0003350238548591733)),(to_sfixed_a(-0.00013194289931561798)),(to_sfixed_a(-1.4456100871029776e-05)),(to_sfixed_a(0.00022180045198183507)),(to_sfixed_a(1.1479239219625015e-05)),(to_sfixed_a(-1.9967503249063157e-05)),(to_sfixed_a(-0.0001944604009622708)),(to_sfixed_a(-0.008844810537993908)),(to_sfixed_a(-0.0002082803111989051)),(to_sfixed_a(-8.562244329368696e-05)),(to_sfixed_a(-4.6525638026650995e-06)),(to_sfixed_a(-8.838360372465104e-05)),(to_sfixed_a(8.775390597293153e-05)),(to_sfixed_a(-1.038067875924753e-05)),(to_sfixed_a(0.0001911595609271899)),(to_sfixed_a(4.119724690099247e-05)),(to_sfixed_a(-0.0001652726496104151)),(to_sfixed_a(5.685393625753932e-05)),(to_sfixed_a(-1.6332866152879433e-06)),(to_sfixed_a(9.169027907773852e-05)),(to_sfixed_a(-6.877214036649093e-05)),(to_sfixed_a(-0.0001487648842157796)),(to_sfixed_a(-0.00016938384214881808)),(to_sfixed_a(4.3349438783479854e-05)),(to_sfixed_a(-4.163246921962127e-05)),(to_sfixed_a(-4.1265488107455894e-05)),(to_sfixed_a(-0.00022369813814293593)),(to_sfixed_a(6.36404802207835e-05)),(to_sfixed_a(2.5421347800147487e-06)),(to_sfixed_a(-0.0002594068937469274)),(to_sfixed_a(0.03890242427587509)),(to_sfixed_a(-5.637784852297045e-05)),(to_sfixed_a(0.04404234513640404)),(to_sfixed_a(0.04810762032866478)),(to_sfixed_a(0.08382581919431686)),(to_sfixed_a(0.03502571955323219)),(to_sfixed_a(0.06907660514116287)),(to_sfixed_a(0.0048457724042236805)),(to_sfixed_a(0.02389080449938774)),(to_sfixed_a(-0.01917085237801075)),(to_sfixed_a(0.0005992625374346972)),(to_sfixed_a(-0.034933026880025864)),(to_sfixed_a(-0.009196680039167404)),(to_sfixed_a(-0.018555225804448128)),(to_sfixed_a(0.00012341247929725796)),(to_sfixed_a(3.4630591017048573e-06)),(to_sfixed_a(-6.558919267263263e-05)),(to_sfixed_a(-8.542474824935198e-05)),(to_sfixed_a(5.7911511248676106e-05)),(to_sfixed_a(3.0118912036414258e-05)),(to_sfixed_a(-0.00031675814534537494)),(to_sfixed_a(-8.521169547748286e-06)),(to_sfixed_a(0.00013017021410632879)),(to_sfixed_a(8.091517520369962e-05)),(to_sfixed_a(-0.0001510914007667452)),(to_sfixed_a(0.00013502778892870992)),(to_sfixed_a(0.00043545971857383847)),(to_sfixed_a(-0.02207726612687111)),(to_sfixed_a(0.013253478333353996)),(to_sfixed_a(0.058231402188539505)),(to_sfixed_a(0.1364811509847641)),(to_sfixed_a(0.005466788541525602)),(to_sfixed_a(0.0051977732218801975)),(to_sfixed_a(0.07033272087574005)),(to_sfixed_a(0.1193663626909256)),(to_sfixed_a(0.0049211434088647366)),(to_sfixed_a(-0.0035395915620028973)),(to_sfixed_a(0.015985306352376938)),(to_sfixed_a(-0.02540731057524681)),(to_sfixed_a(-0.0774737223982811)),(to_sfixed_a(-0.0007211426855064929)),(to_sfixed_a(0.03252384439110756)),(to_sfixed_a(-0.007899337448179722)),(to_sfixed_a(3.992153779108776e-06)),(to_sfixed_a(-0.0004773239779751748)),(to_sfixed_a(-7.554019248345867e-05)),(to_sfixed_a(-0.00023989632609300315)),(to_sfixed_a(0.00013792593381367624)),(to_sfixed_a(6.114385178079829e-05)),(to_sfixed_a(0.00010887996177189052)),(to_sfixed_a(-1.916440851346124e-05)),(to_sfixed_a(-0.0002270678960485384)),(to_sfixed_a(0.000861856562551111)),(to_sfixed_a(-0.04579664021730423)),(to_sfixed_a(-0.012115118093788624)),(to_sfixed_a(-0.10166051238775253)),(to_sfixed_a(0.13482515513896942)),(to_sfixed_a(0.06804143637418747)),(to_sfixed_a(0.05711133033037186)),(to_sfixed_a(0.04076460376381874)),(to_sfixed_a(0.057584285736083984)),(to_sfixed_a(0.04097244516015053)),(to_sfixed_a(0.2053077220916748)),(to_sfixed_a(0.18358521163463593)),(to_sfixed_a(0.03282671794295311)),(to_sfixed_a(-0.14982709288597107)),(to_sfixed_a(-0.06319776922464371)),(to_sfixed_a(-0.362210214138031)),(to_sfixed_a(-0.08083507418632507)),(to_sfixed_a(0.061606742441654205)),(to_sfixed_a(-0.002831418067216873)),(to_sfixed_a(-0.06190493330359459)),(to_sfixed_a(0.0018038098933175206)),(to_sfixed_a(0.00016562097880523652)),(to_sfixed_a(-8.383942622458562e-05)),(to_sfixed_a(-3.14630196953658e-05)),(to_sfixed_a(0.0001288160856347531)),(to_sfixed_a(-6.288349686656147e-05)),(to_sfixed_a(-1.9792347302427515e-05)),(to_sfixed_a(8.223256736528128e-05)),(to_sfixed_a(-4.944071770296432e-05)),(to_sfixed_a(-0.04328230023384094)),(to_sfixed_a(-0.07699614018201828)),(to_sfixed_a(-0.00716425059363246)),(to_sfixed_a(-0.0030027537140995264)),(to_sfixed_a(0.20138226449489594)),(to_sfixed_a(0.20628252625465393)),(to_sfixed_a(0.17187665402889252)),(to_sfixed_a(0.20423242449760437)),(to_sfixed_a(0.19103772938251495)),(to_sfixed_a(0.06824459880590439)),(to_sfixed_a(0.036851461976766586)),(to_sfixed_a(0.06264133751392365)),(to_sfixed_a(-0.1351865977048874)),(to_sfixed_a(-0.033052440732717514)),(to_sfixed_a(-0.2586902976036072)),(to_sfixed_a(0.06127459183335304)),(to_sfixed_a(0.0697999820113182)),(to_sfixed_a(0.1678377091884613)),(to_sfixed_a(0.12006557732820511)),(to_sfixed_a(0.010364130139350891)),(to_sfixed_a(0.010681950487196445)),(to_sfixed_a(0.007339585572481155)),(to_sfixed_a(9.179888002108783e-05)),(to_sfixed_a(0.00018965904018841684)),(to_sfixed_a(-5.7228120567742735e-05)),(to_sfixed_a(-8.55353573570028e-05)),(to_sfixed_a(1.1752080354199279e-05)),(to_sfixed_a(-0.0003360616392455995)),(to_sfixed_a(-0.0552351213991642)),(to_sfixed_a(0.033741142600774765)),(to_sfixed_a(-0.13820800185203552)),(to_sfixed_a(0.13260121643543243)),(to_sfixed_a(0.03514852002263069)),(to_sfixed_a(0.45647236704826355)),(to_sfixed_a(0.0017892435425892472)),(to_sfixed_a(-0.08393023163080215)),(to_sfixed_a(-0.019790804013609886)),(to_sfixed_a(0.033310867846012115)),(to_sfixed_a(0.039400603622198105)),(to_sfixed_a(0.20205627381801605)),(to_sfixed_a(-0.0935598611831665)),(to_sfixed_a(0.17964215576648712)),(to_sfixed_a(-0.11186651140451431)),(to_sfixed_a(-0.2509855031967163)),(to_sfixed_a(-0.19838674366474152)),(to_sfixed_a(0.03077571466565132)),(to_sfixed_a(-0.10571415722370148)),(to_sfixed_a(0.03847919777035713)),(to_sfixed_a(0.0016728321788832545)),(to_sfixed_a(7.19395829946734e-05)),(to_sfixed_a(-0.00022445312060881406)),(to_sfixed_a(0.00011343023652443662)),(to_sfixed_a(-0.00011389212886570022)),(to_sfixed_a(-7.488662231480703e-05)),(to_sfixed_a(0.00014702185580972582)),(to_sfixed_a(0.014152834191918373)),(to_sfixed_a(0.031478311866521835)),(to_sfixed_a(-0.1084209755063057)),(to_sfixed_a(0.016328129917383194)),(to_sfixed_a(-0.05950123071670532)),(to_sfixed_a(0.029292987659573555)),(to_sfixed_a(-0.2278757244348526)),(to_sfixed_a(0.061081767082214355)),(to_sfixed_a(-0.0769888311624527)),(to_sfixed_a(-1.3223899259173777e-05)),(to_sfixed_a(-0.09182246029376984)),(to_sfixed_a(0.1389807164669037)),(to_sfixed_a(0.16817811131477356)),(to_sfixed_a(0.09856107831001282)),(to_sfixed_a(0.10791287571191788)),(to_sfixed_a(0.02791057713329792)),(to_sfixed_a(-0.04171190410852432)),(to_sfixed_a(0.03446929529309273)),(to_sfixed_a(-0.07382512837648392)),(to_sfixed_a(-0.08522894233465195)),(to_sfixed_a(0.1471608430147171)),(to_sfixed_a(0.025873957201838493)),(to_sfixed_a(-0.00013305796892382205)),(to_sfixed_a(-7.270503556355834e-05)),(to_sfixed_a(0.00032932599424384534)),(to_sfixed_a(9.575548028806224e-05)),(to_sfixed_a(5.014971975469962e-05)),(to_sfixed_a(-9.611214773030952e-05)),(to_sfixed_a(-0.0008570587961003184)),(to_sfixed_a(0.025090565904974937)),(to_sfixed_a(0.09066049009561539)),(to_sfixed_a(0.18926270306110382)),(to_sfixed_a(-0.011998314410448074)),(to_sfixed_a(0.05641862377524376)),(to_sfixed_a(0.31392478942871094)),(to_sfixed_a(-0.18525001406669617)),(to_sfixed_a(-0.015824662521481514)),(to_sfixed_a(-0.3295517563819885)),(to_sfixed_a(0.03388894721865654)),(to_sfixed_a(-0.19817721843719482)),(to_sfixed_a(-0.0954718366265297)),(to_sfixed_a(0.11844197660684586)),(to_sfixed_a(0.2832833528518677)),(to_sfixed_a(-0.009953691624104977)),(to_sfixed_a(-0.09416665881872177)),(to_sfixed_a(0.06048703193664551)),(to_sfixed_a(-0.06173420324921608)),(to_sfixed_a(0.0730782076716423)),(to_sfixed_a(0.1561950147151947)),(to_sfixed_a(-2.9786667710141046e-06)),(to_sfixed_a(4.046177491545677e-05)),(to_sfixed_a(-0.00011494549107737839)),(to_sfixed_a(0.00016637169755995274)),(to_sfixed_a(0.00010771750385174528)),(to_sfixed_a(-5.858648000867106e-05)),(to_sfixed_a(0.00019148981664329767)),(to_sfixed_a(-0.002380810445174575)),(to_sfixed_a(-0.03893166780471802)),(to_sfixed_a(0.1941869705915451)),(to_sfixed_a(0.03424539417028427)),(to_sfixed_a(0.08394502103328705)),(to_sfixed_a(-0.02863362431526184)),(to_sfixed_a(0.04739703610539436)),(to_sfixed_a(0.05861463397741318)),(to_sfixed_a(-0.08701782673597336)),(to_sfixed_a(-0.26518282294273376)),(to_sfixed_a(-0.03009316697716713)),(to_sfixed_a(-0.07483396679162979)),(to_sfixed_a(-0.02768641710281372)),(to_sfixed_a(0.05065630376338959)),(to_sfixed_a(0.1535540223121643)),(to_sfixed_a(0.06495677679777145)),(to_sfixed_a(0.05780955031514168)),(to_sfixed_a(-0.031905706971883774)),(to_sfixed_a(0.03726860508322716)),(to_sfixed_a(-0.2777196168899536)),(to_sfixed_a(0.008760022930800915)),(to_sfixed_a(0.06886519491672516)),(to_sfixed_a(0.0001330274244537577)),(to_sfixed_a(0.00016608115402050316)),(to_sfixed_a(-0.00011613788228714839)),(to_sfixed_a(4.767937571159564e-05)),(to_sfixed_a(-0.0001452042633900419)),(to_sfixed_a(0.0610005185008049)),(to_sfixed_a(0.030882300809025764)),(to_sfixed_a(0.2084943652153015)),(to_sfixed_a(0.02518501505255699)),(to_sfixed_a(0.1635316014289856)),(to_sfixed_a(0.14232957363128662)),(to_sfixed_a(0.07535640150308609)),(to_sfixed_a(0.17278815805912018)),(to_sfixed_a(0.05505989491939545)),(to_sfixed_a(-0.012876706197857857)),(to_sfixed_a(-0.16605132818222046)),(to_sfixed_a(0.23371478915214539)),(to_sfixed_a(0.0057477569207549095)),(to_sfixed_a(-0.017852790653705597)),(to_sfixed_a(0.022649377584457397)),(to_sfixed_a(0.07779985666275024)),(to_sfixed_a(0.01914866827428341)),(to_sfixed_a(0.03768140822649002)),(to_sfixed_a(0.09616079926490784)),(to_sfixed_a(0.15776148438453674)),(to_sfixed_a(-0.1507982462644577)),(to_sfixed_a(-0.12576882541179657)),(to_sfixed_a(-0.0001285423495573923)),(to_sfixed_a(1.568447805766482e-05)),(to_sfixed_a(0.000172246087458916)),(to_sfixed_a(-0.00014545161684509367)),(to_sfixed_a(0.0003998780739493668)),(to_sfixed_a(-5.1960389100713655e-05)),(to_sfixed_a(0.00011462176917120814)),(to_sfixed_a(0.14424745738506317)),(to_sfixed_a(0.10568548738956451)),(to_sfixed_a(0.06330152601003647)),(to_sfixed_a(0.18962204456329346)),(to_sfixed_a(0.20870418846607208)),(to_sfixed_a(0.15134014189243317)),(to_sfixed_a(0.04850504547357559)),(to_sfixed_a(-0.08609425276517868)),(to_sfixed_a(0.27910786867141724)),(to_sfixed_a(0.06553985178470612)),(to_sfixed_a(-0.3060428500175476)),(to_sfixed_a(-0.1056511253118515)),(to_sfixed_a(0.5689222812652588)),(to_sfixed_a(0.1950451135635376)),(to_sfixed_a(0.2063814103603363)),(to_sfixed_a(0.14917778968811035)),(to_sfixed_a(-0.29385292530059814)),(to_sfixed_a(-0.010677475482225418)),(to_sfixed_a(-0.16894449293613434)),(to_sfixed_a(-0.2620165944099426)),(to_sfixed_a(0.07179324328899384)),(to_sfixed_a(-5.04462695971597e-05)),(to_sfixed_a(-2.5788878701860085e-05)),(to_sfixed_a(4.532469029072672e-05)),(to_sfixed_a(7.368214573943987e-05)),(to_sfixed_a(-0.00012436967517714947)),(to_sfixed_a(-6.201201176736504e-05)),(to_sfixed_a(5.497694291989319e-05)),(to_sfixed_a(0.08632243424654007)),(to_sfixed_a(-0.08869689702987671)),(to_sfixed_a(-0.3401416838169098)),(to_sfixed_a(-0.20423460006713867)),(to_sfixed_a(-0.17061302065849304)),(to_sfixed_a(0.18841348588466644)),(to_sfixed_a(0.3141796886920929)),(to_sfixed_a(-0.0487915575504303)),(to_sfixed_a(0.16709637641906738)),(to_sfixed_a(0.0794471725821495)),(to_sfixed_a(-0.01940491981804371)),(to_sfixed_a(-0.1564416140317917)),(to_sfixed_a(-0.0051275016739964485)),(to_sfixed_a(-0.2020488828420639)),(to_sfixed_a(-0.020103519782423973)),(to_sfixed_a(0.06645502895116806)),(to_sfixed_a(0.060797542333602905)),(to_sfixed_a(-0.028232503682374954)),(to_sfixed_a(0.1796504110097885)),(to_sfixed_a(0.030545754358172417)),(to_sfixed_a(0.048188626766204834)),(to_sfixed_a(-0.002235487336292863)),(to_sfixed_a(-0.0012480049626901746)),(to_sfixed_a(1.0217093404207844e-05)),(to_sfixed_a(0.0004153370391577482)),(to_sfixed_a(-0.0003074830456171185)),(to_sfixed_a(0.00018920146976597607)),(to_sfixed_a(0.00011694066051859409)),(to_sfixed_a(-0.0013374659465625882)),(to_sfixed_a(0.09859468042850494)),(to_sfixed_a(0.02392793446779251)),(to_sfixed_a(-0.1944165676832199)),(to_sfixed_a(0.00013714376837015152)),(to_sfixed_a(-0.09514984488487244)),(to_sfixed_a(0.002940661273896694)),(to_sfixed_a(0.013220146298408508)),(to_sfixed_a(0.12972740828990936)),(to_sfixed_a(0.1288406103849411)),(to_sfixed_a(-0.11596477031707764)),(to_sfixed_a(0.019729794934391975)),(to_sfixed_a(0.17142614722251892)),(to_sfixed_a(-0.053109075874090195)),(to_sfixed_a(0.09260623157024384)),(to_sfixed_a(-0.22114627063274384)),(to_sfixed_a(0.023535188287496567)),(to_sfixed_a(0.14190684258937836)),(to_sfixed_a(0.013745012693107128)),(to_sfixed_a(-0.10059540718793869)),(to_sfixed_a(-0.08942531794309616)),(to_sfixed_a(0.00028456078143790364)),(to_sfixed_a(6.759937241440639e-05)),(to_sfixed_a(-6.464063335442916e-05)),(to_sfixed_a(0.00016477554163429886)),(to_sfixed_a(-0.00017017238133121282)),(to_sfixed_a(0.00026507300208322704)),(to_sfixed_a(0.00014015339547768235)),(to_sfixed_a(-0.05064806342124939)),(to_sfixed_a(0.09122154861688614)),(to_sfixed_a(-0.11746852844953537)),(to_sfixed_a(-0.12208898365497589)),(to_sfixed_a(-0.15522652864456177)),(to_sfixed_a(-0.18202465772628784)),(to_sfixed_a(-0.3449864387512207)),(to_sfixed_a(0.1382833868265152)),(to_sfixed_a(-0.36691462993621826)),(to_sfixed_a(-0.3468811511993408)),(to_sfixed_a(-0.1654495745897293)),(to_sfixed_a(-0.15323375165462494)),(to_sfixed_a(0.04014718532562256)),(to_sfixed_a(-0.0397137850522995)),(to_sfixed_a(0.05853910371661186)),(to_sfixed_a(0.188277930021286)),(to_sfixed_a(-0.24003472924232483)),(to_sfixed_a(-0.19336995482444763)),(to_sfixed_a(-0.14486567676067352)),(to_sfixed_a(-0.12034922093153)),(to_sfixed_a(-0.052962541580200195)),(to_sfixed_a(2.164673787774518e-06)),(to_sfixed_a(2.1948715129838092e-06)),(to_sfixed_a(0.00010910101264016703)),(to_sfixed_a(-0.00011372726294212043)),(to_sfixed_a(9.640224743634462e-05)),(to_sfixed_a(-0.00015839954721741378)),(to_sfixed_a(0.0009171133278869092)),(to_sfixed_a(-0.09575700759887695)),(to_sfixed_a(-0.19713042676448822)),(to_sfixed_a(-0.10808927565813065)),(to_sfixed_a(-0.04223612695932388)),(to_sfixed_a(-0.005430104210972786)),(to_sfixed_a(0.027408935129642487)),(to_sfixed_a(0.15949681401252747)),(to_sfixed_a(0.041519708931446075)),(to_sfixed_a(0.14356593787670135)),(to_sfixed_a(-0.37907537817955017)),(to_sfixed_a(-0.03503909707069397)),(to_sfixed_a(0.03883685544133186)),(to_sfixed_a(0.06427082419395447)),(to_sfixed_a(-0.07941178232431412)),(to_sfixed_a(-0.017362812533974648)),(to_sfixed_a(0.04368222504854202)),(to_sfixed_a(0.19145572185516357)),(to_sfixed_a(-0.25559067726135254)),(to_sfixed_a(-0.022691717371344566)),(to_sfixed_a(-0.022839633747935295)),(to_sfixed_a(0.04867358133196831)),(to_sfixed_a(-0.01504239346832037)),(to_sfixed_a(3.46801862178836e-05)),(to_sfixed_a(-0.0004105223051737994)),(to_sfixed_a(0.0001092359161702916)),(to_sfixed_a(0.0001397549785906449)),(to_sfixed_a(0.0011253129923716187)),(to_sfixed_a(0.001358525361865759)),(to_sfixed_a(-0.13465090095996857)),(to_sfixed_a(-0.08551681786775589)),(to_sfixed_a(0.13864834606647491)),(to_sfixed_a(0.30637606978416443)),(to_sfixed_a(0.12788672745227814)),(to_sfixed_a(0.3191869854927063)),(to_sfixed_a(0.1852385699748993)),(to_sfixed_a(0.057019732892513275)),(to_sfixed_a(0.10270003974437714)),(to_sfixed_a(-0.0921376496553421)),(to_sfixed_a(0.043940480798482895)),(to_sfixed_a(-0.026960909366607666)),(to_sfixed_a(0.059046097099781036)),(to_sfixed_a(0.14799053966999054)),(to_sfixed_a(-0.042578618973493576)),(to_sfixed_a(-0.18956850469112396)),(to_sfixed_a(0.1019841805100441)),(to_sfixed_a(-0.11259292811155319)),(to_sfixed_a(-0.1513511836528778)),(to_sfixed_a(0.014030327089130878)),(to_sfixed_a(-0.00011923745478270575)),(to_sfixed_a(8.924784197006375e-05)),(to_sfixed_a(0.00016229355242103338)),(to_sfixed_a(-0.00023222492018248886)),(to_sfixed_a(5.162063462194055e-05)),(to_sfixed_a(-2.9698710932279937e-05)),(to_sfixed_a(0.00012681186490226537)),(to_sfixed_a(-0.026900362223386765)),(to_sfixed_a(-0.08006476610898972)),(to_sfixed_a(0.12584559619426727)),(to_sfixed_a(0.06922028958797455)),(to_sfixed_a(-0.253696084022522)),(to_sfixed_a(0.19553004205226898)),(to_sfixed_a(0.16207759082317352)),(to_sfixed_a(0.03036903403699398)),(to_sfixed_a(-0.24555151164531708)),(to_sfixed_a(0.12789495289325714)),(to_sfixed_a(-0.03208323195576668)),(to_sfixed_a(-0.04770027473568916)),(to_sfixed_a(0.04431269317865372)),(to_sfixed_a(0.02297489158809185)),(to_sfixed_a(-0.06244485452771187)),(to_sfixed_a(-0.09278196096420288)),(to_sfixed_a(-0.1749681979417801)),(to_sfixed_a(-0.06223299354314804)),(to_sfixed_a(-0.012674812227487564)),(to_sfixed_a(-0.03994690626859665)),(to_sfixed_a(0.057235438376665115)),(to_sfixed_a(-0.025481106713414192)),(to_sfixed_a(-9.802527347346768e-05)),(to_sfixed_a(-0.0002053165517281741)),(to_sfixed_a(-0.0001821824989747256)),(to_sfixed_a(-1.5625237210770138e-05)),(to_sfixed_a(-7.471370918210596e-05)),(to_sfixed_a(-4.3507639929885045e-05)),(to_sfixed_a(0.01793404296040535)),(to_sfixed_a(0.0027184486389160156)),(to_sfixed_a(0.03901493921875954)),(to_sfixed_a(0.03408067673444748)),(to_sfixed_a(0.040301576256752014)),(to_sfixed_a(-0.096303790807724)),(to_sfixed_a(0.02583850361406803)),(to_sfixed_a(-0.1176682785153389)),(to_sfixed_a(-0.06888938695192337)),(to_sfixed_a(-0.10890021920204163)),(to_sfixed_a(-0.19557324051856995)),(to_sfixed_a(0.24219810962677002)),(to_sfixed_a(0.02036578767001629)),(to_sfixed_a(-0.18125778436660767)),(to_sfixed_a(-0.13958041369915009)),(to_sfixed_a(-0.09243994951248169)),(to_sfixed_a(0.03162984177470207)),(to_sfixed_a(-0.1397714465856552)),(to_sfixed_a(-0.15123344957828522)),(to_sfixed_a(-0.0808444693684578)),(to_sfixed_a(0.21747279167175293)),(to_sfixed_a(7.162959809647873e-05)),(to_sfixed_a(-7.649597682757303e-05)),(to_sfixed_a(3.634066888480447e-05)),(to_sfixed_a(0.00010307905176887289)),(to_sfixed_a(4.484701275941916e-05)),(to_sfixed_a(-6.946035682631191e-06)),(to_sfixed_a(0.000267314026132226)),(to_sfixed_a(-0.0002348503767279908)),(to_sfixed_a(-0.05649681016802788)),(to_sfixed_a(-0.07119841128587723)),(to_sfixed_a(-0.2138209193944931)),(to_sfixed_a(-0.0889916941523552)),(to_sfixed_a(-0.15904545783996582)),(to_sfixed_a(-0.26433607935905457)),(to_sfixed_a(-0.04843030124902725)),(to_sfixed_a(0.015525979921221733)),(to_sfixed_a(0.00029625376919284463)),(to_sfixed_a(0.09961730241775513)),(to_sfixed_a(-0.08988707512617111)),(to_sfixed_a(0.07512310892343521)),(to_sfixed_a(-0.042198602110147476)),(to_sfixed_a(0.11226072907447815)),(to_sfixed_a(-0.06424987316131592)),(to_sfixed_a(-0.07365092635154724)),(to_sfixed_a(-0.0654987245798111)),(to_sfixed_a(0.13355664908885956)),(to_sfixed_a(0.055226318538188934)),(to_sfixed_a(0.007299893070012331)),(to_sfixed_a(-0.1183227151632309)),(to_sfixed_a(-0.00012454920215532184)),(to_sfixed_a(-7.35646317480132e-05)),(to_sfixed_a(-0.00012252926535438746)),(to_sfixed_a(-0.00025664069107733667)),(to_sfixed_a(-0.00012769091699738055)),(to_sfixed_a(-0.00016591584426350892)),(to_sfixed_a(-0.00013153083273209631)),(to_sfixed_a(-0.04668572545051575)),(to_sfixed_a(0.0008091052295640111)),(to_sfixed_a(-0.11823111027479172)),(to_sfixed_a(-0.07708434015512466)),(to_sfixed_a(-0.30190786719322205)),(to_sfixed_a(-0.018463807180523872)),(to_sfixed_a(-0.14008860290050507)),(to_sfixed_a(-0.17285145819187164)),(to_sfixed_a(0.2536349296569824)),(to_sfixed_a(0.3467632234096527)),(to_sfixed_a(0.1259981244802475)),(to_sfixed_a(-0.07850561290979385)),(to_sfixed_a(-0.0396231971681118)),(to_sfixed_a(-0.06724733114242554)),(to_sfixed_a(-0.04374051094055176)),(to_sfixed_a(-0.16764385998249054)),(to_sfixed_a(-0.38938504457473755)),(to_sfixed_a(-0.09311895817518234)),(to_sfixed_a(0.3354151248931885)),(to_sfixed_a(-0.0008336447644978762)),(to_sfixed_a(-0.11661506444215775)),(to_sfixed_a(-0.00030217727180570364)),(to_sfixed_a(-6.275168561842293e-05)),(to_sfixed_a(-7.215433925011894e-06)),(to_sfixed_a(-3.2057007047114894e-05)),(to_sfixed_a(-7.823541818652302e-05)),(to_sfixed_a(-7.106606790330261e-05)),(to_sfixed_a(8.629407966509461e-05)),(to_sfixed_a(-0.00021122870384715497)),(to_sfixed_a(-0.046928729861974716)),(to_sfixed_a(0.00745473662391305)),(to_sfixed_a(-0.2151174247264862)),(to_sfixed_a(-0.13215860724449158)),(to_sfixed_a(-0.0060606542974710464)),(to_sfixed_a(0.09899847954511642)),(to_sfixed_a(-0.028816035017371178)),(to_sfixed_a(0.14081214368343353)),(to_sfixed_a(0.02981039322912693)),(to_sfixed_a(-0.0241754949092865)),(to_sfixed_a(0.10628047585487366)),(to_sfixed_a(0.11190882325172424)),(to_sfixed_a(-0.05252726376056671)),(to_sfixed_a(0.002533236052840948)),(to_sfixed_a(0.02376389130949974)),(to_sfixed_a(-0.0296358410269022)),(to_sfixed_a(-0.031292181462049484)),(to_sfixed_a(-0.15487511456012726)),(to_sfixed_a(-0.006271626800298691)),(to_sfixed_a(-1.0146431122848298e-05)),(to_sfixed_a(2.875497557397466e-05)),(to_sfixed_a(-3.356713932589628e-05)),(to_sfixed_a(-9.549684909870848e-05)),(to_sfixed_a(-0.00023903556575533003)),(to_sfixed_a(9.777572267921641e-05)),(to_sfixed_a(5.625990525004454e-05)),(to_sfixed_a(-6.580712943105027e-05)),(to_sfixed_a(-0.00041055865585803986)),(to_sfixed_a(0.015629244968295097)),(to_sfixed_a(-0.019313830882310867)),(to_sfixed_a(0.06497838348150253)),(to_sfixed_a(0.03969530761241913)),(to_sfixed_a(-0.0028550466522574425)),(to_sfixed_a(0.06644735485315323)),(to_sfixed_a(-0.030908668413758278)),(to_sfixed_a(0.050328340381383896)),(to_sfixed_a(0.13056470453739166)),(to_sfixed_a(0.0044177924282848835)),(to_sfixed_a(-0.03579352796077728)),(to_sfixed_a(0.3007063567638397)),(to_sfixed_a(-0.018318625167012215)),(to_sfixed_a(-0.03799862787127495)),(to_sfixed_a(0.2313663810491562)),(to_sfixed_a(-0.04308691620826721)),(to_sfixed_a(0.21453642845153809)),(to_sfixed_a(-0.007383568212389946)),(to_sfixed_a(0.1624637097120285)),(to_sfixed_a(-2.8471977202570997e-06)),(to_sfixed_a(0.0001586935541126877)),(to_sfixed_a(-0.00010275063687004149)),(to_sfixed_a(5.729604163207114e-05)),(to_sfixed_a(5.854979463038035e-05)),(to_sfixed_a(8.279213216155767e-05)),(to_sfixed_a(-8.996743417810649e-05)),(to_sfixed_a(-9.393491200171411e-05)),(to_sfixed_a(-0.07211201637983322)),(to_sfixed_a(0.0033522050362080336)),(to_sfixed_a(-0.29933226108551025)),(to_sfixed_a(-0.18973524868488312)),(to_sfixed_a(-0.07708225399255753)),(to_sfixed_a(-0.0681142657995224)),(to_sfixed_a(-0.02861202508211136)),(to_sfixed_a(0.18145343661308289)),(to_sfixed_a(0.08561132848262787)),(to_sfixed_a(-0.10087792575359344)),(to_sfixed_a(0.14898893237113953)),(to_sfixed_a(0.07104746997356415)),(to_sfixed_a(0.007864448241889477)),(to_sfixed_a(0.009730542078614235)),(to_sfixed_a(-0.05818244814872742)),(to_sfixed_a(0.1694507896900177)),(to_sfixed_a(-0.005133577156811953)),(to_sfixed_a(0.18001128733158112)),(to_sfixed_a(0.08158402144908905)),(to_sfixed_a(-0.005996671970933676)),(to_sfixed_a(-6.89281223458238e-05)),(to_sfixed_a(-8.444801642326638e-05)),(to_sfixed_a(0.0004473002627491951)),(to_sfixed_a(0.00016271004278678447)),(to_sfixed_a(-5.547650653170422e-05)),(to_sfixed_a(-0.00019547842384781688)),(to_sfixed_a(-0.00020763781503774226)),(to_sfixed_a(-3.211611692677252e-05)),(to_sfixed_a(-0.0002334356540814042)),(to_sfixed_a(-0.037781305611133575)),(to_sfixed_a(-0.18066909909248352)),(to_sfixed_a(-0.1642087996006012)),(to_sfixed_a(-0.15576781332492828)),(to_sfixed_a(0.012751097790896893)),(to_sfixed_a(-0.2542774975299835)),(to_sfixed_a(-0.07287537306547165)),(to_sfixed_a(-0.06870690733194351)),(to_sfixed_a(-0.04162006080150604)),(to_sfixed_a(0.08249829709529877)),(to_sfixed_a(-0.0004611636104527861)),(to_sfixed_a(0.17279614508152008)),(to_sfixed_a(0.0752858892083168)),(to_sfixed_a(0.007058217190206051)),(to_sfixed_a(0.013224725611507893)),(to_sfixed_a(-0.01391254086047411)),(to_sfixed_a(-0.0007348176441155374)),(to_sfixed_a(-0.0014842725358903408)),(to_sfixed_a(-0.002138787182047963)),(to_sfixed_a(0.0001889597624540329)),(to_sfixed_a(0.00014676936552859843)),(to_sfixed_a(0.00015715553308837116)),(to_sfixed_a(7.055084279272705e-05)),(to_sfixed_a(0.00013870580005459487)),(to_sfixed_a(2.2689217075821944e-05)),(to_sfixed_a(-9.590700938133523e-05)),(to_sfixed_a(-0.0003600929630920291)),(to_sfixed_a(7.57170855649747e-05)),(to_sfixed_a(-0.00010682287393137813)),(to_sfixed_a(-9.446278272662312e-05)),(to_sfixed_a(-0.0002521787246223539)),(to_sfixed_a(-6.964921340113506e-05)),(to_sfixed_a(0.0002375917974859476)),(to_sfixed_a(-0.009158694185316563)),(to_sfixed_a(-0.0028822252061218023)),(to_sfixed_a(-0.00041713693644851446)),(to_sfixed_a(-0.010461854748427868)),(to_sfixed_a(-0.08460540324449539)),(to_sfixed_a(-0.0031073852442204952)),(to_sfixed_a(-0.002546908101066947)),(to_sfixed_a(-0.007160363253206015)),(to_sfixed_a(-0.012250948697328568)),(to_sfixed_a(-0.008079725317656994)),(to_sfixed_a(-0.0019427173538133502)),(to_sfixed_a(-0.00014544531586579978)),(to_sfixed_a(-0.00020131752535235137)),(to_sfixed_a(0.00010199384269071743)),(to_sfixed_a(-9.496917482465506e-05)),(to_sfixed_a(0.00018383990391157568)),(to_sfixed_a(-6.762716657249257e-05)),(to_sfixed_a(-5.07950026076287e-05)),(to_sfixed_a(-0.00024136187857948244)),(to_sfixed_a(-0.0002829649893101305)),(to_sfixed_a(0.00011259485472692177)),(to_sfixed_a(0.0002331918221898377)),(to_sfixed_a(5.51520315639209e-06)),(to_sfixed_a(-2.104270606650971e-05)),(to_sfixed_a(-3.366324745002203e-05)),(to_sfixed_a(0.00010304342868039384)),(to_sfixed_a(0.00018203230865765363)),(to_sfixed_a(0.0001512024027761072)),(to_sfixed_a(0.0002964752202387899)),(to_sfixed_a(2.563509769970551e-05)),(to_sfixed_a(-0.00020322170166764408)),(to_sfixed_a(0.00018976465798914433)),(to_sfixed_a(0.00026093574706465006)),(to_sfixed_a(8.848186553223059e-05)),(to_sfixed_a(-1.494535717938561e-05)),(to_sfixed_a(-0.0002943199942819774)),(to_sfixed_a(-0.00011826066474895924)),(to_sfixed_a(-5.4492513299919665e-05)),(to_sfixed_a(-0.0001678004628047347)),(to_sfixed_a(5.822872117278166e-05)),(to_sfixed_a(-0.00025969650596380234)),(to_sfixed_a(7.14767593308352e-05)),(to_sfixed_a(-0.0001035414679790847)),(to_sfixed_a(9.00485465535894e-05)),(to_sfixed_a(0.00022152015299070626)),(to_sfixed_a(7.904231460997835e-05)));

    constant weight_n0_32 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(2.589764108051895e-06)),(to_sfixed_a(-0.0001434392761439085)),(to_sfixed_a(0.00017276150174438953)),(to_sfixed_a(-0.00012160986079834402)),(to_sfixed_a(-0.00022851451649330556)),(to_sfixed_a(-0.0002528642653487623)),(to_sfixed_a(-0.00029124243883416057)),(to_sfixed_a(0.0002182076423196122)),(to_sfixed_a(0.00023309135576710105)),(to_sfixed_a(-6.118967576185241e-06)),(to_sfixed_a(-9.293396578868851e-05)),(to_sfixed_a(-2.1361649487516843e-05)),(to_sfixed_a(-0.00020294632122386247)),(to_sfixed_a(0.0003980742476414889)),(to_sfixed_a(0.00010929234849754721)),(to_sfixed_a(-0.000134915899252519)),(to_sfixed_a(-0.0001758273137966171)),(to_sfixed_a(-0.00010571284656180069)),(to_sfixed_a(0.00011240585445193574)),(to_sfixed_a(-0.00018497528799343854)),(to_sfixed_a(-0.00020356786262709647)),(to_sfixed_a(8.405917469644919e-05)),(to_sfixed_a(-6.8512192228809e-05)),(to_sfixed_a(0.00012722646351903677)),(to_sfixed_a(0.00019960325153078884)),(to_sfixed_a(-3.91539215343073e-05)),(to_sfixed_a(-0.0001940354995895177)),(to_sfixed_a(-0.00011612648813752457)),(to_sfixed_a(-0.00011906869622180238)),(to_sfixed_a(8.608197094872594e-05)),(to_sfixed_a(-4.3695676140487194e-05)),(to_sfixed_a(-0.0003502968465909362)),(to_sfixed_a(-0.00010792538523674011)),(to_sfixed_a(-2.1819765606778674e-05)),(to_sfixed_a(-0.00013922201469540596)),(to_sfixed_a(2.708346187318966e-07)),(to_sfixed_a(3.1502244382863864e-05)),(to_sfixed_a(0.00013564406253863126)),(to_sfixed_a(1.4611168808187358e-05)),(to_sfixed_a(-0.00018418255785945803)),(to_sfixed_a(-3.77290380129125e-05)),(to_sfixed_a(3.325031138956547e-05)),(to_sfixed_a(6.975654741836479e-06)),(to_sfixed_a(0.00010512669541640207)),(to_sfixed_a(-1.4417631064134184e-05)),(to_sfixed_a(0.00038039745413698256)),(to_sfixed_a(-0.00014493399066850543)),(to_sfixed_a(0.0001716376282274723)),(to_sfixed_a(-3.974495120928623e-05)),(to_sfixed_a(0.00035843445220962167)),(to_sfixed_a(-9.86068625934422e-05)),(to_sfixed_a(1.745854751789011e-05)),(to_sfixed_a(2.9187422114773653e-05)),(to_sfixed_a(2.762623807939235e-05)),(to_sfixed_a(-0.00015673354209866375)),(to_sfixed_a(-8.262971277872566e-06)),(to_sfixed_a(-9.967074583983049e-05)),(to_sfixed_a(-0.0003290653112344444)),(to_sfixed_a(7.436699524987489e-05)),(to_sfixed_a(0.00010256393579766154)),(to_sfixed_a(-0.00033678143518045545)),(to_sfixed_a(5.233764386503026e-05)),(to_sfixed_a(-5.3342209866968915e-06)),(to_sfixed_a(-0.00011517074017319828)),(to_sfixed_a(1.172479460365139e-05)),(to_sfixed_a(-6.962127372389659e-05)),(to_sfixed_a(0.00014386222756002098)),(to_sfixed_a(0.00010721399303292856)),(to_sfixed_a(-9.251990377379116e-06)),(to_sfixed_a(0.015440764836966991)),(to_sfixed_a(0.0001115667910198681)),(to_sfixed_a(0.0001298486749874428)),(to_sfixed_a(-0.0001440512714907527)),(to_sfixed_a(-6.788846803829074e-05)),(to_sfixed_a(5.177565981284715e-05)),(to_sfixed_a(-0.00022193403856363147)),(to_sfixed_a(0.0001620194670977071)),(to_sfixed_a(-6.114074494689703e-05)),(to_sfixed_a(7.652006024727598e-05)),(to_sfixed_a(-0.0003529250680003315)),(to_sfixed_a(-7.98465553089045e-05)),(to_sfixed_a(2.3236454580910504e-05)),(to_sfixed_a(0.0003203601227141917)),(to_sfixed_a(0.00014370410644914955)),(to_sfixed_a(-2.7192189008928835e-05)),(to_sfixed_a(1.675618113949895e-05)),(to_sfixed_a(-6.385153392329812e-05)),(to_sfixed_a(6.573526479769498e-05)),(to_sfixed_a(-0.0002613795513752848)),(to_sfixed_a(6.996267620706931e-05)),(to_sfixed_a(0.00011260976316407323)),(to_sfixed_a(-0.0002991393266711384)),(to_sfixed_a(0.05940299108624458)),(to_sfixed_a(-8.068147144513205e-05)),(to_sfixed_a(0.06754381209611893)),(to_sfixed_a(-0.07593285292387009)),(to_sfixed_a(0.015287719666957855)),(to_sfixed_a(-0.1410147249698639)),(to_sfixed_a(0.13851536810398102)),(to_sfixed_a(0.09973737597465515)),(to_sfixed_a(-0.004486073739826679)),(to_sfixed_a(-0.03351910039782524)),(to_sfixed_a(0.07446770370006561)),(to_sfixed_a(0.08589833974838257)),(to_sfixed_a(0.030695827677845955)),(to_sfixed_a(0.06218996271491051)),(to_sfixed_a(-4.098617137060501e-05)),(to_sfixed_a(3.5894783650292084e-05)),(to_sfixed_a(-0.00013913874863646924)),(to_sfixed_a(-5.828905341331847e-05)),(to_sfixed_a(4.5213131670607254e-05)),(to_sfixed_a(-0.00014637834101449698)),(to_sfixed_a(-0.0002735272573772818)),(to_sfixed_a(-3.5891560401069e-05)),(to_sfixed_a(0.0001634296786505729)),(to_sfixed_a(2.3303235138882883e-05)),(to_sfixed_a(-9.897536074277014e-05)),(to_sfixed_a(0.00015959699521772563)),(to_sfixed_a(-0.000622364750597626)),(to_sfixed_a(-0.09428201615810394)),(to_sfixed_a(-0.035811085253953934)),(to_sfixed_a(0.08641970157623291)),(to_sfixed_a(0.04247445613145828)),(to_sfixed_a(-0.10517636686563492)),(to_sfixed_a(-0.08448796719312668)),(to_sfixed_a(-0.2522713243961334)),(to_sfixed_a(0.21382588148117065)),(to_sfixed_a(-0.13803064823150635)),(to_sfixed_a(-0.06989958137273788)),(to_sfixed_a(-0.20261667668819427)),(to_sfixed_a(-0.12288523465394974)),(to_sfixed_a(0.0685390830039978)),(to_sfixed_a(0.0289777759462595)),(to_sfixed_a(0.027185767889022827)),(to_sfixed_a(0.006032662466168404)),(to_sfixed_a(0.00012911620433442295)),(to_sfixed_a(-0.0013718530535697937)),(to_sfixed_a(-0.00013232500350568444)),(to_sfixed_a(2.161957490898203e-05)),(to_sfixed_a(-5.4787724366178736e-05)),(to_sfixed_a(0.00024540306185372174)),(to_sfixed_a(-0.00012025439355056733)),(to_sfixed_a(-0.00014866601850371808)),(to_sfixed_a(0.00010235208901576698)),(to_sfixed_a(-0.000524758652318269)),(to_sfixed_a(-0.14309333264827728)),(to_sfixed_a(-0.006706268992275)),(to_sfixed_a(-0.09363085776567459)),(to_sfixed_a(0.04548060894012451)),(to_sfixed_a(0.021371306851506233)),(to_sfixed_a(-0.005435141734778881)),(to_sfixed_a(-0.0030606435611844063)),(to_sfixed_a(0.19480471312999725)),(to_sfixed_a(0.1744859665632248)),(to_sfixed_a(-0.05803268030285835)),(to_sfixed_a(-0.05774126201868057)),(to_sfixed_a(-0.016682041808962822)),(to_sfixed_a(-0.11281926929950714)),(to_sfixed_a(0.17308840155601501)),(to_sfixed_a(0.2554265558719635)),(to_sfixed_a(0.1320902407169342)),(to_sfixed_a(0.10423523932695389)),(to_sfixed_a(-0.002168591134250164)),(to_sfixed_a(0.041446857154369354)),(to_sfixed_a(0.0005255045252852142)),(to_sfixed_a(-0.0001563978148624301)),(to_sfixed_a(-7.192078192019835e-05)),(to_sfixed_a(7.267255568876863e-05)),(to_sfixed_a(8.686073124408722e-05)),(to_sfixed_a(0.0001427860406693071)),(to_sfixed_a(0.0002935251977760345)),(to_sfixed_a(5.4496504162671044e-05)),(to_sfixed_a(-0.00019364373292773962)),(to_sfixed_a(-0.13786770403385162)),(to_sfixed_a(-0.11885369569063187)),(to_sfixed_a(-0.14588072896003723)),(to_sfixed_a(-0.03581538796424866)),(to_sfixed_a(-0.2292720377445221)),(to_sfixed_a(0.27559584379196167)),(to_sfixed_a(0.25202447175979614)),(to_sfixed_a(0.26825615763664246)),(to_sfixed_a(0.14269934594631195)),(to_sfixed_a(-0.04746202751994133)),(to_sfixed_a(0.11987106502056122)),(to_sfixed_a(0.14439362287521362)),(to_sfixed_a(-0.11393433064222336)),(to_sfixed_a(-0.21622289717197418)),(to_sfixed_a(0.08430170267820358)),(to_sfixed_a(0.13085752725601196)),(to_sfixed_a(-0.17962424457073212)),(to_sfixed_a(0.07321402430534363)),(to_sfixed_a(0.07980527728796005)),(to_sfixed_a(0.001697380794212222)),(to_sfixed_a(0.0026553585194051266)),(to_sfixed_a(2.7206311642657965e-05)),(to_sfixed_a(7.130185258574784e-05)),(to_sfixed_a(0.0001658687397139147)),(to_sfixed_a(-0.00013146636774763465)),(to_sfixed_a(4.382199404062703e-05)),(to_sfixed_a(0.0001084384712157771)),(to_sfixed_a(-9.420670539839193e-05)),(to_sfixed_a(-0.04933329299092293)),(to_sfixed_a(-0.22249950468540192)),(to_sfixed_a(-0.032687410712242126)),(to_sfixed_a(-0.0040446179918944836)),(to_sfixed_a(0.09853166341781616)),(to_sfixed_a(0.18877851963043213)),(to_sfixed_a(-0.0173850916326046)),(to_sfixed_a(0.07434115558862686)),(to_sfixed_a(-0.08764202147722244)),(to_sfixed_a(0.04258757829666138)),(to_sfixed_a(0.3991721570491791)),(to_sfixed_a(0.009281668812036514)),(to_sfixed_a(-0.05509011447429657)),(to_sfixed_a(0.12893199920654297)),(to_sfixed_a(-0.4507445693016052)),(to_sfixed_a(0.08170993626117706)),(to_sfixed_a(-0.07721653580665588)),(to_sfixed_a(-0.00784184131771326)),(to_sfixed_a(-0.15760545432567596)),(to_sfixed_a(-0.050627704709768295)),(to_sfixed_a(-0.009589401073753834)),(to_sfixed_a(0.000242047623032704)),(to_sfixed_a(-0.0003161122731398791)),(to_sfixed_a(6.796023808419704e-05)),(to_sfixed_a(-0.00014395029575098306)),(to_sfixed_a(2.3327202143264003e-05)),(to_sfixed_a(-3.107385782641359e-05)),(to_sfixed_a(-0.018306216225028038)),(to_sfixed_a(0.028363699093461037)),(to_sfixed_a(-0.06988635659217834)),(to_sfixed_a(0.06268413364887238)),(to_sfixed_a(0.019830897450447083)),(to_sfixed_a(0.025401026010513306)),(to_sfixed_a(-0.07987931370735168)),(to_sfixed_a(-0.13932690024375916)),(to_sfixed_a(-0.1016930565237999)),(to_sfixed_a(-0.12919187545776367)),(to_sfixed_a(-0.236967995762825)),(to_sfixed_a(-0.10888451337814331)),(to_sfixed_a(-0.24833276867866516)),(to_sfixed_a(-0.23178631067276)),(to_sfixed_a(-0.06512026488780975)),(to_sfixed_a(-0.12959721684455872)),(to_sfixed_a(0.021440895274281502)),(to_sfixed_a(0.04063611477613449)),(to_sfixed_a(-0.3879053592681885)),(to_sfixed_a(-0.02124856226146221)),(to_sfixed_a(-0.19188712537288666)),(to_sfixed_a(0.013029411435127258)),(to_sfixed_a(0.00015772551705595106)),(to_sfixed_a(0.00018368876772001386)),(to_sfixed_a(-0.0001857886090874672)),(to_sfixed_a(-1.3396414942690171e-05)),(to_sfixed_a(-2.6904364858637564e-05)),(to_sfixed_a(-0.00011225149501115084)),(to_sfixed_a(-0.0028621158562600613)),(to_sfixed_a(-0.0858345702290535)),(to_sfixed_a(-0.03833940252661705)),(to_sfixed_a(-0.14242948591709137)),(to_sfixed_a(-0.010159142315387726)),(to_sfixed_a(0.13247227668762207)),(to_sfixed_a(-0.02959500066936016)),(to_sfixed_a(0.021533025428652763)),(to_sfixed_a(-0.03991219028830528)),(to_sfixed_a(-0.03852704539895058)),(to_sfixed_a(-0.2503407895565033)),(to_sfixed_a(0.0388832613825798)),(to_sfixed_a(0.16721542179584503)),(to_sfixed_a(0.2683942914009094)),(to_sfixed_a(0.02688984014093876)),(to_sfixed_a(0.1330782175064087)),(to_sfixed_a(-0.022596541792154312)),(to_sfixed_a(-0.04050667583942413)),(to_sfixed_a(0.015130724757909775)),(to_sfixed_a(-0.0389418788254261)),(to_sfixed_a(-0.10237722098827362)),(to_sfixed_a(8.067620365181938e-05)),(to_sfixed_a(-0.00013410981046035886)),(to_sfixed_a(-0.00013853158452548087)),(to_sfixed_a(-0.00019333753152750432)),(to_sfixed_a(-0.0002113699883921072)),(to_sfixed_a(0.0001059755522874184)),(to_sfixed_a(0.00017641960585024208)),(to_sfixed_a(-0.008087065070867538)),(to_sfixed_a(-0.03726969286799431)),(to_sfixed_a(0.02897948957979679)),(to_sfixed_a(0.23516185581684113)),(to_sfixed_a(0.3917222023010254)),(to_sfixed_a(0.17875303328037262)),(to_sfixed_a(0.25357913970947266)),(to_sfixed_a(-0.22762571275234222)),(to_sfixed_a(0.10638141632080078)),(to_sfixed_a(0.15260405838489532)),(to_sfixed_a(-0.18381306529045105)),(to_sfixed_a(-0.0894593670964241)),(to_sfixed_a(-0.10878970474004745)),(to_sfixed_a(0.07321377098560333)),(to_sfixed_a(0.1022929847240448)),(to_sfixed_a(0.18446442484855652)),(to_sfixed_a(-0.24465593695640564)),(to_sfixed_a(-0.031019283458590508)),(to_sfixed_a(-0.10109210014343262)),(to_sfixed_a(-0.07466411590576172)),(to_sfixed_a(-0.050881922245025635)),(to_sfixed_a(-0.07274985313415527)),(to_sfixed_a(4.387934677652083e-05)),(to_sfixed_a(-0.00015760568203404546)),(to_sfixed_a(7.083137461449951e-05)),(to_sfixed_a(0.0001601028343429789)),(to_sfixed_a(-6.057776772649959e-05)),(to_sfixed_a(-0.007221960928291082)),(to_sfixed_a(-0.11567354947328568)),(to_sfixed_a(0.09036403149366379)),(to_sfixed_a(0.1620536893606186)),(to_sfixed_a(0.11863264441490173)),(to_sfixed_a(0.048704370856285095)),(to_sfixed_a(-0.21678657829761505)),(to_sfixed_a(-0.039918504655361176)),(to_sfixed_a(0.026310406625270844)),(to_sfixed_a(-0.1805085390806198)),(to_sfixed_a(-0.1381259709596634)),(to_sfixed_a(0.07032277435064316)),(to_sfixed_a(-0.16423293948173523)),(to_sfixed_a(0.04474879801273346)),(to_sfixed_a(-0.21630991995334625)),(to_sfixed_a(-0.20281198620796204)),(to_sfixed_a(0.08112015575170517)),(to_sfixed_a(-0.022543897852301598)),(to_sfixed_a(-0.012425053864717484)),(to_sfixed_a(-0.005381404887884855)),(to_sfixed_a(0.03133666142821312)),(to_sfixed_a(-0.0035106269642710686)),(to_sfixed_a(3.5403703805059195e-05)),(to_sfixed_a(-5.02465127283358e-06)),(to_sfixed_a(0.00022873308626003563)),(to_sfixed_a(-0.00026025951956398785)),(to_sfixed_a(3.490993185550906e-05)),(to_sfixed_a(-0.00010160644887946546)),(to_sfixed_a(-0.0002716233138926327)),(to_sfixed_a(0.004980041645467281)),(to_sfixed_a(-0.11926020681858063)),(to_sfixed_a(0.12169419229030609)),(to_sfixed_a(0.07735291123390198)),(to_sfixed_a(0.07360547035932541)),(to_sfixed_a(0.25897565484046936)),(to_sfixed_a(-0.03707878664135933)),(to_sfixed_a(0.1814797818660736)),(to_sfixed_a(-0.08838150650262833)),(to_sfixed_a(0.07513174414634705)),(to_sfixed_a(0.09501276165246964)),(to_sfixed_a(0.30701544880867004)),(to_sfixed_a(-0.03916981443762779)),(to_sfixed_a(-0.42488551139831543)),(to_sfixed_a(-0.28669479489326477)),(to_sfixed_a(-0.18149220943450928)),(to_sfixed_a(0.03078218549489975)),(to_sfixed_a(-0.0005634701810777187)),(to_sfixed_a(0.10207848995923996)),(to_sfixed_a(0.08273891359567642)),(to_sfixed_a(0.11438696086406708)),(to_sfixed_a(6.504291377495974e-05)),(to_sfixed_a(-0.00040226170676760375)),(to_sfixed_a(2.537224099796731e-05)),(to_sfixed_a(-6.179865158628672e-05)),(to_sfixed_a(-0.0004129692679271102)),(to_sfixed_a(-9.144790965365246e-05)),(to_sfixed_a(-5.0833816203521565e-05)),(to_sfixed_a(-0.08145427703857422)),(to_sfixed_a(0.29592886567115784)),(to_sfixed_a(0.2998674213886261)),(to_sfixed_a(0.1473691314458847)),(to_sfixed_a(0.057267963886260986)),(to_sfixed_a(-0.034952301532030106)),(to_sfixed_a(0.030639395117759705)),(to_sfixed_a(0.09616692364215851)),(to_sfixed_a(0.15544842183589935)),(to_sfixed_a(0.23057842254638672)),(to_sfixed_a(0.13038477301597595)),(to_sfixed_a(0.12747427821159363)),(to_sfixed_a(0.1592312604188919)),(to_sfixed_a(0.02760910987854004)),(to_sfixed_a(0.05047251656651497)),(to_sfixed_a(-0.04977641999721527)),(to_sfixed_a(-0.15017452836036682)),(to_sfixed_a(-0.023495325818657875)),(to_sfixed_a(-0.07386118173599243)),(to_sfixed_a(0.1803218573331833)),(to_sfixed_a(0.0735110491514206)),(to_sfixed_a(-0.002075615106150508)),(to_sfixed_a(-0.0028840978629887104)),(to_sfixed_a(-0.000110713837784715)),(to_sfixed_a(0.00017447583377361298)),(to_sfixed_a(2.0649193174904212e-05)),(to_sfixed_a(-0.00017630266665946692)),(to_sfixed_a(-2.3837961634853855e-05)),(to_sfixed_a(-0.000428132334491238)),(to_sfixed_a(0.016524052247405052)),(to_sfixed_a(-0.1374868005514145)),(to_sfixed_a(0.08251402527093887)),(to_sfixed_a(-0.01763956807553768)),(to_sfixed_a(0.1572428196668625)),(to_sfixed_a(0.14708425104618073)),(to_sfixed_a(-0.05010148882865906)),(to_sfixed_a(-0.0956963449716568)),(to_sfixed_a(0.03182687610387802)),(to_sfixed_a(0.22811667621135712)),(to_sfixed_a(0.1163419708609581)),(to_sfixed_a(0.24148915708065033)),(to_sfixed_a(0.031119193881750107)),(to_sfixed_a(0.22131307423114777)),(to_sfixed_a(0.24461044371128082)),(to_sfixed_a(0.05293119698762894)),(to_sfixed_a(-0.051134347915649414)),(to_sfixed_a(0.07004071772098541)),(to_sfixed_a(-0.11537499725818634)),(to_sfixed_a(-0.04796300455927849)),(to_sfixed_a(0.0003336480294819921)),(to_sfixed_a(5.161946319276467e-05)),(to_sfixed_a(-0.0001322456228081137)),(to_sfixed_a(3.580813790904358e-05)),(to_sfixed_a(0.0002256254811072722)),(to_sfixed_a(0.00014530261978507042)),(to_sfixed_a(0.00029291133978404105)),(to_sfixed_a(-0.011320228688418865)),(to_sfixed_a(-0.0954727753996849)),(to_sfixed_a(-0.11153594404459)),(to_sfixed_a(-0.2319220006465912)),(to_sfixed_a(-0.18083813786506653)),(to_sfixed_a(-0.16536399722099304)),(to_sfixed_a(-0.025138305500149727)),(to_sfixed_a(-0.09427409619092941)),(to_sfixed_a(0.015101495198905468)),(to_sfixed_a(-0.18445737659931183)),(to_sfixed_a(0.09646584093570709)),(to_sfixed_a(0.16917982697486877)),(to_sfixed_a(-0.0036745723336935043)),(to_sfixed_a(0.18971988558769226)),(to_sfixed_a(-0.06368666887283325)),(to_sfixed_a(-0.24166826903820038)),(to_sfixed_a(0.15751902759075165)),(to_sfixed_a(0.018056286498904228)),(to_sfixed_a(-0.05006202682852745)),(to_sfixed_a(-0.21420380473136902)),(to_sfixed_a(-0.2077312022447586)),(to_sfixed_a(-0.0001473867305321619)),(to_sfixed_a(1.68967671925202e-05)),(to_sfixed_a(6.613508594455197e-05)),(to_sfixed_a(0.00010672663484001532)),(to_sfixed_a(3.373820072738454e-05)),(to_sfixed_a(0.0006284762057475746)),(to_sfixed_a(0.00419491296634078)),(to_sfixed_a(-0.03473835811018944)),(to_sfixed_a(0.028673024848103523)),(to_sfixed_a(0.09957192838191986)),(to_sfixed_a(-0.012849811464548111)),(to_sfixed_a(0.013295860961079597)),(to_sfixed_a(0.08442194014787674)),(to_sfixed_a(-0.3204008638858795)),(to_sfixed_a(0.01735297590494156)),(to_sfixed_a(0.06520681083202362)),(to_sfixed_a(0.013196642510592937)),(to_sfixed_a(0.10777821391820908)),(to_sfixed_a(0.09010849893093109)),(to_sfixed_a(-0.055630315095186234)),(to_sfixed_a(-0.1479761302471161)),(to_sfixed_a(0.022365843877196312)),(to_sfixed_a(0.13145828247070312)),(to_sfixed_a(0.06074976176023483)),(to_sfixed_a(0.16756777465343475)),(to_sfixed_a(0.13976797461509705)),(to_sfixed_a(0.020937198773026466)),(to_sfixed_a(-0.002118652453646064)),(to_sfixed_a(0.0011910126777365804)),(to_sfixed_a(-0.00018352946790400892)),(to_sfixed_a(-1.9635130229289643e-05)),(to_sfixed_a(-0.0001854794390965253)),(to_sfixed_a(0.0002967939944937825)),(to_sfixed_a(0.0027318557258695364)),(to_sfixed_a(0.003971211612224579)),(to_sfixed_a(0.043963853269815445)),(to_sfixed_a(-0.03903884440660477)),(to_sfixed_a(0.07597287744283676)),(to_sfixed_a(0.05484018102288246)),(to_sfixed_a(0.1747598648071289)),(to_sfixed_a(0.035453710705041885)),(to_sfixed_a(0.03642283007502556)),(to_sfixed_a(-0.03823558986186981)),(to_sfixed_a(0.048074424266815186)),(to_sfixed_a(-0.07861354202032089)),(to_sfixed_a(-0.09785307198762894)),(to_sfixed_a(0.2347615361213684)),(to_sfixed_a(-0.13481475412845612)),(to_sfixed_a(-0.062405407428741455)),(to_sfixed_a(0.04340699687600136)),(to_sfixed_a(-0.00790938176214695)),(to_sfixed_a(0.26176393032073975)),(to_sfixed_a(0.019539320841431618)),(to_sfixed_a(0.059296805411577225)),(to_sfixed_a(0.01890646666288376)),(to_sfixed_a(-6.084756751079112e-05)),(to_sfixed_a(-8.96686760825105e-05)),(to_sfixed_a(-0.00020632980158552527)),(to_sfixed_a(-0.00010008040408138186)),(to_sfixed_a(-5.768576738773845e-05)),(to_sfixed_a(-9.67984669841826e-05)),(to_sfixed_a(-0.00018520107551012188)),(to_sfixed_a(-0.037031449377536774)),(to_sfixed_a(-0.23195362091064453)),(to_sfixed_a(-0.047297582030296326)),(to_sfixed_a(0.159199059009552)),(to_sfixed_a(0.004895062185823917)),(to_sfixed_a(0.07380408048629761)),(to_sfixed_a(-0.04222428426146507)),(to_sfixed_a(-0.10310903191566467)),(to_sfixed_a(-0.004522316623479128)),(to_sfixed_a(0.1901821494102478)),(to_sfixed_a(-0.07645919919013977)),(to_sfixed_a(0.1916980743408203)),(to_sfixed_a(0.18494316935539246)),(to_sfixed_a(0.05840786173939705)),(to_sfixed_a(-0.27362775802612305)),(to_sfixed_a(0.08206894993782043)),(to_sfixed_a(0.17602220177650452)),(to_sfixed_a(0.022754890844225883)),(to_sfixed_a(0.10707405209541321)),(to_sfixed_a(-0.1926620602607727)),(to_sfixed_a(0.13006675243377686)),(to_sfixed_a(0.03468632698059082)),(to_sfixed_a(-0.00015819915279280394)),(to_sfixed_a(-0.00017982478311751038)),(to_sfixed_a(-0.00016840992611832917)),(to_sfixed_a(4.596372673404403e-05)),(to_sfixed_a(0.00024037202820181847)),(to_sfixed_a(0.00017291450058110058)),(to_sfixed_a(0.07742426544427872)),(to_sfixed_a(0.001290846150368452)),(to_sfixed_a(0.11563131213188171)),(to_sfixed_a(-0.012296071276068687)),(to_sfixed_a(-0.05341227352619171)),(to_sfixed_a(0.1506214290857315)),(to_sfixed_a(0.052194468677043915)),(to_sfixed_a(-0.03963275998830795)),(to_sfixed_a(-0.1443156749010086)),(to_sfixed_a(-0.018560854718089104)),(to_sfixed_a(0.08951643109321594)),(to_sfixed_a(0.013214148581027985)),(to_sfixed_a(0.09877745807170868)),(to_sfixed_a(0.006434533279389143)),(to_sfixed_a(0.000310048257233575)),(to_sfixed_a(-0.032375890761613846)),(to_sfixed_a(-0.12830482423305511)),(to_sfixed_a(0.15510213375091553)),(to_sfixed_a(0.009984559379518032)),(to_sfixed_a(-0.07122134417295456)),(to_sfixed_a(0.18038484454154968)),(to_sfixed_a(-0.0001805193314794451)),(to_sfixed_a(-2.9910384910181165e-05)),(to_sfixed_a(-1.3889638466935139e-05)),(to_sfixed_a(-6.421317721105879e-06)),(to_sfixed_a(0.00013160538219381124)),(to_sfixed_a(7.592196925543249e-05)),(to_sfixed_a(-7.025873856036924e-07)),(to_sfixed_a(0.0001931682782014832)),(to_sfixed_a(0.011064654216170311)),(to_sfixed_a(0.07348048686981201)),(to_sfixed_a(-0.0983906015753746)),(to_sfixed_a(-0.001965261297300458)),(to_sfixed_a(0.047350749373435974)),(to_sfixed_a(-0.362234503030777)),(to_sfixed_a(0.011651811189949512)),(to_sfixed_a(0.031338583678007126)),(to_sfixed_a(-0.050010327249765396)),(to_sfixed_a(0.10038862377405167)),(to_sfixed_a(0.07733022421598434)),(to_sfixed_a(-0.13101226091384888)),(to_sfixed_a(-0.05501218140125275)),(to_sfixed_a(-0.32142478227615356)),(to_sfixed_a(0.31518280506134033)),(to_sfixed_a(-0.15462587773799896)),(to_sfixed_a(0.051822468638420105)),(to_sfixed_a(-0.04434122517704964)),(to_sfixed_a(0.002729987958446145)),(to_sfixed_a(0.0966009721159935)),(to_sfixed_a(0.07375118136405945)),(to_sfixed_a(3.755549755624088e-07)),(to_sfixed_a(-0.0001803044433472678)),(to_sfixed_a(5.8998608437832445e-05)),(to_sfixed_a(-0.0001852225832408294)),(to_sfixed_a(3.5930734156863764e-05)),(to_sfixed_a(8.771824650466442e-05)),(to_sfixed_a(-0.0001468061818741262)),(to_sfixed_a(-0.03533115237951279)),(to_sfixed_a(-0.00019487836107145995)),(to_sfixed_a(-0.01038985513150692)),(to_sfixed_a(0.11941518634557724)),(to_sfixed_a(0.15650002658367157)),(to_sfixed_a(0.10667537152767181)),(to_sfixed_a(0.1005769670009613)),(to_sfixed_a(0.18015913665294647)),(to_sfixed_a(0.25731390714645386)),(to_sfixed_a(0.16258203983306885)),(to_sfixed_a(0.1235722005367279)),(to_sfixed_a(-0.00783667154610157)),(to_sfixed_a(-0.2004621922969818)),(to_sfixed_a(-0.07390686869621277)),(to_sfixed_a(0.154449462890625)),(to_sfixed_a(0.1711592674255371)),(to_sfixed_a(0.06538457423448563)),(to_sfixed_a(0.049614548683166504)),(to_sfixed_a(0.1875150203704834)),(to_sfixed_a(-0.0010546606499701738)),(to_sfixed_a(-0.006810266990214586)),(to_sfixed_a(7.33394845155999e-05)),(to_sfixed_a(0.000244278518948704)),(to_sfixed_a(-0.00014613034727517515)),(to_sfixed_a(-2.5840650778263807e-05)),(to_sfixed_a(2.376963857386727e-05)),(to_sfixed_a(-0.0001628230238566175)),(to_sfixed_a(-5.739982225350104e-05)),(to_sfixed_a(3.228764035156928e-05)),(to_sfixed_a(-0.11189757287502289)),(to_sfixed_a(0.02421584539115429)),(to_sfixed_a(0.005641013849526644)),(to_sfixed_a(0.053367286920547485)),(to_sfixed_a(0.02450387366116047)),(to_sfixed_a(0.46036070585250854)),(to_sfixed_a(0.13178329169750214)),(to_sfixed_a(0.19517122209072113)),(to_sfixed_a(-0.08839356154203415)),(to_sfixed_a(-0.0087073789909482)),(to_sfixed_a(0.0781116783618927)),(to_sfixed_a(0.015856992453336716)),(to_sfixed_a(0.0958237424492836)),(to_sfixed_a(0.009986547753214836)),(to_sfixed_a(-0.061470404267311096)),(to_sfixed_a(-0.0029459355864673853)),(to_sfixed_a(0.03974022716283798)),(to_sfixed_a(0.027897492051124573)),(to_sfixed_a(0.005091212689876556)),(to_sfixed_a(9.059945296030492e-05)),(to_sfixed_a(-5.3109779400983825e-05)),(to_sfixed_a(0.00013870472321286798)),(to_sfixed_a(-0.00010923163790721446)),(to_sfixed_a(-0.00010058362386189401)),(to_sfixed_a(6.0655314882751554e-05)),(to_sfixed_a(-0.00017567910254001617)),(to_sfixed_a(0.00020146789029240608)),(to_sfixed_a(0.00011215486301807687)),(to_sfixed_a(-0.02796495519578457)),(to_sfixed_a(-0.15460383892059326)),(to_sfixed_a(-0.023878125473856926)),(to_sfixed_a(0.011998915113508701)),(to_sfixed_a(0.07218564301729202)),(to_sfixed_a(0.0719129666686058)),(to_sfixed_a(-0.07262138277292252)),(to_sfixed_a(0.03905637562274933)),(to_sfixed_a(0.08450096100568771)),(to_sfixed_a(-0.019264891743659973)),(to_sfixed_a(-0.09264260530471802)),(to_sfixed_a(0.10673155635595322)),(to_sfixed_a(-0.06644532084465027)),(to_sfixed_a(-0.19865472614765167)),(to_sfixed_a(-0.07323294878005981)),(to_sfixed_a(-0.021494600921869278)),(to_sfixed_a(0.1738327443599701)),(to_sfixed_a(0.003377046901732683)),(to_sfixed_a(0.12039678543806076)),(to_sfixed_a(-4.888023340754444e-06)),(to_sfixed_a(-5.284519829729106e-06)),(to_sfixed_a(-0.00019424255879130214)),(to_sfixed_a(8.591001824242994e-05)),(to_sfixed_a(0.00010691994975786656)),(to_sfixed_a(0.00011339305638102815)),(to_sfixed_a(-0.00015656827599741518)),(to_sfixed_a(-0.0002539922425057739)),(to_sfixed_a(0.020157162100076675)),(to_sfixed_a(-0.025260047987103462)),(to_sfixed_a(0.08262445032596588)),(to_sfixed_a(0.25757497549057007)),(to_sfixed_a(-0.09017838537693024)),(to_sfixed_a(0.12645772099494934)),(to_sfixed_a(0.007353881374001503)),(to_sfixed_a(0.0796312689781189)),(to_sfixed_a(0.19950659573078156)),(to_sfixed_a(0.04919160157442093)),(to_sfixed_a(-0.13538607954978943)),(to_sfixed_a(-0.009196851402521133)),(to_sfixed_a(0.15833650529384613)),(to_sfixed_a(-0.09778513014316559)),(to_sfixed_a(0.13914687931537628)),(to_sfixed_a(0.17777687311172485)),(to_sfixed_a(-0.0007299963035620749)),(to_sfixed_a(0.16835671663284302)),(to_sfixed_a(0.055375102907419205)),(to_sfixed_a(-0.007890784181654453)),(to_sfixed_a(-9.06101122382097e-05)),(to_sfixed_a(-0.00014369368727784604)),(to_sfixed_a(-5.8608689869288355e-05)),(to_sfixed_a(1.782455001375638e-05)),(to_sfixed_a(2.1515554180950858e-05)),(to_sfixed_a(0.00010298092820448801)),(to_sfixed_a(-6.90920787747018e-05)),(to_sfixed_a(-0.0002257009909953922)),(to_sfixed_a(0.0001879468181869015)),(to_sfixed_a(-0.0072603123262524605)),(to_sfixed_a(0.05068746581673622)),(to_sfixed_a(0.023728495463728905)),(to_sfixed_a(0.23169279098510742)),(to_sfixed_a(0.16643160581588745)),(to_sfixed_a(0.10716293007135391)),(to_sfixed_a(0.005175813566893339)),(to_sfixed_a(0.06476879119873047)),(to_sfixed_a(-0.006156292278319597)),(to_sfixed_a(0.12505152821540833)),(to_sfixed_a(0.07203979790210724)),(to_sfixed_a(-0.4642889201641083)),(to_sfixed_a(-0.158610001206398)),(to_sfixed_a(-0.00987773947417736)),(to_sfixed_a(-0.029090186581015587)),(to_sfixed_a(-0.10825307667255402)),(to_sfixed_a(-0.0012445731554180384)),(to_sfixed_a(-0.004305812064558268)),(to_sfixed_a(-0.004199300426989794)),(to_sfixed_a(0.00016555105685256422)),(to_sfixed_a(1.9747782062040642e-05)),(to_sfixed_a(-5.5661515943938866e-05)),(to_sfixed_a(0.00020368928380776197)),(to_sfixed_a(-4.8071349738165736e-05)),(to_sfixed_a(-3.704552727867849e-05)),(to_sfixed_a(-8.247635560110211e-05)),(to_sfixed_a(0.00010714621748775244)),(to_sfixed_a(8.957678073784336e-05)),(to_sfixed_a(0.00034998581395484507)),(to_sfixed_a(0.00040030243690125644)),(to_sfixed_a(-0.0002711682172957808)),(to_sfixed_a(-9.955957648344338e-05)),(to_sfixed_a(0.0001004358273348771)),(to_sfixed_a(-0.06354519724845886)),(to_sfixed_a(0.0020249024964869022)),(to_sfixed_a(-0.0008215576526708901)),(to_sfixed_a(-0.052091438323259354)),(to_sfixed_a(-0.045115210115909576)),(to_sfixed_a(-0.017081422731280327)),(to_sfixed_a(0.014209304004907608)),(to_sfixed_a(-0.05136284604668617)),(to_sfixed_a(-0.07189937680959702)),(to_sfixed_a(-0.007716489490121603)),(to_sfixed_a(-0.0008297229069285095)),(to_sfixed_a(6.34976095170714e-05)),(to_sfixed_a(0.00022241460101213306)),(to_sfixed_a(-7.608256419189274e-05)),(to_sfixed_a(0.00021503058087546378)),(to_sfixed_a(0.00013601176033262163)),(to_sfixed_a(0.00017735797155182809)),(to_sfixed_a(-0.00011968802573392168)),(to_sfixed_a(-7.121761882444844e-05)),(to_sfixed_a(-0.00011507284216349944)),(to_sfixed_a(0.00021410673798527569)),(to_sfixed_a(-7.337035640375689e-05)),(to_sfixed_a(-6.723785918438807e-05)),(to_sfixed_a(0.000152700231410563)),(to_sfixed_a(-7.673478830838576e-05)),(to_sfixed_a(8.061859261943027e-05)),(to_sfixed_a(0.00011097933747805655)),(to_sfixed_a(-6.395915261236951e-05)),(to_sfixed_a(-8.655201236251742e-05)),(to_sfixed_a(-0.00014654493134003133)),(to_sfixed_a(6.0447015130193904e-05)),(to_sfixed_a(-0.00023346887610387057)),(to_sfixed_a(0.00028582336381077766)),(to_sfixed_a(-1.8387077943771146e-05)),(to_sfixed_a(-2.4483540983055718e-05)),(to_sfixed_a(0.00018526424537412822)),(to_sfixed_a(-0.00011318333417875692)),(to_sfixed_a(0.0002573724777903408)),(to_sfixed_a(8.448809967376292e-05)),(to_sfixed_a(-0.00016856346337590367)),(to_sfixed_a(3.415666287764907e-05)),(to_sfixed_a(-0.00017359404591843486)),(to_sfixed_a(5.842382233822718e-05)),(to_sfixed_a(-5.354394670575857e-05)),(to_sfixed_a(-8.868020813679323e-05)),(to_sfixed_a(-0.00022418401204049587)));

    constant weight_n0_33 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-3.320176256238483e-05)),(to_sfixed_a(0.00020626223704311997)),(to_sfixed_a(4.234688822180033e-05)),(to_sfixed_a(0.00011335566523484886)),(to_sfixed_a(-5.57231942366343e-05)),(to_sfixed_a(-4.090759466635063e-05)),(to_sfixed_a(8.460634853690863e-05)),(to_sfixed_a(4.4686689193440543e-07)),(to_sfixed_a(-2.171545202145353e-05)),(to_sfixed_a(-0.0001786990906111896)),(to_sfixed_a(1.9565579350455664e-05)),(to_sfixed_a(-0.00012467059423215687)),(to_sfixed_a(-0.00011221855675103143)),(to_sfixed_a(2.6124618557332724e-07)),(to_sfixed_a(3.298676892882213e-05)),(to_sfixed_a(0.0001224229927174747)),(to_sfixed_a(-2.665121246536728e-05)),(to_sfixed_a(4.369204179965891e-05)),(to_sfixed_a(-0.000148417180753313)),(to_sfixed_a(0.0003220373473595828)),(to_sfixed_a(4.833815182792023e-05)),(to_sfixed_a(0.00016950326971709728)),(to_sfixed_a(0.00015094055561348796)),(to_sfixed_a(-0.0002565581235103309)),(to_sfixed_a(-2.49940603680443e-06)),(to_sfixed_a(-5.191807940718718e-05)),(to_sfixed_a(-7.739226566627622e-05)),(to_sfixed_a(0.00011368651030352339)),(to_sfixed_a(-2.9579794500023127e-05)),(to_sfixed_a(0.00016957965272013098)),(to_sfixed_a(-0.00022938716574572027)),(to_sfixed_a(-0.00021302129607647657)),(to_sfixed_a(-0.00021364974963944405)),(to_sfixed_a(-3.92031179217156e-05)),(to_sfixed_a(0.00012335578503552824)),(to_sfixed_a(0.00013860661420039833)),(to_sfixed_a(0.00013309608038980514)),(to_sfixed_a(1.9272591089247726e-05)),(to_sfixed_a(0.00015503492613788694)),(to_sfixed_a(-0.0002048520400421694)),(to_sfixed_a(-0.0004416059819050133)),(to_sfixed_a(7.999538502190262e-05)),(to_sfixed_a(0.00015055878611747175)),(to_sfixed_a(0.00026532739866524935)),(to_sfixed_a(-8.183743193512782e-05)),(to_sfixed_a(-0.00014253452536650002)),(to_sfixed_a(-6.73527320032008e-05)),(to_sfixed_a(-0.00018883949087467045)),(to_sfixed_a(-0.0002248612727271393)),(to_sfixed_a(-9.51245783653576e-06)),(to_sfixed_a(-0.00021723246027249843)),(to_sfixed_a(5.733905709348619e-06)),(to_sfixed_a(-0.0004993689362891018)),(to_sfixed_a(0.0002483213902451098)),(to_sfixed_a(5.585920007433742e-05)),(to_sfixed_a(-0.00019399287702981383)),(to_sfixed_a(-6.294460774824984e-08)),(to_sfixed_a(9.984085045289248e-05)),(to_sfixed_a(-0.00019158096984028816)),(to_sfixed_a(-9.472779493080452e-05)),(to_sfixed_a(-5.911655898671597e-05)),(to_sfixed_a(-0.00024350930470973253)),(to_sfixed_a(-0.00012591000995598733)),(to_sfixed_a(-7.791679672664031e-05)),(to_sfixed_a(0.00013933645095676184)),(to_sfixed_a(-0.00034379313001409173)),(to_sfixed_a(-0.0001402619236614555)),(to_sfixed_a(-0.00014747884415555745)),(to_sfixed_a(0.00013884651707485318)),(to_sfixed_a(0.026482049375772476)),(to_sfixed_a(0.0001521910453448072)),(to_sfixed_a(0.00021567557996604592)),(to_sfixed_a(-7.73978463257663e-05)),(to_sfixed_a(0.00010119854414369911)),(to_sfixed_a(0.0001579806412337348)),(to_sfixed_a(-5.740662891184911e-05)),(to_sfixed_a(1.4844427823845763e-05)),(to_sfixed_a(-4.229397018207237e-05)),(to_sfixed_a(0.00014527815801557153)),(to_sfixed_a(0.00011702490883180872)),(to_sfixed_a(-0.0001625852019060403)),(to_sfixed_a(-8.787225851847325e-06)),(to_sfixed_a(-0.0001387900992995128)),(to_sfixed_a(3.136352097499184e-05)),(to_sfixed_a(-2.3981592676136643e-05)),(to_sfixed_a(-3.6937832192052156e-05)),(to_sfixed_a(-0.0001076961780199781)),(to_sfixed_a(0.00020851557201240212)),(to_sfixed_a(3.455948535702191e-05)),(to_sfixed_a(-0.0002814959443639964)),(to_sfixed_a(-6.965469219721854e-05)),(to_sfixed_a(0.00013080240751150995)),(to_sfixed_a(-0.03729808330535889)),(to_sfixed_a(-8.058820094447583e-05)),(to_sfixed_a(-0.042418815195560455)),(to_sfixed_a(0.043658655136823654)),(to_sfixed_a(-0.17509445548057556)),(to_sfixed_a(-0.10849184542894363)),(to_sfixed_a(-0.08575934916734695)),(to_sfixed_a(-0.0612458810210228)),(to_sfixed_a(0.003520858706906438)),(to_sfixed_a(-0.04366172477602959)),(to_sfixed_a(0.12814444303512573)),(to_sfixed_a(0.12806262075901031)),(to_sfixed_a(0.04195259511470795)),(to_sfixed_a(0.0853230357170105)),(to_sfixed_a(-7.935360372357536e-06)),(to_sfixed_a(0.00016695998783688992)),(to_sfixed_a(9.62526974035427e-05)),(to_sfixed_a(-0.00020338835020083934)),(to_sfixed_a(-0.00018868375627789646)),(to_sfixed_a(-0.00014389835996553302)),(to_sfixed_a(0.00011270945105934516)),(to_sfixed_a(-0.0001697393017821014)),(to_sfixed_a(7.419112807838246e-05)),(to_sfixed_a(-0.0001288921048399061)),(to_sfixed_a(-0.00012627204705495387)),(to_sfixed_a(0.00010245924931950867)),(to_sfixed_a(-0.0009678601054474711)),(to_sfixed_a(0.023656409233808517)),(to_sfixed_a(-0.0018601736519485712)),(to_sfixed_a(-0.04892222583293915)),(to_sfixed_a(-0.010515243746340275)),(to_sfixed_a(-0.024149825796484947)),(to_sfixed_a(-0.148515984416008)),(to_sfixed_a(-0.21767085790634155)),(to_sfixed_a(-0.0747813954949379)),(to_sfixed_a(-0.19696687161922455)),(to_sfixed_a(-0.08625050634145737)),(to_sfixed_a(-0.09030117094516754)),(to_sfixed_a(0.007269750349223614)),(to_sfixed_a(0.013132489286363125)),(to_sfixed_a(0.01892920583486557)),(to_sfixed_a(-0.02746289037168026)),(to_sfixed_a(-0.0033369315788149834)),(to_sfixed_a(-0.00010107544221682474)),(to_sfixed_a(-0.0017777306493371725)),(to_sfixed_a(-0.00022518700279761106)),(to_sfixed_a(2.4218488761107437e-05)),(to_sfixed_a(0.00012453646922949702)),(to_sfixed_a(-7.293685484910384e-05)),(to_sfixed_a(0.00010875576845137402)),(to_sfixed_a(-0.0001292639208259061)),(to_sfixed_a(-5.822159891977208e-06)),(to_sfixed_a(-0.0013064314844086766)),(to_sfixed_a(0.03115016035735607)),(to_sfixed_a(-0.006408087443560362)),(to_sfixed_a(0.12405948340892792)),(to_sfixed_a(0.04668688401579857)),(to_sfixed_a(-0.031677860766649246)),(to_sfixed_a(-0.12514673173427582)),(to_sfixed_a(-0.010977436788380146)),(to_sfixed_a(-0.05511119216680527)),(to_sfixed_a(0.012925227172672749)),(to_sfixed_a(-0.02663337253034115)),(to_sfixed_a(0.06588665395975113)),(to_sfixed_a(0.056876957416534424)),(to_sfixed_a(0.1652776449918747)),(to_sfixed_a(0.0070565794594585896)),(to_sfixed_a(-0.08315035700798035)),(to_sfixed_a(-0.023549100384116173)),(to_sfixed_a(0.02266114391386509)),(to_sfixed_a(-0.0004557082720566541)),(to_sfixed_a(0.05347435548901558)),(to_sfixed_a(-0.0009752217447385192)),(to_sfixed_a(-0.0004001148627139628)),(to_sfixed_a(4.40935036749579e-05)),(to_sfixed_a(0.0002793400199152529)),(to_sfixed_a(-0.0001430659758625552)),(to_sfixed_a(9.781355038285255e-05)),(to_sfixed_a(6.997327727731317e-05)),(to_sfixed_a(-6.355749064823613e-05)),(to_sfixed_a(-0.00033386365976184607)),(to_sfixed_a(0.03284706175327301)),(to_sfixed_a(-0.06498569250106812)),(to_sfixed_a(0.08814915269613266)),(to_sfixed_a(-0.07543295621871948)),(to_sfixed_a(0.06942091882228851)),(to_sfixed_a(0.1453583538532257)),(to_sfixed_a(0.15117715299129486)),(to_sfixed_a(0.04840913042426109)),(to_sfixed_a(-0.1123947948217392)),(to_sfixed_a(-0.13328982889652252)),(to_sfixed_a(0.1502576321363449)),(to_sfixed_a(0.18500544130802155)),(to_sfixed_a(0.01893104612827301)),(to_sfixed_a(-0.12240415811538696)),(to_sfixed_a(-0.004127637483179569)),(to_sfixed_a(0.08119688928127289)),(to_sfixed_a(-0.08628514409065247)),(to_sfixed_a(-0.02583800069987774)),(to_sfixed_a(0.10305601358413696)),(to_sfixed_a(-0.0012522978940978646)),(to_sfixed_a(-0.0017722531920298934)),(to_sfixed_a(-0.003051512874662876)),(to_sfixed_a(-3.399734850972891e-05)),(to_sfixed_a(7.021654164418578e-05)),(to_sfixed_a(-0.00024927029153332114)),(to_sfixed_a(6.909895455464721e-05)),(to_sfixed_a(0.00013673448120243847)),(to_sfixed_a(-2.0376544853206724e-05)),(to_sfixed_a(0.02480965666472912)),(to_sfixed_a(-0.05735347792506218)),(to_sfixed_a(0.024489259347319603)),(to_sfixed_a(-0.005327625200152397)),(to_sfixed_a(0.0981426015496254)),(to_sfixed_a(0.0112910782918334)),(to_sfixed_a(0.05684739351272583)),(to_sfixed_a(-0.04123882204294205)),(to_sfixed_a(-0.31519803404808044)),(to_sfixed_a(0.1339910328388214)),(to_sfixed_a(0.2609637677669525)),(to_sfixed_a(0.023560943081974983)),(to_sfixed_a(-0.020847579464316368)),(to_sfixed_a(-0.10062995553016663)),(to_sfixed_a(-0.041323695331811905)),(to_sfixed_a(-0.17708277702331543)),(to_sfixed_a(0.023600321263074875)),(to_sfixed_a(-0.12286150455474854)),(to_sfixed_a(0.026132341474294662)),(to_sfixed_a(0.012499538250267506)),(to_sfixed_a(0.004442824516445398)),(to_sfixed_a(0.00011330875713611022)),(to_sfixed_a(-4.963629908161238e-05)),(to_sfixed_a(0.0001922155061038211)),(to_sfixed_a(2.3886104827397503e-05)),(to_sfixed_a(-0.00033258143230341375)),(to_sfixed_a(-7.276071119122207e-05)),(to_sfixed_a(-0.027988966554403305)),(to_sfixed_a(0.05307381600141525)),(to_sfixed_a(0.012592049315571785)),(to_sfixed_a(0.1818832904100418)),(to_sfixed_a(-0.18543991446495056)),(to_sfixed_a(0.040073197335004807)),(to_sfixed_a(0.07496237754821777)),(to_sfixed_a(-0.046972908079624176)),(to_sfixed_a(-0.16073206067085266)),(to_sfixed_a(0.18941083550453186)),(to_sfixed_a(0.26217204332351685)),(to_sfixed_a(0.15773652493953705)),(to_sfixed_a(-0.0786285474896431)),(to_sfixed_a(-0.07562515139579773)),(to_sfixed_a(-0.16573679447174072)),(to_sfixed_a(-0.31270936131477356)),(to_sfixed_a(-0.11448230594396591)),(to_sfixed_a(-0.05327434465289116)),(to_sfixed_a(-0.04941850155591965)),(to_sfixed_a(-0.010676269419491291)),(to_sfixed_a(-0.05366731807589531)),(to_sfixed_a(0.07669105380773544)),(to_sfixed_a(0.00014910339086782187)),(to_sfixed_a(3.733090125024319e-05)),(to_sfixed_a(-8.189355139620602e-05)),(to_sfixed_a(-0.0001521117374068126)),(to_sfixed_a(-0.00019833586702588946)),(to_sfixed_a(-5.9060927014797926e-05)),(to_sfixed_a(-0.00023794254229869694)),(to_sfixed_a(-0.04561794921755791)),(to_sfixed_a(-0.013312757015228271)),(to_sfixed_a(0.0013546458212658763)),(to_sfixed_a(0.025566881522536278)),(to_sfixed_a(-0.027034824714064598)),(to_sfixed_a(-0.20454953610897064)),(to_sfixed_a(0.0994325801730156)),(to_sfixed_a(-0.03415681794285774)),(to_sfixed_a(0.10717999935150146)),(to_sfixed_a(0.1984003782272339)),(to_sfixed_a(0.23890119791030884)),(to_sfixed_a(0.027936050668358803)),(to_sfixed_a(-0.010230564512312412)),(to_sfixed_a(-0.2662663161754608)),(to_sfixed_a(0.13436102867126465)),(to_sfixed_a(-0.09972500056028366)),(to_sfixed_a(-0.07852798700332642)),(to_sfixed_a(0.09753797948360443)),(to_sfixed_a(0.10603451728820801)),(to_sfixed_a(0.34116846323013306)),(to_sfixed_a(2.2492482457892038e-05)),(to_sfixed_a(0.00047078888746909797)),(to_sfixed_a(-4.5023680286249146e-05)),(to_sfixed_a(-0.0001220154226757586)),(to_sfixed_a(-0.00012106877693440765)),(to_sfixed_a(-0.0001745067856973037)),(to_sfixed_a(-0.0001637902169022709)),(to_sfixed_a(0.002387670800089836)),(to_sfixed_a(0.011555960401892662)),(to_sfixed_a(-0.17221283912658691)),(to_sfixed_a(-0.0007138987421058118)),(to_sfixed_a(-0.10700614750385284)),(to_sfixed_a(-0.22380448877811432)),(to_sfixed_a(0.1862535923719406)),(to_sfixed_a(0.3492991626262665)),(to_sfixed_a(-0.03691992908716202)),(to_sfixed_a(0.045483339577913284)),(to_sfixed_a(0.22382839024066925)),(to_sfixed_a(-0.15818020701408386)),(to_sfixed_a(-0.24283716082572937)),(to_sfixed_a(0.04930886626243591)),(to_sfixed_a(0.25736817717552185)),(to_sfixed_a(0.1228606179356575)),(to_sfixed_a(-0.08586964011192322)),(to_sfixed_a(0.0194181390106678)),(to_sfixed_a(-0.10413076728582382)),(to_sfixed_a(-0.20854437351226807)),(to_sfixed_a(0.08010285347700119)),(to_sfixed_a(0.0060285525396466255)),(to_sfixed_a(6.741341348970309e-05)),(to_sfixed_a(7.782904867781326e-05)),(to_sfixed_a(0.00011684927449095994)),(to_sfixed_a(-0.0001721802109386772)),(to_sfixed_a(-1.2861794857599307e-05)),(to_sfixed_a(-0.011010128073394299)),(to_sfixed_a(-0.019386162981390953)),(to_sfixed_a(-0.08083939552307129)),(to_sfixed_a(-0.048588115721940994)),(to_sfixed_a(0.21622276306152344)),(to_sfixed_a(0.12414642423391342)),(to_sfixed_a(-0.02656400017440319)),(to_sfixed_a(-0.006649858318269253)),(to_sfixed_a(0.2895413935184479)),(to_sfixed_a(0.21494485437870026)),(to_sfixed_a(-0.2556138038635254)),(to_sfixed_a(-0.3270900249481201)),(to_sfixed_a(0.0019807443022727966)),(to_sfixed_a(0.2238772213459015)),(to_sfixed_a(0.15714780986309052)),(to_sfixed_a(0.19351288676261902)),(to_sfixed_a(0.14574748277664185)),(to_sfixed_a(-0.0011080449912697077)),(to_sfixed_a(-2.642559411469847e-05)),(to_sfixed_a(0.014637188985943794)),(to_sfixed_a(-0.019423052668571472)),(to_sfixed_a(-0.07552646845579147)),(to_sfixed_a(-2.7155578209203668e-05)),(to_sfixed_a(-7.047737744869664e-05)),(to_sfixed_a(0.00014731950068380684)),(to_sfixed_a(0.00020268683147151023)),(to_sfixed_a(2.171758569602389e-05)),(to_sfixed_a(0.0003104649658780545)),(to_sfixed_a(-0.00023587190662510693)),(to_sfixed_a(0.06605423986911774)),(to_sfixed_a(-0.11139979213476181)),(to_sfixed_a(-0.10396900773048401)),(to_sfixed_a(0.11163749545812607)),(to_sfixed_a(0.043507881462574005)),(to_sfixed_a(-0.12591080367565155)),(to_sfixed_a(-0.1558179408311844)),(to_sfixed_a(0.15972213447093964)),(to_sfixed_a(0.148818239569664)),(to_sfixed_a(-0.3841722309589386)),(to_sfixed_a(-0.16597966849803925)),(to_sfixed_a(-0.14250479638576508)),(to_sfixed_a(0.34301725029945374)),(to_sfixed_a(-0.3781462609767914)),(to_sfixed_a(-0.03092154674232006)),(to_sfixed_a(-0.22447195649147034)),(to_sfixed_a(0.18252599239349365)),(to_sfixed_a(0.12039253860712051)),(to_sfixed_a(0.16215632855892181)),(to_sfixed_a(0.14946894347667694)),(to_sfixed_a(-0.14222843945026398)),(to_sfixed_a(-0.0002088916371576488)),(to_sfixed_a(-5.22498412465211e-05)),(to_sfixed_a(7.260566235345323e-06)),(to_sfixed_a(4.8351601435570046e-05)),(to_sfixed_a(0.00018346557044424117)),(to_sfixed_a(-2.9492723115254194e-05)),(to_sfixed_a(-0.00013387942453846335)),(to_sfixed_a(0.06968086957931519)),(to_sfixed_a(-0.12933409214019775)),(to_sfixed_a(-0.06134568899869919)),(to_sfixed_a(-0.3177449703216553)),(to_sfixed_a(-0.1785557121038437)),(to_sfixed_a(-0.12848792970180511)),(to_sfixed_a(-0.06336959451436996)),(to_sfixed_a(0.25342532992362976)),(to_sfixed_a(0.09545409679412842)),(to_sfixed_a(-0.3361538052558899)),(to_sfixed_a(0.2646827697753906)),(to_sfixed_a(0.3179202675819397)),(to_sfixed_a(-0.05070051923394203)),(to_sfixed_a(0.037243179976940155)),(to_sfixed_a(-0.02366812527179718)),(to_sfixed_a(-0.20101939141750336)),(to_sfixed_a(-0.004886047914624214)),(to_sfixed_a(0.03312086686491966)),(to_sfixed_a(-0.01948951743543148)),(to_sfixed_a(-0.30247822403907776)),(to_sfixed_a(-0.04626155272126198)),(to_sfixed_a(0.0004079253994859755)),(to_sfixed_a(-0.00014365864626597613)),(to_sfixed_a(0.0003240200167056173)),(to_sfixed_a(0.0001764375192578882)),(to_sfixed_a(-0.00017726424266584218)),(to_sfixed_a(9.643840894568712e-05)),(to_sfixed_a(-8.051403710851446e-05)),(to_sfixed_a(0.00017029624723363668)),(to_sfixed_a(0.006623373366892338)),(to_sfixed_a(0.12426529824733734)),(to_sfixed_a(-0.12021064013242722)),(to_sfixed_a(0.038942787796258926)),(to_sfixed_a(-0.22172223031520844)),(to_sfixed_a(0.11430633068084717)),(to_sfixed_a(0.17691200971603394)),(to_sfixed_a(0.18004237115383148)),(to_sfixed_a(0.20492297410964966)),(to_sfixed_a(-0.08079227805137634)),(to_sfixed_a(-0.1082909032702446)),(to_sfixed_a(-0.06921429187059402)),(to_sfixed_a(0.006335573270916939)),(to_sfixed_a(-0.06683731824159622)),(to_sfixed_a(-0.00915964413434267)),(to_sfixed_a(0.08168469369411469)),(to_sfixed_a(-0.0023592032957822084)),(to_sfixed_a(-0.07154854387044907)),(to_sfixed_a(-0.10290678590536118)),(to_sfixed_a(-0.12979988753795624)),(to_sfixed_a(0.00042272169957868755)),(to_sfixed_a(0.00031824232428334653)),(to_sfixed_a(0.0001696034159976989)),(to_sfixed_a(-4.724943210021593e-05)),(to_sfixed_a(-0.00019485711527522653)),(to_sfixed_a(0.0002063749561784789)),(to_sfixed_a(9.830180351855233e-05)),(to_sfixed_a(-0.09236299246549606)),(to_sfixed_a(0.2964903712272644)),(to_sfixed_a(0.02013995312154293)),(to_sfixed_a(0.3089197278022766)),(to_sfixed_a(0.06523758172988892)),(to_sfixed_a(0.14575642347335815)),(to_sfixed_a(0.02320033498108387)),(to_sfixed_a(-0.039542440325021744)),(to_sfixed_a(-0.24082982540130615)),(to_sfixed_a(-0.38018831610679626)),(to_sfixed_a(-0.009570026770234108)),(to_sfixed_a(-0.15566423535346985)),(to_sfixed_a(-0.17325903475284576)),(to_sfixed_a(0.2066013664007187)),(to_sfixed_a(-0.07020985335111618)),(to_sfixed_a(0.07087689638137817)),(to_sfixed_a(-0.053478579968214035)),(to_sfixed_a(-0.05026025325059891)),(to_sfixed_a(-0.06438365578651428)),(to_sfixed_a(-0.08408305048942566)),(to_sfixed_a(-0.09660346806049347)),(to_sfixed_a(0.0004158385854680091)),(to_sfixed_a(0.00016247591702267528)),(to_sfixed_a(-7.065842510201037e-05)),(to_sfixed_a(2.924594264186453e-05)),(to_sfixed_a(0.00022079143673181534)),(to_sfixed_a(-0.00015372819325421005)),(to_sfixed_a(-0.0008756523602642119)),(to_sfixed_a(-0.09506651014089584)),(to_sfixed_a(-0.22049222886562347)),(to_sfixed_a(-0.3385869860649109)),(to_sfixed_a(-0.03828989714384079)),(to_sfixed_a(-0.08501880615949631)),(to_sfixed_a(0.111969493329525)),(to_sfixed_a(-0.08181123435497284)),(to_sfixed_a(0.15883402526378632)),(to_sfixed_a(0.058025062084198)),(to_sfixed_a(0.27289900183677673)),(to_sfixed_a(0.016604473814368248)),(to_sfixed_a(-0.1312999725341797)),(to_sfixed_a(0.06068481504917145)),(to_sfixed_a(-0.0006359754479490221)),(to_sfixed_a(0.062062498182058334)),(to_sfixed_a(0.08279695361852646)),(to_sfixed_a(0.04059295728802681)),(to_sfixed_a(-0.2336675524711609)),(to_sfixed_a(-0.06075901538133621)),(to_sfixed_a(0.05749012529850006)),(to_sfixed_a(-0.06863896548748016)),(to_sfixed_a(-0.0015523299807682633)),(to_sfixed_a(-0.00015915239055175334)),(to_sfixed_a(-2.5703784558572806e-06)),(to_sfixed_a(5.365890683606267e-05)),(to_sfixed_a(0.00016420324391219765)),(to_sfixed_a(-0.0011363350786268711)),(to_sfixed_a(-0.000859367020893842)),(to_sfixed_a(-0.0097538772970438)),(to_sfixed_a(-0.13590431213378906)),(to_sfixed_a(0.10108472406864166)),(to_sfixed_a(-0.13752101361751556)),(to_sfixed_a(0.07570706307888031)),(to_sfixed_a(0.009914057329297066)),(to_sfixed_a(-0.0017948949243873358)),(to_sfixed_a(0.006326089613139629)),(to_sfixed_a(0.1644914746284485)),(to_sfixed_a(0.0725165605545044)),(to_sfixed_a(0.15842007100582123)),(to_sfixed_a(-0.0251007117331028)),(to_sfixed_a(-0.10393897444009781)),(to_sfixed_a(0.015864094719290733)),(to_sfixed_a(0.2548043727874756)),(to_sfixed_a(0.321184903383255)),(to_sfixed_a(0.11675352603197098)),(to_sfixed_a(0.07088932394981384)),(to_sfixed_a(-0.01317583303898573)),(to_sfixed_a(-0.007591592613607645)),(to_sfixed_a(-6.85801642248407e-05)),(to_sfixed_a(3.1907471566228196e-05)),(to_sfixed_a(9.395951929036528e-05)),(to_sfixed_a(-0.00024803754058666527)),(to_sfixed_a(5.0536174967419356e-05)),(to_sfixed_a(-8.774175512371585e-05)),(to_sfixed_a(-0.00010524096433073282)),(to_sfixed_a(0.03561824560165405)),(to_sfixed_a(-0.04417188838124275)),(to_sfixed_a(0.15044988691806793)),(to_sfixed_a(0.018239231780171394)),(to_sfixed_a(0.1939723640680313)),(to_sfixed_a(0.034076083451509476)),(to_sfixed_a(-0.08106677234172821)),(to_sfixed_a(0.01417980995029211)),(to_sfixed_a(-0.19136296212673187)),(to_sfixed_a(0.13015031814575195)),(to_sfixed_a(0.1855199933052063)),(to_sfixed_a(0.02365162782371044)),(to_sfixed_a(-0.10044983774423599)),(to_sfixed_a(0.09150830656290054)),(to_sfixed_a(0.03159298002719879)),(to_sfixed_a(0.009994210675358772)),(to_sfixed_a(0.20546197891235352)),(to_sfixed_a(-0.015345829539000988)),(to_sfixed_a(-0.30701300501823425)),(to_sfixed_a(-0.06858176738023758)),(to_sfixed_a(-0.04582514986395836)),(to_sfixed_a(0.014645291492342949)),(to_sfixed_a(0.000228230856009759)),(to_sfixed_a(-0.00016778135614003986)),(to_sfixed_a(0.00011119562259409577)),(to_sfixed_a(-0.00010396140714874491)),(to_sfixed_a(3.6566001654136926e-05)),(to_sfixed_a(-0.00012282833631616086)),(to_sfixed_a(-0.10759031772613525)),(to_sfixed_a(0.0012672959128394723)),(to_sfixed_a(-0.07046038657426834)),(to_sfixed_a(0.08421697467565536)),(to_sfixed_a(0.0007777499267831445)),(to_sfixed_a(0.18979205191135406)),(to_sfixed_a(-0.06731338053941727)),(to_sfixed_a(0.4008682072162628)),(to_sfixed_a(-0.029336797073483467)),(to_sfixed_a(0.03531724959611893)),(to_sfixed_a(0.05364220216870308)),(to_sfixed_a(-0.1535843461751938)),(to_sfixed_a(0.011614824645221233)),(to_sfixed_a(-0.020520461723208427)),(to_sfixed_a(0.1425265520811081)),(to_sfixed_a(0.1786748617887497)),(to_sfixed_a(0.06447850912809372)),(to_sfixed_a(-0.09345323592424393)),(to_sfixed_a(0.020658783614635468)),(to_sfixed_a(-0.01703077368438244)),(to_sfixed_a(-0.010718753561377525)),(to_sfixed_a(8.765058737481013e-05)),(to_sfixed_a(3.386045864317566e-05)),(to_sfixed_a(8.864166011335328e-05)),(to_sfixed_a(0.00026925330166704953)),(to_sfixed_a(0.0002813022874761373)),(to_sfixed_a(-0.0001128909716499038)),(to_sfixed_a(6.159289478091523e-05)),(to_sfixed_a(0.0002489185717422515)),(to_sfixed_a(0.014178465120494366)),(to_sfixed_a(0.10506469756364822)),(to_sfixed_a(-0.034802984446287155)),(to_sfixed_a(0.02092389389872551)),(to_sfixed_a(-0.24850071966648102)),(to_sfixed_a(0.07298602908849716)),(to_sfixed_a(0.07798899710178375)),(to_sfixed_a(-0.10571154952049255)),(to_sfixed_a(-0.10332021117210388)),(to_sfixed_a(-0.11649785190820694)),(to_sfixed_a(-0.09085571020841599)),(to_sfixed_a(-0.21603234112262726)),(to_sfixed_a(-0.15666750073432922)),(to_sfixed_a(0.10154970735311508)),(to_sfixed_a(-0.1887323558330536)),(to_sfixed_a(0.04566310718655586)),(to_sfixed_a(-0.03105500526726246)),(to_sfixed_a(-0.17459671199321747)),(to_sfixed_a(-0.007005732506513596)),(to_sfixed_a(-0.05667901411652565)),(to_sfixed_a(-0.022594798356294632)),(to_sfixed_a(-8.333107689395547e-05)),(to_sfixed_a(1.309394974668976e-05)),(to_sfixed_a(0.00023335246078204364)),(to_sfixed_a(-0.00016972121375147253)),(to_sfixed_a(1.1453144907136448e-05)),(to_sfixed_a(-8.179802534868941e-05)),(to_sfixed_a(-1.8620681657921523e-05)),(to_sfixed_a(-0.004402644000947475)),(to_sfixed_a(2.9799728508805856e-05)),(to_sfixed_a(-0.062350593507289886)),(to_sfixed_a(-0.10108086466789246)),(to_sfixed_a(-0.15954959392547607)),(to_sfixed_a(-0.26333433389663696)),(to_sfixed_a(0.015075293369591236)),(to_sfixed_a(-0.27796807885169983)),(to_sfixed_a(-0.07306621223688126)),(to_sfixed_a(-0.030909547582268715)),(to_sfixed_a(0.13967782258987427)),(to_sfixed_a(-0.07397949695587158)),(to_sfixed_a(-0.10646868497133255)),(to_sfixed_a(-0.12980717420578003)),(to_sfixed_a(0.05987562611699104)),(to_sfixed_a(0.06833244115114212)),(to_sfixed_a(0.2693159282207489)),(to_sfixed_a(0.06857199966907501)),(to_sfixed_a(-0.004988408647477627)),(to_sfixed_a(8.116262324620038e-05)),(to_sfixed_a(0.0012435032986104488)),(to_sfixed_a(0.00023155026428867131)),(to_sfixed_a(0.00016314847744069993)),(to_sfixed_a(-0.00024946441408246756)),(to_sfixed_a(-0.00011559456470422447)),(to_sfixed_a(-4.4085343688493595e-05)),(to_sfixed_a(-0.0002512720529921353)),(to_sfixed_a(0.00022574805188924074)),(to_sfixed_a(0.00026802808861248195)),(to_sfixed_a(-0.059310995042324066)),(to_sfixed_a(-0.18980740010738373)),(to_sfixed_a(-0.10021552443504333)),(to_sfixed_a(0.0844636932015419)),(to_sfixed_a(-0.045756421983242035)),(to_sfixed_a(-0.2853037118911743)),(to_sfixed_a(-0.24424996972084045)),(to_sfixed_a(-0.09981080144643784)),(to_sfixed_a(-0.0179641954600811)),(to_sfixed_a(0.06836207956075668)),(to_sfixed_a(0.023264681920409203)),(to_sfixed_a(0.027682499960064888)),(to_sfixed_a(0.10708136111497879)),(to_sfixed_a(-0.036742307245731354)),(to_sfixed_a(-0.056061942130327225)),(to_sfixed_a(0.024906722828745842)),(to_sfixed_a(0.007925606332719326)),(to_sfixed_a(-0.006582255940884352)),(to_sfixed_a(0.0057002645917236805)),(to_sfixed_a(0.0001049917918862775)),(to_sfixed_a(-9.90582429949427e-06)),(to_sfixed_a(5.46347328054253e-05)),(to_sfixed_a(-4.9192633014172316e-05)),(to_sfixed_a(-0.00011890979658346623)),(to_sfixed_a(-0.0001558194198878482)),(to_sfixed_a(-0.00023888178111519665)),(to_sfixed_a(2.7352863980922848e-05)),(to_sfixed_a(0.00010981447121594101)),(to_sfixed_a(0.019739432260394096)),(to_sfixed_a(0.1063503548502922)),(to_sfixed_a(-0.024134932085871696)),(to_sfixed_a(0.15803810954093933)),(to_sfixed_a(0.009125441312789917)),(to_sfixed_a(-0.010904519818723202)),(to_sfixed_a(-0.09678726643323898)),(to_sfixed_a(0.09757666289806366)),(to_sfixed_a(0.02107452228665352)),(to_sfixed_a(0.20634374022483826)),(to_sfixed_a(0.08074028044939041)),(to_sfixed_a(-0.003422666108235717)),(to_sfixed_a(0.013860217295587063)),(to_sfixed_a(-0.07782334834337234)),(to_sfixed_a(-0.17962203919887543)),(to_sfixed_a(0.07375858724117279)),(to_sfixed_a(-0.003953675273805857)),(to_sfixed_a(0.005144242197275162)),(to_sfixed_a(-0.008168576285243034)),(to_sfixed_a(-8.065568545134738e-05)),(to_sfixed_a(5.098223118693568e-05)),(to_sfixed_a(4.644127329811454e-05)),(to_sfixed_a(1.4527739949699026e-05)),(to_sfixed_a(-0.0003333195927552879)),(to_sfixed_a(1.7614676835364662e-05)),(to_sfixed_a(7.309197098948061e-05)),(to_sfixed_a(0.00011654686386464164)),(to_sfixed_a(0.010407908819615841)),(to_sfixed_a(0.03265632688999176)),(to_sfixed_a(0.04249238595366478)),(to_sfixed_a(-0.028032127767801285)),(to_sfixed_a(0.0008819757495075464)),(to_sfixed_a(-0.1974126249551773)),(to_sfixed_a(-0.08812791109085083)),(to_sfixed_a(0.0038263017777353525)),(to_sfixed_a(-0.010914653539657593)),(to_sfixed_a(0.012163319624960423)),(to_sfixed_a(-0.05324752256274223)),(to_sfixed_a(-0.11824353784322739)),(to_sfixed_a(-0.12424761056900024)),(to_sfixed_a(-0.15030108392238617)),(to_sfixed_a(-0.05201084911823273)),(to_sfixed_a(-0.06427236646413803)),(to_sfixed_a(-0.003837121417745948)),(to_sfixed_a(-0.029589267447590828)),(to_sfixed_a(-0.009873666800558567)),(to_sfixed_a(-0.0049257124774158)),(to_sfixed_a(0.000146375474287197)),(to_sfixed_a(2.733863948378712e-05)),(to_sfixed_a(3.4790537029039115e-05)),(to_sfixed_a(-2.0283805497456342e-05)),(to_sfixed_a(0.00020074886560905725)),(to_sfixed_a(-2.754856541287154e-05)),(to_sfixed_a(-0.00020948951714672148)),(to_sfixed_a(9.161651541944593e-05)),(to_sfixed_a(4.0935385186458007e-05)),(to_sfixed_a(-0.08344212919473648)),(to_sfixed_a(0.02592557854950428)),(to_sfixed_a(0.04008553549647331)),(to_sfixed_a(0.013142501004040241)),(to_sfixed_a(0.18382740020751953)),(to_sfixed_a(0.0629594698548317)),(to_sfixed_a(-0.08116243034601212)),(to_sfixed_a(0.14909346401691437)),(to_sfixed_a(-0.04755023121833801)),(to_sfixed_a(0.04036759212613106)),(to_sfixed_a(0.045316632837057114)),(to_sfixed_a(-0.25341325998306274)),(to_sfixed_a(-0.008395558223128319)),(to_sfixed_a(-0.008330662734806538)),(to_sfixed_a(-0.17313505709171295)),(to_sfixed_a(-0.18270717561244965)),(to_sfixed_a(-0.00041163747664541006)),(to_sfixed_a(-0.0013655382208526134)),(to_sfixed_a(-0.0018307806458324194)),(to_sfixed_a(2.4216531528509222e-05)),(to_sfixed_a(-5.4036023357184604e-05)),(to_sfixed_a(-3.4368746128166094e-05)),(to_sfixed_a(-6.74107504892163e-05)),(to_sfixed_a(0.00010250561899738386)),(to_sfixed_a(-0.00023269763914868236)),(to_sfixed_a(4.313584940973669e-05)),(to_sfixed_a(-0.0002531373465899378)),(to_sfixed_a(-3.901176751242019e-05)),(to_sfixed_a(0.0009987056255340576)),(to_sfixed_a(0.001038354472257197)),(to_sfixed_a(-7.529029244324192e-05)),(to_sfixed_a(-3.9990532968658954e-05)),(to_sfixed_a(0.0001885115634649992)),(to_sfixed_a(-0.17014780640602112)),(to_sfixed_a(-0.0039326841942965984)),(to_sfixed_a(-0.0011852941242977977)),(to_sfixed_a(-0.12424057722091675)),(to_sfixed_a(0.004544905852526426)),(to_sfixed_a(0.0029495658818632364)),(to_sfixed_a(0.001900032046250999)),(to_sfixed_a(-0.1324819177389145)),(to_sfixed_a(-0.17415444552898407)),(to_sfixed_a(0.0028495744336396456)),(to_sfixed_a(0.000435639958595857)),(to_sfixed_a(-5.153358506504446e-05)),(to_sfixed_a(-0.00021071876108180732)),(to_sfixed_a(-0.00016026235243771225)),(to_sfixed_a(-0.00015334298950619996)),(to_sfixed_a(0.00024385142023675144)),(to_sfixed_a(-0.00018194981385022402)),(to_sfixed_a(2.9861459552193992e-05)),(to_sfixed_a(-0.00016907521057873964)),(to_sfixed_a(-0.00011176317639183253)),(to_sfixed_a(0.00012042924208799377)),(to_sfixed_a(0.0001237071555806324)),(to_sfixed_a(5.5098600569181144e-05)),(to_sfixed_a(0.00014837371418252587)),(to_sfixed_a(-0.0001461473439121619)),(to_sfixed_a(-0.00014543446013703942)),(to_sfixed_a(-0.00013237792882137)),(to_sfixed_a(-0.00022756152611691505)),(to_sfixed_a(0.00016816053539514542)),(to_sfixed_a(5.950056220171973e-05)),(to_sfixed_a(-0.000107483436295297)),(to_sfixed_a(5.231095929048024e-05)),(to_sfixed_a(8.947041351348162e-05)),(to_sfixed_a(-5.420112574938685e-05)),(to_sfixed_a(0.00029895250918343663)),(to_sfixed_a(-6.584506627405062e-05)),(to_sfixed_a(0.00021054985700175166)),(to_sfixed_a(9.309273445978761e-05)),(to_sfixed_a(-0.00013889017282053828)),(to_sfixed_a(-0.00020181034051347524)),(to_sfixed_a(9.320170647697523e-05)),(to_sfixed_a(-7.62125346227549e-05)),(to_sfixed_a(5.704915747628547e-05)),(to_sfixed_a(-0.0001961267553269863)),(to_sfixed_a(-9.207769835484214e-06)),(to_sfixed_a(-3.5624525480670854e-05)));

    constant weight_n0_34 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(-8.82572348928079e-05)),(to_sfixed_a(1.8203309082309715e-05)),(to_sfixed_a(0.0002462588017806411)),(to_sfixed_a(-1.1754000297514722e-05)),(to_sfixed_a(8.316994353663176e-05)),(to_sfixed_a(-9.445509203942493e-05)),(to_sfixed_a(-3.769485829252517e-06)),(to_sfixed_a(0.00038743377081118524)),(to_sfixed_a(-0.00023959418467711657)),(to_sfixed_a(-0.00013469092664308846)),(to_sfixed_a(-0.0001697690604487434)),(to_sfixed_a(8.540867565898225e-05)),(to_sfixed_a(0.000144315417855978)),(to_sfixed_a(-6.180385389598086e-05)),(to_sfixed_a(-6.503280746983364e-05)),(to_sfixed_a(0.00026734487619251013)),(to_sfixed_a(-7.001664926065132e-05)),(to_sfixed_a(0.0001008655090117827)),(to_sfixed_a(-0.00010283359733875841)),(to_sfixed_a(-9.96431554085575e-05)),(to_sfixed_a(-0.0001861931523308158)),(to_sfixed_a(0.00024923047749325633)),(to_sfixed_a(0.00025221583200618625)),(to_sfixed_a(-0.00014388297859113663)),(to_sfixed_a(0.0002464482095092535)),(to_sfixed_a(-3.769869726966135e-05)),(to_sfixed_a(-2.1318390281521715e-05)),(to_sfixed_a(8.650815289001912e-05)),(to_sfixed_a(5.004610284231603e-05)),(to_sfixed_a(-3.497244688333012e-05)),(to_sfixed_a(1.4954932339605875e-05)),(to_sfixed_a(-5.917781527386978e-05)),(to_sfixed_a(0.00016155806952156126)),(to_sfixed_a(5.382459676184226e-06)),(to_sfixed_a(-3.446214032010175e-05)),(to_sfixed_a(-5.711643825634383e-05)),(to_sfixed_a(-8.19609995232895e-05)),(to_sfixed_a(-2.6341102056903765e-05)),(to_sfixed_a(4.6390516217797995e-05)),(to_sfixed_a(-0.0002171070664189756)),(to_sfixed_a(5.716604573535733e-05)),(to_sfixed_a(0.00027158530429005623)),(to_sfixed_a(-0.0001954545296030119)),(to_sfixed_a(0.0001288895873585716)),(to_sfixed_a(6.882230809424073e-05)),(to_sfixed_a(5.5945998610695824e-05)),(to_sfixed_a(0.0001777630386641249)),(to_sfixed_a(-0.0001997380459215492)),(to_sfixed_a(-3.5046945413341746e-05)),(to_sfixed_a(9.652676089899614e-05)),(to_sfixed_a(3.6006411392008886e-05)),(to_sfixed_a(4.1716093619470485e-06)),(to_sfixed_a(0.00017442538228351623)),(to_sfixed_a(-8.174126560334116e-05)),(to_sfixed_a(0.00012844866432715207)),(to_sfixed_a(3.114791979896836e-05)),(to_sfixed_a(0.00012637866893783212)),(to_sfixed_a(5.7507197197992355e-05)),(to_sfixed_a(0.00018104798800777644)),(to_sfixed_a(0.00020627093908842653)),(to_sfixed_a(5.413536564446986e-05)),(to_sfixed_a(-3.3932345104403794e-05)),(to_sfixed_a(0.00015978579176589847)),(to_sfixed_a(-2.9954218916827813e-05)),(to_sfixed_a(4.057597470819019e-05)),(to_sfixed_a(-2.7761439923779108e-05)),(to_sfixed_a(0.000241165587794967)),(to_sfixed_a(-0.00013025416410528123)),(to_sfixed_a(9.302333637606353e-05)),(to_sfixed_a(-0.02873297780752182)),(to_sfixed_a(6.136661249911413e-05)),(to_sfixed_a(0.00011872733739437535)),(to_sfixed_a(9.266405868402217e-06)),(to_sfixed_a(0.00012858725676778704)),(to_sfixed_a(6.270670564845204e-05)),(to_sfixed_a(8.73270837473683e-05)),(to_sfixed_a(0.00018283443932887167)),(to_sfixed_a(7.14191555744037e-05)),(to_sfixed_a(-4.957253622706048e-05)),(to_sfixed_a(0.00048513736692257226)),(to_sfixed_a(0.00018446701869834214)),(to_sfixed_a(0.00015562820772174746)),(to_sfixed_a(4.875044396612793e-05)),(to_sfixed_a(-5.683152994606644e-05)),(to_sfixed_a(-1.1652413377305493e-05)),(to_sfixed_a(9.983817290049046e-05)),(to_sfixed_a(-4.4779844756703824e-05)),(to_sfixed_a(-0.00014862777607049793)),(to_sfixed_a(0.00020498734374996275)),(to_sfixed_a(0.0001236903917742893)),(to_sfixed_a(7.991636812221259e-05)),(to_sfixed_a(-7.576032203360228e-06)),(to_sfixed_a(0.04831165447831154)),(to_sfixed_a(-0.00023457745555788279)),(to_sfixed_a(0.054647281765937805)),(to_sfixed_a(-0.025623155757784843)),(to_sfixed_a(0.0732036754488945)),(to_sfixed_a(0.05270499736070633)),(to_sfixed_a(0.09980852901935577)),(to_sfixed_a(0.17402751743793488)),(to_sfixed_a(-0.013974525034427643)),(to_sfixed_a(0.16411800682544708)),(to_sfixed_a(-0.12688368558883667)),(to_sfixed_a(-0.08729236572980881)),(to_sfixed_a(-0.01699436642229557)),(to_sfixed_a(-0.03451834246516228)),(to_sfixed_a(6.626189133385196e-05)),(to_sfixed_a(8.565034659113735e-05)),(to_sfixed_a(-9.02005413081497e-05)),(to_sfixed_a(-0.0001019686897052452)),(to_sfixed_a(0.00021044351160526276)),(to_sfixed_a(-0.00011841873492812738)),(to_sfixed_a(-0.00025709636975079775)),(to_sfixed_a(-0.0001098373977583833)),(to_sfixed_a(2.8957440008525737e-05)),(to_sfixed_a(-6.355899677146226e-05)),(to_sfixed_a(3.274892515037209e-05)),(to_sfixed_a(4.996838470106013e-06)),(to_sfixed_a(0.001239487319253385)),(to_sfixed_a(-0.04695524647831917)),(to_sfixed_a(0.025547632947564125)),(to_sfixed_a(0.07277921587228775)),(to_sfixed_a(-0.242929607629776)),(to_sfixed_a(-0.11514008045196533)),(to_sfixed_a(0.2361040562391281)),(to_sfixed_a(0.08070625364780426)),(to_sfixed_a(0.10927731543779373)),(to_sfixed_a(0.2940632104873657)),(to_sfixed_a(0.3332069516181946)),(to_sfixed_a(0.03144285827875137)),(to_sfixed_a(-0.049981698393821716)),(to_sfixed_a(0.024216603487730026)),(to_sfixed_a(-0.01736045442521572)),(to_sfixed_a(-0.1349487602710724)),(to_sfixed_a(-0.04175374284386635)),(to_sfixed_a(0.0001069547506631352)),(to_sfixed_a(0.0006868471973575652)),(to_sfixed_a(-8.233397238655016e-05)),(to_sfixed_a(8.483812052872963e-06)),(to_sfixed_a(-0.00011262127372901887)),(to_sfixed_a(-9.268052963307127e-06)),(to_sfixed_a(-0.00020271427638363093)),(to_sfixed_a(-0.00015282738604582846)),(to_sfixed_a(-1.001712735160254e-05)),(to_sfixed_a(-4.021831409772858e-05)),(to_sfixed_a(-0.06468971818685532)),(to_sfixed_a(0.008854739367961884)),(to_sfixed_a(-0.01827158033847809)),(to_sfixed_a(0.03487249091267586)),(to_sfixed_a(-0.15442301332950592)),(to_sfixed_a(-0.08899430930614471)),(to_sfixed_a(0.1794530153274536)),(to_sfixed_a(0.05364637449383736)),(to_sfixed_a(0.3221901059150696)),(to_sfixed_a(0.3193114101886749)),(to_sfixed_a(0.23531709611415863)),(to_sfixed_a(0.06777464598417282)),(to_sfixed_a(-0.11350873857736588)),(to_sfixed_a(0.07489147782325745)),(to_sfixed_a(-0.004568919539451599)),(to_sfixed_a(-0.0016728364862501621)),(to_sfixed_a(-0.09842196106910706)),(to_sfixed_a(0.0013726847246289253)),(to_sfixed_a(-0.012665082700550556)),(to_sfixed_a(0.002580928383395076)),(to_sfixed_a(9.628544648876414e-05)),(to_sfixed_a(-7.926363468868658e-05)),(to_sfixed_a(0.00026244239415973425)),(to_sfixed_a(5.407561911852099e-05)),(to_sfixed_a(2.6855230316868983e-05)),(to_sfixed_a(7.403325525956461e-06)),(to_sfixed_a(-7.137688953662291e-06)),(to_sfixed_a(0.00016836656141094863)),(to_sfixed_a(-0.06475140154361725)),(to_sfixed_a(-0.06704606860876083)),(to_sfixed_a(-0.13115832209587097)),(to_sfixed_a(-0.12103359401226044)),(to_sfixed_a(-0.15159255266189575)),(to_sfixed_a(0.3498294949531555)),(to_sfixed_a(0.290958046913147)),(to_sfixed_a(0.04910518601536751)),(to_sfixed_a(0.2030821442604065)),(to_sfixed_a(0.13208448886871338)),(to_sfixed_a(0.04476664587855339)),(to_sfixed_a(0.156744122505188)),(to_sfixed_a(0.06402429193258286)),(to_sfixed_a(-0.20973283052444458)),(to_sfixed_a(-0.054341334849596024)),(to_sfixed_a(-0.10133137553930283)),(to_sfixed_a(0.12023799121379852)),(to_sfixed_a(0.09785519540309906)),(to_sfixed_a(0.03773988410830498)),(to_sfixed_a(0.0028292564675211906)),(to_sfixed_a(0.0028361622244119644)),(to_sfixed_a(0.0013224383583292365)),(to_sfixed_a(-0.00021526828641071916)),(to_sfixed_a(-0.0001380104513373226)),(to_sfixed_a(-0.00013889861293137074)),(to_sfixed_a(-5.063740536570549e-05)),(to_sfixed_a(-0.00026018277276307344)),(to_sfixed_a(-0.00014376474427990615)),(to_sfixed_a(-0.027296463027596474)),(to_sfixed_a(-0.04145296663045883)),(to_sfixed_a(-0.10883836448192596)),(to_sfixed_a(0.15999922156333923)),(to_sfixed_a(0.1322227567434311)),(to_sfixed_a(0.3887496292591095)),(to_sfixed_a(-0.035315509885549545)),(to_sfixed_a(-0.23675888776779175)),(to_sfixed_a(0.09121537953615189)),(to_sfixed_a(-0.18890070915222168)),(to_sfixed_a(0.11813008785247803)),(to_sfixed_a(0.04165979474782944)),(to_sfixed_a(0.08753149211406708)),(to_sfixed_a(0.15288884937763214)),(to_sfixed_a(0.3862465023994446)),(to_sfixed_a(0.07779204845428467)),(to_sfixed_a(-0.27669790387153625)),(to_sfixed_a(0.002007882809266448)),(to_sfixed_a(-0.03767571225762367)),(to_sfixed_a(-0.007830284535884857)),(to_sfixed_a(0.003029701765626669)),(to_sfixed_a(-3.256453783251345e-05)),(to_sfixed_a(-0.0002539419801905751)),(to_sfixed_a(-6.6874340518552344e-06)),(to_sfixed_a(0.00010562109673628584)),(to_sfixed_a(-0.00018464720051269978)),(to_sfixed_a(-0.00018197015742771327)),(to_sfixed_a(0.029152149334549904)),(to_sfixed_a(-0.10250464826822281)),(to_sfixed_a(-0.006465062033385038)),(to_sfixed_a(0.06473474949598312)),(to_sfixed_a(-0.19110122323036194)),(to_sfixed_a(0.05412956699728966)),(to_sfixed_a(0.3604489266872406)),(to_sfixed_a(-0.1557917594909668)),(to_sfixed_a(-0.2733123302459717)),(to_sfixed_a(0.08128976076841354)),(to_sfixed_a(-0.15968672931194305)),(to_sfixed_a(0.3663398325443268)),(to_sfixed_a(-0.00431346520781517)),(to_sfixed_a(0.1029479131102562)),(to_sfixed_a(0.07628174871206284)),(to_sfixed_a(0.09008952230215073)),(to_sfixed_a(0.27112892270088196)),(to_sfixed_a(0.10078506916761398)),(to_sfixed_a(-0.04986388981342316)),(to_sfixed_a(0.14868609607219696)),(to_sfixed_a(0.11533964425325394)),(to_sfixed_a(0.016723329201340675)),(to_sfixed_a(-3.0144627089612186e-05)),(to_sfixed_a(-0.0002484588185325265)),(to_sfixed_a(-0.00028039992321282625)),(to_sfixed_a(7.633002678630874e-05)),(to_sfixed_a(8.739367331145331e-05)),(to_sfixed_a(-0.0002577236155048013)),(to_sfixed_a(-0.0019483116921037436)),(to_sfixed_a(-0.02863944135606289)),(to_sfixed_a(0.03263188526034355)),(to_sfixed_a(-0.11077747493982315)),(to_sfixed_a(-0.04949130862951279)),(to_sfixed_a(-0.07555872946977615)),(to_sfixed_a(0.30828434228897095)),(to_sfixed_a(0.2638789713382721)),(to_sfixed_a(0.05155729129910469)),(to_sfixed_a(0.04243630915880203)),(to_sfixed_a(-0.1360289752483368)),(to_sfixed_a(0.3770749270915985)),(to_sfixed_a(0.028905440121889114)),(to_sfixed_a(0.17989562451839447)),(to_sfixed_a(0.07218275964260101)),(to_sfixed_a(-0.2039022445678711)),(to_sfixed_a(-0.20251326262950897)),(to_sfixed_a(-0.025716397911310196)),(to_sfixed_a(0.18721242249011993)),(to_sfixed_a(0.13425412774085999)),(to_sfixed_a(-0.011488810181617737)),(to_sfixed_a(-6.475250847870484e-05)),(to_sfixed_a(-5.0538026698632166e-05)),(to_sfixed_a(-6.976692384341732e-05)),(to_sfixed_a(1.5145344150369056e-05)),(to_sfixed_a(-4.158377487328835e-05)),(to_sfixed_a(9.208938718074933e-05)),(to_sfixed_a(9.562447667121887e-05)),(to_sfixed_a(0.010991767980158329)),(to_sfixed_a(0.002469389932230115)),(to_sfixed_a(0.195283442735672)),(to_sfixed_a(0.06259558349847794)),(to_sfixed_a(0.19801166653633118)),(to_sfixed_a(-0.047413576394319534)),(to_sfixed_a(0.1409243941307068)),(to_sfixed_a(-0.30328676104545593)),(to_sfixed_a(-0.14094699919223785)),(to_sfixed_a(-0.22164572775363922)),(to_sfixed_a(0.2589260935783386)),(to_sfixed_a(-0.024164345115423203)),(to_sfixed_a(0.22257600724697113)),(to_sfixed_a(0.06687722355127335)),(to_sfixed_a(-0.04791047424077988)),(to_sfixed_a(0.016755636781454086)),(to_sfixed_a(0.04602816700935364)),(to_sfixed_a(-0.05401041731238365)),(to_sfixed_a(0.043793339282274246)),(to_sfixed_a(-0.19180777668952942)),(to_sfixed_a(0.0989367887377739)),(to_sfixed_a(0.003462923923507333)),(to_sfixed_a(-8.938307473727036e-06)),(to_sfixed_a(0.00026711076498031616)),(to_sfixed_a(-0.0003117866290267557)),(to_sfixed_a(0.00011368070408934727)),(to_sfixed_a(-2.555290166128543e-06)),(to_sfixed_a(-0.03494463115930557)),(to_sfixed_a(0.054843366146087646)),(to_sfixed_a(0.046854496002197266)),(to_sfixed_a(0.06490899622440338)),(to_sfixed_a(0.0029757481534034014)),(to_sfixed_a(-0.030476462095975876)),(to_sfixed_a(-0.10019876062870026)),(to_sfixed_a(-0.03302069380879402)),(to_sfixed_a(-0.03056558594107628)),(to_sfixed_a(-0.09287760406732559)),(to_sfixed_a(0.17662963271141052)),(to_sfixed_a(-0.031572744250297546)),(to_sfixed_a(0.03306341543793678)),(to_sfixed_a(-0.0030935194808989763)),(to_sfixed_a(0.05317390710115433)),(to_sfixed_a(0.05289237201213837)),(to_sfixed_a(-0.02354745753109455)),(to_sfixed_a(0.005836424417793751)),(to_sfixed_a(0.157302588224411)),(to_sfixed_a(-0.01953013613820076)),(to_sfixed_a(-0.188542902469635)),(to_sfixed_a(-0.0748453140258789)),(to_sfixed_a(-3.180869316565804e-05)),(to_sfixed_a(-0.00024031769135035574)),(to_sfixed_a(-5.760676140198484e-05)),(to_sfixed_a(-0.00020459819643292576)),(to_sfixed_a(-9.578950994182378e-05)),(to_sfixed_a(5.614344627247192e-05)),(to_sfixed_a(-0.0001226829190272838)),(to_sfixed_a(-0.04603379964828491)),(to_sfixed_a(0.13387691974639893)),(to_sfixed_a(0.08885631710290909)),(to_sfixed_a(0.013060878962278366)),(to_sfixed_a(0.029006628319621086)),(to_sfixed_a(-0.21854902803897858)),(to_sfixed_a(-0.12601657211780548)),(to_sfixed_a(0.06916269659996033)),(to_sfixed_a(0.101469986140728)),(to_sfixed_a(-0.09041465818881989)),(to_sfixed_a(0.09743347018957138)),(to_sfixed_a(0.18448254466056824)),(to_sfixed_a(-0.0058603896759450436)),(to_sfixed_a(-0.0317230261862278)),(to_sfixed_a(0.33086127042770386)),(to_sfixed_a(0.06235295906662941)),(to_sfixed_a(-0.006676380056887865)),(to_sfixed_a(0.01879231631755829)),(to_sfixed_a(-0.040762174874544144)),(to_sfixed_a(0.03220660611987114)),(to_sfixed_a(0.012379618361592293)),(to_sfixed_a(-0.00010877431486733258)),(to_sfixed_a(0.00017999298870563507)),(to_sfixed_a(0.0001944681425811723)),(to_sfixed_a(1.6907746612560004e-05)),(to_sfixed_a(-1.3360370758164208e-05)),(to_sfixed_a(-3.5505239793565124e-05)),(to_sfixed_a(-0.00014235432900022715)),(to_sfixed_a(0.06075885519385338)),(to_sfixed_a(0.08825115114450455)),(to_sfixed_a(0.2326866090297699)),(to_sfixed_a(0.11490431427955627)),(to_sfixed_a(-0.049646131694316864)),(to_sfixed_a(0.025026442483067513)),(to_sfixed_a(-0.03617095574736595)),(to_sfixed_a(0.09636319428682327)),(to_sfixed_a(-0.06957514584064484)),(to_sfixed_a(-1.6652026033625589e-06)),(to_sfixed_a(-0.027942858636379242)),(to_sfixed_a(0.13444958627223969)),(to_sfixed_a(-0.12542884051799774)),(to_sfixed_a(0.014490281231701374)),(to_sfixed_a(-0.058968909084796906)),(to_sfixed_a(0.0906587615609169)),(to_sfixed_a(0.010973842814564705)),(to_sfixed_a(-0.02748027630150318)),(to_sfixed_a(0.06129835173487663)),(to_sfixed_a(0.01765337772667408)),(to_sfixed_a(0.06492459774017334)),(to_sfixed_a(0.0036575712729245424)),(to_sfixed_a(0.0044291336089372635)),(to_sfixed_a(-0.00012120314931962639)),(to_sfixed_a(-3.3107698982348666e-05)),(to_sfixed_a(-5.698743188986555e-05)),(to_sfixed_a(-1.3772742022410966e-05)),(to_sfixed_a(-9.221530490322039e-05)),(to_sfixed_a(0.001743473345413804)),(to_sfixed_a(0.17008058726787567)),(to_sfixed_a(0.006419460289180279)),(to_sfixed_a(0.09931452572345734)),(to_sfixed_a(-0.052940886467695236)),(to_sfixed_a(-0.23390372097492218)),(to_sfixed_a(-0.03152807056903839)),(to_sfixed_a(0.04164842888712883)),(to_sfixed_a(-0.05023786798119545)),(to_sfixed_a(-0.08897493779659271)),(to_sfixed_a(0.011130531318485737)),(to_sfixed_a(-0.060825053602457047)),(to_sfixed_a(-0.34998998045921326)),(to_sfixed_a(0.02569674700498581)),(to_sfixed_a(0.1376599818468094)),(to_sfixed_a(0.0762835443019867)),(to_sfixed_a(0.039015818387269974)),(to_sfixed_a(-0.12606407701969147)),(to_sfixed_a(-0.003134318860247731)),(to_sfixed_a(-0.027676871046423912)),(to_sfixed_a(-0.019543366506695747)),(to_sfixed_a(7.919922609289642e-06)),(to_sfixed_a(9.608526306692511e-05)),(to_sfixed_a(2.183215292461682e-05)),(to_sfixed_a(5.682626215275377e-05)),(to_sfixed_a(-0.00012281279487069696)),(to_sfixed_a(0.00025324951275251806)),(to_sfixed_a(0.00032801320776343346)),(to_sfixed_a(0.02343016117811203)),(to_sfixed_a(0.1123499944806099)),(to_sfixed_a(0.016210224479436874)),(to_sfixed_a(0.12677372992038727)),(to_sfixed_a(-0.1599269062280655)),(to_sfixed_a(0.1735956221818924)),(to_sfixed_a(0.022607002407312393)),(to_sfixed_a(-0.2055586725473404)),(to_sfixed_a(-0.13815516233444214)),(to_sfixed_a(0.14119303226470947)),(to_sfixed_a(0.033250756561756134)),(to_sfixed_a(-0.05974534526467323)),(to_sfixed_a(-0.26696690917015076)),(to_sfixed_a(0.19412407279014587)),(to_sfixed_a(0.0290987491607666)),(to_sfixed_a(0.13952331244945526)),(to_sfixed_a(-0.03416077420115471)),(to_sfixed_a(-0.01622546650469303)),(to_sfixed_a(-0.011700299568474293)),(to_sfixed_a(-0.07550361752510071)),(to_sfixed_a(0.004081662744283676)),(to_sfixed_a(0.0002771352883428335)),(to_sfixed_a(7.2706238825048786e-06)),(to_sfixed_a(0.00012977400911040604)),(to_sfixed_a(-0.00024855704396031797)),(to_sfixed_a(7.949527207529172e-05)),(to_sfixed_a(5.3503852541325614e-05)),(to_sfixed_a(0.0025370034854859114)),(to_sfixed_a(0.010410089045763016)),(to_sfixed_a(0.02366134710609913)),(to_sfixed_a(0.008997534401714802)),(to_sfixed_a(-0.1222863420844078)),(to_sfixed_a(0.00581109756603837)),(to_sfixed_a(-0.17265582084655762)),(to_sfixed_a(-0.08040039986371994)),(to_sfixed_a(0.1386273056268692)),(to_sfixed_a(-0.11506524682044983)),(to_sfixed_a(-0.015225746668875217)),(to_sfixed_a(-0.04212841019034386)),(to_sfixed_a(-0.17963725328445435)),(to_sfixed_a(-0.1258951723575592)),(to_sfixed_a(0.21359451115131378)),(to_sfixed_a(0.11633287370204926)),(to_sfixed_a(-0.0017612648662179708)),(to_sfixed_a(0.17016145586967468)),(to_sfixed_a(0.1065862700343132)),(to_sfixed_a(0.06020290404558182)),(to_sfixed_a(-0.0640861839056015)),(to_sfixed_a(0.09035584330558777)),(to_sfixed_a(-0.005634885281324387)),(to_sfixed_a(-0.00011697873560478911)),(to_sfixed_a(-8.063539667091391e-07)),(to_sfixed_a(8.73347744345665e-05)),(to_sfixed_a(0.00019366668129805475)),(to_sfixed_a(0.0021186843514442444)),(to_sfixed_a(0.0025957238394767046)),(to_sfixed_a(0.032141413539648056)),(to_sfixed_a(0.009728864766657352)),(to_sfixed_a(-0.08554144948720932)),(to_sfixed_a(-0.14864566922187805)),(to_sfixed_a(0.013134266249835491)),(to_sfixed_a(-0.02710714004933834)),(to_sfixed_a(0.013018274679780006)),(to_sfixed_a(-0.024296436458826065)),(to_sfixed_a(-0.15674154460430145)),(to_sfixed_a(-0.02877386473119259)),(to_sfixed_a(-0.07182876020669937)),(to_sfixed_a(0.053315792232751846)),(to_sfixed_a(-0.045346830040216446)),(to_sfixed_a(0.12300878763198853)),(to_sfixed_a(-0.08442674577236176)),(to_sfixed_a(0.121673084795475)),(to_sfixed_a(0.1211804747581482)),(to_sfixed_a(-0.08724111318588257)),(to_sfixed_a(-0.17731167376041412)),(to_sfixed_a(-0.018358446657657623)),(to_sfixed_a(0.00027181149926036596)),(to_sfixed_a(7.506613474106416e-05)),(to_sfixed_a(2.5705485313665122e-05)),(to_sfixed_a(3.2589287002338096e-05)),(to_sfixed_a(-1.1744531548174564e-05)),(to_sfixed_a(-0.00010773645772133023)),(to_sfixed_a(6.309125456027687e-05)),(to_sfixed_a(-0.0006731604225933552)),(to_sfixed_a(-0.0012744998093694448)),(to_sfixed_a(-0.17260698974132538)),(to_sfixed_a(-0.29613035917282104)),(to_sfixed_a(-0.08727958798408508)),(to_sfixed_a(0.08661136776208878)),(to_sfixed_a(-0.03098464570939541)),(to_sfixed_a(0.19391174614429474)),(to_sfixed_a(0.03759711608290672)),(to_sfixed_a(0.059156570583581924)),(to_sfixed_a(-0.17822477221488953)),(to_sfixed_a(0.24548742175102234)),(to_sfixed_a(0.20280945301055908)),(to_sfixed_a(0.260099858045578)),(to_sfixed_a(0.17791466414928436)),(to_sfixed_a(0.2004663646221161)),(to_sfixed_a(0.2680543065071106)),(to_sfixed_a(0.04181119054555893)),(to_sfixed_a(-0.14268679916858673)),(to_sfixed_a(-0.03924514353275299)),(to_sfixed_a(0.05414824187755585)),(to_sfixed_a(0.0026676193810999393)),(to_sfixed_a(0.00012956939463037997)),(to_sfixed_a(-0.00023289656382985413)),(to_sfixed_a(-0.00011195868137292564)),(to_sfixed_a(0.00015199236804619431)),(to_sfixed_a(0.0001253080554306507)),(to_sfixed_a(5.8699391956906766e-05)),(to_sfixed_a(0.0008909716852940619)),(to_sfixed_a(-0.0037925569340586662)),(to_sfixed_a(-0.046207740902900696)),(to_sfixed_a(-0.10489504039287567)),(to_sfixed_a(-0.15580162405967712)),(to_sfixed_a(-0.17329294979572296)),(to_sfixed_a(-0.22127659618854523)),(to_sfixed_a(0.07644560933113098)),(to_sfixed_a(0.0094583285972476)),(to_sfixed_a(0.2065931111574173)),(to_sfixed_a(0.2476678490638733)),(to_sfixed_a(0.1175297349691391)),(to_sfixed_a(-0.029564637690782547)),(to_sfixed_a(-0.05989053100347519)),(to_sfixed_a(0.10831031203269958)),(to_sfixed_a(0.16190756857395172)),(to_sfixed_a(0.023891400545835495)),(to_sfixed_a(-0.04913540557026863)),(to_sfixed_a(0.037790052592754364)),(to_sfixed_a(0.009117105975747108)),(to_sfixed_a(-0.09551562368869781)),(to_sfixed_a(-4.841382906306535e-05)),(to_sfixed_a(9.856148608378135e-06)),(to_sfixed_a(2.5578036002116278e-05)),(to_sfixed_a(0.00018035453103948385)),(to_sfixed_a(3.097969454302074e-07)),(to_sfixed_a(0.00011975429515587166)),(to_sfixed_a(5.2527273510349914e-05)),(to_sfixed_a(6.636950274696574e-05)),(to_sfixed_a(-0.037209149450063705)),(to_sfixed_a(-0.03156067430973053)),(to_sfixed_a(-0.27865123748779297)),(to_sfixed_a(0.2936984896659851)),(to_sfixed_a(0.00872021447867155)),(to_sfixed_a(0.09747698158025742)),(to_sfixed_a(-0.19298993051052094)),(to_sfixed_a(0.24288904666900635)),(to_sfixed_a(-0.07072034478187561)),(to_sfixed_a(-0.10107100009918213)),(to_sfixed_a(-0.13703222572803497)),(to_sfixed_a(0.18871526420116425)),(to_sfixed_a(0.12679733335971832)),(to_sfixed_a(0.16029170155525208)),(to_sfixed_a(0.1629333347082138)),(to_sfixed_a(0.18646065890789032)),(to_sfixed_a(0.014949637465178967)),(to_sfixed_a(0.072471022605896)),(to_sfixed_a(0.04801400005817413)),(to_sfixed_a(0.04075966402888298)),(to_sfixed_a(0.06183795630931854)),(to_sfixed_a(-0.0001426608068868518)),(to_sfixed_a(-5.6161377870012075e-05)),(to_sfixed_a(-4.6737513912376016e-05)),(to_sfixed_a(0.00017022498650476336)),(to_sfixed_a(-0.0001043895972543396)),(to_sfixed_a(-0.00011231517419219017)),(to_sfixed_a(5.73874385736417e-05)),(to_sfixed_a(-0.01310705952346325)),(to_sfixed_a(-0.0017653737450018525)),(to_sfixed_a(0.04737546294927597)),(to_sfixed_a(0.39137810468673706)),(to_sfixed_a(-0.014829814434051514)),(to_sfixed_a(-0.10605539381504059)),(to_sfixed_a(0.02612663432955742)),(to_sfixed_a(0.10680824518203735)),(to_sfixed_a(0.04581147059798241)),(to_sfixed_a(0.04379052296280861)),(to_sfixed_a(-0.14352205395698547)),(to_sfixed_a(-0.1282610297203064)),(to_sfixed_a(-0.06637676805257797)),(to_sfixed_a(0.011774025857448578)),(to_sfixed_a(-0.028104247525334358)),(to_sfixed_a(-0.015372782945632935)),(to_sfixed_a(0.29798251390457153)),(to_sfixed_a(0.10109852999448776)),(to_sfixed_a(-0.21862071752548218)),(to_sfixed_a(0.0007103574462234974)),(to_sfixed_a(0.030185271054506302)),(to_sfixed_a(0.0001308481878368184)),(to_sfixed_a(-9.128437523031607e-05)),(to_sfixed_a(0.00010015119187301025)),(to_sfixed_a(-0.00015082801110111177)),(to_sfixed_a(0.00021003533038310707)),(to_sfixed_a(-7.316830306081101e-05)),(to_sfixed_a(-0.000271448923740536)),(to_sfixed_a(-0.0004212800704408437)),(to_sfixed_a(0.036951787769794464)),(to_sfixed_a(0.020491180941462517)),(to_sfixed_a(-0.101023830473423)),(to_sfixed_a(-0.03140052780508995)),(to_sfixed_a(0.0776955857872963)),(to_sfixed_a(-0.0088008102029562)),(to_sfixed_a(-0.06803110241889954)),(to_sfixed_a(-0.08835390955209732)),(to_sfixed_a(0.05051247775554657)),(to_sfixed_a(-0.037823986262083054)),(to_sfixed_a(-0.037543896585702896)),(to_sfixed_a(0.053493428975343704)),(to_sfixed_a(-0.15073001384735107)),(to_sfixed_a(-0.09510762244462967)),(to_sfixed_a(-0.12167669087648392)),(to_sfixed_a(0.013028956018388271)),(to_sfixed_a(-0.028965376317501068)),(to_sfixed_a(-0.018980909138917923)),(to_sfixed_a(-0.0017271337565034628)),(to_sfixed_a(-5.223428888712078e-05)),(to_sfixed_a(-0.00010469312110217288)),(to_sfixed_a(9.092795517062768e-05)),(to_sfixed_a(0.00020024807599838823)),(to_sfixed_a(0.00010836917499545962)),(to_sfixed_a(-6.899714935570955e-05)),(to_sfixed_a(-4.7858284233370796e-05)),(to_sfixed_a(2.822863098117523e-05)),(to_sfixed_a(-0.0004062283842358738)),(to_sfixed_a(0.013230407610535622)),(to_sfixed_a(-0.002151066903024912)),(to_sfixed_a(-0.05941149592399597)),(to_sfixed_a(-0.028506722301244736)),(to_sfixed_a(-0.07231637835502625)),(to_sfixed_a(-0.04832589998841286)),(to_sfixed_a(-0.07009827345609665)),(to_sfixed_a(0.04352465271949768)),(to_sfixed_a(-0.16967275738716125)),(to_sfixed_a(-0.0444134920835495)),(to_sfixed_a(0.004782574716955423)),(to_sfixed_a(-0.2728830873966217)),(to_sfixed_a(-0.2135871946811676)),(to_sfixed_a(-0.017094623297452927)),(to_sfixed_a(0.007563436403870583)),(to_sfixed_a(-0.04716477543115616)),(to_sfixed_a(-0.3419141173362732)),(to_sfixed_a(0.005525572691112757)),(to_sfixed_a(-0.25217634439468384)),(to_sfixed_a(-2.545898678363301e-05)),(to_sfixed_a(-1.2677409358730074e-05)),(to_sfixed_a(2.549789314798545e-05)),(to_sfixed_a(-7.460491906385869e-05)),(to_sfixed_a(2.793501698761247e-05)),(to_sfixed_a(-6.402565873031563e-07)),(to_sfixed_a(0.00010492804722161964)),(to_sfixed_a(5.2270839660195634e-05)),(to_sfixed_a(-0.04631797596812248)),(to_sfixed_a(-0.03020639345049858)),(to_sfixed_a(-0.19202692806720734)),(to_sfixed_a(-0.04393446817994118)),(to_sfixed_a(0.06423083692789078)),(to_sfixed_a(0.1559796780347824)),(to_sfixed_a(0.01287910994142294)),(to_sfixed_a(-0.0072944508865475655)),(to_sfixed_a(-0.05934688448905945)),(to_sfixed_a(-0.07759847491979599)),(to_sfixed_a(-0.08377248048782349)),(to_sfixed_a(-0.0772584080696106)),(to_sfixed_a(0.08292289823293686)),(to_sfixed_a(-0.02121976763010025)),(to_sfixed_a(-0.0031499930191785097)),(to_sfixed_a(-0.2782745361328125)),(to_sfixed_a(0.005802174564450979)),(to_sfixed_a(-0.27401599287986755)),(to_sfixed_a(-0.1231689453125)),(to_sfixed_a(0.011850825510919094)),(to_sfixed_a(-6.870767538202927e-05)),(to_sfixed_a(7.182348326750798e-06)),(to_sfixed_a(-0.00011366981198079884)),(to_sfixed_a(6.771496555302292e-05)),(to_sfixed_a(-8.667397924000397e-05)),(to_sfixed_a(-6.326151196844876e-05)),(to_sfixed_a(-1.7397565898136236e-05)),(to_sfixed_a(0.00019213331688661128)),(to_sfixed_a(-0.00017198498244397342)),(to_sfixed_a(-0.01786726340651512)),(to_sfixed_a(-0.1161731481552124)),(to_sfixed_a(-0.10642290115356445)),(to_sfixed_a(-0.11815112084150314)),(to_sfixed_a(-0.0631486251950264)),(to_sfixed_a(-0.21643444895744324)),(to_sfixed_a(0.024571746587753296)),(to_sfixed_a(-0.005879649892449379)),(to_sfixed_a(-0.03184497356414795)),(to_sfixed_a(0.015191017650067806)),(to_sfixed_a(-0.002613103948533535)),(to_sfixed_a(-0.09422408789396286)),(to_sfixed_a(0.0355994738638401)),(to_sfixed_a(0.009081951342523098)),(to_sfixed_a(-0.05329563841223717)),(to_sfixed_a(0.18699268996715546)),(to_sfixed_a(0.0005750391283072531)),(to_sfixed_a(0.006334299687296152)),(to_sfixed_a(0.006554936058819294)),(to_sfixed_a(9.496403072262183e-05)),(to_sfixed_a(0.0003769296745304018)),(to_sfixed_a(4.421743142302148e-05)),(to_sfixed_a(0.00015034529496915638)),(to_sfixed_a(-0.00013269427290651947)),(to_sfixed_a(-0.00012628748663701117)),(to_sfixed_a(7.424484647344798e-05)),(to_sfixed_a(-4.695082225225633e-06)),(to_sfixed_a(4.582779365591705e-05)),(to_sfixed_a(-0.0008630690863355994)),(to_sfixed_a(-0.0007313894457183778)),(to_sfixed_a(3.29461254295893e-05)),(to_sfixed_a(6.62191814626567e-05)),(to_sfixed_a(0.0005066730664111674)),(to_sfixed_a(0.05628981813788414)),(to_sfixed_a(0.007109944708645344)),(to_sfixed_a(0.0016936756437644362)),(to_sfixed_a(0.045818571001291275)),(to_sfixed_a(-0.04313244670629501)),(to_sfixed_a(-0.022182181477546692)),(to_sfixed_a(-0.06393956393003464)),(to_sfixed_a(0.040498506277799606)),(to_sfixed_a(0.06459994614124298)),(to_sfixed_a(0.015588314272463322)),(to_sfixed_a(0.00495017459616065)),(to_sfixed_a(1.2309817066125106e-05)),(to_sfixed_a(1.1333412658132147e-05)),(to_sfixed_a(-0.00026062389952130616)),(to_sfixed_a(-0.000387116422643885)),(to_sfixed_a(-0.00013605646381620318)),(to_sfixed_a(0.000205707605346106)),(to_sfixed_a(-8.434318442596123e-05)),(to_sfixed_a(0.0002549214696045965)),(to_sfixed_a(0.000330889830365777)),(to_sfixed_a(5.3402352932607755e-05)),(to_sfixed_a(0.00017938348173629493)),(to_sfixed_a(0.00017732100968714803)),(to_sfixed_a(1.0503343219170347e-05)),(to_sfixed_a(0.00017989524349104613)),(to_sfixed_a(0.0003108694509137422)),(to_sfixed_a(5.7935190852731466e-05)),(to_sfixed_a(0.00028126456891186535)),(to_sfixed_a(0.00011204813199583441)),(to_sfixed_a(-0.000154643232235685)),(to_sfixed_a(2.3854758183006197e-05)),(to_sfixed_a(-4.446151797310449e-05)),(to_sfixed_a(0.000433913228334859)),(to_sfixed_a(0.00015279659419320524)),(to_sfixed_a(0.0001366765209240839)),(to_sfixed_a(0.000302442058455199)),(to_sfixed_a(0.00011503748100949451)),(to_sfixed_a(-0.00021746079437434673)),(to_sfixed_a(-0.000174495653482154)),(to_sfixed_a(0.0001437674800399691)),(to_sfixed_a(9.099706949200481e-05)),(to_sfixed_a(-0.00025936454767361283)),(to_sfixed_a(2.841899731720332e-05)),(to_sfixed_a(-0.0001707281480776146)),(to_sfixed_a(8.746905223233625e-05)),(to_sfixed_a(0.00021324244153220206)));

    constant weight_n0_35 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(9.062876051757485e-05)),(to_sfixed_a(-0.000148109276778996)),(to_sfixed_a(-0.00013275073433760554)),(to_sfixed_a(-1.618426358618308e-05)),(to_sfixed_a(-6.188327097333968e-05)),(to_sfixed_a(0.00012871739454567432)),(to_sfixed_a(0.00015802336565684527)),(to_sfixed_a(-3.325511352159083e-05)),(to_sfixed_a(0.0002885019057430327)),(to_sfixed_a(0.0002269537653774023)),(to_sfixed_a(-2.610689307402936e-06)),(to_sfixed_a(-8.108275505946949e-05)),(to_sfixed_a(-6.383093568729237e-05)),(to_sfixed_a(-0.00019907066598534584)),(to_sfixed_a(-0.00010634636419126764)),(to_sfixed_a(-0.00016194504860322922)),(to_sfixed_a(-0.0001830048713600263)),(to_sfixed_a(-6.543695781147107e-05)),(to_sfixed_a(9.991461411118507e-05)),(to_sfixed_a(0.00021572531841229647)),(to_sfixed_a(-0.00010736856347648427)),(to_sfixed_a(-0.00024265347747132182)),(to_sfixed_a(-2.105149360431824e-05)),(to_sfixed_a(-3.409985583857633e-05)),(to_sfixed_a(-0.000123854391858913)),(to_sfixed_a(3.111913247266784e-05)),(to_sfixed_a(0.00012527989747468382)),(to_sfixed_a(5.524312655325048e-05)),(to_sfixed_a(5.683406925527379e-05)),(to_sfixed_a(-7.273205847013742e-05)),(to_sfixed_a(7.697943510720506e-05)),(to_sfixed_a(-0.0002123538579326123)),(to_sfixed_a(0.00011533971701283008)),(to_sfixed_a(5.3203420975478366e-05)),(to_sfixed_a(-7.052686851238832e-05)),(to_sfixed_a(-0.00030455656815320253)),(to_sfixed_a(2.7103051252197474e-05)),(to_sfixed_a(0.0002042550768237561)),(to_sfixed_a(5.7805547839961946e-05)),(to_sfixed_a(-0.00010528980783419684)),(to_sfixed_a(1.1696547517203726e-05)),(to_sfixed_a(3.294291309430264e-05)),(to_sfixed_a(-0.00030495994724333286)),(to_sfixed_a(-0.00013078803021926433)),(to_sfixed_a(-7.298071068362333e-06)),(to_sfixed_a(3.58204088115599e-05)),(to_sfixed_a(6.382119318004698e-05)),(to_sfixed_a(-0.0001289801875827834)),(to_sfixed_a(-0.00014282586926128715)),(to_sfixed_a(4.2306186514906585e-05)),(to_sfixed_a(7.036341412458569e-05)),(to_sfixed_a(0.00013557127385865897)),(to_sfixed_a(1.8470898794475943e-05)),(to_sfixed_a(0.00019866431830450892)),(to_sfixed_a(0.0001383641647407785)),(to_sfixed_a(-6.606139504583552e-05)),(to_sfixed_a(6.19251950411126e-05)),(to_sfixed_a(-0.0004644119180738926)),(to_sfixed_a(-0.0001162965054390952)),(to_sfixed_a(1.7842870875028893e-05)),(to_sfixed_a(4.546178752207197e-05)),(to_sfixed_a(-3.7623340176651254e-06)),(to_sfixed_a(0.00021474128880072385)),(to_sfixed_a(0.0001310324587393552)),(to_sfixed_a(-0.00017703072808217257)),(to_sfixed_a(-5.941180279478431e-05)),(to_sfixed_a(1.4697012375108898e-05)),(to_sfixed_a(1.9234001058521244e-07)),(to_sfixed_a(0.00011766995157813653)),(to_sfixed_a(-0.035616371780633926)),(to_sfixed_a(0.00013759435387328267)),(to_sfixed_a(0.00034687298466451466)),(to_sfixed_a(-4.024149529868737e-05)),(to_sfixed_a(-0.00014218577416613698)),(to_sfixed_a(8.582227019360289e-05)),(to_sfixed_a(-0.00010861296323128045)),(to_sfixed_a(0.0001922921946970746)),(to_sfixed_a(1.701648761809338e-05)),(to_sfixed_a(9.545517968945205e-05)),(to_sfixed_a(0.00012533064000308514)),(to_sfixed_a(-0.00044169038301333785)),(to_sfixed_a(-0.00030591050744988024)),(to_sfixed_a(-1.4418484170164447e-05)),(to_sfixed_a(6.597619358217344e-05)),(to_sfixed_a(9.35654024942778e-05)),(to_sfixed_a(0.00022968862322159111)),(to_sfixed_a(0.0001243526057805866)),(to_sfixed_a(0.00024982247850857675)),(to_sfixed_a(0.0001553614711156115)),(to_sfixed_a(-0.00023007688287179917)),(to_sfixed_a(-5.466554284794256e-05)),(to_sfixed_a(4.4619941036216915e-05)),(to_sfixed_a(0.032352015376091)),(to_sfixed_a(-4.081604856764898e-05)),(to_sfixed_a(0.03682651370763779)),(to_sfixed_a(0.02993047423660755)),(to_sfixed_a(0.03183991461992264)),(to_sfixed_a(0.018515318632125854)),(to_sfixed_a(0.045577019453048706)),(to_sfixed_a(-0.025806808844208717)),(to_sfixed_a(0.009628570638597012)),(to_sfixed_a(-0.09047248959541321)),(to_sfixed_a(0.06942758709192276)),(to_sfixed_a(-0.07423418015241623)),(to_sfixed_a(-0.0016073834849521518)),(to_sfixed_a(-0.0034198062494397163)),(to_sfixed_a(-5.573764155997196e-06)),(to_sfixed_a(-8.674577838974074e-05)),(to_sfixed_a(-0.00022368351346813142)),(to_sfixed_a(1.1520835869305301e-05)),(to_sfixed_a(-0.0002592217642813921)),(to_sfixed_a(0.0001770038070390001)),(to_sfixed_a(0.00012434128439053893)),(to_sfixed_a(-8.37125026009744e-06)),(to_sfixed_a(0.00019872441771440208)),(to_sfixed_a(9.291060268878937e-05)),(to_sfixed_a(-0.0001654896914260462)),(to_sfixed_a(-9.854313975665718e-05)),(to_sfixed_a(0.0002199467271566391)),(to_sfixed_a(-0.005612611770629883)),(to_sfixed_a(0.025920245796442032)),(to_sfixed_a(0.049214087426662445)),(to_sfixed_a(0.2096690833568573)),(to_sfixed_a(0.06316259503364563)),(to_sfixed_a(0.0587693452835083)),(to_sfixed_a(0.041210055351257324)),(to_sfixed_a(-0.14181344211101532)),(to_sfixed_a(-0.020131710916757584)),(to_sfixed_a(-0.0677284300327301)),(to_sfixed_a(-0.19660775363445282)),(to_sfixed_a(-0.021384742110967636)),(to_sfixed_a(0.011016763746738434)),(to_sfixed_a(-0.004675441887229681)),(to_sfixed_a(0.03450296074151993)),(to_sfixed_a(0.054458219558000565)),(to_sfixed_a(-0.00016619292728137225)),(to_sfixed_a(0.00035776966251432896)),(to_sfixed_a(-0.00020756959565915167)),(to_sfixed_a(-0.00014379186904989183)),(to_sfixed_a(-0.00022766370966564864)),(to_sfixed_a(-0.00017353483417537063)),(to_sfixed_a(-9.711613529361784e-05)),(to_sfixed_a(0.00021692995505873114)),(to_sfixed_a(5.6096843763953075e-05)),(to_sfixed_a(0.0010037869215011597)),(to_sfixed_a(-0.029530677944421768)),(to_sfixed_a(-0.015045526437461376)),(to_sfixed_a(-0.03713976964354515)),(to_sfixed_a(0.07438945770263672)),(to_sfixed_a(0.07268674671649933)),(to_sfixed_a(0.0068653360940515995)),(to_sfixed_a(0.16125167906284332)),(to_sfixed_a(0.1549442559480667)),(to_sfixed_a(-0.12808053195476532)),(to_sfixed_a(0.06405133008956909)),(to_sfixed_a(0.16041551530361176)),(to_sfixed_a(0.28507569432258606)),(to_sfixed_a(-0.10970904678106308)),(to_sfixed_a(-0.05511665716767311)),(to_sfixed_a(-0.0090376827865839)),(to_sfixed_a(0.06445523351430893)),(to_sfixed_a(0.17609770596027374)),(to_sfixed_a(0.003127256641164422)),(to_sfixed_a(0.029075242578983307)),(to_sfixed_a(0.0026456185150891542)),(to_sfixed_a(-0.00018210694543085992)),(to_sfixed_a(-0.00011837971396744251)),(to_sfixed_a(0.0001444131921743974)),(to_sfixed_a(0.00021446544269565493)),(to_sfixed_a(-0.00011501425615279004)),(to_sfixed_a(-0.00027713956660591066)),(to_sfixed_a(0.00023049963056109846)),(to_sfixed_a(-0.0004422779311425984)),(to_sfixed_a(-0.026342013850808144)),(to_sfixed_a(-0.02182878367602825)),(to_sfixed_a(-0.046566084027290344)),(to_sfixed_a(0.0919690728187561)),(to_sfixed_a(0.03286700323224068)),(to_sfixed_a(0.17574463784694672)),(to_sfixed_a(0.18561211228370667)),(to_sfixed_a(0.07077830284833908)),(to_sfixed_a(0.007424721959978342)),(to_sfixed_a(0.0014402579981833696)),(to_sfixed_a(-0.13994693756103516)),(to_sfixed_a(0.09736280143260956)),(to_sfixed_a(0.08115837723016739)),(to_sfixed_a(-0.029217099770903587)),(to_sfixed_a(-0.017588822171092033)),(to_sfixed_a(0.07072935253381729)),(to_sfixed_a(0.20048180222511292)),(to_sfixed_a(0.4713997542858124)),(to_sfixed_a(0.24519386887550354)),(to_sfixed_a(-0.003517819568514824)),(to_sfixed_a(-0.004430384375154972)),(to_sfixed_a(-0.004463774152100086)),(to_sfixed_a(0.00020641613809857517)),(to_sfixed_a(-7.0174181018956e-05)),(to_sfixed_a(-0.00020963513816241175)),(to_sfixed_a(5.480271647684276e-05)),(to_sfixed_a(0.0001879082847153768)),(to_sfixed_a(-3.4215860068798065e-05)),(to_sfixed_a(0.013427800498902798)),(to_sfixed_a(0.04542751982808113)),(to_sfixed_a(-0.1675015091896057)),(to_sfixed_a(-0.29770427942276)),(to_sfixed_a(-0.12454425543546677)),(to_sfixed_a(-0.11847042292356491)),(to_sfixed_a(0.008920280262827873)),(to_sfixed_a(-0.13899412751197815)),(to_sfixed_a(0.00816324632614851)),(to_sfixed_a(-0.04693219065666199)),(to_sfixed_a(0.07068974524736404)),(to_sfixed_a(0.031362470239400864)),(to_sfixed_a(0.2426666021347046)),(to_sfixed_a(-0.18144024908542633)),(to_sfixed_a(0.14216060936450958)),(to_sfixed_a(0.584881067276001)),(to_sfixed_a(0.06335508078336716)),(to_sfixed_a(-0.04785444214940071)),(to_sfixed_a(-0.06764055043458939)),(to_sfixed_a(-0.02505354955792427)),(to_sfixed_a(-0.0059943851083517075)),(to_sfixed_a(5.429066368378699e-05)),(to_sfixed_a(2.555697392381262e-05)),(to_sfixed_a(-0.00010956451296806335)),(to_sfixed_a(0.00018976135470438749)),(to_sfixed_a(0.00024878946715034544)),(to_sfixed_a(1.3095447002342553e-06)),(to_sfixed_a(0.0057904478162527084)),(to_sfixed_a(0.0338442400097847)),(to_sfixed_a(-0.07457667589187622)),(to_sfixed_a(-0.09627904742956161)),(to_sfixed_a(0.20802132785320282)),(to_sfixed_a(0.22331024706363678)),(to_sfixed_a(0.11651966720819473)),(to_sfixed_a(-0.022246617823839188)),(to_sfixed_a(-0.14061859250068665)),(to_sfixed_a(0.16144488751888275)),(to_sfixed_a(0.06920226663351059)),(to_sfixed_a(0.028637384995818138)),(to_sfixed_a(-0.4597623646259308)),(to_sfixed_a(-0.1450687050819397)),(to_sfixed_a(-0.0764351636171341)),(to_sfixed_a(-0.12146110832691193)),(to_sfixed_a(-0.1175616905093193)),(to_sfixed_a(-0.002066462766379118)),(to_sfixed_a(0.07361232489347458)),(to_sfixed_a(-0.12268023937940598)),(to_sfixed_a(-0.08367535471916199)),(to_sfixed_a(0.07327312231063843)),(to_sfixed_a(0.00012231980508659035)),(to_sfixed_a(0.00018200477643404156)),(to_sfixed_a(-1.4782847756578121e-05)),(to_sfixed_a(3.930210368707776e-05)),(to_sfixed_a(-0.00014354093582369387)),(to_sfixed_a(0.00019818372675217688)),(to_sfixed_a(-0.0007252951618283987)),(to_sfixed_a(-0.05670234188437462)),(to_sfixed_a(0.013288356363773346)),(to_sfixed_a(0.08935817331075668)),(to_sfixed_a(-0.03658558428287506)),(to_sfixed_a(0.06083736941218376)),(to_sfixed_a(-0.1153487041592598)),(to_sfixed_a(-0.01339772529900074)),(to_sfixed_a(-0.27615639567375183)),(to_sfixed_a(0.00046439841389656067)),(to_sfixed_a(-0.08581564575433731)),(to_sfixed_a(-0.03033786080777645)),(to_sfixed_a(-0.00776295643299818)),(to_sfixed_a(0.07100845873355865)),(to_sfixed_a(-0.1525123417377472)),(to_sfixed_a(-0.016392456367611885)),(to_sfixed_a(-0.03951917216181755)),(to_sfixed_a(-0.029815305024385452)),(to_sfixed_a(0.17030908167362213)),(to_sfixed_a(-0.01877477392554283)),(to_sfixed_a(-0.0065632350742816925)),(to_sfixed_a(8.626408089185134e-05)),(to_sfixed_a(-0.00012153737770859152)),(to_sfixed_a(0.00011107634054496884)),(to_sfixed_a(-0.0002229135570814833)),(to_sfixed_a(0.00016095205501187593)),(to_sfixed_a(0.00016002310439944267)),(to_sfixed_a(0.0002344518870813772)),(to_sfixed_a(-0.010553708299994469)),(to_sfixed_a(0.02602844126522541)),(to_sfixed_a(0.09492171555757523)),(to_sfixed_a(0.06518951803445816)),(to_sfixed_a(0.04768291488289833)),(to_sfixed_a(0.1657814234495163)),(to_sfixed_a(0.2171633094549179)),(to_sfixed_a(-0.00159633404109627)),(to_sfixed_a(-0.15103952586650848)),(to_sfixed_a(0.11455602943897247)),(to_sfixed_a(0.07404616475105286)),(to_sfixed_a(-0.1558917611837387)),(to_sfixed_a(-0.18771901726722717)),(to_sfixed_a(0.03894402086734772)),(to_sfixed_a(-0.03650370240211487)),(to_sfixed_a(0.0755511224269867)),(to_sfixed_a(0.051699817180633545)),(to_sfixed_a(-0.05742698162794113)),(to_sfixed_a(-0.0088883051648736)),(to_sfixed_a(0.15350298583507538)),(to_sfixed_a(0.051326051354408264)),(to_sfixed_a(-0.01840570569038391)),(to_sfixed_a(0.00021539966110140085)),(to_sfixed_a(-0.00026666276971809566)),(to_sfixed_a(-0.00020393339218571782)),(to_sfixed_a(8.340071508428082e-05)),(to_sfixed_a(-0.00016860202595125884)),(to_sfixed_a(-0.03169861063361168)),(to_sfixed_a(0.06792168319225311)),(to_sfixed_a(0.061084046959877014)),(to_sfixed_a(0.07803920656442642)),(to_sfixed_a(-0.09098010510206223)),(to_sfixed_a(-0.004031778313219547)),(to_sfixed_a(0.10575473308563232)),(to_sfixed_a(0.030562834814190865)),(to_sfixed_a(0.07396964728832245)),(to_sfixed_a(0.09626869112253189)),(to_sfixed_a(-0.12837441265583038)),(to_sfixed_a(-0.14254365861415863)),(to_sfixed_a(-0.10101769119501114)),(to_sfixed_a(0.16724088788032532)),(to_sfixed_a(0.15112313628196716)),(to_sfixed_a(-0.1495646983385086)),(to_sfixed_a(-0.09760576486587524)),(to_sfixed_a(-0.14821180701255798)),(to_sfixed_a(-0.061352167278528214)),(to_sfixed_a(-0.2142803817987442)),(to_sfixed_a(0.05526040866971016)),(to_sfixed_a(-0.02268979884684086)),(to_sfixed_a(-0.00013669395411852747)),(to_sfixed_a(2.040213621512521e-05)),(to_sfixed_a(1.0832871339516714e-05)),(to_sfixed_a(0.00011738756438717246)),(to_sfixed_a(2.1874595404369757e-05)),(to_sfixed_a(1.918507769005373e-05)),(to_sfixed_a(4.756358976010233e-05)),(to_sfixed_a(-0.09337735176086426)),(to_sfixed_a(0.04056740179657936)),(to_sfixed_a(0.07163326442241669)),(to_sfixed_a(-0.08272732049226761)),(to_sfixed_a(0.03354959189891815)),(to_sfixed_a(0.11372610181570053)),(to_sfixed_a(-0.16265101730823517)),(to_sfixed_a(-0.14765988290309906)),(to_sfixed_a(0.15044768154621124)),(to_sfixed_a(0.30868253111839294)),(to_sfixed_a(-0.1372194141149521)),(to_sfixed_a(0.05055040493607521)),(to_sfixed_a(-0.11654053628444672)),(to_sfixed_a(-0.01458723470568657)),(to_sfixed_a(0.13578826189041138)),(to_sfixed_a(0.15035684406757355)),(to_sfixed_a(0.15102308988571167)),(to_sfixed_a(-0.11355002224445343)),(to_sfixed_a(0.014030421152710915)),(to_sfixed_a(-0.01235441118478775)),(to_sfixed_a(-0.1547495275735855)),(to_sfixed_a(-0.00017481736722402275)),(to_sfixed_a(0.0001878371404018253)),(to_sfixed_a(-0.0001274446549359709)),(to_sfixed_a(-0.0004415680014062673)),(to_sfixed_a(7.549837027909234e-05)),(to_sfixed_a(0.00011589863424887881)),(to_sfixed_a(-0.0002648905210662633)),(to_sfixed_a(0.02089528925716877)),(to_sfixed_a(0.022796090692281723)),(to_sfixed_a(0.11460471898317337)),(to_sfixed_a(0.06150548905134201)),(to_sfixed_a(0.2165834605693817)),(to_sfixed_a(-0.1518218219280243)),(to_sfixed_a(-0.00017208440112881362)),(to_sfixed_a(-0.047265633940696716)),(to_sfixed_a(-0.02093140408396721)),(to_sfixed_a(0.470389187335968)),(to_sfixed_a(-0.11864116787910461)),(to_sfixed_a(0.04882889986038208)),(to_sfixed_a(-0.16392821073532104)),(to_sfixed_a(0.05374367535114288)),(to_sfixed_a(0.0318443737924099)),(to_sfixed_a(-0.05301814526319504)),(to_sfixed_a(-0.02093994803726673)),(to_sfixed_a(-0.08838430047035217)),(to_sfixed_a(-0.02927263081073761)),(to_sfixed_a(-0.03702929615974426)),(to_sfixed_a(0.042851775884628296)),(to_sfixed_a(0.0007960947696119547)),(to_sfixed_a(0.000624359177891165)),(to_sfixed_a(0.00035679011489264667)),(to_sfixed_a(-0.00022827716020401567)),(to_sfixed_a(-1.3133984793967102e-05)),(to_sfixed_a(-0.00031442393083125353)),(to_sfixed_a(-5.4410429584095255e-06)),(to_sfixed_a(-0.0005710511468350887)),(to_sfixed_a(-0.2072313129901886)),(to_sfixed_a(-0.10011883080005646)),(to_sfixed_a(0.1381145864725113)),(to_sfixed_a(-0.1325111836194992)),(to_sfixed_a(-0.38063162565231323)),(to_sfixed_a(0.11711133271455765)),(to_sfixed_a(0.0241530928760767)),(to_sfixed_a(-0.12622250616550446)),(to_sfixed_a(0.09092655032873154)),(to_sfixed_a(-0.47171419858932495)),(to_sfixed_a(0.09401512891054153)),(to_sfixed_a(0.10266885906457901)),(to_sfixed_a(0.1286969631910324)),(to_sfixed_a(-0.009618307463824749)),(to_sfixed_a(0.05553469434380531)),(to_sfixed_a(-0.025064408779144287)),(to_sfixed_a(0.15575635433197021)),(to_sfixed_a(0.12887151539325714)),(to_sfixed_a(0.27928152680397034)),(to_sfixed_a(0.013180899433791637)),(to_sfixed_a(0.0002719186304602772)),(to_sfixed_a(-0.00017100537661463022)),(to_sfixed_a(1.0516911970626097e-05)),(to_sfixed_a(5.5829128541518e-05)),(to_sfixed_a(-3.232923972973367e-06)),(to_sfixed_a(0.00025914813159033656)),(to_sfixed_a(-0.00012352908379398286)),(to_sfixed_a(0.017562810331583023)),(to_sfixed_a(-0.047477565705776215)),(to_sfixed_a(-0.00546477735042572)),(to_sfixed_a(-0.016454575583338737)),(to_sfixed_a(-0.16022007167339325)),(to_sfixed_a(0.004102595616132021)),(to_sfixed_a(-0.03943076729774475)),(to_sfixed_a(-0.02617098204791546)),(to_sfixed_a(0.0307554192841053)),(to_sfixed_a(-0.3416389524936676)),(to_sfixed_a(-0.14278864860534668)),(to_sfixed_a(-0.09910870343446732)),(to_sfixed_a(-0.00717378593981266)),(to_sfixed_a(0.10086967796087265)),(to_sfixed_a(0.041518718004226685)),(to_sfixed_a(0.03412879630923271)),(to_sfixed_a(-0.0331602580845356)),(to_sfixed_a(-0.09500216692686081)),(to_sfixed_a(0.025955766439437866)),(to_sfixed_a(0.1369408518075943)),(to_sfixed_a(0.14379577338695526)),(to_sfixed_a(0.0003685190458782017)),(to_sfixed_a(0.00024945830227807164)),(to_sfixed_a(-0.00012640828208532184)),(to_sfixed_a(0.000213250721571967)),(to_sfixed_a(-0.0001985821727430448)),(to_sfixed_a(-0.0002024487912422046)),(to_sfixed_a(0.00019966342370025814)),(to_sfixed_a(0.04225275665521622)),(to_sfixed_a(0.04719846695661545)),(to_sfixed_a(0.12827429175376892)),(to_sfixed_a(-0.029149705544114113)),(to_sfixed_a(-0.06153135374188423)),(to_sfixed_a(-0.05421239882707596)),(to_sfixed_a(0.08024347573518753)),(to_sfixed_a(0.29926466941833496)),(to_sfixed_a(-0.09335380792617798)),(to_sfixed_a(-0.03990792855620384)),(to_sfixed_a(-0.04759536311030388)),(to_sfixed_a(0.1357099860906601)),(to_sfixed_a(-0.007312118075788021)),(to_sfixed_a(-0.05445511266589165)),(to_sfixed_a(-0.17799267172813416)),(to_sfixed_a(-0.21613530814647675)),(to_sfixed_a(-0.13105668127536774)),(to_sfixed_a(0.06578356772661209)),(to_sfixed_a(-0.0855443924665451)),(to_sfixed_a(-0.004069230053573847)),(to_sfixed_a(0.09488257765769958)),(to_sfixed_a(-0.012650753371417522)),(to_sfixed_a(2.984627462865319e-05)),(to_sfixed_a(-8.599031571066007e-05)),(to_sfixed_a(0.00011014730989700183)),(to_sfixed_a(-0.00017679658776614815)),(to_sfixed_a(0.0006384681328199804)),(to_sfixed_a(0.0005968979676254094)),(to_sfixed_a(0.034064121544361115)),(to_sfixed_a(0.0928850769996643)),(to_sfixed_a(-0.03155157342553139)),(to_sfixed_a(0.32037773728370667)),(to_sfixed_a(-0.10012207180261612)),(to_sfixed_a(-0.179775670170784)),(to_sfixed_a(0.144120454788208)),(to_sfixed_a(-0.3008531332015991)),(to_sfixed_a(0.09739670902490616)),(to_sfixed_a(-0.12781335413455963)),(to_sfixed_a(-0.29837578535079956)),(to_sfixed_a(-0.19905798137187958)),(to_sfixed_a(-0.17431576550006866)),(to_sfixed_a(0.08020913600921631)),(to_sfixed_a(-0.2334292232990265)),(to_sfixed_a(-0.43918105959892273)),(to_sfixed_a(-0.1733304262161255)),(to_sfixed_a(0.08238445222377777)),(to_sfixed_a(0.23615007102489471)),(to_sfixed_a(0.008689300157129765)),(to_sfixed_a(6.465818296419457e-05)),(to_sfixed_a(3.972254489781335e-05)),(to_sfixed_a(-4.226947930874303e-05)),(to_sfixed_a(-0.00017611625662539154)),(to_sfixed_a(0.0004968621069565415)),(to_sfixed_a(-9.023796155815944e-05)),(to_sfixed_a(-0.00010421157639939338)),(to_sfixed_a(0.012780360877513885)),(to_sfixed_a(0.144815132021904)),(to_sfixed_a(0.04143647477030754)),(to_sfixed_a(0.09637759625911713)),(to_sfixed_a(0.22010886669158936)),(to_sfixed_a(0.057703908532857895)),(to_sfixed_a(-0.3471035659313202)),(to_sfixed_a(-0.09691240638494492)),(to_sfixed_a(-0.14938554167747498)),(to_sfixed_a(0.18093818426132202)),(to_sfixed_a(-0.11911381036043167)),(to_sfixed_a(-0.23104047775268555)),(to_sfixed_a(0.08100878447294235)),(to_sfixed_a(0.269060879945755)),(to_sfixed_a(-0.02759772539138794)),(to_sfixed_a(-0.19752711057662964)),(to_sfixed_a(-0.22711844742298126)),(to_sfixed_a(-0.07538950443267822)),(to_sfixed_a(0.08094379305839539)),(to_sfixed_a(-0.1056891456246376)),(to_sfixed_a(-0.021490657702088356)),(to_sfixed_a(0.008191976696252823)),(to_sfixed_a(0.0001827729429351166)),(to_sfixed_a(-0.0003262547543272376)),(to_sfixed_a(-0.0003596260503400117)),(to_sfixed_a(-0.00010247050522593781)),(to_sfixed_a(-0.00013352074893191457)),(to_sfixed_a(0.00010573495092103258)),(to_sfixed_a(0.07736217230558395)),(to_sfixed_a(-0.0026038577780127525)),(to_sfixed_a(0.05121344327926636)),(to_sfixed_a(-0.03101346269249916)),(to_sfixed_a(-0.0002366645639995113)),(to_sfixed_a(0.03435685858130455)),(to_sfixed_a(-0.16440653800964355)),(to_sfixed_a(-0.14281044900417328)),(to_sfixed_a(0.023744385689496994)),(to_sfixed_a(0.055639516562223434)),(to_sfixed_a(-0.12015572190284729)),(to_sfixed_a(-0.24640712141990662)),(to_sfixed_a(-0.26736047863960266)),(to_sfixed_a(-0.11122220009565353)),(to_sfixed_a(0.058916591107845306)),(to_sfixed_a(0.02044004015624523)),(to_sfixed_a(0.09868761897087097)),(to_sfixed_a(0.08566023409366608)),(to_sfixed_a(0.04503311961889267)),(to_sfixed_a(0.030257603153586388)),(to_sfixed_a(0.09492176026105881)),(to_sfixed_a(-1.562076977279503e-05)),(to_sfixed_a(-3.2063635444501415e-05)),(to_sfixed_a(0.0001658085238886997)),(to_sfixed_a(-4.1983905248343945e-05)),(to_sfixed_a(0.0001819436438381672)),(to_sfixed_a(-0.00024130685778800398)),(to_sfixed_a(3.082347757299431e-05)),(to_sfixed_a(9.916789167618845e-06)),(to_sfixed_a(0.05790366977453232)),(to_sfixed_a(0.004942577797919512)),(to_sfixed_a(0.008425166830420494)),(to_sfixed_a(0.24725188314914703)),(to_sfixed_a(-0.18168610334396362)),(to_sfixed_a(-0.016056498512625694)),(to_sfixed_a(-0.048449207097291946)),(to_sfixed_a(0.01634281314909458)),(to_sfixed_a(0.10532398521900177)),(to_sfixed_a(-0.11391294002532959)),(to_sfixed_a(0.02065260335803032)),(to_sfixed_a(0.009934481233358383)),(to_sfixed_a(-0.08229481428861618)),(to_sfixed_a(0.1148582324385643)),(to_sfixed_a(-0.18955323100090027)),(to_sfixed_a(-0.1509300321340561)),(to_sfixed_a(-0.15721625089645386)),(to_sfixed_a(0.13582751154899597)),(to_sfixed_a(-0.22825098037719727)),(to_sfixed_a(-0.15593458712100983)),(to_sfixed_a(0.021038323640823364)),(to_sfixed_a(-5.157292616786435e-05)),(to_sfixed_a(-4.972638635081239e-05)),(to_sfixed_a(-5.1829309086315334e-05)),(to_sfixed_a(6.987567758187652e-05)),(to_sfixed_a(0.0003365794545970857)),(to_sfixed_a(-9.18037912924774e-05)),(to_sfixed_a(9.527585643809289e-05)),(to_sfixed_a(0.028957147151231766)),(to_sfixed_a(0.00013908298569731414)),(to_sfixed_a(-0.12483326345682144)),(to_sfixed_a(0.15707668662071228)),(to_sfixed_a(-0.057645734399557114)),(to_sfixed_a(-0.1247016191482544)),(to_sfixed_a(-0.1217479258775711)),(to_sfixed_a(0.03094884194433689)),(to_sfixed_a(-0.12451212853193283)),(to_sfixed_a(-0.3006700277328491)),(to_sfixed_a(0.001978556625545025)),(to_sfixed_a(-0.06518350541591644)),(to_sfixed_a(0.08698909729719162)),(to_sfixed_a(0.1696780025959015)),(to_sfixed_a(-0.12200365215539932)),(to_sfixed_a(-0.019991468638181686)),(to_sfixed_a(0.21282006800174713)),(to_sfixed_a(0.10486137121915817)),(to_sfixed_a(0.348757266998291)),(to_sfixed_a(-0.0005465284339152277)),(to_sfixed_a(0.021448493003845215)),(to_sfixed_a(2.1120695237186737e-05)),(to_sfixed_a(5.6056065659504384e-05)),(to_sfixed_a(-0.00015660005738027394)),(to_sfixed_a(0.00018200595513917506)),(to_sfixed_a(-0.00020207725174259394)),(to_sfixed_a(3.636549536167877e-06)),(to_sfixed_a(-5.812084964418318e-06)),(to_sfixed_a(-0.00022432625701185316)),(to_sfixed_a(-0.07002268731594086)),(to_sfixed_a(-0.15149106085300446)),(to_sfixed_a(-0.08293747901916504)),(to_sfixed_a(0.12027843296527863)),(to_sfixed_a(0.010537040419876575)),(to_sfixed_a(-0.25051629543304443)),(to_sfixed_a(0.043897707015275955)),(to_sfixed_a(-0.024169402197003365)),(to_sfixed_a(-0.025708744302392006)),(to_sfixed_a(0.005914923269301653)),(to_sfixed_a(-0.04572217911481857)),(to_sfixed_a(-0.1584823876619339)),(to_sfixed_a(-0.009422963485121727)),(to_sfixed_a(-0.18979261815547943)),(to_sfixed_a(-0.10255863517522812)),(to_sfixed_a(0.021959958598017693)),(to_sfixed_a(-0.013242008164525032)),(to_sfixed_a(-0.023013757541775703)),(to_sfixed_a(-0.0024909251369535923)),(to_sfixed_a(9.359773684991524e-05)),(to_sfixed_a(-4.179256939096376e-05)),(to_sfixed_a(-0.00017290280084125698)),(to_sfixed_a(0.00012335117207840085)),(to_sfixed_a(0.00012982331099919975)),(to_sfixed_a(-7.57697198423557e-05)),(to_sfixed_a(-0.00019390825764276087)),(to_sfixed_a(-3.364944495842792e-05)),(to_sfixed_a(-6.30793219897896e-05)),(to_sfixed_a(-0.029495511204004288)),(to_sfixed_a(0.09244713187217712)),(to_sfixed_a(-0.010347392410039902)),(to_sfixed_a(-0.17068536579608917)),(to_sfixed_a(-0.0024239381309598684)),(to_sfixed_a(0.05877894163131714)),(to_sfixed_a(0.11001550406217575)),(to_sfixed_a(-0.12919482588768005)),(to_sfixed_a(0.042361751198768616)),(to_sfixed_a(0.17441056668758392)),(to_sfixed_a(0.0329921580851078)),(to_sfixed_a(-0.0876849815249443)),(to_sfixed_a(-0.3074156939983368)),(to_sfixed_a(0.009901588782668114)),(to_sfixed_a(-0.04159209504723549)),(to_sfixed_a(-0.07430718839168549)),(to_sfixed_a(0.1340421438217163)),(to_sfixed_a(-0.007865720428526402)),(to_sfixed_a(0.10975135117769241)),(to_sfixed_a(7.593585178256035e-05)),(to_sfixed_a(5.442845213110559e-05)),(to_sfixed_a(0.00015526937204413116)),(to_sfixed_a(-0.00026320110191591084)),(to_sfixed_a(0.0002979027049150318)),(to_sfixed_a(-3.759237006306648e-05)),(to_sfixed_a(-6.118362944107503e-05)),(to_sfixed_a(2.3534701540484093e-05)),(to_sfixed_a(-0.011577471159398556)),(to_sfixed_a(0.03407776355743408)),(to_sfixed_a(-0.048423729836940765)),(to_sfixed_a(0.06563232094049454)),(to_sfixed_a(0.13786709308624268)),(to_sfixed_a(0.0019461262272670865)),(to_sfixed_a(0.05389423668384552)),(to_sfixed_a(-0.020264126360416412)),(to_sfixed_a(-0.08478625863790512)),(to_sfixed_a(0.015290710143744946)),(to_sfixed_a(-0.011502218432724476)),(to_sfixed_a(-0.03470984846353531)),(to_sfixed_a(-0.11035323888063431)),(to_sfixed_a(0.0972815752029419)),(to_sfixed_a(-0.02123936451971531)),(to_sfixed_a(0.043152716010808945)),(to_sfixed_a(-0.012827766127884388)),(to_sfixed_a(0.10422168672084808)),(to_sfixed_a(0.049246691167354584)),(to_sfixed_a(-0.00324833020567894)),(to_sfixed_a(-7.779573206789792e-05)),(to_sfixed_a(-7.012178684817627e-05)),(to_sfixed_a(-6.999916513450444e-05)),(to_sfixed_a(-0.00025290960911661386)),(to_sfixed_a(-1.7877402569865808e-05)),(to_sfixed_a(-8.338969200849533e-05)),(to_sfixed_a(-0.00020583107834681869)),(to_sfixed_a(-0.0001284525787923485)),(to_sfixed_a(-2.4140301320585422e-05)),(to_sfixed_a(-0.0014958492247387767)),(to_sfixed_a(-0.02828865870833397)),(to_sfixed_a(-0.05215238779783249)),(to_sfixed_a(-0.16840173304080963)),(to_sfixed_a(-0.012633557431399822)),(to_sfixed_a(0.10622277110815048)),(to_sfixed_a(0.036666687577962875)),(to_sfixed_a(0.17908114194869995)),(to_sfixed_a(0.0052010295912623405)),(to_sfixed_a(-0.08528666198253632)),(to_sfixed_a(-0.15040266513824463)),(to_sfixed_a(0.16611257195472717)),(to_sfixed_a(-0.0021323177497833967)),(to_sfixed_a(-0.006891870405524969)),(to_sfixed_a(-0.0649334192276001)),(to_sfixed_a(-0.04259553179144859)),(to_sfixed_a(-0.0006233849562704563)),(to_sfixed_a(0.004011609125882387)),(to_sfixed_a(0.00420718127861619)),(to_sfixed_a(-8.317150786751881e-05)),(to_sfixed_a(-9.823772415984422e-05)),(to_sfixed_a(0.00035731293610297143)),(to_sfixed_a(0.0001931161095853895)),(to_sfixed_a(4.0358645492233336e-05)),(to_sfixed_a(0.00025702061248011887)),(to_sfixed_a(-7.452417048625648e-05)),(to_sfixed_a(-0.00013053606380708516)),(to_sfixed_a(-7.029085827525705e-05)),(to_sfixed_a(0.00025576187181286514)),(to_sfixed_a(0.00030387972947210073)),(to_sfixed_a(0.00012443153536878526)),(to_sfixed_a(0.0001050061036949046)),(to_sfixed_a(0.00045425863936543465)),(to_sfixed_a(0.0036203449126333)),(to_sfixed_a(-0.004953399766236544)),(to_sfixed_a(-0.0010828896192833781)),(to_sfixed_a(0.0055136894807219505)),(to_sfixed_a(-0.19214744865894318)),(to_sfixed_a(-0.013861503452062607)),(to_sfixed_a(-0.01580815576016903)),(to_sfixed_a(0.0033836751244962215)),(to_sfixed_a(-0.003690349403768778)),(to_sfixed_a(-0.012237644754350185)),(to_sfixed_a(-0.0029953133780509233)),(to_sfixed_a(0.00023795294691808522)),(to_sfixed_a(-0.0003176607715431601)),(to_sfixed_a(-6.853693048469722e-05)),(to_sfixed_a(0.00019721098942682147)),(to_sfixed_a(0.0001464368251617998)),(to_sfixed_a(0.0001284962781937793)),(to_sfixed_a(-0.00015345861902460456)),(to_sfixed_a(-8.886046998668462e-05)),(to_sfixed_a(-0.0003773548232857138)),(to_sfixed_a(1.2870068530901335e-05)),(to_sfixed_a(-0.00017120222037192434)),(to_sfixed_a(0.00041025527752935886)),(to_sfixed_a(-7.14433190296404e-05)),(to_sfixed_a(-0.0001050099017447792)),(to_sfixed_a(2.966802094306331e-05)),(to_sfixed_a(1.5440056813531555e-05)),(to_sfixed_a(9.646523540141061e-05)),(to_sfixed_a(-0.00017526741430629045)),(to_sfixed_a(0.00024104535987135023)),(to_sfixed_a(-0.00011617781274253502)),(to_sfixed_a(-0.00018190366972703487)),(to_sfixed_a(-0.00027563809999264777)),(to_sfixed_a(-0.00021165057842154056)),(to_sfixed_a(-0.00015719549264758825)),(to_sfixed_a(0.00018552850815467536)),(to_sfixed_a(-6.345423025777563e-05)),(to_sfixed_a(-6.68216816848144e-05)),(to_sfixed_a(-5.986582254990935e-05)),(to_sfixed_a(0.00011724401701940224)),(to_sfixed_a(7.98763066995889e-05)),(to_sfixed_a(-2.371428763581207e-06)),(to_sfixed_a(-0.00014794888556934893)),(to_sfixed_a(0.00010621990804793313)),(to_sfixed_a(0.0002129068598151207)),(to_sfixed_a(7.4148723797407e-05)));

    constant weight_n0_36 : sfixed_bus_array(784 downto 0) := ((to_sfixed_a(0.0)),(to_sfixed_a(0.00031424424378201365)),(to_sfixed_a(0.0002694699796847999)),(to_sfixed_a(-0.000265035341726616)),(to_sfixed_a(-8.486809383612126e-05)),(to_sfixed_a(0.00016792021051514894)),(to_sfixed_a(0.0003482877218630165)),(to_sfixed_a(3.4651922760531306e-05)),(to_sfixed_a(9.069435327546671e-05)),(to_sfixed_a(0.00012134513235650957)),(to_sfixed_a(-0.00021198503964114934)),(to_sfixed_a(-0.00018805508443620056)),(to_sfixed_a(8.329401680384763e-06)),(to_sfixed_a(0.00013671908527612686)),(to_sfixed_a(4.034560697618872e-05)),(to_sfixed_a(0.000137848561280407)),(to_sfixed_a(-0.0002227544755442068)),(to_sfixed_a(4.986625935998745e-05)),(to_sfixed_a(-4.844412615057081e-05)),(to_sfixed_a(0.0001010095511446707)),(to_sfixed_a(9.367070742882788e-05)),(to_sfixed_a(5.567608695855597e-06)),(to_sfixed_a(0.00011565551540115848)),(to_sfixed_a(-9.899590804707259e-05)),(to_sfixed_a(-1.0389187082182616e-05)),(to_sfixed_a(-4.886868191533722e-05)),(to_sfixed_a(0.0003041209129150957)),(to_sfixed_a(0.0003535287396516651)),(to_sfixed_a(0.00024848684552125633)),(to_sfixed_a(-0.00023467856226488948)),(to_sfixed_a(4.8436490033054724e-05)),(to_sfixed_a(-3.712849775183713e-06)),(to_sfixed_a(-0.00011363402882125229)),(to_sfixed_a(3.9301547076320276e-05)),(to_sfixed_a(2.4100885639199987e-05)),(to_sfixed_a(0.00017851762822829187)),(to_sfixed_a(-6.845731695648283e-05)),(to_sfixed_a(-5.4161126172402874e-05)),(to_sfixed_a(-0.0003522353363223374)),(to_sfixed_a(-8.448553126072511e-05)),(to_sfixed_a(2.713081266847439e-05)),(to_sfixed_a(4.87634570163209e-05)),(to_sfixed_a(-0.00011683047341648489)),(to_sfixed_a(-9.193293954012915e-05)),(to_sfixed_a(0.0003555284929461777)),(to_sfixed_a(0.00014595183893106878)),(to_sfixed_a(-0.00011370726133463904)),(to_sfixed_a(0.0001588845334481448)),(to_sfixed_a(0.00033973462996073067)),(to_sfixed_a(-0.0001309294457314536)),(to_sfixed_a(-6.822559225838631e-05)),(to_sfixed_a(7.837956218281761e-05)),(to_sfixed_a(0.00017846828268375248)),(to_sfixed_a(-7.837217708583921e-06)),(to_sfixed_a(-4.1691870137583464e-05)),(to_sfixed_a(0.00010093110176967457)),(to_sfixed_a(7.867241220083088e-05)),(to_sfixed_a(-9.889203647617251e-05)),(to_sfixed_a(0.0003290297172497958)),(to_sfixed_a(-6.72194582875818e-05)),(to_sfixed_a(0.00019423365301918238)),(to_sfixed_a(0.00011737523891497403)),(to_sfixed_a(-5.014779162593186e-05)),(to_sfixed_a(0.00010366425703978166)),(to_sfixed_a(0.00016034282452892512)),(to_sfixed_a(-4.1510840674163774e-05)),(to_sfixed_a(-0.0001820637844502926)),(to_sfixed_a(0.00017934902280103415)),(to_sfixed_a(-0.00014626915799453855)),(to_sfixed_a(0.00013234518701210618)),(to_sfixed_a(0.015846578404307365)),(to_sfixed_a(1.869006700871978e-05)),(to_sfixed_a(7.70308033679612e-05)),(to_sfixed_a(-0.0001445914531359449)),(to_sfixed_a(-8.656309364596382e-05)),(to_sfixed_a(-0.00020138302352279425)),(to_sfixed_a(-3.8958751247264445e-05)),(to_sfixed_a(0.00011567707406356931)),(to_sfixed_a(4.3929579987889156e-05)),(to_sfixed_a(0.00022307151812128723)),(to_sfixed_a(-1.2815149602829479e-05)),(to_sfixed_a(0.00010755992116173729)),(to_sfixed_a(2.4729630240472034e-05)),(to_sfixed_a(-3.082940384047106e-05)),(to_sfixed_a(-3.6524315873975866e-06)),(to_sfixed_a(-0.0001312699750997126)),(to_sfixed_a(0.00024372634652536362)),(to_sfixed_a(-0.0001285907783312723)),(to_sfixed_a(-0.00019211573817301542)),(to_sfixed_a(-8.649774827063084e-05)),(to_sfixed_a(9.962152398657054e-05)),(to_sfixed_a(3.130575714749284e-05)),(to_sfixed_a(-0.00010859522444661707)),(to_sfixed_a(0.030818412080407143)),(to_sfixed_a(-2.1668649424100295e-05)),(to_sfixed_a(0.035009823739528656)),(to_sfixed_a(0.015125089325010777)),(to_sfixed_a(0.04050071910023689)),(to_sfixed_a(-0.014347623102366924)),(to_sfixed_a(0.003564863232895732)),(to_sfixed_a(-0.022557226940989494)),(to_sfixed_a(-0.0024103608448058367)),(to_sfixed_a(0.049587756395339966)),(to_sfixed_a(0.0013451420236378908)),(to_sfixed_a(0.045414187014102936)),(to_sfixed_a(0.0073984949849545956)),(to_sfixed_a(0.01502532884478569)),(to_sfixed_a(0.00019090110436081886)),(to_sfixed_a(5.150130527908914e-05)),(to_sfixed_a(0.0001558007497806102)),(to_sfixed_a(9.177173342322931e-05)),(to_sfixed_a(8.593391248723492e-05)),(to_sfixed_a(6.229264545254409e-05)),(to_sfixed_a(0.0002922892745118588)),(to_sfixed_a(-7.588968583149835e-05)),(to_sfixed_a(-0.00013470888370648026)),(to_sfixed_a(-2.686236439330969e-05)),(to_sfixed_a(-9.565136133460328e-05)),(to_sfixed_a(8.242845069617033e-06)),(to_sfixed_a(0.0002503058931324631)),(to_sfixed_a(0.02043864130973816)),(to_sfixed_a(0.009730469435453415)),(to_sfixed_a(0.04163171350955963)),(to_sfixed_a(-0.17075400054454803)),(to_sfixed_a(-0.07687877118587494)),(to_sfixed_a(-0.033803343772888184)),(to_sfixed_a(-0.04796620085835457)),(to_sfixed_a(0.012631249614059925)),(to_sfixed_a(-0.004459437448531389)),(to_sfixed_a(0.0737391859292984)),(to_sfixed_a(0.1470678597688675)),(to_sfixed_a(0.028901556506752968)),(to_sfixed_a(-0.021148277446627617)),(to_sfixed_a(0.019142942503094673)),(to_sfixed_a(0.02730490453541279)),(to_sfixed_a(-0.009179343469440937)),(to_sfixed_a(-1.7383190424880013e-05)),(to_sfixed_a(0.0015480199363082647)),(to_sfixed_a(9.30005990085192e-05)),(to_sfixed_a(3.3029955375241116e-05)),(to_sfixed_a(0.0001270411885343492)),(to_sfixed_a(0.00021890809875912964)),(to_sfixed_a(-1.8087501302943565e-05)),(to_sfixed_a(-6.746016879333183e-05)),(to_sfixed_a(-0.00014105137961450964)),(to_sfixed_a(0.0007092932937666774)),(to_sfixed_a(0.02074708230793476)),(to_sfixed_a(-0.008028407581150532)),(to_sfixed_a(0.07616481184959412)),(to_sfixed_a(-0.023425012826919556)),(to_sfixed_a(0.0009552279370836914)),(to_sfixed_a(0.04288429394364357)),(to_sfixed_a(0.007065703626722097)),(to_sfixed_a(-0.03912671282887459)),(to_sfixed_a(-0.0781133696436882)),(to_sfixed_a(0.03765111044049263)),(to_sfixed_a(-0.034542448818683624)),(to_sfixed_a(-0.11093224585056305)),(to_sfixed_a(-0.018059011548757553)),(to_sfixed_a(-0.16250523924827576)),(to_sfixed_a(0.057628083974123)),(to_sfixed_a(-0.10741754621267319)),(to_sfixed_a(0.017158325761556625)),(to_sfixed_a(0.0037349797785282135)),(to_sfixed_a(0.03363623842597008)),(to_sfixed_a(-0.0018335197819396853)),(to_sfixed_a(-0.00014303289935924113)),(to_sfixed_a(-0.0001293532841373235)),(to_sfixed_a(0.0001658113906159997)),(to_sfixed_a(-3.673828132377821e-06)),(to_sfixed_a(-0.0001625986333237961)),(to_sfixed_a(-5.60849548492115e-05)),(to_sfixed_a(-0.00024805188877508044)),(to_sfixed_a(0.00028092769207432866)),(to_sfixed_a(0.023560646921396255)),(to_sfixed_a(-0.04752209410071373)),(to_sfixed_a(0.08131477981805801)),(to_sfixed_a(-0.0927279144525528)),(to_sfixed_a(0.08931402117013931)),(to_sfixed_a(-0.12611296772956848)),(to_sfixed_a(-0.13338764011859894)),(to_sfixed_a(-0.06544560194015503)),(to_sfixed_a(-0.11115392297506332)),(to_sfixed_a(0.06356688588857651)),(to_sfixed_a(-0.23137861490249634)),(to_sfixed_a(-0.027430908754467964)),(to_sfixed_a(0.008609906770288944)),(to_sfixed_a(0.04937785491347313)),(to_sfixed_a(0.13631509244441986)),(to_sfixed_a(0.06536249816417694)),(to_sfixed_a(-0.01130281575024128)),(to_sfixed_a(-0.0737706646323204)),(to_sfixed_a(0.0863923728466034)),(to_sfixed_a(-0.00655896682292223)),(to_sfixed_a(-0.007721601985394955)),(to_sfixed_a(-0.0026083264965564013)),(to_sfixed_a(0.00017931639740709215)),(to_sfixed_a(0.0001334047265117988)),(to_sfixed_a(1.622094259801088e-06)),(to_sfixed_a(-5.677935769199394e-05)),(to_sfixed_a(0.00017062283586710691)),(to_sfixed_a(-0.0001057116242009215)),(to_sfixed_a(-0.05304324999451637)),(to_sfixed_a(-0.029799124225974083)),(to_sfixed_a(0.0669381245970726)),(to_sfixed_a(0.09388559311628342)),(to_sfixed_a(-0.0626121386885643)),(to_sfixed_a(0.06319733709096909)),(to_sfixed_a(0.08612173050642014)),(to_sfixed_a(-0.09278891980648041)),(to_sfixed_a(-0.014801681973040104)),(to_sfixed_a(-0.22121308743953705)),(to_sfixed_a(-0.2033265233039856)),(to_sfixed_a(-0.2029494196176529)),(to_sfixed_a(-0.010171499103307724)),(to_sfixed_a(-0.11212141811847687)),(to_sfixed_a(-0.2011241614818573)),(to_sfixed_a(0.30278587341308594)),(to_sfixed_a(0.020996227860450745)),(to_sfixed_a(-0.0712059885263443)),(to_sfixed_a(-0.0004365210188552737)),(to_sfixed_a(0.015416920185089111)),(to_sfixed_a(0.005420309491455555)),(to_sfixed_a(-0.00013882074563298374)),(to_sfixed_a(6.508298247354105e-05)),(to_sfixed_a(7.723978342255577e-05)),(to_sfixed_a(0.00017295742873102427)),(to_sfixed_a(0.00011440987145761028)),(to_sfixed_a(0.00013424758799374104)),(to_sfixed_a(-0.0009553000563755631)),(to_sfixed_a(-0.01755272038280964)),(to_sfixed_a(-0.04961804300546646)),(to_sfixed_a(0.005295753013342619)),(to_sfixed_a(-0.16710767149925232)),(to_sfixed_a(0.07463064044713974)),(to_sfixed_a(-0.222280815243721)),(to_sfixed_a(0.06672609597444534)),(to_sfixed_a(-0.07864115387201309)),(to_sfixed_a(0.018781930208206177)),(to_sfixed_a(0.03877149522304535)),(to_sfixed_a(-0.05392494425177574)),(to_sfixed_a(-0.28850653767585754)),(to_sfixed_a(-0.10952064394950867)),(to_sfixed_a(-0.08778389543294907)),(to_sfixed_a(0.024909986183047295)),(to_sfixed_a(0.06940849125385284)),(to_sfixed_a(0.0005707707605324686)),(to_sfixed_a(0.33049508929252625)),(to_sfixed_a(0.30546215176582336)),(to_sfixed_a(-0.03191136196255684)),(to_sfixed_a(0.13444116711616516)),(to_sfixed_a(-0.00010185020073549822)),(to_sfixed_a(9.4386181444861e-05)),(to_sfixed_a(0.00013864434731658548)),(to_sfixed_a(-0.00013523046800401062)),(to_sfixed_a(5.578134732786566e-05)),(to_sfixed_a(-0.0002387118001934141)),(to_sfixed_a(0.002001167042180896)),(to_sfixed_a(0.08492323011159897)),(to_sfixed_a(0.009107181802392006)),(to_sfixed_a(-0.05505486950278282)),(to_sfixed_a(0.014870290644466877)),(to_sfixed_a(-0.04073600471019745)),(to_sfixed_a(-0.1086367517709732)),(to_sfixed_a(-0.18611331284046173)),(to_sfixed_a(-0.6185534596443176)),(to_sfixed_a(-0.08906549960374832)),(to_sfixed_a(0.03522461652755737)),(to_sfixed_a(0.13297387957572937)),(to_sfixed_a(-0.07946416735649109)),(to_sfixed_a(-0.11281570047140121)),(to_sfixed_a(-0.32684841752052307)),(to_sfixed_a(0.04183969274163246)),(to_sfixed_a(0.1045260801911354)),(to_sfixed_a(-0.1254514902830124)),(to_sfixed_a(0.09989741444587708)),(to_sfixed_a(0.21005956828594208)),(to_sfixed_a(0.11268991231918335)),(to_sfixed_a(-1.179227069769695e-06)),(to_sfixed_a(6.67685380904004e-05)),(to_sfixed_a(0.00017282327462453395)),(to_sfixed_a(0.00010696062236092985)),(to_sfixed_a(0.00013409717939794064)),(to_sfixed_a(-0.00023053477343637496)),(to_sfixed_a(0.00021050506620667875)),(to_sfixed_a(-0.005899271462112665)),(to_sfixed_a(-0.06031855195760727)),(to_sfixed_a(0.17161662876605988)),(to_sfixed_a(0.042796120047569275)),(to_sfixed_a(0.010669095441699028)),(to_sfixed_a(0.14755289256572723)),(to_sfixed_a(-0.03889171779155731)),(to_sfixed_a(0.05398840457201004)),(to_sfixed_a(-0.15015269815921783)),(to_sfixed_a(-0.11008233577013016)),(to_sfixed_a(0.24438294768333435)),(to_sfixed_a(-0.03655137121677399)),(to_sfixed_a(0.04820484295487404)),(to_sfixed_a(-0.1044662669301033)),(to_sfixed_a(-0.040474653244018555)),(to_sfixed_a(0.012828600592911243)),(to_sfixed_a(-0.3138067126274109)),(to_sfixed_a(0.10622821003198624)),(to_sfixed_a(-0.09256172180175781)),(to_sfixed_a(0.1279442310333252)),(to_sfixed_a(-0.039395302534103394)),(to_sfixed_a(-0.022299541160464287)),(to_sfixed_a(-8.887228614185005e-05)),(to_sfixed_a(-0.0001200874030473642)),(to_sfixed_a(0.00027176993899047375)),(to_sfixed_a(0.00014276975707616657)),(to_sfixed_a(0.0001103757822420448)),(to_sfixed_a(-0.019660264253616333)),(to_sfixed_a(0.020427586510777473)),(to_sfixed_a(0.008329185657203197)),(to_sfixed_a(0.1730598360300064)),(to_sfixed_a(0.2760225534439087)),(to_sfixed_a(0.22397641837596893)),(to_sfixed_a(0.27075982093811035)),(to_sfixed_a(0.02436225302517414)),(to_sfixed_a(0.10455435514450073)),(to_sfixed_a(-0.049584876745939255)),(to_sfixed_a(-0.10699085146188736)),(to_sfixed_a(-0.059420377016067505)),(to_sfixed_a(0.1311654895544052)),(to_sfixed_a(0.18079419434070587)),(to_sfixed_a(-0.11709260940551758)),(to_sfixed_a(0.1468966156244278)),(to_sfixed_a(-0.0017167243640869856)),(to_sfixed_a(-0.08911654353141785)),(to_sfixed_a(-0.11620558798313141)),(to_sfixed_a(-0.10987038165330887)),(to_sfixed_a(-0.014129852876067162)),(to_sfixed_a(-0.11890698224306107)),(to_sfixed_a(4.035948222735897e-05)),(to_sfixed_a(0.00013597364886663854)),(to_sfixed_a(6.270927406148985e-05)),(to_sfixed_a(8.440350939054042e-05)),(to_sfixed_a(0.00013829283125232905)),(to_sfixed_a(0.00031092195422388613)),(to_sfixed_a(-4.162755431025289e-06)),(to_sfixed_a(0.04419245943427086)),(to_sfixed_a(0.09450766444206238)),(to_sfixed_a(-0.17399539053440094)),(to_sfixed_a(0.07707252353429794)),(to_sfixed_a(-0.0760088637471199)),(to_sfixed_a(-0.047055140137672424)),(to_sfixed_a(-0.2629384696483612)),(to_sfixed_a(-0.18377496302127838)),(to_sfixed_a(0.3281697630882263)),(to_sfixed_a(0.09379842877388)),(to_sfixed_a(-0.01884714514017105)),(to_sfixed_a(-0.08629918843507767)),(to_sfixed_a(-0.27908894419670105)),(to_sfixed_a(-0.16476984322071075)),(to_sfixed_a(-0.08356615900993347)),(to_sfixed_a(-0.029391439631581306)),(to_sfixed_a(0.13373932242393494)),(to_sfixed_a(-0.16520603001117706)),(to_sfixed_a(-0.1611817181110382)),(to_sfixed_a(0.03100133314728737)),(to_sfixed_a(0.050047434866428375)),(to_sfixed_a(-3.7982823414495215e-05)),(to_sfixed_a(0.00020954498904757202)),(to_sfixed_a(-0.00018052443920169026)),(to_sfixed_a(0.0001384935312671587)),(to_sfixed_a(2.416666802673717e-06)),(to_sfixed_a(0.00030006689485162497)),(to_sfixed_a(0.0002969179768115282)),(to_sfixed_a(-0.008589588105678558)),(to_sfixed_a(-0.28623637557029724)),(to_sfixed_a(-0.33233901858329773)),(to_sfixed_a(-0.2920602560043335)),(to_sfixed_a(-0.008787398226559162)),(to_sfixed_a(0.07286802679300308)),(to_sfixed_a(0.17136071622371674)),(to_sfixed_a(-0.16571353375911713)),(to_sfixed_a(-0.041884198784828186)),(to_sfixed_a(0.1012805849313736)),(to_sfixed_a(0.025111904367804527)),(to_sfixed_a(0.07253863662481308)),(to_sfixed_a(0.1140674501657486)),(to_sfixed_a(-0.13371995091438293)),(to_sfixed_a(0.0723714828491211)),(to_sfixed_a(-0.10901133716106415)),(to_sfixed_a(-0.0714629590511322)),(to_sfixed_a(0.09521596133708954)),(to_sfixed_a(-0.09365516155958176)),(to_sfixed_a(-0.04256637394428253)),(to_sfixed_a(0.0380689799785614)),(to_sfixed_a(-0.0009940601885318756)),(to_sfixed_a(-9.48470551520586e-05)),(to_sfixed_a(-0.0002448020095471293)),(to_sfixed_a(-2.9621904104715213e-05)),(to_sfixed_a(0.00010960645886370912)),(to_sfixed_a(-3.721311441040598e-05)),(to_sfixed_a(0.0001071592778316699)),(to_sfixed_a(-0.001987676601856947)),(to_sfixed_a(0.10279069095849991)),(to_sfixed_a(-0.01666453666985035)),(to_sfixed_a(0.09258385747671127)),(to_sfixed_a(0.07932820171117783)),(to_sfixed_a(0.1900816261768341)),(to_sfixed_a(-0.08443696796894073)),(to_sfixed_a(-0.18833550810813904)),(to_sfixed_a(-0.15377672016620636)),(to_sfixed_a(-0.4285418391227722)),(to_sfixed_a(0.022250164300203323)),(to_sfixed_a(0.007005214691162109)),(to_sfixed_a(0.07645364105701447)),(to_sfixed_a(0.06132746487855911)),(to_sfixed_a(-0.12504693865776062)),(to_sfixed_a(0.09357050061225891)),(to_sfixed_a(-0.07273638248443604)),(to_sfixed_a(-0.1075301244854927)),(to_sfixed_a(-0.013628276064991951)),(to_sfixed_a(-0.09299767017364502)),(to_sfixed_a(-0.08022445440292358)),(to_sfixed_a(-0.0001697802363196388)),(to_sfixed_a(-6.640559149673209e-05)),(to_sfixed_a(-3.724032922036713e-06)),(to_sfixed_a(0.00020569664775393903)),(to_sfixed_a(4.616955266101286e-05)),(to_sfixed_a(1.9333627278683707e-05)),(to_sfixed_a(8.337569306604564e-05)),(to_sfixed_a(0.07671436667442322)),(to_sfixed_a(-0.039712850004434586)),(to_sfixed_a(-0.05506132170557976)),(to_sfixed_a(-0.19055385887622833)),(to_sfixed_a(0.09447810053825378)),(to_sfixed_a(-0.10790002346038818)),(to_sfixed_a(-0.10105305165052414)),(to_sfixed_a(0.03350131958723068)),(to_sfixed_a(-0.2865872085094452)),(to_sfixed_a(-0.26594963669776917)),(to_sfixed_a(0.18689344823360443)),(to_sfixed_a(0.021537823602557182)),(to_sfixed_a(0.05429196357727051)),(to_sfixed_a(-0.09289032220840454)),(to_sfixed_a(0.02940160036087036)),(to_sfixed_a(-0.07543246448040009)),(to_sfixed_a(0.17661042511463165)),(to_sfixed_a(0.10108614712953568)),(to_sfixed_a(0.021009132266044617)),(to_sfixed_a(-0.04313071072101593)),(to_sfixed_a(-0.00824267603456974)),(to_sfixed_a(-3.59198274964001e-05)),(to_sfixed_a(4.9436996050644666e-05)),(to_sfixed_a(0.00010012042184825987)),(to_sfixed_a(2.843487345671747e-05)),(to_sfixed_a(4.0487189835403115e-05)),(to_sfixed_a(-2.9843686206731945e-05)),(to_sfixed_a(-0.0012031844817101955)),(to_sfixed_a(-0.08197052031755447)),(to_sfixed_a(-0.16230209171772003)),(to_sfixed_a(-0.055466074496507645)),(to_sfixed_a(-0.05754358321428299)),(to_sfixed_a(0.06469656527042389)),(to_sfixed_a(0.09934751689434052)),(to_sfixed_a(0.12236618250608444)),(to_sfixed_a(-0.024517040699720383)),(to_sfixed_a(0.1257968246936798)),(to_sfixed_a(0.13469301164150238)),(to_sfixed_a(-0.029915794730186462)),(to_sfixed_a(0.046074677258729935)),(to_sfixed_a(0.14263589680194855)),(to_sfixed_a(-0.11531415581703186)),(to_sfixed_a(-0.24264484643936157)),(to_sfixed_a(0.03432602062821388)),(to_sfixed_a(0.31329163908958435)),(to_sfixed_a(0.22726194560527802)),(to_sfixed_a(0.09648571908473969)),(to_sfixed_a(-0.04343944787979126)),(to_sfixed_a(0.039401132613420486)),(to_sfixed_a(0.002484922530129552)),(to_sfixed_a(-3.9400369132636115e-05)),(to_sfixed_a(-4.218116737320088e-05)),(to_sfixed_a(5.812918607261963e-05)),(to_sfixed_a(-5.7858200307236984e-05)),(to_sfixed_a(-0.0008559307898394763)),(to_sfixed_a(-0.0016876491717994213)),(to_sfixed_a(-0.06515036523342133)),(to_sfixed_a(-0.06952890753746033)),(to_sfixed_a(0.00205044518224895)),(to_sfixed_a(0.02908722124993801)),(to_sfixed_a(0.2515430450439453)),(to_sfixed_a(0.14288823306560516)),(to_sfixed_a(0.0453847274184227)),(to_sfixed_a(-0.20956936478614807)),(to_sfixed_a(-0.08457377552986145)),(to_sfixed_a(0.02355487085878849)),(to_sfixed_a(0.1408759206533432)),(to_sfixed_a(0.034162137657403946)),(to_sfixed_a(-0.13546328246593475)),(to_sfixed_a(-0.31773799657821655)),(to_sfixed_a(0.05705868825316429)),(to_sfixed_a(0.038756195455789566)),(to_sfixed_a(-0.05571659654378891)),(to_sfixed_a(-0.1873294711112976)),(to_sfixed_a(-0.2867854833602905)),(to_sfixed_a(-0.02929459698498249)),(to_sfixed_a(-3.7415327824419364e-05)),(to_sfixed_a(8.524853001290467e-06)),(to_sfixed_a(0.00020071813196409494)),(to_sfixed_a(0.00014490280591417104)),(to_sfixed_a(2.944307379948441e-05)),(to_sfixed_a(-0.00019528152188286185)),(to_sfixed_a(6.567870150320232e-05)),(to_sfixed_a(0.0025400235317647457)),(to_sfixed_a(-0.006456168368458748)),(to_sfixed_a(0.017648490145802498)),(to_sfixed_a(-0.049996476620435715)),(to_sfixed_a(-0.13078488409519196)),(to_sfixed_a(-0.047439564019441605)),(to_sfixed_a(0.15932705998420715)),(to_sfixed_a(0.04618912190198898)),(to_sfixed_a(-0.06786841154098511)),(to_sfixed_a(-0.079686738550663)),(to_sfixed_a(-0.074649378657341)),(to_sfixed_a(0.016032053157687187)),(to_sfixed_a(-0.19238194823265076)),(to_sfixed_a(-0.04136090353131294)),(to_sfixed_a(0.25781795382499695)),(to_sfixed_a(0.08813707530498505)),(to_sfixed_a(0.25082698464393616)),(to_sfixed_a(0.0066245500929653645)),(to_sfixed_a(-0.10267887264490128)),(to_sfixed_a(0.02177899330854416)),(to_sfixed_a(0.050412699580192566)),(to_sfixed_a(-0.023907382041215897)),(to_sfixed_a(-0.00017651075904723257)),(to_sfixed_a(-6.243404641281813e-06)),(to_sfixed_a(-0.00020983275317121297)),(to_sfixed_a(-3.533784911269322e-05)),(to_sfixed_a(3.481415205897065e-06)),(to_sfixed_a(0.00021083014144096524)),(to_sfixed_a(0.008305365219712257)),(to_sfixed_a(-0.007221548818051815)),(to_sfixed_a(-0.13959656655788422)),(to_sfixed_a(-0.03709132969379425)),(to_sfixed_a(-0.15257921814918518)),(to_sfixed_a(-0.1275075078010559)),(to_sfixed_a(-0.12879911065101624)),(to_sfixed_a(0.11662749201059341)),(to_sfixed_a(0.10081692039966583)),(to_sfixed_a(-0.05436611548066139)),(to_sfixed_a(0.04087338596582413)),(to_sfixed_a(-0.2482473999261856)),(to_sfixed_a(0.025065764784812927)),(to_sfixed_a(0.04455975815653801)),(to_sfixed_a(-0.03643093258142471)),(to_sfixed_a(0.0351611003279686)),(to_sfixed_a(0.011541258543729782)),(to_sfixed_a(-0.2535924017429352)),(to_sfixed_a(-0.2030743509531021)),(to_sfixed_a(0.07196179777383804)),(to_sfixed_a(-0.15889780223369598)),(to_sfixed_a(-9.901681187329814e-05)),(to_sfixed_a(2.819359360728413e-05)),(to_sfixed_a(3.582973295124248e-05)),(to_sfixed_a(0.00032096379436552525)),(to_sfixed_a(-0.00017217331333085895)),(to_sfixed_a(5.436172796180472e-05)),(to_sfixed_a(-0.0002156387345166877)),(to_sfixed_a(4.166732196608791e-06)),(to_sfixed_a(0.034779492765665054)),(to_sfixed_a(0.04921070858836174)),(to_sfixed_a(-0.2123032659292221)),(to_sfixed_a(0.018472984433174133)),(to_sfixed_a(0.044072821736335754)),(to_sfixed_a(-0.06256858259439468)),(to_sfixed_a(-0.0012793118366971612)),(to_sfixed_a(0.3489546477794647)),(to_sfixed_a(0.06075180694460869)),(to_sfixed_a(-0.004493484739214182)),(to_sfixed_a(-0.2252625674009323)),(to_sfixed_a(-0.10987751930952072)),(to_sfixed_a(-0.005108116194605827)),(to_sfixed_a(-0.01984139159321785)),(to_sfixed_a(0.4026002287864685)),(to_sfixed_a(-0.24497947096824646)),(to_sfixed_a(-0.2075992077589035)),(to_sfixed_a(0.01289727259427309)),(to_sfixed_a(-0.06437888741493225)),(to_sfixed_a(-0.09606292843818665)),(to_sfixed_a(-0.04784626513719559)),(to_sfixed_a(0.00022431985416915268)),(to_sfixed_a(0.00021874844969715923)),(to_sfixed_a(-6.30518261459656e-05)),(to_sfixed_a(0.0001686378091108054)),(to_sfixed_a(3.9509595808340237e-05)),(to_sfixed_a(-0.00032608062610961497)),(to_sfixed_a(2.232629958598409e-05)),(to_sfixed_a(-0.08846824616193771)),(to_sfixed_a(-0.0015697136987000704)),(to_sfixed_a(-0.03112010471522808)),(to_sfixed_a(0.20414157211780548)),(to_sfixed_a(-0.0141939427703619)),(to_sfixed_a(0.08076047152280807)),(to_sfixed_a(0.015398778021335602)),(to_sfixed_a(0.07575934380292892)),(to_sfixed_a(0.04646960645914078)),(to_sfixed_a(0.08509595692157745)),(to_sfixed_a(-0.029774032533168793)),(to_sfixed_a(-0.10424510389566422)),(to_sfixed_a(-0.04999883472919464)),(to_sfixed_a(0.07954595237970352)),(to_sfixed_a(-0.021363340318202972)),(to_sfixed_a(-0.21617361903190613)),(to_sfixed_a(-0.2615976929664612)),(to_sfixed_a(-0.012325955554842949)),(to_sfixed_a(-0.06064538657665253)),(to_sfixed_a(0.000460107228718698)),(to_sfixed_a(0.08283963799476624)),(to_sfixed_a(-4.643779175239615e-05)),(to_sfixed_a(0.00011289336543995887)),(to_sfixed_a(0.00015507993521168828)),(to_sfixed_a(3.208002817700617e-05)),(to_sfixed_a(-7.862881466280669e-05)),(to_sfixed_a(4.8118334234459326e-05)),(to_sfixed_a(0.00018651795107871294)),(to_sfixed_a(-0.00026241305749863386)),(to_sfixed_a(0.030295029282569885)),(to_sfixed_a(0.08132651448249817)),(to_sfixed_a(-0.005566726438701153)),(to_sfixed_a(0.14002031087875366)),(to_sfixed_a(0.09122613817453384)),(to_sfixed_a(0.08528723567724228)),(to_sfixed_a(0.06888504326343536)),(to_sfixed_a(0.06078638136386871)),(to_sfixed_a(0.026209501549601555)),(to_sfixed_a(-0.07290918380022049)),(to_sfixed_a(-0.16868053376674652)),(to_sfixed_a(0.02014540694653988)),(to_sfixed_a(-0.15973082184791565)),(to_sfixed_a(-0.07166661322116852)),(to_sfixed_a(-0.23145881295204163)),(to_sfixed_a(0.06316483020782471)),(to_sfixed_a(0.005690003279596567)),(to_sfixed_a(0.10823506861925125)),(to_sfixed_a(-0.00047286663902923465)),(to_sfixed_a(1.3993870197737124e-05)),(to_sfixed_a(-0.00014925967843737453)),(to_sfixed_a(3.439943247940391e-05)),(to_sfixed_a(-0.00016501314530614763)),(to_sfixed_a(2.999956086569e-05)),(to_sfixed_a(0.0002584054309409112)),(to_sfixed_a(-6.316047074506059e-05)),(to_sfixed_a(-0.0002941639395430684)),(to_sfixed_a(-0.00018109005759470165)),(to_sfixed_a(0.021465463563799858)),(to_sfixed_a(-0.06775542348623276)),(to_sfixed_a(0.08716654032468796)),(to_sfixed_a(0.13616713881492615)),(to_sfixed_a(0.07787284255027771)),(to_sfixed_a(-0.020046377554535866)),(to_sfixed_a(-0.16439764201641083)),(to_sfixed_a(0.08015695959329605)),(to_sfixed_a(0.019333569332957268)),(to_sfixed_a(-0.16434946656227112)),(to_sfixed_a(-0.223136305809021)),(to_sfixed_a(-0.39373958110809326)),(to_sfixed_a(0.055130671709775925)),(to_sfixed_a(0.05015916749835014)),(to_sfixed_a(-0.10722585022449493)),(to_sfixed_a(-0.042538270354270935)),(to_sfixed_a(0.015593932941555977)),(to_sfixed_a(-0.007023069076240063)),(to_sfixed_a(0.021560154855251312)),(to_sfixed_a(-0.00019676813099067658)),(to_sfixed_a(-7.740101864328608e-05)),(to_sfixed_a(0.0001343186158919707)),(to_sfixed_a(0.00025402806932106614)),(to_sfixed_a(0.000128896368551068)),(to_sfixed_a(0.00015134969726204872)),(to_sfixed_a(-0.00019667491142172366)),(to_sfixed_a(0.00011758596519939601)),(to_sfixed_a(0.025150662288069725)),(to_sfixed_a(0.04479619115591049)),(to_sfixed_a(0.10487376898527145)),(to_sfixed_a(0.20264899730682373)),(to_sfixed_a(0.00712551036849618)),(to_sfixed_a(0.14702534675598145)),(to_sfixed_a(0.29742926359176636)),(to_sfixed_a(0.2133646160364151)),(to_sfixed_a(-0.020087607204914093)),(to_sfixed_a(0.022087113931775093)),(to_sfixed_a(0.07320687919855118)),(to_sfixed_a(-0.3142896890640259)),(to_sfixed_a(0.11573982983827591)),(to_sfixed_a(-0.018907396122813225)),(to_sfixed_a(0.0910559892654419)),(to_sfixed_a(0.14250941574573517)),(to_sfixed_a(-0.002447272650897503)),(to_sfixed_a(0.042918235063552856)),(to_sfixed_a(0.008847476914525032)),(to_sfixed_a(-0.00035842577926814556)),(to_sfixed_a(3.0716328183189034e-05)),(to_sfixed_a(-0.00013163259427528828)),(to_sfixed_a(-0.00012576371955219656)),(to_sfixed_a(-0.0002548191696405411)),(to_sfixed_a(7.037272735033184e-05)),(to_sfixed_a(-6.546684016939253e-05)),(to_sfixed_a(2.3438167772837915e-05)),(to_sfixed_a(-4.37917624367401e-05)),(to_sfixed_a(0.00011488056043162942)),(to_sfixed_a(-0.0601184256374836)),(to_sfixed_a(0.06339297443628311)),(to_sfixed_a(0.06316977739334106)),(to_sfixed_a(-0.011800582520663738)),(to_sfixed_a(0.02565780095756054)),(to_sfixed_a(0.11650180071592331)),(to_sfixed_a(0.16824041306972504)),(to_sfixed_a(-0.17383095622062683)),(to_sfixed_a(-0.16403962671756744)),(to_sfixed_a(0.01044321246445179)),(to_sfixed_a(0.039898861199617386)),(to_sfixed_a(0.2432948350906372)),(to_sfixed_a(-0.022722618654370308)),(to_sfixed_a(-0.002825530245900154)),(to_sfixed_a(0.024920091032981873)),(to_sfixed_a(0.0987178161740303)),(to_sfixed_a(0.0003241840749979019)),(to_sfixed_a(0.0042738099582493305)),(to_sfixed_a(0.0045082829892635345)),(to_sfixed_a(0.0002755149616859853)),(to_sfixed_a(0.0001728791103232652)),(to_sfixed_a(-0.0003080469905398786)),(to_sfixed_a(-7.993719191290438e-05)),(to_sfixed_a(0.00024336742353625596)),(to_sfixed_a(-0.00010091933654621243)),(to_sfixed_a(-0.0001600650284672156)),(to_sfixed_a(-0.00012906844494864345)),(to_sfixed_a(3.995216957264347e-06)),(to_sfixed_a(-0.0007056161994114518)),(to_sfixed_a(-0.0009981272742152214)),(to_sfixed_a(0.00010548056161496788)),(to_sfixed_a(-4.6717213990632445e-05)),(to_sfixed_a(-7.001517951721326e-05)),(to_sfixed_a(0.1011510118842125)),(to_sfixed_a(-0.001671159639954567)),(to_sfixed_a(-0.0007968945428729057)),(to_sfixed_a(0.06829197704792023)),(to_sfixed_a(0.007292653899639845)),(to_sfixed_a(-0.013617271557450294)),(to_sfixed_a(-0.08027315139770508)),(to_sfixed_a(0.07986258715391159)),(to_sfixed_a(0.09918459504842758)),(to_sfixed_a(-0.0036869405303150415)),(to_sfixed_a(0.000770356273278594)),(to_sfixed_a(-0.00010288838529959321)),(to_sfixed_a(-9.040503209689632e-05)),(to_sfixed_a(-6.9704897214251105e-06)),(to_sfixed_a(-4.350560266175307e-05)),(to_sfixed_a(5.481170228449628e-05)),(to_sfixed_a(-0.00015142980555538088)),(to_sfixed_a(0.00030370260355994105)),(to_sfixed_a(-0.000391979148844257)),(to_sfixed_a(-6.003363159834407e-05)),(to_sfixed_a(0.00022814670228399336)),(to_sfixed_a(-0.00032972119515761733)),(to_sfixed_a(-0.00034368489286862314)),(to_sfixed_a(0.00010933009616564959)),(to_sfixed_a(9.362814307678491e-05)),(to_sfixed_a(0.00013228601892478764)),(to_sfixed_a(-6.628158735111356e-05)),(to_sfixed_a(-0.0001586509752087295)),(to_sfixed_a(8.096050441963598e-05)),(to_sfixed_a(7.699763227719814e-05)),(to_sfixed_a(-0.0001445846282877028)),(to_sfixed_a(0.00012175209121778607)),(to_sfixed_a(-0.00017590635980013758)),(to_sfixed_a(0.00012997294834349304)),(to_sfixed_a(-9.569364920025691e-05)),(to_sfixed_a(-0.0001198393729282543)),(to_sfixed_a(5.5578333558514714e-05)),(to_sfixed_a(0.00010342238965677097)),(to_sfixed_a(6.970308731979458e-06)),(to_sfixed_a(8.206020720535889e-05)),(to_sfixed_a(-7.074181485222653e-05)),(to_sfixed_a(-0.00011835682380478829)),(to_sfixed_a(4.183677810942754e-05)),(to_sfixed_a(2.604131395855802e-06)),(to_sfixed_a(0.00014284589269664139)),(to_sfixed_a(0.0001067443226929754)));


    constant weight_n1_0 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.26857462525367737)),(to_sfixed_a(0.15818241238594055)),(to_sfixed_a(-0.09932118654251099)),(to_sfixed_a(0.05585562810301781)),(to_sfixed_a(-0.27512967586517334)),(to_sfixed_a(0.13638116419315338)),(to_sfixed_a(-0.09296657890081406)),(to_sfixed_a(0.37282323837280273)),(to_sfixed_a(-0.051479991525411606)),(to_sfixed_a(0.0160475242882967)),(to_sfixed_a(-0.09117770940065384)),(to_sfixed_a(0.05607093870639801)),(to_sfixed_a(-0.006856780033558607)),(to_sfixed_a(0.017905578017234802)),(to_sfixed_a(-0.13606004416942596)),(to_sfixed_a(0.08857106417417526)),(to_sfixed_a(0.021214909851551056)),(to_sfixed_a(-0.03554689139127731)),(to_sfixed_a(0.12546369433403015)),(to_sfixed_a(-0.034939348697662354)),(to_sfixed_a(0.017086323350667953)),(to_sfixed_a(-0.04089096188545227)),(to_sfixed_a(0.03259311616420746)),(to_sfixed_a(-0.050422560423612595)),(to_sfixed_a(0.02862045168876648)),(to_sfixed_a(-0.028437357395887375)),(to_sfixed_a(0.11800219863653183)),(to_sfixed_a(-0.10884242504835129)),(to_sfixed_a(0.027524899691343307)),(to_sfixed_a(-0.027564655989408493)),(to_sfixed_a(0.030370092019438744)),(to_sfixed_a(-0.031228313222527504)),(to_sfixed_a(0.07185275107622147)),(to_sfixed_a(-0.12782397866249084)),(to_sfixed_a(0.08902892470359802)),(to_sfixed_a(0.061225052922964096)),(to_sfixed_a(-0.13357798755168915)),(to_sfixed_a(0.09745524078607559)));

    constant weight_n1_1 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.11653158813714981)),(to_sfixed_a(-0.16737987101078033)),(to_sfixed_a(0.1952148973941803)),(to_sfixed_a(0.3540059030056)),(to_sfixed_a(0.09454912692308426)),(to_sfixed_a(-0.26575082540512085)),(to_sfixed_a(-0.14997558295726776)),(to_sfixed_a(0.13294170796871185)),(to_sfixed_a(-0.12724949419498444)),(to_sfixed_a(0.030200498178601265)),(to_sfixed_a(-0.014742099680006504)),(to_sfixed_a(0.08816825598478317)),(to_sfixed_a(-0.09772039204835892)),(to_sfixed_a(0.10576991736888885)),(to_sfixed_a(0.0485399067401886)),(to_sfixed_a(-0.012724384665489197)),(to_sfixed_a(0.01232899073511362)),(to_sfixed_a(0.06273873150348663)),(to_sfixed_a(0.13095198571681976)),(to_sfixed_a(0.1252007782459259)),(to_sfixed_a(-0.0389835424721241)),(to_sfixed_a(0.03918081894516945)),(to_sfixed_a(-0.07045861333608627)),(to_sfixed_a(-0.07181385904550552)),(to_sfixed_a(0.056487083435058594)),(to_sfixed_a(-0.018197134137153625)),(to_sfixed_a(0.01888197846710682)),(to_sfixed_a(-0.08307944238185883)),(to_sfixed_a(-0.0491032712161541)),(to_sfixed_a(-0.15943187475204468)),(to_sfixed_a(-0.019068164750933647)),(to_sfixed_a(0.014393425546586514)),(to_sfixed_a(0.1169649064540863)),(to_sfixed_a(-0.11605530232191086)),(to_sfixed_a(0.16043850779533386)),(to_sfixed_a(0.03865216299891472)),(to_sfixed_a(0.0975082591176033)),(to_sfixed_a(0.014351104386150837)));

    constant weight_n1_2 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.039211712777614594)),(to_sfixed_a(2.4149998353095725e-05)),(to_sfixed_a(-4.231023194734007e-05)),(to_sfixed_a(-1.185695145977661e-05)),(to_sfixed_a(-1.4452069081016816e-05)),(to_sfixed_a(-3.951803591917269e-05)),(to_sfixed_a(7.372170512098819e-05)),(to_sfixed_a(-7.3499772952345666e-06)),(to_sfixed_a(-3.990705863543553e-06)),(to_sfixed_a(2.3116277588997036e-05)),(to_sfixed_a(-2.346436849620659e-05)),(to_sfixed_a(-9.685069926490542e-06)),(to_sfixed_a(-7.106752309482545e-05)),(to_sfixed_a(-4.840418478124775e-05)),(to_sfixed_a(-1.4213788745109923e-05)),(to_sfixed_a(-1.4970097254263237e-05)),(to_sfixed_a(5.715493534808047e-05)),(to_sfixed_a(-2.844909431587439e-05)),(to_sfixed_a(-1.2832385436922777e-05)),(to_sfixed_a(-9.829067494138144e-06)),(to_sfixed_a(-9.57935208134586e-06)),(to_sfixed_a(-3.175942038069479e-05)),(to_sfixed_a(1.721599073789548e-05)),(to_sfixed_a(2.0218833014951088e-05)),(to_sfixed_a(-8.399247599299997e-05)),(to_sfixed_a(-2.2315662135952152e-05)),(to_sfixed_a(-5.894893911317922e-05)),(to_sfixed_a(-6.0945283621549606e-05)),(to_sfixed_a(-4.3846910557476804e-05)),(to_sfixed_a(6.356229278026149e-05)),(to_sfixed_a(3.9660830225329846e-05)),(to_sfixed_a(-7.071408617775887e-05)),(to_sfixed_a(-2.6008628992713057e-05)),(to_sfixed_a(-1.5890735085122287e-05)),(to_sfixed_a(6.496573041658849e-05)),(to_sfixed_a(-4.4153930502943695e-05)),(to_sfixed_a(5.595977199845947e-05)),(to_sfixed_a(8.240571332862601e-05)));

    constant weight_n1_3 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.3379265069961548)),(to_sfixed_a(0.16886776685714722)),(to_sfixed_a(0.14295214414596558)),(to_sfixed_a(-0.10420683771371841)),(to_sfixed_a(0.0981055349111557)),(to_sfixed_a(0.024965625256299973)),(to_sfixed_a(-0.0814669281244278)),(to_sfixed_a(0.038729432970285416)),(to_sfixed_a(-0.06920734792947769)),(to_sfixed_a(0.17118120193481445)),(to_sfixed_a(0.011932230554521084)),(to_sfixed_a(-0.011460971087217331)),(to_sfixed_a(0.02570553869009018)),(to_sfixed_a(0.00027774961199611425)),(to_sfixed_a(0.06925780326128006)),(to_sfixed_a(-0.006529553327709436)),(to_sfixed_a(0.01880149357020855)),(to_sfixed_a(0.08185700327157974)),(to_sfixed_a(-0.003691137069836259)),(to_sfixed_a(0.06619725376367569)),(to_sfixed_a(-0.013248084113001823)),(to_sfixed_a(-0.023897798731923103)),(to_sfixed_a(-0.026968074962496758)),(to_sfixed_a(0.044933341443538666)),(to_sfixed_a(0.03138574957847595)),(to_sfixed_a(-0.023528164252638817)),(to_sfixed_a(0.0906636044383049)),(to_sfixed_a(0.028517525643110275)),(to_sfixed_a(-0.05360987037420273)),(to_sfixed_a(-0.02265637181699276)),(to_sfixed_a(-0.010809159837663174)),(to_sfixed_a(0.010148060508072376)),(to_sfixed_a(0.03270250931382179)),(to_sfixed_a(-0.17746861279010773)),(to_sfixed_a(-0.0822485014796257)),(to_sfixed_a(0.020584480836987495)),(to_sfixed_a(-0.0035666662734001875)),(to_sfixed_a(0.04482071101665497)));

    constant weight_n1_4 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.11215491592884064)),(to_sfixed_a(3.8331174437189475e-05)),(to_sfixed_a(2.697216405067593e-05)),(to_sfixed_a(-5.037014852860011e-05)),(to_sfixed_a(7.1922281676961575e-06)),(to_sfixed_a(1.849016007327009e-05)),(to_sfixed_a(1.5477848137379624e-05)),(to_sfixed_a(-1.1789345080615021e-05)),(to_sfixed_a(-1.1727777746273205e-05)),(to_sfixed_a(1.0654444849933498e-05)),(to_sfixed_a(-3.258040305809118e-05)),(to_sfixed_a(-2.6578052711556666e-05)),(to_sfixed_a(-2.3767170205246657e-05)),(to_sfixed_a(-7.70648148318287e-06)),(to_sfixed_a(-2.1684249077225104e-05)),(to_sfixed_a(5.474382487591356e-05)),(to_sfixed_a(3.757014201255515e-05)),(to_sfixed_a(4.3609790623122535e-07)),(to_sfixed_a(-4.8048834287328646e-05)),(to_sfixed_a(-2.902816731875646e-06)),(to_sfixed_a(-3.7866549973841757e-05)),(to_sfixed_a(-2.624066110001877e-05)),(to_sfixed_a(7.463905831173179e-07)),(to_sfixed_a(4.0195867768488824e-05)),(to_sfixed_a(9.222715561918449e-06)),(to_sfixed_a(1.3247809874883387e-05)),(to_sfixed_a(-4.7853507567197084e-05)),(to_sfixed_a(-9.02125975699164e-05)),(to_sfixed_a(2.4754443074925803e-05)),(to_sfixed_a(3.2475480111315846e-05)),(to_sfixed_a(5.570216671912931e-05)),(to_sfixed_a(-7.17601869837381e-05)),(to_sfixed_a(-4.802000694326125e-05)),(to_sfixed_a(0.0001426732778782025)),(to_sfixed_a(2.9226728656794876e-05)),(to_sfixed_a(2.7689118724083528e-05)),(to_sfixed_a(-5.115023668622598e-05)),(to_sfixed_a(6.744180427631363e-05)));

    constant weight_n1_5 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.050697844475507736)),(to_sfixed_a(0.015035470016300678)),(to_sfixed_a(-0.007022355683147907)),(to_sfixed_a(0.0059525067918002605)),(to_sfixed_a(0.004136690869927406)),(to_sfixed_a(0.06668811291456223)),(to_sfixed_a(-0.004012113902717829)),(to_sfixed_a(0.031852614134550095)),(to_sfixed_a(-0.0020002599339932203)),(to_sfixed_a(-0.009257077239453793)),(to_sfixed_a(0.026583164930343628)),(to_sfixed_a(0.0009079622686840594)),(to_sfixed_a(0.01956120692193508)),(to_sfixed_a(0.01813969388604164)),(to_sfixed_a(0.006271607708185911)),(to_sfixed_a(-0.002843568567186594)),(to_sfixed_a(-0.013166356831789017)),(to_sfixed_a(-0.015075779519975185)),(to_sfixed_a(-0.006709179375320673)),(to_sfixed_a(-0.001612727646715939)),(to_sfixed_a(-0.0013017579913139343)),(to_sfixed_a(-0.020032577216625214)),(to_sfixed_a(0.058552175760269165)),(to_sfixed_a(-0.029722347855567932)),(to_sfixed_a(0.006953700911253691)),(to_sfixed_a(-0.010933692567050457)),(to_sfixed_a(-0.0035803159698843956)),(to_sfixed_a(-0.00796044897288084)),(to_sfixed_a(0.010197357274591923)),(to_sfixed_a(-0.02198655530810356)),(to_sfixed_a(-0.008931138552725315)),(to_sfixed_a(-0.013845750130712986)),(to_sfixed_a(-0.05660836026072502)),(to_sfixed_a(0.014847858808934689)),(to_sfixed_a(-0.08114135265350342)),(to_sfixed_a(-0.01505602803081274)),(to_sfixed_a(-0.01899748295545578)),(to_sfixed_a(-0.036082714796066284)));

    constant weight_n1_6 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.015744978561997414)),(to_sfixed_a(1.1420460396038834e-05)),(to_sfixed_a(6.359732196870027e-06)),(to_sfixed_a(-1.4991082935011946e-06)),(to_sfixed_a(-7.021556666586548e-05)),(to_sfixed_a(-3.2109048220263503e-07)),(to_sfixed_a(0.00010045590897789225)),(to_sfixed_a(-5.781998697784729e-05)),(to_sfixed_a(-6.2685016928298865e-06)),(to_sfixed_a(1.2368000170681626e-06)),(to_sfixed_a(-4.5137461711419746e-05)),(to_sfixed_a(-3.534622737788595e-05)),(to_sfixed_a(1.269530002900865e-05)),(to_sfixed_a(-4.819002060685307e-05)),(to_sfixed_a(7.034498412394896e-05)),(to_sfixed_a(1.521240938018309e-05)),(to_sfixed_a(1.0336617378925439e-05)),(to_sfixed_a(-2.102018697769381e-05)),(to_sfixed_a(-1.6076963902378338e-06)),(to_sfixed_a(-8.429053195868619e-06)),(to_sfixed_a(-3.8116215819172794e-06)),(to_sfixed_a(3.8080219383118674e-05)),(to_sfixed_a(-4.123781400267035e-05)),(to_sfixed_a(9.082672477234155e-05)),(to_sfixed_a(-7.065742101985961e-05)),(to_sfixed_a(-4.198877650196664e-05)),(to_sfixed_a(-2.6362376956967637e-05)),(to_sfixed_a(6.411064532585442e-05)),(to_sfixed_a(-5.405781848821789e-06)),(to_sfixed_a(2.9930761229479685e-05)),(to_sfixed_a(-0.0001303711615037173)),(to_sfixed_a(2.7766142011387274e-05)),(to_sfixed_a(0.00014115730300545692)),(to_sfixed_a(4.312702367315069e-05)),(to_sfixed_a(1.6441811467871048e-08)),(to_sfixed_a(0.00013068935368210077)),(to_sfixed_a(-9.98249597614631e-05)),(to_sfixed_a(-7.287285825441359e-06)));

    constant weight_n1_7 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.07947754859924316)),(to_sfixed_a(-3.9332720916718245e-05)),(to_sfixed_a(6.478033174062148e-05)),(to_sfixed_a(-1.42151620821096e-05)),(to_sfixed_a(-4.708571941591799e-05)),(to_sfixed_a(2.1217962057562545e-05)),(to_sfixed_a(-2.3111675545806065e-05)),(to_sfixed_a(4.419219840201549e-05)),(to_sfixed_a(3.0494502425426617e-06)),(to_sfixed_a(1.4397675840882584e-05)),(to_sfixed_a(-3.9267284591915086e-05)),(to_sfixed_a(-8.811485713522416e-06)),(to_sfixed_a(-5.3398201998788863e-05)),(to_sfixed_a(-5.9789326769532636e-05)),(to_sfixed_a(-5.6618882808834314e-06)),(to_sfixed_a(4.041564170620404e-05)),(to_sfixed_a(-2.067320565402042e-05)),(to_sfixed_a(4.214725413476117e-05)),(to_sfixed_a(-4.305940365156857e-06)),(to_sfixed_a(1.95164539036341e-05)),(to_sfixed_a(2.0994031729060225e-05)),(to_sfixed_a(2.90724328806391e-05)),(to_sfixed_a(8.495446309098043e-06)),(to_sfixed_a(4.8654808779247105e-05)),(to_sfixed_a(-2.079859041259624e-05)),(to_sfixed_a(-8.382088708458468e-06)),(to_sfixed_a(-7.356279093073681e-05)),(to_sfixed_a(-6.3737229538674e-06)),(to_sfixed_a(6.079428203520365e-05)),(to_sfixed_a(3.5715929698199034e-05)),(to_sfixed_a(5.308543222781736e-06)),(to_sfixed_a(2.598266746645095e-06)),(to_sfixed_a(1.0225084224657621e-05)),(to_sfixed_a(3.4669188607949764e-05)),(to_sfixed_a(1.7385860701324418e-05)),(to_sfixed_a(-9.735272215039004e-06)),(to_sfixed_a(1.4547736100212205e-05)),(to_sfixed_a(7.007097156019881e-05)));

    constant weight_n1_8 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.04679664969444275)),(to_sfixed_a(-3.133989230263978e-05)),(to_sfixed_a(3.1207148367684567e-06)),(to_sfixed_a(4.990431625628844e-05)),(to_sfixed_a(-4.333142896939535e-06)),(to_sfixed_a(1.8687775082071312e-05)),(to_sfixed_a(3.90123859688174e-05)),(to_sfixed_a(-1.320640734547851e-07)),(to_sfixed_a(-3.845479295705445e-05)),(to_sfixed_a(6.525398202938959e-05)),(to_sfixed_a(1.515791973361047e-05)),(to_sfixed_a(3.859485877910629e-05)),(to_sfixed_a(-4.871340934187174e-05)),(to_sfixed_a(5.342719305190258e-05)),(to_sfixed_a(-3.205979510312318e-06)),(to_sfixed_a(-1.4558981092704926e-05)),(to_sfixed_a(-1.340911603620043e-05)),(to_sfixed_a(-4.320687730796635e-05)),(to_sfixed_a(-7.016912422841415e-05)),(to_sfixed_a(-4.435560913407244e-05)),(to_sfixed_a(-4.9873237003339455e-05)),(to_sfixed_a(-2.4782602849882096e-05)),(to_sfixed_a(-7.261850259965286e-05)),(to_sfixed_a(3.257264324929565e-05)),(to_sfixed_a(2.7724406663764967e-06)),(to_sfixed_a(-2.435583337501157e-05)),(to_sfixed_a(6.111434777267277e-05)),(to_sfixed_a(-4.523115785559639e-05)),(to_sfixed_a(6.932188989594579e-05)),(to_sfixed_a(3.659737922134809e-05)),(to_sfixed_a(2.9598912078654394e-05)),(to_sfixed_a(4.85837554151658e-05)),(to_sfixed_a(-1.3019831385463476e-05)),(to_sfixed_a(1.9494453226798214e-05)),(to_sfixed_a(5.829525980516337e-05)),(to_sfixed_a(9.614016016712412e-05)),(to_sfixed_a(4.512126179179177e-05)),(to_sfixed_a(-1.4355097846419085e-05)));

    constant weight_n1_9 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.13859863579273224)),(to_sfixed_a(2.8186377676320262e-06)),(to_sfixed_a(-5.143622911418788e-05)),(to_sfixed_a(2.0338846297818236e-05)),(to_sfixed_a(-5.7547887990949675e-05)),(to_sfixed_a(3.095579450018704e-05)),(to_sfixed_a(2.1011258013459155e-06)),(to_sfixed_a(-8.561214053770527e-05)),(to_sfixed_a(9.28775807551574e-06)),(to_sfixed_a(1.1634942893579137e-05)),(to_sfixed_a(1.9620350940385833e-05)),(to_sfixed_a(8.701080514583737e-05)),(to_sfixed_a(4.403571438160725e-05)),(to_sfixed_a(-2.3286225768970326e-05)),(to_sfixed_a(1.7820631910581142e-05)),(to_sfixed_a(4.140750752412714e-05)),(to_sfixed_a(3.292912515462376e-05)),(to_sfixed_a(7.113526953617111e-05)),(to_sfixed_a(1.0266438948747236e-05)),(to_sfixed_a(8.03855000413023e-05)),(to_sfixed_a(6.994355771894334e-06)),(to_sfixed_a(-5.533502553589642e-05)),(to_sfixed_a(3.922747509932378e-06)),(to_sfixed_a(1.6358163179575058e-07)),(to_sfixed_a(-4.5814176701242104e-05)),(to_sfixed_a(7.545742118963972e-05)),(to_sfixed_a(1.1007704415533226e-05)),(to_sfixed_a(2.048036731139291e-05)),(to_sfixed_a(-6.596747425646754e-06)),(to_sfixed_a(7.627205923199654e-05)),(to_sfixed_a(6.529536040034145e-05)),(to_sfixed_a(-4.019200423499569e-05)),(to_sfixed_a(7.89731930126436e-05)),(to_sfixed_a(5.6300767028005794e-05)),(to_sfixed_a(-9.482368477620184e-05)),(to_sfixed_a(-7.042314973659813e-05)),(to_sfixed_a(-0.00014334460138343275)),(to_sfixed_a(7.453082798747346e-05)));

    constant weight_n1_10 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.17103831470012665)),(to_sfixed_a(0.0614740364253521)),(to_sfixed_a(0.0006711016758345068)),(to_sfixed_a(-0.025853773579001427)),(to_sfixed_a(-0.038828276097774506)),(to_sfixed_a(0.005968389101326466)),(to_sfixed_a(-0.05593744292855263)),(to_sfixed_a(0.008937756530940533)),(to_sfixed_a(0.11350423097610474)),(to_sfixed_a(-0.10846909880638123)),(to_sfixed_a(0.02403467707335949)),(to_sfixed_a(0.040796466171741486)),(to_sfixed_a(-0.0962071567773819)),(to_sfixed_a(0.021514827385544777)),(to_sfixed_a(-0.02442052960395813)),(to_sfixed_a(0.08134536445140839)),(to_sfixed_a(0.0236167274415493)),(to_sfixed_a(0.016735034063458443)),(to_sfixed_a(-0.04444570094347)),(to_sfixed_a(-0.05264649540185928)),(to_sfixed_a(-0.03281961753964424)),(to_sfixed_a(-0.05315263569355011)),(to_sfixed_a(0.034936923533678055)),(to_sfixed_a(0.0201769657433033)),(to_sfixed_a(-0.05612295866012573)),(to_sfixed_a(-0.02113477885723114)),(to_sfixed_a(0.013476909138262272)),(to_sfixed_a(-0.14845694601535797)),(to_sfixed_a(0.0006540837930515409)),(to_sfixed_a(-0.007310713641345501)),(to_sfixed_a(0.13859446346759796)),(to_sfixed_a(0.10219548642635345)),(to_sfixed_a(0.020377367734909058)),(to_sfixed_a(0.0616360679268837)),(to_sfixed_a(-0.08567667752504349)),(to_sfixed_a(0.04238154739141464)),(to_sfixed_a(-0.056573301553726196)),(to_sfixed_a(-0.04883790388703346)));

    constant weight_n1_11 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.11341952532529831)),(to_sfixed_a(-0.026317300274968147)),(to_sfixed_a(0.0409589558839798)),(to_sfixed_a(0.03191305696964264)),(to_sfixed_a(-0.040321458131074905)),(to_sfixed_a(-0.11767902970314026)),(to_sfixed_a(0.0181435439735651)),(to_sfixed_a(-0.004268655553460121)),(to_sfixed_a(0.028239089995622635)),(to_sfixed_a(0.055681515485048294)),(to_sfixed_a(-0.034894876182079315)),(to_sfixed_a(-0.039741892367601395)),(to_sfixed_a(-0.06331753730773926)),(to_sfixed_a(-0.144149050116539)),(to_sfixed_a(-0.06954652070999146)),(to_sfixed_a(0.024052636697888374)),(to_sfixed_a(-0.03521512448787689)),(to_sfixed_a(0.10069277882575989)),(to_sfixed_a(0.0014001692179590464)),(to_sfixed_a(0.035027388483285904)),(to_sfixed_a(0.017579125240445137)),(to_sfixed_a(-0.2330130785703659)),(to_sfixed_a(-0.043469756841659546)),(to_sfixed_a(0.02332572638988495)),(to_sfixed_a(0.09242324531078339)),(to_sfixed_a(-0.041768841445446014)),(to_sfixed_a(0.04586224630475044)),(to_sfixed_a(-0.10828771442174911)),(to_sfixed_a(0.0007045158999972045)),(to_sfixed_a(-0.0778326541185379)),(to_sfixed_a(0.04657679796218872)),(to_sfixed_a(-0.02362852357327938)),(to_sfixed_a(-0.23534852266311646)),(to_sfixed_a(0.04642012342810631)),(to_sfixed_a(0.056198980659246445)),(to_sfixed_a(-0.13656072318553925)),(to_sfixed_a(0.23521552979946136)),(to_sfixed_a(0.15305617451667786)));

    constant weight_n1_12 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.2920524775981903)),(to_sfixed_a(0.03501550480723381)),(to_sfixed_a(-0.002417318057268858)),(to_sfixed_a(-0.021824073046445847)),(to_sfixed_a(0.017649631947278976)),(to_sfixed_a(0.0048333145678043365)),(to_sfixed_a(0.005597617942839861)),(to_sfixed_a(-0.023650407791137695)),(to_sfixed_a(0.0506531298160553)),(to_sfixed_a(0.04199686273932457)),(to_sfixed_a(-0.036798976361751556)),(to_sfixed_a(-0.013894523493945599)),(to_sfixed_a(0.004769275896251202)),(to_sfixed_a(0.07394711673259735)),(to_sfixed_a(0.010715867392718792)),(to_sfixed_a(0.00821800995618105)),(to_sfixed_a(-0.03664388880133629)),(to_sfixed_a(-0.0076658520847558975)),(to_sfixed_a(0.027281934395432472)),(to_sfixed_a(-0.008547087199985981)),(to_sfixed_a(0.02250680699944496)),(to_sfixed_a(0.0299187283962965)),(to_sfixed_a(-0.002334908116608858)),(to_sfixed_a(-0.012529107742011547)),(to_sfixed_a(0.08033888041973114)),(to_sfixed_a(0.049621231853961945)),(to_sfixed_a(-0.11581474542617798)),(to_sfixed_a(0.10583952069282532)),(to_sfixed_a(-0.021658213809132576)),(to_sfixed_a(0.0024980963207781315)),(to_sfixed_a(0.11425088346004486)),(to_sfixed_a(0.04996525123715401)),(to_sfixed_a(-0.07764647156000137)),(to_sfixed_a(-0.08274644613265991)),(to_sfixed_a(-0.017955681309103966)),(to_sfixed_a(-0.098851278424263)),(to_sfixed_a(-0.029629837721586227)),(to_sfixed_a(-0.006459848955273628)));

    constant weight_n1_13 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.014934713020920753)),(to_sfixed_a(1.4530212865793146e-05)),(to_sfixed_a(1.3598315490526147e-05)),(to_sfixed_a(9.089058039535303e-06)),(to_sfixed_a(1.5541914763161913e-05)),(to_sfixed_a(4.235604501445778e-05)),(to_sfixed_a(-4.803050401847031e-09)),(to_sfixed_a(-3.95621573261451e-05)),(to_sfixed_a(2.150761974917259e-05)),(to_sfixed_a(-4.616214027919341e-06)),(to_sfixed_a(-1.0909316188190132e-05)),(to_sfixed_a(4.1650600905995816e-05)),(to_sfixed_a(4.361571427580202e-06)),(to_sfixed_a(6.839739216957241e-05)),(to_sfixed_a(8.55863545439206e-05)),(to_sfixed_a(3.781135819735937e-05)),(to_sfixed_a(-3.616501635406166e-05)),(to_sfixed_a(7.721572728769388e-06)),(to_sfixed_a(1.3436238077702e-05)),(to_sfixed_a(1.221490583702689e-05)),(to_sfixed_a(4.599786552716978e-05)),(to_sfixed_a(4.245980017003603e-05)),(to_sfixed_a(-5.6801975006237626e-05)),(to_sfixed_a(4.585271381074563e-05)),(to_sfixed_a(-4.3401661969255656e-05)),(to_sfixed_a(1.3239232430350967e-05)),(to_sfixed_a(-0.00011260768224019557)),(to_sfixed_a(-1.988045551115647e-05)),(to_sfixed_a(7.069456478348002e-05)),(to_sfixed_a(-9.573467650625389e-06)),(to_sfixed_a(-6.757337541785091e-05)),(to_sfixed_a(-9.067940482054837e-06)),(to_sfixed_a(-6.288174336077645e-05)),(to_sfixed_a(-0.00010406968794995919)),(to_sfixed_a(-4.470314524951391e-05)),(to_sfixed_a(3.6941735743312165e-05)),(to_sfixed_a(2.167256570828613e-05)),(to_sfixed_a(1.3042786122241523e-05)));

    constant weight_n1_14 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.13107313215732574)),(to_sfixed_a(-2.2140882720123045e-05)),(to_sfixed_a(-3.0082868761382997e-05)),(to_sfixed_a(6.567626314790687e-06)),(to_sfixed_a(2.150773798348382e-05)),(to_sfixed_a(-1.4039650523045566e-05)),(to_sfixed_a(-2.6031932065961882e-05)),(to_sfixed_a(4.023025758215226e-05)),(to_sfixed_a(1.3357777788769454e-05)),(to_sfixed_a(1.9364173567737453e-05)),(to_sfixed_a(5.801308361697011e-05)),(to_sfixed_a(2.4718117856536992e-05)),(to_sfixed_a(6.28880225121975e-05)),(to_sfixed_a(1.1884176274179481e-05)),(to_sfixed_a(1.5964275007718243e-05)),(to_sfixed_a(9.388769103679806e-05)),(to_sfixed_a(-1.4434684999287128e-05)),(to_sfixed_a(4.5737331674899906e-05)),(to_sfixed_a(-8.308610995300114e-05)),(to_sfixed_a(0.00013881881022825837)),(to_sfixed_a(-5.884081110707484e-05)),(to_sfixed_a(0.00010356376878917217)),(to_sfixed_a(-9.10647286218591e-05)),(to_sfixed_a(-1.2864459677075502e-05)),(to_sfixed_a(1.083550614566775e-06)),(to_sfixed_a(-1.8740369341685437e-05)),(to_sfixed_a(1.9797087588813156e-05)),(to_sfixed_a(-3.281267709098756e-05)),(to_sfixed_a(-3.153168290737085e-05)),(to_sfixed_a(3.0346604944497813e-06)),(to_sfixed_a(-3.6627293411584105e-06)),(to_sfixed_a(8.164777682395652e-05)),(to_sfixed_a(1.2592829534696648e-06)),(to_sfixed_a(-0.00016151474846992642)),(to_sfixed_a(-3.17012527375482e-05)),(to_sfixed_a(5.3305309847928584e-05)),(to_sfixed_a(1.393083221046254e-05)),(to_sfixed_a(2.0613038941519335e-05)));

    constant weight_n1_15 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.015202323906123638)),(to_sfixed_a(-0.02352963015437126)),(to_sfixed_a(0.025957437232136726)),(to_sfixed_a(0.3061273396015167)),(to_sfixed_a(0.048959676176309586)),(to_sfixed_a(0.22984431684017181)),(to_sfixed_a(-0.11880534142255783)),(to_sfixed_a(-0.17512862384319305)),(to_sfixed_a(0.0008002542890608311)),(to_sfixed_a(0.004522469826042652)),(to_sfixed_a(0.10902024060487747)),(to_sfixed_a(0.09125497192144394)),(to_sfixed_a(0.014196276664733887)),(to_sfixed_a(-0.050648946315050125)),(to_sfixed_a(-0.012354864738881588)),(to_sfixed_a(0.04260382428765297)),(to_sfixed_a(0.0725390836596489)),(to_sfixed_a(-0.09840375930070877)),(to_sfixed_a(0.13160580396652222)),(to_sfixed_a(-0.0255353432148695)),(to_sfixed_a(-0.1083298996090889)),(to_sfixed_a(0.013997605070471764)),(to_sfixed_a(-0.0404827781021595)),(to_sfixed_a(0.08997572958469391)),(to_sfixed_a(0.04456348344683647)),(to_sfixed_a(0.1287689208984375)),(to_sfixed_a(0.09198031574487686)),(to_sfixed_a(0.095248743891716)),(to_sfixed_a(-0.1458067148923874)),(to_sfixed_a(-0.0601942203938961)),(to_sfixed_a(-0.07245971262454987)),(to_sfixed_a(0.06619004905223846)),(to_sfixed_a(-0.024960199370980263)),(to_sfixed_a(0.08997520804405212)),(to_sfixed_a(-0.1819012612104416)),(to_sfixed_a(0.17305707931518555)),(to_sfixed_a(0.07605673372745514)),(to_sfixed_a(0.1577741652727127)));

    constant weight_n1_16 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.017475103959441185)),(to_sfixed_a(3.172887591063045e-05)),(to_sfixed_a(-2.5790039217099547e-05)),(to_sfixed_a(3.528831803123467e-05)),(to_sfixed_a(-4.421017729328014e-05)),(to_sfixed_a(5.670318569173105e-05)),(to_sfixed_a(8.310656994581223e-06)),(to_sfixed_a(7.342788649111753e-06)),(to_sfixed_a(-3.7691675970563665e-05)),(to_sfixed_a(3.383087459951639e-05)),(to_sfixed_a(-7.754666148684919e-05)),(to_sfixed_a(5.190007505007088e-05)),(to_sfixed_a(-2.4373068299610168e-05)),(to_sfixed_a(9.929191264745896e-07)),(to_sfixed_a(5.3616069635609165e-05)),(to_sfixed_a(-3.813704097410664e-05)),(to_sfixed_a(9.97560073301429e-06)),(to_sfixed_a(-5.184283963899361e-06)),(to_sfixed_a(-4.6812081563984975e-05)),(to_sfixed_a(1.648104989726562e-05)),(to_sfixed_a(3.1124185625230893e-05)),(to_sfixed_a(-1.9053964933846146e-05)),(to_sfixed_a(6.214872701093554e-05)),(to_sfixed_a(-1.9368333596503362e-05)),(to_sfixed_a(4.7312416427303106e-05)),(to_sfixed_a(1.1834777978947386e-05)),(to_sfixed_a(5.65147365705343e-06)),(to_sfixed_a(0.00011306261149002239)),(to_sfixed_a(-2.7716032491298392e-06)),(to_sfixed_a(-3.719871983776102e-06)),(to_sfixed_a(3.2487627322552726e-05)),(to_sfixed_a(-0.00011334140435792506)),(to_sfixed_a(3.337083398946561e-05)),(to_sfixed_a(-1.8217155229649507e-05)),(to_sfixed_a(-3.657582783489488e-05)),(to_sfixed_a(-4.844179056817666e-05)),(to_sfixed_a(6.244388350751251e-05)),(to_sfixed_a(4.74773914902471e-05)));

    constant weight_n1_17 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.0537727065384388)),(to_sfixed_a(-0.08204742521047592)),(to_sfixed_a(-0.06005287915468216)),(to_sfixed_a(0.0735192820429802)),(to_sfixed_a(-0.13016249239444733)),(to_sfixed_a(-0.016805002465844154)),(to_sfixed_a(0.05877940356731415)),(to_sfixed_a(-0.006903945934027433)),(to_sfixed_a(0.23488624393939972)),(to_sfixed_a(0.012688315473496914)),(to_sfixed_a(0.151970773935318)),(to_sfixed_a(-0.06357371062040329)),(to_sfixed_a(0.05499701946973801)),(to_sfixed_a(0.08942292630672455)),(to_sfixed_a(0.050369929522275925)),(to_sfixed_a(0.09305092692375183)),(to_sfixed_a(-0.15917854011058807)),(to_sfixed_a(-0.0848456546664238)),(to_sfixed_a(0.06381462514400482)),(to_sfixed_a(0.22983798384666443)),(to_sfixed_a(0.07247018814086914)),(to_sfixed_a(-0.16501854360103607)),(to_sfixed_a(0.11710082739591599)),(to_sfixed_a(0.17672866582870483)),(to_sfixed_a(0.1357259452342987)),(to_sfixed_a(0.12570247054100037)),(to_sfixed_a(0.18784934282302856)),(to_sfixed_a(-0.08817286789417267)),(to_sfixed_a(-0.2600935995578766)),(to_sfixed_a(0.18642134964466095)),(to_sfixed_a(0.10146913677453995)),(to_sfixed_a(-0.07884285598993301)),(to_sfixed_a(-0.02237175963819027)),(to_sfixed_a(0.09940338134765625)),(to_sfixed_a(0.2051762342453003)),(to_sfixed_a(-0.08147265017032623)),(to_sfixed_a(0.026116836816072464)),(to_sfixed_a(-0.0248823594301939)));

    constant weight_n1_18 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.3387475609779358)),(to_sfixed_a(0.0024274757597595453)),(to_sfixed_a(-0.0055298395454883575)),(to_sfixed_a(-0.044792693108320236)),(to_sfixed_a(-0.0387197881937027)),(to_sfixed_a(-0.05853961035609245)),(to_sfixed_a(0.021882900968194008)),(to_sfixed_a(-0.02764962427318096)),(to_sfixed_a(-0.033059198409318924)),(to_sfixed_a(-0.002233870793133974)),(to_sfixed_a(-0.025641929358243942)),(to_sfixed_a(-0.034686580300331116)),(to_sfixed_a(-0.040365319699048996)),(to_sfixed_a(-0.02291906252503395)),(to_sfixed_a(0.038523975759744644)),(to_sfixed_a(0.07094667851924896)),(to_sfixed_a(-0.010684475302696228)),(to_sfixed_a(0.07148140668869019)),(to_sfixed_a(0.022285571321845055)),(to_sfixed_a(0.03772582486271858)),(to_sfixed_a(-0.020542137324810028)),(to_sfixed_a(0.020144859328866005)),(to_sfixed_a(-0.012900346890091896)),(to_sfixed_a(-0.004108199384063482)),(to_sfixed_a(-0.038626622408628464)),(to_sfixed_a(0.022806620225310326)),(to_sfixed_a(0.024955814704298973)),(to_sfixed_a(-0.013200457207858562)),(to_sfixed_a(0.08242509514093399)),(to_sfixed_a(0.04301447421312332)),(to_sfixed_a(0.05456922948360443)),(to_sfixed_a(-0.039809197187423706)),(to_sfixed_a(0.02875654771924019)),(to_sfixed_a(-0.05503278970718384)),(to_sfixed_a(0.03412732109427452)),(to_sfixed_a(0.04942793399095535)),(to_sfixed_a(0.011432480998337269)),(to_sfixed_a(0.01405561063438654)));

    constant weight_n1_19 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.009435213170945644)),(to_sfixed_a(-2.5920289772329852e-05)),(to_sfixed_a(1.6719879567972384e-05)),(to_sfixed_a(-1.88440262718359e-05)),(to_sfixed_a(4.790538514498621e-05)),(to_sfixed_a(9.964627679437399e-05)),(to_sfixed_a(5.9968893765471876e-05)),(to_sfixed_a(3.888646824634634e-05)),(to_sfixed_a(1.0224235666100867e-05)),(to_sfixed_a(-3.2365638617193326e-05)),(to_sfixed_a(3.84001832571812e-05)),(to_sfixed_a(-1.149012769019464e-05)),(to_sfixed_a(5.756412065238692e-05)),(to_sfixed_a(-0.00011372340668458492)),(to_sfixed_a(1.9437029550317675e-05)),(to_sfixed_a(2.0609704733942635e-06)),(to_sfixed_a(5.897384471609257e-05)),(to_sfixed_a(1.891100396278489e-06)),(to_sfixed_a(3.5076329368166625e-05)),(to_sfixed_a(4.380163591122255e-05)),(to_sfixed_a(1.6776975826360285e-05)),(to_sfixed_a(6.600220513064414e-05)),(to_sfixed_a(-1.6750347640481777e-05)),(to_sfixed_a(4.372330295154825e-05)),(to_sfixed_a(5.387702799453109e-07)),(to_sfixed_a(4.9363781727151945e-05)),(to_sfixed_a(6.01743595325388e-05)),(to_sfixed_a(3.5220335121266544e-05)),(to_sfixed_a(-5.095193046145141e-06)),(to_sfixed_a(-9.858630619419273e-06)),(to_sfixed_a(6.990307156229392e-05)),(to_sfixed_a(3.461899177636951e-05)),(to_sfixed_a(-4.557673310046084e-05)),(to_sfixed_a(6.321540422504768e-05)),(to_sfixed_a(2.836689782270696e-05)),(to_sfixed_a(4.903970693703741e-05)),(to_sfixed_a(2.9268212529132143e-05)),(to_sfixed_a(-4.8875604989007115e-05)));

    constant weight_n1_20 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.016156548634171486)),(to_sfixed_a(-1.0837058653123677e-05)),(to_sfixed_a(1.2692167729255743e-05)),(to_sfixed_a(-2.7813159249490127e-05)),(to_sfixed_a(4.7979456212488e-06)),(to_sfixed_a(-9.650644642533734e-06)),(to_sfixed_a(3.4928299896819226e-07)),(to_sfixed_a(2.023770139203407e-05)),(to_sfixed_a(1.834616341511719e-05)),(to_sfixed_a(-3.031984078916139e-06)),(to_sfixed_a(-2.847695031960029e-05)),(to_sfixed_a(-1.640959453652613e-05)),(to_sfixed_a(-1.2779550161212683e-05)),(to_sfixed_a(-4.1904422687366605e-05)),(to_sfixed_a(5.474931822391227e-05)),(to_sfixed_a(2.804094947350677e-05)),(to_sfixed_a(-5.388021236285567e-05)),(to_sfixed_a(4.207202073303051e-05)),(to_sfixed_a(3.381960777915083e-05)),(to_sfixed_a(-9.629229316487908e-05)),(to_sfixed_a(1.8610047845868394e-05)),(to_sfixed_a(-1.980873457796406e-05)),(to_sfixed_a(2.497848072380293e-05)),(to_sfixed_a(-6.818756810389459e-05)),(to_sfixed_a(-5.0430160627001897e-05)),(to_sfixed_a(-1.4618382920161821e-05)),(to_sfixed_a(-3.649169593700208e-05)),(to_sfixed_a(-0.00011295972217340022)),(to_sfixed_a(-0.00010907367686741054)),(to_sfixed_a(1.5424697267008014e-05)),(to_sfixed_a(-1.1284837455605157e-05)),(to_sfixed_a(-6.850846693851054e-05)),(to_sfixed_a(2.0531746486085467e-05)),(to_sfixed_a(-3.331353946123272e-05)),(to_sfixed_a(-4.446764705789974e-06)),(to_sfixed_a(-2.4965031116153114e-05)),(to_sfixed_a(1.0520142495806795e-05)),(to_sfixed_a(4.297954001231119e-05)));

    constant weight_n1_21 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.08488751947879791)),(to_sfixed_a(-0.020529722794890404)),(to_sfixed_a(-0.01853235997259617)),(to_sfixed_a(0.011093569919466972)),(to_sfixed_a(-0.00963394995778799)),(to_sfixed_a(-0.009139927104115486)),(to_sfixed_a(0.0070523424074053764)),(to_sfixed_a(0.0006077342550270259)),(to_sfixed_a(-0.0060120983980596066)),(to_sfixed_a(-0.012668251991271973)),(to_sfixed_a(-0.013077937066555023)),(to_sfixed_a(-0.010562249459326267)),(to_sfixed_a(0.0066162901930511)),(to_sfixed_a(-0.018595939502120018)),(to_sfixed_a(-0.006859954446554184)),(to_sfixed_a(0.010857721790671349)),(to_sfixed_a(0.010170870460569859)),(to_sfixed_a(0.02267252840101719)),(to_sfixed_a(0.022155610844492912)),(to_sfixed_a(0.0003730496682692319)),(to_sfixed_a(-0.0048335250467062)),(to_sfixed_a(-0.02047053724527359)),(to_sfixed_a(0.00574149563908577)),(to_sfixed_a(0.0011244899360463023)),(to_sfixed_a(-0.010817439295351505)),(to_sfixed_a(0.014260541647672653)),(to_sfixed_a(0.016751041635870934)),(to_sfixed_a(0.004489622078835964)),(to_sfixed_a(-0.014937720261514187)),(to_sfixed_a(0.027436671778559685)),(to_sfixed_a(-0.01443813182413578)),(to_sfixed_a(0.024904325604438782)),(to_sfixed_a(-0.027660798281431198)),(to_sfixed_a(0.060921818017959595)),(to_sfixed_a(0.03192202374339104)),(to_sfixed_a(-0.019927339628338814)),(to_sfixed_a(-0.009106406010687351)),(to_sfixed_a(0.043623361736536026)));

    constant weight_n1_22 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.3388829529285431)),(to_sfixed_a(0.06306254863739014)),(to_sfixed_a(-0.018247975036501884)),(to_sfixed_a(0.03590216860175133)),(to_sfixed_a(-0.020651960745453835)),(to_sfixed_a(-0.08568773418664932)),(to_sfixed_a(-0.04015800356864929)),(to_sfixed_a(-0.019480496644973755)),(to_sfixed_a(0.027028487995266914)),(to_sfixed_a(-0.034305471926927567)),(to_sfixed_a(0.0039274548180401325)),(to_sfixed_a(-0.05321979895234108)),(to_sfixed_a(-0.00013266783207654953)),(to_sfixed_a(0.04884318634867668)),(to_sfixed_a(-0.03205883130431175)),(to_sfixed_a(0.04282161220908165)),(to_sfixed_a(0.06464540213346481)),(to_sfixed_a(-0.06791651993989944)),(to_sfixed_a(0.06039780005812645)),(to_sfixed_a(0.0048140776343643665)),(to_sfixed_a(-0.0719352588057518)),(to_sfixed_a(0.04713510721921921)),(to_sfixed_a(-0.027387501671910286)),(to_sfixed_a(-0.032816462218761444)),(to_sfixed_a(-0.03368411213159561)),(to_sfixed_a(-0.03883130103349686)),(to_sfixed_a(-0.06563253700733185)),(to_sfixed_a(0.1437264382839203)),(to_sfixed_a(0.019028550013899803)),(to_sfixed_a(-0.11508702486753464)),(to_sfixed_a(0.029440855607390404)),(to_sfixed_a(-0.1737305372953415)),(to_sfixed_a(-0.05599354952573776)),(to_sfixed_a(0.003721206448972225)),(to_sfixed_a(-0.07292850315570831)),(to_sfixed_a(-0.004272350575774908)),(to_sfixed_a(0.16978232562541962)),(to_sfixed_a(0.14072251319885254)));

    constant weight_n1_23 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.056550316512584686)),(to_sfixed_a(0.0449211485683918)),(to_sfixed_a(-0.030508941039443016)),(to_sfixed_a(0.1516026109457016)),(to_sfixed_a(0.03930116072297096)),(to_sfixed_a(0.10340327769517899)),(to_sfixed_a(-0.09394613653421402)),(to_sfixed_a(-0.05316054821014404)),(to_sfixed_a(-0.003112674690783024)),(to_sfixed_a(0.012571916915476322)),(to_sfixed_a(0.04554963856935501)),(to_sfixed_a(0.0371282622218132)),(to_sfixed_a(0.02268599532544613)),(to_sfixed_a(-0.005893521476536989)),(to_sfixed_a(-0.0016376242274418473)),(to_sfixed_a(0.03731324523687363)),(to_sfixed_a(0.002526202006265521)),(to_sfixed_a(0.004861832596361637)),(to_sfixed_a(-0.004817882552742958)),(to_sfixed_a(-0.04363107681274414)),(to_sfixed_a(-0.10020943731069565)),(to_sfixed_a(-0.02396233193576336)),(to_sfixed_a(-0.04851171746850014)),(to_sfixed_a(0.04124967381358147)),(to_sfixed_a(0.03072277456521988)),(to_sfixed_a(0.06056436523795128)),(to_sfixed_a(0.0024369489401578903)),(to_sfixed_a(-0.02203507162630558)),(to_sfixed_a(0.020647209137678146)),(to_sfixed_a(0.005436315201222897)),(to_sfixed_a(-0.04950582608580589)),(to_sfixed_a(0.024004587903618813)),(to_sfixed_a(0.01738583669066429)),(to_sfixed_a(-0.0030787745490670204)),(to_sfixed_a(-0.023057792335748672)),(to_sfixed_a(0.023140501230955124)),(to_sfixed_a(0.022840334102511406)),(to_sfixed_a(0.035981565713882446)));

    constant weight_n1_24 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.19301003217697144)),(to_sfixed_a(-0.08251790702342987)),(to_sfixed_a(0.003770522540435195)),(to_sfixed_a(0.11204762011766434)),(to_sfixed_a(-0.001243185717612505)),(to_sfixed_a(0.03264708071947098)),(to_sfixed_a(-0.09348401427268982)),(to_sfixed_a(0.01337931677699089)),(to_sfixed_a(-0.020748762413859367)),(to_sfixed_a(0.09647747874259949)),(to_sfixed_a(0.05486660078167915)),(to_sfixed_a(0.08404608815908432)),(to_sfixed_a(0.00650600902736187)),(to_sfixed_a(-0.0943351536989212)),(to_sfixed_a(0.023348968476057053)),(to_sfixed_a(-0.12768979370594025)),(to_sfixed_a(-0.0835750475525856)),(to_sfixed_a(-0.06101038306951523)),(to_sfixed_a(0.07830838114023209)),(to_sfixed_a(-0.053954754024744034)),(to_sfixed_a(-0.07084871083498001)),(to_sfixed_a(-0.03486349806189537)),(to_sfixed_a(0.046172041445970535)),(to_sfixed_a(0.058099523186683655)),(to_sfixed_a(0.06421691179275513)),(to_sfixed_a(-0.005437719635665417)),(to_sfixed_a(-0.031151944771409035)),(to_sfixed_a(0.045289650559425354)),(to_sfixed_a(-0.15294359624385834)),(to_sfixed_a(-0.017683226615190506)),(to_sfixed_a(-0.07156246155500412)),(to_sfixed_a(-0.04347074031829834)),(to_sfixed_a(-0.01558687910437584)),(to_sfixed_a(0.002036845311522484)),(to_sfixed_a(-0.01487888302654028)),(to_sfixed_a(-0.05039219930768013)),(to_sfixed_a(-0.03567424789071083)),(to_sfixed_a(-0.1966315656900406)));

    constant weight_n1_25 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.010163313709199429)),(to_sfixed_a(1.2898179193143733e-05)),(to_sfixed_a(-1.0600236919344752e-06)),(to_sfixed_a(5.459773092297837e-05)),(to_sfixed_a(5.515712473425083e-05)),(to_sfixed_a(-3.396939791855402e-05)),(to_sfixed_a(-2.893924101954326e-05)),(to_sfixed_a(-3.980580731877126e-05)),(to_sfixed_a(-1.7427390048396774e-05)),(to_sfixed_a(-4.002129571745172e-06)),(to_sfixed_a(4.6797333197901025e-05)),(to_sfixed_a(-2.2756286853109486e-05)),(to_sfixed_a(5.3070874855620787e-05)),(to_sfixed_a(6.559685425600037e-05)),(to_sfixed_a(-2.16426433325978e-05)),(to_sfixed_a(2.2228065063245595e-05)),(to_sfixed_a(6.672349172731629e-06)),(to_sfixed_a(1.4202535567164887e-05)),(to_sfixed_a(6.167924584588036e-05)),(to_sfixed_a(2.344448603253113e-06)),(to_sfixed_a(-4.158891533734277e-05)),(to_sfixed_a(3.4999837225768715e-05)),(to_sfixed_a(1.1655652997433208e-05)),(to_sfixed_a(1.2754225281241816e-05)),(to_sfixed_a(-0.0001065957112587057)),(to_sfixed_a(-4.324758629081771e-05)),(to_sfixed_a(5.0717433623503894e-05)),(to_sfixed_a(1.766321474860888e-05)),(to_sfixed_a(-2.3439546566805802e-05)),(to_sfixed_a(4.362399340607226e-05)),(to_sfixed_a(-1.0852242667169776e-05)),(to_sfixed_a(-7.76855358708417e-06)),(to_sfixed_a(7.476705650333315e-05)),(to_sfixed_a(2.8469379685702734e-05)),(to_sfixed_a(2.847196810762398e-05)),(to_sfixed_a(-7.71917257225141e-06)),(to_sfixed_a(0.0001657532120589167)),(to_sfixed_a(-1.3389705600275192e-05)));

    constant weight_n1_26 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.0329965315759182)),(to_sfixed_a(-9.062649041879922e-05)),(to_sfixed_a(-0.002058528596535325)),(to_sfixed_a(-0.005019751843065023)),(to_sfixed_a(0.011407322250306606)),(to_sfixed_a(0.005671403836458921)),(to_sfixed_a(0.013461073860526085)),(to_sfixed_a(0.013788748532533646)),(to_sfixed_a(-0.013404661789536476)),(to_sfixed_a(0.002446400932967663)),(to_sfixed_a(0.023130428045988083)),(to_sfixed_a(-0.008108756504952908)),(to_sfixed_a(0.011350600980222225)),(to_sfixed_a(0.02682788297533989)),(to_sfixed_a(-0.0034642554819583893)),(to_sfixed_a(-0.01153501681983471)),(to_sfixed_a(0.020764490589499474)),(to_sfixed_a(-0.022120937705039978)),(to_sfixed_a(-0.01843954063951969)),(to_sfixed_a(0.009535438381135464)),(to_sfixed_a(-0.009312060661613941)),(to_sfixed_a(-0.007188678253442049)),(to_sfixed_a(0.018942443653941154)),(to_sfixed_a(-0.01691923849284649)),(to_sfixed_a(-0.015326433815062046)),(to_sfixed_a(-0.009579800069332123)),(to_sfixed_a(0.019484343007206917)),(to_sfixed_a(-0.036345914006233215)),(to_sfixed_a(0.0035756740253418684)),(to_sfixed_a(0.007985001429915428)),(to_sfixed_a(0.01699298433959484)),(to_sfixed_a(-0.00042654338176362216)),(to_sfixed_a(-0.021779607981443405)),(to_sfixed_a(0.02008412964642048)),(to_sfixed_a(0.0017966337036341429)),(to_sfixed_a(-0.0040507023222744465)),(to_sfixed_a(0.012073630467057228)),(to_sfixed_a(0.037682197988033295)));

    constant weight_n1_27 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.02159428969025612)),(to_sfixed_a(-0.014393184334039688)),(to_sfixed_a(0.008365826681256294)),(to_sfixed_a(0.0035537080839276314)),(to_sfixed_a(0.004869292490184307)),(to_sfixed_a(-0.020336203277111053)),(to_sfixed_a(-0.007681902498006821)),(to_sfixed_a(-0.012311539612710476)),(to_sfixed_a(-0.006020972039550543)),(to_sfixed_a(-0.006949135102331638)),(to_sfixed_a(0.030094359070062637)),(to_sfixed_a(-0.0039281644858419895)),(to_sfixed_a(-0.00407027080655098)),(to_sfixed_a(-0.00831606611609459)),(to_sfixed_a(0.007891851477324963)),(to_sfixed_a(0.02703656256198883)),(to_sfixed_a(0.008740690536797047)),(to_sfixed_a(0.016362076625227928)),(to_sfixed_a(-0.007794732693582773)),(to_sfixed_a(0.02467302605509758)),(to_sfixed_a(-0.025755755603313446)),(to_sfixed_a(0.007268762681633234)),(to_sfixed_a(0.009031897410750389)),(to_sfixed_a(-0.002296414691954851)),(to_sfixed_a(0.0216505229473114)),(to_sfixed_a(-0.02662508189678192)),(to_sfixed_a(-0.022067934274673462)),(to_sfixed_a(-0.015787839889526367)),(to_sfixed_a(0.012669256888329983)),(to_sfixed_a(-0.005016736686229706)),(to_sfixed_a(-0.009141343645751476)),(to_sfixed_a(-0.017870984971523285)),(to_sfixed_a(-0.002690694760531187)),(to_sfixed_a(-0.008945876732468605)),(to_sfixed_a(-0.014038554392755032)),(to_sfixed_a(0.006788910366594791)),(to_sfixed_a(0.011806518770754337)),(to_sfixed_a(0.0029020707588642836)));

    constant weight_n1_28 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.011202746070921421)),(to_sfixed_a(2.0296545699238777e-05)),(to_sfixed_a(-2.6980862458003685e-05)),(to_sfixed_a(1.985494418477174e-05)),(to_sfixed_a(-3.5252526231488446e-06)),(to_sfixed_a(-3.0463997973129153e-05)),(to_sfixed_a(-2.5120089048868977e-05)),(to_sfixed_a(2.9635508326464333e-05)),(to_sfixed_a(1.796440665202681e-05)),(to_sfixed_a(-4.17538576584775e-05)),(to_sfixed_a(-2.742660626608995e-06)),(to_sfixed_a(-4.0443283069180325e-05)),(to_sfixed_a(-2.0109671822865494e-05)),(to_sfixed_a(4.653645009966567e-05)),(to_sfixed_a(5.736068851547316e-05)),(to_sfixed_a(5.3261803259374574e-05)),(to_sfixed_a(4.668645851779729e-05)),(to_sfixed_a(-4.837666710955091e-05)),(to_sfixed_a(-2.56992152571911e-05)),(to_sfixed_a(2.9374834412010387e-05)),(to_sfixed_a(4.287116098566912e-05)),(to_sfixed_a(-3.7841371522517875e-05)),(to_sfixed_a(-4.188726961729117e-05)),(to_sfixed_a(6.002026202622801e-05)),(to_sfixed_a(3.827758337138221e-05)),(to_sfixed_a(1.4391062904905993e-05)),(to_sfixed_a(-4.373728734208271e-05)),(to_sfixed_a(-5.662022522301413e-05)),(to_sfixed_a(-3.647309131338261e-05)),(to_sfixed_a(-2.7613883503363468e-05)),(to_sfixed_a(5.6151493481593207e-05)),(to_sfixed_a(-4.490287392400205e-05)),(to_sfixed_a(3.2180623747990467e-06)),(to_sfixed_a(2.550003773649223e-05)),(to_sfixed_a(6.744553684256971e-05)),(to_sfixed_a(-8.888895536074415e-06)),(to_sfixed_a(-3.1962626962922513e-05)),(to_sfixed_a(8.762521611060947e-05)));

    constant weight_n1_29 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.41458073258399963)),(to_sfixed_a(0.0496169812977314)),(to_sfixed_a(-0.09348423779010773)),(to_sfixed_a(-0.06423758715391159)),(to_sfixed_a(-0.056709885597229004)),(to_sfixed_a(-0.028395043686032295)),(to_sfixed_a(-0.07823291420936584)),(to_sfixed_a(-0.08101323992013931)),(to_sfixed_a(0.03184331953525543)),(to_sfixed_a(-0.017670053988695145)),(to_sfixed_a(0.08884914219379425)),(to_sfixed_a(0.09264938533306122)),(to_sfixed_a(-0.06004953756928444)),(to_sfixed_a(0.011180934496223927)),(to_sfixed_a(0.029058970510959625)),(to_sfixed_a(-0.27775058150291443)),(to_sfixed_a(-0.04640975221991539)),(to_sfixed_a(-0.09134308248758316)),(to_sfixed_a(-0.10197075456380844)),(to_sfixed_a(-0.05831557884812355)),(to_sfixed_a(0.03168844059109688)),(to_sfixed_a(-0.09096752107143402)),(to_sfixed_a(0.04497425630688667)),(to_sfixed_a(0.001022822572849691)),(to_sfixed_a(0.096289724111557)),(to_sfixed_a(-0.1656755656003952)),(to_sfixed_a(0.057180941104888916)),(to_sfixed_a(0.06149530038237572)),(to_sfixed_a(-0.028992680832743645)),(to_sfixed_a(-0.02861592173576355)),(to_sfixed_a(-0.16682828962802887)),(to_sfixed_a(0.1214914619922638)),(to_sfixed_a(-0.09630978852510452)),(to_sfixed_a(-0.13230551779270172)),(to_sfixed_a(0.12290908396244049)),(to_sfixed_a(-0.008306160569190979)),(to_sfixed_a(0.041780050843954086)),(to_sfixed_a(0.011248485185205936)));

    constant weight_n1_30 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.02053939551115036)),(to_sfixed_a(2.8517195460153744e-05)),(to_sfixed_a(3.480026498436928e-05)),(to_sfixed_a(1.0416860277473461e-05)),(to_sfixed_a(3.834104791167192e-05)),(to_sfixed_a(1.9546798284864053e-05)),(to_sfixed_a(-3.474478216958232e-05)),(to_sfixed_a(-2.7014390070689842e-05)),(to_sfixed_a(-2.231075086456258e-05)),(to_sfixed_a(4.063319465785753e-06)),(to_sfixed_a(1.201015584229026e-05)),(to_sfixed_a(6.61985836813983e-07)),(to_sfixed_a(1.8664168237592094e-05)),(to_sfixed_a(-2.710166882025078e-05)),(to_sfixed_a(-4.159766831435263e-05)),(to_sfixed_a(-6.539830792462453e-05)),(to_sfixed_a(-2.562947520345915e-05)),(to_sfixed_a(3.0177488952176645e-05)),(to_sfixed_a(-4.023610472358996e-06)),(to_sfixed_a(-1.0215784413958318e-06)),(to_sfixed_a(-3.347160236444324e-05)),(to_sfixed_a(7.043007826723624e-06)),(to_sfixed_a(6.12858566455543e-05)),(to_sfixed_a(-0.00011171379446750507)),(to_sfixed_a(2.8180404115119018e-05)),(to_sfixed_a(2.6096322471858002e-05)),(to_sfixed_a(-4.549518052954227e-05)),(to_sfixed_a(-2.7726371627068147e-05)),(to_sfixed_a(-8.485346188535914e-05)),(to_sfixed_a(5.00196692883037e-05)),(to_sfixed_a(-1.2899876310257241e-05)),(to_sfixed_a(-2.2137639462016523e-05)),(to_sfixed_a(1.4004352806296083e-06)),(to_sfixed_a(1.7627871784497984e-05)),(to_sfixed_a(3.823037332040258e-05)),(to_sfixed_a(3.8139809475978836e-05)),(to_sfixed_a(5.151443838258274e-05)),(to_sfixed_a(6.3091119955061e-06)));

    constant weight_n1_31 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.09969425946474075)),(to_sfixed_a(0.02652564086019993)),(to_sfixed_a(0.009515817277133465)),(to_sfixed_a(0.00795727875083685)),(to_sfixed_a(0.024598848074674606)),(to_sfixed_a(-0.03224800154566765)),(to_sfixed_a(0.06432005017995834)),(to_sfixed_a(0.023707177489995956)),(to_sfixed_a(0.018295006826519966)),(to_sfixed_a(0.07519587129354477)),(to_sfixed_a(0.12931033968925476)),(to_sfixed_a(-0.038277167826890945)),(to_sfixed_a(-0.0067866044119000435)),(to_sfixed_a(0.048066262155771255)),(to_sfixed_a(0.06508086621761322)),(to_sfixed_a(-0.04784635454416275)),(to_sfixed_a(0.06611470878124237)),(to_sfixed_a(0.017964407801628113)),(to_sfixed_a(0.04861770570278168)),(to_sfixed_a(-0.029589783400297165)),(to_sfixed_a(-0.11960361897945404)),(to_sfixed_a(-0.024361642077565193)),(to_sfixed_a(0.09739729017019272)),(to_sfixed_a(0.0037093795835971832)),(to_sfixed_a(0.03514132648706436)),(to_sfixed_a(0.019491203129291534)),(to_sfixed_a(-0.13953617215156555)),(to_sfixed_a(0.008575394749641418)),(to_sfixed_a(0.011234205216169357)),(to_sfixed_a(0.030775075778365135)),(to_sfixed_a(0.038455672562122345)),(to_sfixed_a(-0.08407005667686462)),(to_sfixed_a(-0.10178883373737335)),(to_sfixed_a(0.01745462231338024)),(to_sfixed_a(0.08732061833143234)),(to_sfixed_a(0.10064733773469925)),(to_sfixed_a(-0.06719191372394562)),(to_sfixed_a(-0.012944987043738365)));

    constant weight_n1_32 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.20669777691364288)),(to_sfixed_a(-2.7330992452334613e-05)),(to_sfixed_a(-2.1414934963104315e-05)),(to_sfixed_a(-2.7258252885076217e-05)),(to_sfixed_a(3.1445066269952804e-05)),(to_sfixed_a(-8.48708805278875e-05)),(to_sfixed_a(4.9175077947438695e-06)),(to_sfixed_a(-1.6701200365787372e-05)),(to_sfixed_a(-2.60975521086948e-05)),(to_sfixed_a(-1.4275540252128849e-06)),(to_sfixed_a(1.5401845303131267e-05)),(to_sfixed_a(3.3881107810884714e-05)),(to_sfixed_a(-1.5610527043463662e-05)),(to_sfixed_a(2.606187990750186e-05)),(to_sfixed_a(-0.00011214752157684416)),(to_sfixed_a(0.00011702156189130619)),(to_sfixed_a(4.263222581357695e-05)),(to_sfixed_a(-7.475245365640149e-05)),(to_sfixed_a(1.1118473594251554e-05)),(to_sfixed_a(-1.0623281241350924e-06)),(to_sfixed_a(6.586474773939699e-05)),(to_sfixed_a(3.3793341572163627e-05)),(to_sfixed_a(1.5652187357773073e-05)),(to_sfixed_a(4.0455466660205275e-05)),(to_sfixed_a(9.18121531867655e-06)),(to_sfixed_a(9.558304736856371e-05)),(to_sfixed_a(6.689759175060317e-05)),(to_sfixed_a(-1.9595139747252688e-05)),(to_sfixed_a(-5.260952457319945e-05)),(to_sfixed_a(1.7078269593184814e-05)),(to_sfixed_a(-9.312208931078203e-06)),(to_sfixed_a(-0.0001648550241952762)),(to_sfixed_a(4.629913019016385e-05)),(to_sfixed_a(3.007261966558872e-06)),(to_sfixed_a(7.600748358527198e-05)),(to_sfixed_a(2.322045293112751e-05)),(to_sfixed_a(5.1824452384607866e-05)),(to_sfixed_a(2.2970916688791476e-06)));

    constant weight_n1_33 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.07146091759204865)),(to_sfixed_a(-4.058091508341022e-05)),(to_sfixed_a(-4.4755415729014203e-07)),(to_sfixed_a(-4.341354269854492e-06)),(to_sfixed_a(1.9883545974153094e-06)),(to_sfixed_a(-8.674481250636745e-06)),(to_sfixed_a(-4.128240107093006e-06)),(to_sfixed_a(-6.0098449466750026e-05)),(to_sfixed_a(2.6090741812367924e-05)),(to_sfixed_a(5.397655968408799e-06)),(to_sfixed_a(9.496440725342836e-06)),(to_sfixed_a(9.889603825286031e-05)),(to_sfixed_a(1.8012256987276487e-05)),(to_sfixed_a(6.120403850218281e-05)),(to_sfixed_a(1.2748158724207315e-06)),(to_sfixed_a(-4.852853817283176e-05)),(to_sfixed_a(-1.087601140170591e-05)),(to_sfixed_a(2.1138996089575812e-05)),(to_sfixed_a(1.8851364075089805e-05)),(to_sfixed_a(9.845355816651136e-05)),(to_sfixed_a(-1.561674253025558e-05)),(to_sfixed_a(1.2296522982069291e-05)),(to_sfixed_a(-5.581289951805957e-05)),(to_sfixed_a(-5.042244083597325e-05)),(to_sfixed_a(3.0406619771383703e-05)),(to_sfixed_a(6.471824599429965e-05)),(to_sfixed_a(4.139247721468564e-06)),(to_sfixed_a(4.8274159780703485e-05)),(to_sfixed_a(-2.6610887289280072e-05)),(to_sfixed_a(-4.271467332728207e-05)),(to_sfixed_a(2.4350589228561148e-05)),(to_sfixed_a(2.2336433175951242e-05)),(to_sfixed_a(2.773332926153671e-05)),(to_sfixed_a(1.6469633919768967e-05)),(to_sfixed_a(5.982703805784695e-05)),(to_sfixed_a(-9.1788297140738e-06)),(to_sfixed_a(-1.5460687791346572e-05)),(to_sfixed_a(3.462222593952902e-05)));

    constant weight_n1_34 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.00856279581785202)),(to_sfixed_a(1.065331252902979e-05)),(to_sfixed_a(2.8276310331420973e-05)),(to_sfixed_a(-3.489614027785137e-05)),(to_sfixed_a(-1.8776745491777547e-05)),(to_sfixed_a(1.2638794032682199e-05)),(to_sfixed_a(-2.6175648599746637e-05)),(to_sfixed_a(7.146974439820042e-06)),(to_sfixed_a(5.4250227549346164e-05)),(to_sfixed_a(-1.5343050108640455e-05)),(to_sfixed_a(-2.8624112019315362e-05)),(to_sfixed_a(-1.1095442459918559e-05)),(to_sfixed_a(1.3680629308510106e-05)),(to_sfixed_a(1.2981249710719567e-05)),(to_sfixed_a(4.36340706073679e-05)),(to_sfixed_a(5.9929454437224194e-05)),(to_sfixed_a(-3.5885987017536536e-05)),(to_sfixed_a(4.792472464032471e-05)),(to_sfixed_a(4.3739219108829275e-05)),(to_sfixed_a(1.5416278984048404e-05)),(to_sfixed_a(1.3456181591209315e-07)),(to_sfixed_a(-5.578310810960829e-05)),(to_sfixed_a(-4.877989340457134e-05)),(to_sfixed_a(7.578723852930125e-06)),(to_sfixed_a(-9.168501128442585e-05)),(to_sfixed_a(-0.00010503115481697023)),(to_sfixed_a(-3.4502738799346844e-06)),(to_sfixed_a(3.203453525202349e-05)),(to_sfixed_a(-9.164263246930204e-06)),(to_sfixed_a(-0.0001390495744999498)),(to_sfixed_a(4.335137873567874e-06)),(to_sfixed_a(-3.336522786412388e-05)),(to_sfixed_a(-3.96502400690224e-05)),(to_sfixed_a(-9.476151171838865e-05)),(to_sfixed_a(3.5764063795795664e-05)),(to_sfixed_a(2.1843565264134668e-05)),(to_sfixed_a(8.406141205341555e-07)),(to_sfixed_a(-8.386159606743604e-05)));

    constant weight_n1_35 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.0266406387090683)),(to_sfixed_a(0.18162676692008972)),(to_sfixed_a(0.13585342466831207)),(to_sfixed_a(0.04895550385117531)),(to_sfixed_a(-0.12388446182012558)),(to_sfixed_a(0.0016504505183547735)),(to_sfixed_a(0.122244693338871)),(to_sfixed_a(-0.04715784266591072)),(to_sfixed_a(0.04462355002760887)),(to_sfixed_a(-0.11232420057058334)),(to_sfixed_a(-0.011965760961174965)),(to_sfixed_a(0.20884670317173004)),(to_sfixed_a(0.06653088331222534)),(to_sfixed_a(-0.08450433611869812)),(to_sfixed_a(-0.05941226705908775)),(to_sfixed_a(0.017335068434476852)),(to_sfixed_a(-0.1435462087392807)),(to_sfixed_a(-0.1081174910068512)),(to_sfixed_a(-0.02101902849972248)),(to_sfixed_a(-0.004354189150035381)),(to_sfixed_a(0.14611941576004028)),(to_sfixed_a(-0.005805212073028088)),(to_sfixed_a(-0.00012123692431487143)),(to_sfixed_a(-0.10473925620317459)),(to_sfixed_a(-0.02164047583937645)),(to_sfixed_a(0.09106216579675674)),(to_sfixed_a(0.09423872828483582)),(to_sfixed_a(-0.0495414212346077)),(to_sfixed_a(0.25307950377464294)),(to_sfixed_a(0.03747854009270668)),(to_sfixed_a(-0.13939811289310455)),(to_sfixed_a(0.08381381630897522)),(to_sfixed_a(0.18265843391418457)),(to_sfixed_a(0.11421693861484528)),(to_sfixed_a(0.02418593131005764)),(to_sfixed_a(0.09258756786584854)),(to_sfixed_a(0.09186826646327972)),(to_sfixed_a(-0.028416495770215988)));

    constant weight_n1_36 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.1969679594039917)),(to_sfixed_a(-0.023562146350741386)),(to_sfixed_a(0.04813019931316376)),(to_sfixed_a(-0.018805375322699547)),(to_sfixed_a(-0.09569092094898224)),(to_sfixed_a(-0.03342907130718231)),(to_sfixed_a(-0.04546603932976723)),(to_sfixed_a(-0.051499564200639725)),(to_sfixed_a(-0.1274101287126541)),(to_sfixed_a(-0.0829262062907219)),(to_sfixed_a(-0.01686328835785389)),(to_sfixed_a(-0.17458882927894592)),(to_sfixed_a(-0.18324129283428192)),(to_sfixed_a(-0.09665994346141815)),(to_sfixed_a(0.05041399970650673)),(to_sfixed_a(-0.04245014116168022)),(to_sfixed_a(-0.14277544617652893)),(to_sfixed_a(-0.06258630007505417)),(to_sfixed_a(-0.14937861263751984)),(to_sfixed_a(-0.06661131232976913)),(to_sfixed_a(-0.1402312070131302)),(to_sfixed_a(0.004864975810050964)),(to_sfixed_a(0.052382539957761765)),(to_sfixed_a(-0.10487286746501923)),(to_sfixed_a(0.05524652078747749)),(to_sfixed_a(0.032155510038137436)),(to_sfixed_a(-0.07688811421394348)),(to_sfixed_a(0.05077815800905228)),(to_sfixed_a(-0.10355206578969955)),(to_sfixed_a(0.2109440714120865)),(to_sfixed_a(0.0680193230509758)),(to_sfixed_a(-0.09365606307983398)),(to_sfixed_a(0.17317543923854828)),(to_sfixed_a(-0.14829854667186737)),(to_sfixed_a(0.12366043776273727)),(to_sfixed_a(0.08200504630804062)),(to_sfixed_a(0.06406833231449127)),(to_sfixed_a(-0.03026602976024151)));

    constant weight_n1_37 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.21724003553390503)),(to_sfixed_a(-0.0830828920006752)),(to_sfixed_a(0.12312456220388412)),(to_sfixed_a(-0.11865510791540146)),(to_sfixed_a(-0.07917425781488419)),(to_sfixed_a(0.05279242619872093)),(to_sfixed_a(0.11145859211683273)),(to_sfixed_a(-0.01838619075715542)),(to_sfixed_a(-0.007057107053697109)),(to_sfixed_a(-0.0621245838701725)),(to_sfixed_a(-0.037252675741910934)),(to_sfixed_a(-0.05990028753876686)),(to_sfixed_a(0.15777328610420227)),(to_sfixed_a(0.010463882237672806)),(to_sfixed_a(0.11425227671861649)),(to_sfixed_a(0.24053162336349487)),(to_sfixed_a(0.1770331859588623)),(to_sfixed_a(-0.045516613870859146)),(to_sfixed_a(0.04325200617313385)),(to_sfixed_a(-0.014030414633452892)),(to_sfixed_a(-0.05067521333694458)),(to_sfixed_a(0.092072993516922)),(to_sfixed_a(-0.11903581023216248)),(to_sfixed_a(-0.026314137503504753)),(to_sfixed_a(0.002687961794435978)),(to_sfixed_a(-0.05045778676867485)),(to_sfixed_a(0.083379827439785)),(to_sfixed_a(0.045749861747026443)),(to_sfixed_a(-0.07632926106452942)),(to_sfixed_a(0.10182711482048035)),(to_sfixed_a(-0.017802515998482704)),(to_sfixed_a(0.1311885118484497)),(to_sfixed_a(-0.0557418018579483)),(to_sfixed_a(-0.06105785444378853)),(to_sfixed_a(-0.020344581454992294)),(to_sfixed_a(0.07985810935497284)),(to_sfixed_a(-0.0006487221689894795)),(to_sfixed_a(-0.07559531182050705)));

    constant weight_n1_38 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.07529427856206894)),(to_sfixed_a(1.257499388884753e-05)),(to_sfixed_a(-1.7508273231214844e-05)),(to_sfixed_a(-4.036695827380754e-05)),(to_sfixed_a(4.92162726004608e-05)),(to_sfixed_a(-4.9153506552102044e-05)),(to_sfixed_a(3.178022234351374e-05)),(to_sfixed_a(-2.9284952688612975e-05)),(to_sfixed_a(3.423225280130282e-05)),(to_sfixed_a(-4.121899837628007e-05)),(to_sfixed_a(-1.0566311203774603e-07)),(to_sfixed_a(7.622778412041953e-06)),(to_sfixed_a(1.4071826626604889e-05)),(to_sfixed_a(1.7301103071076795e-05)),(to_sfixed_a(7.243552681757137e-05)),(to_sfixed_a(-2.3565198716823943e-05)),(to_sfixed_a(-1.4556328096659854e-05)),(to_sfixed_a(6.261483940761536e-05)),(to_sfixed_a(1.2447236258594785e-05)),(to_sfixed_a(-6.673907046206295e-05)),(to_sfixed_a(-4.33251989306882e-05)),(to_sfixed_a(6.989594112383202e-05)),(to_sfixed_a(-2.6877280106418766e-05)),(to_sfixed_a(-1.4323519280878827e-05)),(to_sfixed_a(2.775857319647912e-05)),(to_sfixed_a(8.298218745039776e-06)),(to_sfixed_a(-2.2407612050301395e-06)),(to_sfixed_a(-1.1878253644681536e-05)),(to_sfixed_a(6.939073500689119e-05)),(to_sfixed_a(-1.4122284483164549e-05)),(to_sfixed_a(2.3754339053994045e-05)),(to_sfixed_a(3.900226511177607e-05)),(to_sfixed_a(3.439900683588348e-05)),(to_sfixed_a(-1.531933776277583e-05)),(to_sfixed_a(-4.359484955784865e-05)),(to_sfixed_a(-8.412573515670374e-05)),(to_sfixed_a(6.216629117261618e-05)),(to_sfixed_a(-8.668027294334024e-05)));

    constant weight_n1_39 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.005447335075587034)),(to_sfixed_a(0.03176552429795265)),(to_sfixed_a(0.011874721385538578)),(to_sfixed_a(0.08859079331159592)),(to_sfixed_a(0.031830959022045135)),(to_sfixed_a(-0.020778479054570198)),(to_sfixed_a(0.017186889424920082)),(to_sfixed_a(-0.12079209834337234)),(to_sfixed_a(-0.0073029357008636)),(to_sfixed_a(-0.12838466465473175)),(to_sfixed_a(-0.07314012944698334)),(to_sfixed_a(-0.10089340806007385)),(to_sfixed_a(0.08662039786577225)),(to_sfixed_a(0.04296726733446121)),(to_sfixed_a(0.09789104014635086)),(to_sfixed_a(0.006262415088713169)),(to_sfixed_a(-0.10590158402919769)),(to_sfixed_a(0.058560024946928024)),(to_sfixed_a(-0.14494550228118896)),(to_sfixed_a(0.025425666943192482)),(to_sfixed_a(0.15769317746162415)),(to_sfixed_a(-0.01877489872276783)),(to_sfixed_a(0.1201431080698967)),(to_sfixed_a(0.07266348600387573)),(to_sfixed_a(-0.06436872482299805)),(to_sfixed_a(-0.12440609186887741)),(to_sfixed_a(0.08756478130817413)),(to_sfixed_a(0.14958156645298004)),(to_sfixed_a(-0.05129335820674896)),(to_sfixed_a(-0.12455559521913528)),(to_sfixed_a(0.07112924009561539)),(to_sfixed_a(0.03057227097451687)),(to_sfixed_a(0.07679451256990433)),(to_sfixed_a(0.04209667071700096)),(to_sfixed_a(-0.10879042744636536)),(to_sfixed_a(-0.013581089675426483)),(to_sfixed_a(0.04278257489204407)),(to_sfixed_a(0.16500958800315857)));

    constant weight_n1_40 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.19035765528678894)),(to_sfixed_a(0.0712362602353096)),(to_sfixed_a(-0.0474146232008934)),(to_sfixed_a(0.011187578551471233)),(to_sfixed_a(0.08258998394012451)),(to_sfixed_a(-0.04196404293179512)),(to_sfixed_a(0.09632021933794022)),(to_sfixed_a(-0.045297134667634964)),(to_sfixed_a(0.09210360050201416)),(to_sfixed_a(-0.06220036372542381)),(to_sfixed_a(-0.058583248406648636)),(to_sfixed_a(-0.06593438237905502)),(to_sfixed_a(-0.023179957643151283)),(to_sfixed_a(0.018090257421135902)),(to_sfixed_a(-0.0012808497995138168)),(to_sfixed_a(0.11071993410587311)),(to_sfixed_a(-0.09738405793905258)),(to_sfixed_a(-0.17397870123386383)),(to_sfixed_a(0.06015748530626297)),(to_sfixed_a(-0.12033428996801376)),(to_sfixed_a(-0.08908093720674515)),(to_sfixed_a(-0.0004710886860266328)),(to_sfixed_a(0.0523342527449131)),(to_sfixed_a(-0.04938710480928421)),(to_sfixed_a(-0.06273023039102554)),(to_sfixed_a(0.09302904456853867)),(to_sfixed_a(-0.06309803575277328)),(to_sfixed_a(0.07426442205905914)),(to_sfixed_a(-0.005050717853009701)),(to_sfixed_a(-0.13057921826839447)),(to_sfixed_a(0.21305492520332336)),(to_sfixed_a(0.08631724864244461)),(to_sfixed_a(-0.15073128044605255)),(to_sfixed_a(-0.08080693334341049)),(to_sfixed_a(-0.015099374577403069)),(to_sfixed_a(-0.20545001327991486)),(to_sfixed_a(-0.057075198739767075)),(to_sfixed_a(0.12315377593040466)));

    constant weight_n1_41 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.07074088603258133)),(to_sfixed_a(-1.1136384273413569e-05)),(to_sfixed_a(2.3032807803247124e-06)),(to_sfixed_a(6.21457802481018e-05)),(to_sfixed_a(-1.0603248483675998e-05)),(to_sfixed_a(-1.8114766135113314e-05)),(to_sfixed_a(2.1356945580919273e-05)),(to_sfixed_a(3.881518932757899e-05)),(to_sfixed_a(1.56582027557306e-05)),(to_sfixed_a(-6.788881728425622e-05)),(to_sfixed_a(3.079372618230991e-05)),(to_sfixed_a(-1.1915567483811174e-05)),(to_sfixed_a(2.7830241378978826e-05)),(to_sfixed_a(4.340694795246236e-05)),(to_sfixed_a(6.432284408219857e-06)),(to_sfixed_a(1.843018617364578e-05)),(to_sfixed_a(1.4763693798158783e-05)),(to_sfixed_a(-2.2628935766988434e-05)),(to_sfixed_a(-4.58344875369221e-05)),(to_sfixed_a(-4.291859295335598e-05)),(to_sfixed_a(-7.232828465930652e-06)),(to_sfixed_a(-3.6274843296268955e-05)),(to_sfixed_a(-7.693447696510702e-05)),(to_sfixed_a(1.9655594769574236e-06)),(to_sfixed_a(2.6932051696348935e-05)),(to_sfixed_a(-2.9416185498121195e-05)),(to_sfixed_a(-3.31504998030141e-05)),(to_sfixed_a(-1.1903231097676326e-05)),(to_sfixed_a(2.3050004529068246e-05)),(to_sfixed_a(5.124485323904082e-05)),(to_sfixed_a(-3.44292311638128e-05)),(to_sfixed_a(3.55052288796287e-05)),(to_sfixed_a(1.3040909834671766e-05)),(to_sfixed_a(7.2811981226550415e-06)),(to_sfixed_a(-8.288447133963928e-06)),(to_sfixed_a(-7.267398905241862e-05)),(to_sfixed_a(-6.591018063772935e-06)),(to_sfixed_a(1.5874169548624195e-05)));

    constant weight_n1_42 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.016628872603178024)),(to_sfixed_a(-3.116691732429899e-05)),(to_sfixed_a(1.990583405131474e-05)),(to_sfixed_a(1.2032897757308092e-05)),(to_sfixed_a(-2.409979424555786e-05)),(to_sfixed_a(1.5213465303531848e-05)),(to_sfixed_a(-1.68857368407771e-05)),(to_sfixed_a(-1.9488830730551854e-05)),(to_sfixed_a(6.446055340347812e-05)),(to_sfixed_a(-6.814537482568994e-05)),(to_sfixed_a(-6.222318461368559e-06)),(to_sfixed_a(-3.7548696127487347e-05)),(to_sfixed_a(-8.193397661671042e-06)),(to_sfixed_a(-2.3281685571419075e-05)),(to_sfixed_a(-1.9495873857522383e-05)),(to_sfixed_a(3.0426259399973787e-05)),(to_sfixed_a(-1.4297259440354537e-05)),(to_sfixed_a(-3.755724537768401e-05)),(to_sfixed_a(-1.2580611837620381e-05)),(to_sfixed_a(-3.76414718630258e-05)),(to_sfixed_a(1.8566755898064002e-05)),(to_sfixed_a(5.849020817549899e-05)),(to_sfixed_a(-6.003387534292415e-05)),(to_sfixed_a(8.549684935132973e-06)),(to_sfixed_a(-9.480377229920123e-06)),(to_sfixed_a(-1.3130812476447318e-05)),(to_sfixed_a(2.4400285383308074e-06)),(to_sfixed_a(-1.7738451788318343e-05)),(to_sfixed_a(3.9057620597304776e-05)),(to_sfixed_a(-1.049397724273149e-05)),(to_sfixed_a(-1.702739973552525e-05)),(to_sfixed_a(4.5709813889516226e-07)),(to_sfixed_a(7.967960300447885e-06)),(to_sfixed_a(-5.195047560846433e-05)),(to_sfixed_a(5.618398790829815e-05)),(to_sfixed_a(-0.00011629271466517821)),(to_sfixed_a(-8.128946319629904e-06)),(to_sfixed_a(-8.360447100130841e-05)));

    constant weight_n1_43 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.04591955617070198)),(to_sfixed_a(-0.006019068881869316)),(to_sfixed_a(0.024652767926454544)),(to_sfixed_a(0.017296945676207542)),(to_sfixed_a(0.04804329574108124)),(to_sfixed_a(-0.027763977646827698)),(to_sfixed_a(-0.008599646389484406)),(to_sfixed_a(0.057126160711050034)),(to_sfixed_a(0.006229812279343605)),(to_sfixed_a(-0.005852032452821732)),(to_sfixed_a(0.009643700905144215)),(to_sfixed_a(0.007807569578289986)),(to_sfixed_a(-0.013624398037791252)),(to_sfixed_a(0.025606930255889893)),(to_sfixed_a(-0.0029661175794899464)),(to_sfixed_a(-0.014068392105400562)),(to_sfixed_a(-0.037053145468235016)),(to_sfixed_a(0.011286848224699497)),(to_sfixed_a(0.0034929097164422274)),(to_sfixed_a(0.04228723421692848)),(to_sfixed_a(0.009666410274803638)),(to_sfixed_a(0.00280143809504807)),(to_sfixed_a(0.018840203061699867)),(to_sfixed_a(0.02021194063127041)),(to_sfixed_a(0.01404003519564867)),(to_sfixed_a(-0.024166306480765343)),(to_sfixed_a(0.018169119954109192)),(to_sfixed_a(0.030653493478894234)),(to_sfixed_a(0.0357915498316288)),(to_sfixed_a(-0.0243237167596817)),(to_sfixed_a(-0.01969417929649353)),(to_sfixed_a(-0.04793092980980873)),(to_sfixed_a(-0.01237817108631134)),(to_sfixed_a(-0.042249999940395355)),(to_sfixed_a(0.02081766165792942)),(to_sfixed_a(0.025766318663954735)),(to_sfixed_a(0.01245255209505558)),(to_sfixed_a(-0.00986251700669527)));

    constant weight_n1_44 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.31902381777763367)),(to_sfixed_a(-0.13066089153289795)),(to_sfixed_a(-0.1932963877916336)),(to_sfixed_a(-0.005310842301696539)),(to_sfixed_a(0.08940067887306213)),(to_sfixed_a(0.010344060137867928)),(to_sfixed_a(-0.09279582649469376)),(to_sfixed_a(0.034155577421188354)),(to_sfixed_a(0.041580237448215485)),(to_sfixed_a(-0.08445735275745392)),(to_sfixed_a(-0.07952895015478134)),(to_sfixed_a(-0.03987893834710121)),(to_sfixed_a(-0.004737135488539934)),(to_sfixed_a(0.05098966509103775)),(to_sfixed_a(0.02454468235373497)),(to_sfixed_a(-0.16849656403064728)),(to_sfixed_a(0.12362257391214371)),(to_sfixed_a(0.034282926470041275)),(to_sfixed_a(-0.08480673283338547)),(to_sfixed_a(0.11479376256465912)),(to_sfixed_a(-0.17924655973911285)),(to_sfixed_a(-0.06336116790771484)),(to_sfixed_a(-0.018005408346652985)),(to_sfixed_a(0.0721311941742897)),(to_sfixed_a(0.02525591105222702)),(to_sfixed_a(-0.21789856255054474)),(to_sfixed_a(0.14568409323692322)),(to_sfixed_a(0.11774767935276031)),(to_sfixed_a(-0.02313559129834175)),(to_sfixed_a(0.1842147260904312)),(to_sfixed_a(0.056712206453084946)),(to_sfixed_a(-0.0871763601899147)),(to_sfixed_a(-0.09078650921583176)),(to_sfixed_a(-0.1119469478726387)),(to_sfixed_a(0.016146454960107803)),(to_sfixed_a(0.02442394196987152)),(to_sfixed_a(0.04883508384227753)),(to_sfixed_a(0.04966847226023674)));

    constant weight_n1_45 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.3637908399105072)),(to_sfixed_a(-0.27260637283325195)),(to_sfixed_a(0.24570417404174805)),(to_sfixed_a(-0.2552320063114166)),(to_sfixed_a(-0.015071036294102669)),(to_sfixed_a(0.10524673759937286)),(to_sfixed_a(-0.027073057368397713)),(to_sfixed_a(0.04720490798354149)),(to_sfixed_a(0.08305120468139648)),(to_sfixed_a(-0.09043554961681366)),(to_sfixed_a(0.052276767790317535)),(to_sfixed_a(0.11976628750562668)),(to_sfixed_a(0.2147028148174286)),(to_sfixed_a(-0.13471294939517975)),(to_sfixed_a(0.14680492877960205)),(to_sfixed_a(-0.05424348637461662)),(to_sfixed_a(-0.1813412308692932)),(to_sfixed_a(-0.09707316756248474)),(to_sfixed_a(0.03933604434132576)),(to_sfixed_a(-0.20822370052337646)),(to_sfixed_a(-0.22619445621967316)),(to_sfixed_a(-0.21064379811286926)),(to_sfixed_a(0.0593440942466259)),(to_sfixed_a(0.017107142135500908)),(to_sfixed_a(-0.002487629884853959)),(to_sfixed_a(-0.02539048157632351)),(to_sfixed_a(0.09067685902118683)),(to_sfixed_a(0.19321851432323456)),(to_sfixed_a(0.06425876915454865)),(to_sfixed_a(-0.24372194707393646)),(to_sfixed_a(0.052608758211135864)),(to_sfixed_a(-0.10943981260061264)),(to_sfixed_a(0.12083129584789276)),(to_sfixed_a(0.04761389642953873)),(to_sfixed_a(0.11842193454504013)),(to_sfixed_a(-0.010431399568915367)),(to_sfixed_a(-0.05165313184261322)),(to_sfixed_a(0.10119504481554031)));

    constant weight_n1_46 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.003668233286589384)),(to_sfixed_a(0.04517177864909172)),(to_sfixed_a(-0.0030414476059377193)),(to_sfixed_a(-0.06320370733737946)),(to_sfixed_a(0.1397736519575119)),(to_sfixed_a(0.01422558818012476)),(to_sfixed_a(0.020823026075959206)),(to_sfixed_a(-0.000540149980224669)),(to_sfixed_a(-0.15058748424053192)),(to_sfixed_a(-0.059634730219841)),(to_sfixed_a(0.11421829462051392)),(to_sfixed_a(0.07754401862621307)),(to_sfixed_a(-0.0798465758562088)),(to_sfixed_a(0.022587725892663002)),(to_sfixed_a(0.073069728910923)),(to_sfixed_a(0.057980943471193314)),(to_sfixed_a(0.02662649378180504)),(to_sfixed_a(-0.02519812062382698)),(to_sfixed_a(-0.03421357646584511)),(to_sfixed_a(0.017690692096948624)),(to_sfixed_a(0.02040327712893486)),(to_sfixed_a(0.005865143612027168)),(to_sfixed_a(0.0546991229057312)),(to_sfixed_a(-0.06983654201030731)),(to_sfixed_a(-0.013366534374654293)),(to_sfixed_a(0.06980616599321365)),(to_sfixed_a(0.06934813410043716)),(to_sfixed_a(-0.05272345989942551)),(to_sfixed_a(-0.03806633874773979)),(to_sfixed_a(0.033846404403448105)),(to_sfixed_a(0.010210301727056503)),(to_sfixed_a(0.023337559774518013)),(to_sfixed_a(-0.10210350900888443)),(to_sfixed_a(0.0245202649384737)),(to_sfixed_a(0.1335236132144928)),(to_sfixed_a(-0.0774962529540062)),(to_sfixed_a(0.11462164670228958)),(to_sfixed_a(0.09108658879995346)));

    constant weight_n1_47 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.008255274035036564)),(to_sfixed_a(-1.7454147382522933e-05)),(to_sfixed_a(-3.652965460787527e-05)),(to_sfixed_a(-1.2472884009184781e-05)),(to_sfixed_a(-6.926149217179045e-05)),(to_sfixed_a(-5.9510613937163725e-05)),(to_sfixed_a(8.844373951433226e-06)),(to_sfixed_a(5.076039815321565e-05)),(to_sfixed_a(-3.756415389943868e-05)),(to_sfixed_a(-6.673573079751804e-05)),(to_sfixed_a(-0.00010963603563141078)),(to_sfixed_a(-8.509698091074824e-06)),(to_sfixed_a(-2.2087799152359366e-05)),(to_sfixed_a(3.166804162901826e-05)),(to_sfixed_a(-1.000483644020278e-05)),(to_sfixed_a(1.902916847029701e-05)),(to_sfixed_a(-2.629732625791803e-05)),(to_sfixed_a(7.502786320401356e-05)),(to_sfixed_a(2.4789980670902878e-05)),(to_sfixed_a(8.349100426130462e-06)),(to_sfixed_a(6.815762026235461e-05)),(to_sfixed_a(-8.141465514199808e-05)),(to_sfixed_a(-6.065577053959714e-06)),(to_sfixed_a(-7.613841444253922e-05)),(to_sfixed_a(-1.6098356354632415e-05)),(to_sfixed_a(-4.5091004722053185e-05)),(to_sfixed_a(-3.5670422221301123e-05)),(to_sfixed_a(3.704526989167789e-06)),(to_sfixed_a(-0.0001567739964229986)),(to_sfixed_a(-5.4356432883651e-06)),(to_sfixed_a(-2.3046659407555126e-05)),(to_sfixed_a(7.839973841328174e-05)),(to_sfixed_a(-2.3308683012146503e-05)),(to_sfixed_a(4.462726428755559e-05)),(to_sfixed_a(8.890311437426135e-05)),(to_sfixed_a(-1.175810848508263e-05)),(to_sfixed_a(2.419724660285283e-05)),(to_sfixed_a(-1.8489887224859558e-05)));

    constant weight_n1_48 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.0865718200802803)),(to_sfixed_a(0.05380266159772873)),(to_sfixed_a(-0.03508531674742699)),(to_sfixed_a(-0.027473723515868187)),(to_sfixed_a(0.05875749513506889)),(to_sfixed_a(0.01581818424165249)),(to_sfixed_a(-0.04746084660291672)),(to_sfixed_a(0.007051297463476658)),(to_sfixed_a(0.007614086382091045)),(to_sfixed_a(-0.05781165510416031)),(to_sfixed_a(0.05471361428499222)),(to_sfixed_a(-0.08766044676303864)),(to_sfixed_a(0.04486279934644699)),(to_sfixed_a(0.01739463582634926)),(to_sfixed_a(-0.0024155813734978437)),(to_sfixed_a(0.023940715938806534)),(to_sfixed_a(-0.11536595225334167)),(to_sfixed_a(-0.014375580474734306)),(to_sfixed_a(0.13369916379451752)),(to_sfixed_a(-0.07562269270420074)),(to_sfixed_a(-0.03691559657454491)),(to_sfixed_a(0.0987640768289566)),(to_sfixed_a(-0.018896419554948807)),(to_sfixed_a(0.015363910235464573)),(to_sfixed_a(-0.03959064930677414)),(to_sfixed_a(0.06605804711580276)),(to_sfixed_a(0.025451350957155228)),(to_sfixed_a(0.006133111659437418)),(to_sfixed_a(0.13998708128929138)),(to_sfixed_a(-0.1363014578819275)),(to_sfixed_a(-0.05189758166670799)),(to_sfixed_a(-0.02145485207438469)),(to_sfixed_a(-0.05682006850838661)),(to_sfixed_a(0.02733294852077961)),(to_sfixed_a(0.06266630440950394)),(to_sfixed_a(0.06621068716049194)),(to_sfixed_a(0.019259633496403694)),(to_sfixed_a(-0.036333631724119186)));

    constant weight_n1_49 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.06879878044128418)),(to_sfixed_a(-0.02184416353702545)),(to_sfixed_a(-0.05555183067917824)),(to_sfixed_a(0.10928759723901749)),(to_sfixed_a(0.1257307082414627)),(to_sfixed_a(0.012817745096981525)),(to_sfixed_a(-0.029825789853930473)),(to_sfixed_a(0.0021621997002512217)),(to_sfixed_a(0.0856555700302124)),(to_sfixed_a(0.03673386573791504)),(to_sfixed_a(-0.046070635318756104)),(to_sfixed_a(0.11104404181241989)),(to_sfixed_a(0.039827313274145126)),(to_sfixed_a(-0.03551766276359558)),(to_sfixed_a(0.01550880167633295)),(to_sfixed_a(-0.10853254050016403)),(to_sfixed_a(0.11559148877859116)),(to_sfixed_a(0.08091959357261658)),(to_sfixed_a(-0.014973100274801254)),(to_sfixed_a(-0.08364160358905792)),(to_sfixed_a(0.023800693452358246)),(to_sfixed_a(0.00010039465996669605)),(to_sfixed_a(-0.13145548105239868)),(to_sfixed_a(-0.13312044739723206)),(to_sfixed_a(0.017449427396059036)),(to_sfixed_a(0.14481452107429504)),(to_sfixed_a(0.2771148383617401)),(to_sfixed_a(-0.06971599161624908)),(to_sfixed_a(-0.15377067029476166)),(to_sfixed_a(-0.07743644714355469)),(to_sfixed_a(0.04837915301322937)),(to_sfixed_a(0.009075003676116467)),(to_sfixed_a(0.09165150672197342)),(to_sfixed_a(0.10190025717020035)),(to_sfixed_a(-0.020522378385066986)),(to_sfixed_a(0.01584729738533497)),(to_sfixed_a(-0.07755915075540543)),(to_sfixed_a(0.003117790212854743)));

    constant weight_n1_50 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.046556148678064346)),(to_sfixed_a(-0.0045740543864667416)),(to_sfixed_a(0.00624446477741003)),(to_sfixed_a(-0.0009423682931810617)),(to_sfixed_a(-0.010138963349163532)),(to_sfixed_a(0.003856709459796548)),(to_sfixed_a(0.003176681697368622)),(to_sfixed_a(-0.00930843222886324)),(to_sfixed_a(-0.0012746058637276292)),(to_sfixed_a(0.000237318774452433)),(to_sfixed_a(-0.0033976167906075716)),(to_sfixed_a(0.007011029869318008)),(to_sfixed_a(0.0021447420585900545)),(to_sfixed_a(0.010356724262237549)),(to_sfixed_a(0.0036268215626478195)),(to_sfixed_a(-0.003588844323530793)),(to_sfixed_a(0.005706583149731159)),(to_sfixed_a(0.007534582633525133)),(to_sfixed_a(-0.008864904753863811)),(to_sfixed_a(0.006672775838524103)),(to_sfixed_a(0.002503161784261465)),(to_sfixed_a(0.00959249958395958)),(to_sfixed_a(0.001847867970354855)),(to_sfixed_a(-0.00967900175601244)),(to_sfixed_a(0.0020734071731567383)),(to_sfixed_a(-0.006500616203993559)),(to_sfixed_a(-0.00558808958157897)),(to_sfixed_a(-0.006173222791403532)),(to_sfixed_a(-0.006481187883764505)),(to_sfixed_a(0.006462775636464357)),(to_sfixed_a(0.003601294243708253)),(to_sfixed_a(-0.004404537845402956)),(to_sfixed_a(0.0007996528293006122)),(to_sfixed_a(-0.005978450644761324)),(to_sfixed_a(-0.003051137551665306)),(to_sfixed_a(-0.001424587913788855)),(to_sfixed_a(0.01193538960069418)),(to_sfixed_a(0.008373433724045753)));

    constant weight_n1_51 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.028812238946557045)),(to_sfixed_a(7.187318260548636e-06)),(to_sfixed_a(6.378349553415319e-06)),(to_sfixed_a(5.5306973081314936e-05)),(to_sfixed_a(4.25440157414414e-05)),(to_sfixed_a(3.384747469681315e-05)),(to_sfixed_a(-2.550808130763471e-05)),(to_sfixed_a(2.664199928403832e-05)),(to_sfixed_a(7.215738878585398e-05)),(to_sfixed_a(4.132587946514832e-06)),(to_sfixed_a(9.393978217531185e-08)),(to_sfixed_a(-0.00019051962590310723)),(to_sfixed_a(-4.024009103886783e-05)),(to_sfixed_a(1.2579783287947066e-05)),(to_sfixed_a(-4.9817859689937904e-05)),(to_sfixed_a(-3.8456513721030205e-05)),(to_sfixed_a(3.178180122631602e-05)),(to_sfixed_a(7.058263872750103e-05)),(to_sfixed_a(2.5159633878502063e-05)),(to_sfixed_a(-8.972010255092755e-05)),(to_sfixed_a(9.030304499901831e-05)),(to_sfixed_a(8.282008639071137e-05)),(to_sfixed_a(-0.00011355707101756707)),(to_sfixed_a(-6.450121145462617e-05)),(to_sfixed_a(-5.058685565018095e-05)),(to_sfixed_a(6.446316547226161e-05)),(to_sfixed_a(-4.2950374336214736e-05)),(to_sfixed_a(0.00010296962136635557)),(to_sfixed_a(-2.5168330921587767e-06)),(to_sfixed_a(-6.476483395090327e-05)),(to_sfixed_a(-3.180062412866391e-05)),(to_sfixed_a(-1.4555011148331687e-05)),(to_sfixed_a(-3.062988616875373e-05)),(to_sfixed_a(-4.541494854493067e-05)),(to_sfixed_a(8.579315181123093e-05)),(to_sfixed_a(3.725360511452891e-05)),(to_sfixed_a(5.547815453610383e-05)),(to_sfixed_a(0.00011295845615677536)));

    constant weight_n1_52 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.09906929731369019)),(to_sfixed_a(-0.013828490860760212)),(to_sfixed_a(0.03232914209365845)),(to_sfixed_a(0.0012734465999528766)),(to_sfixed_a(-0.045018866658210754)),(to_sfixed_a(0.020669279620051384)),(to_sfixed_a(0.018014784902334213)),(to_sfixed_a(-0.029787147417664528)),(to_sfixed_a(-0.015921344980597496)),(to_sfixed_a(0.013763039372861385)),(to_sfixed_a(0.007778429426252842)),(to_sfixed_a(-0.0012704102555289865)),(to_sfixed_a(-0.014625107869505882)),(to_sfixed_a(-0.003916620276868343)),(to_sfixed_a(0.004620376508682966)),(to_sfixed_a(0.03086179308593273)),(to_sfixed_a(0.050294701009988785)),(to_sfixed_a(0.00923096388578415)),(to_sfixed_a(-0.005462046712636948)),(to_sfixed_a(0.030839044600725174)),(to_sfixed_a(0.004049544222652912)),(to_sfixed_a(0.0029380584601312876)),(to_sfixed_a(0.020242616534233093)),(to_sfixed_a(-0.0032254555262625217)),(to_sfixed_a(0.005735295824706554)),(to_sfixed_a(-0.013185480609536171)),(to_sfixed_a(-0.036168910562992096)),(to_sfixed_a(0.015001952648162842)),(to_sfixed_a(0.02360905148088932)),(to_sfixed_a(0.009613418951630592)),(to_sfixed_a(0.0467267669737339)),(to_sfixed_a(-0.050084274262189865)),(to_sfixed_a(0.01643509976565838)),(to_sfixed_a(-0.0257077869027853)),(to_sfixed_a(-0.004352719988673925)),(to_sfixed_a(-0.04816149175167084)),(to_sfixed_a(0.029103856533765793)),(to_sfixed_a(0.02643240988254547)));

    constant weight_n1_53 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.1588367074728012)),(to_sfixed_a(0.00392673397436738)),(to_sfixed_a(0.015412647277116776)),(to_sfixed_a(0.008701098151504993)),(to_sfixed_a(0.0019151346059516072)),(to_sfixed_a(-0.0629575103521347)),(to_sfixed_a(0.0048899720422923565)),(to_sfixed_a(-0.017888857051730156)),(to_sfixed_a(-0.03479403257369995)),(to_sfixed_a(-0.006186309736222029)),(to_sfixed_a(0.07444296777248383)),(to_sfixed_a(-0.04322582855820656)),(to_sfixed_a(0.03301096707582474)),(to_sfixed_a(-0.00961823109537363)),(to_sfixed_a(-0.09236541390419006)),(to_sfixed_a(-0.12522797286510468)),(to_sfixed_a(-0.13288401067256927)),(to_sfixed_a(0.049091726541519165)),(to_sfixed_a(0.125693678855896)),(to_sfixed_a(-0.13603445887565613)),(to_sfixed_a(-0.01544299628585577)),(to_sfixed_a(0.11120094358921051)),(to_sfixed_a(0.22091946005821228)),(to_sfixed_a(0.05834302678704262)),(to_sfixed_a(0.02883720025420189)),(to_sfixed_a(0.1726359724998474)),(to_sfixed_a(0.09974091500043869)),(to_sfixed_a(-0.0008951641502790153)),(to_sfixed_a(0.04969292879104614)),(to_sfixed_a(0.008089719340205193)),(to_sfixed_a(-0.06984858959913254)),(to_sfixed_a(-0.10471175611019135)),(to_sfixed_a(-0.16862592101097107)),(to_sfixed_a(-0.009859182871878147)),(to_sfixed_a(0.0016617468791082501)),(to_sfixed_a(0.04378673434257507)),(to_sfixed_a(0.030847325921058655)),(to_sfixed_a(0.1198035255074501)));

    constant weight_n1_54 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.06439045071601868)),(to_sfixed_a(-0.0221538245677948)),(to_sfixed_a(0.04477155581116676)),(to_sfixed_a(-0.010537512600421906)),(to_sfixed_a(-0.06680066138505936)),(to_sfixed_a(0.005808650981634855)),(to_sfixed_a(0.05626033991575241)),(to_sfixed_a(-0.05405452102422714)),(to_sfixed_a(-0.05554937943816185)),(to_sfixed_a(0.008701354265213013)),(to_sfixed_a(-0.02520664408802986)),(to_sfixed_a(-0.010151025839149952)),(to_sfixed_a(-0.0022329981438815594)),(to_sfixed_a(0.028753094375133514)),(to_sfixed_a(0.011840506456792355)),(to_sfixed_a(0.13305820524692535)),(to_sfixed_a(0.03856610506772995)),(to_sfixed_a(0.04712958633899689)),(to_sfixed_a(0.07668253779411316)),(to_sfixed_a(-0.014897888526320457)),(to_sfixed_a(0.016705287620425224)),(to_sfixed_a(0.14449690282344818)),(to_sfixed_a(0.02117280475795269)),(to_sfixed_a(-0.0032565398141741753)),(to_sfixed_a(0.037255339324474335)),(to_sfixed_a(0.009827584028244019)),(to_sfixed_a(-0.0125424824655056)),(to_sfixed_a(-0.09012318402528763)),(to_sfixed_a(-0.053176749497652054)),(to_sfixed_a(-0.005178491584956646)),(to_sfixed_a(-0.07197076827287674)),(to_sfixed_a(-0.10460113734006882)),(to_sfixed_a(0.038315463811159134)),(to_sfixed_a(-0.011927434243261814)),(to_sfixed_a(-0.02097705751657486)),(to_sfixed_a(-0.06491109728813171)),(to_sfixed_a(-0.012887990102171898)),(to_sfixed_a(-0.01913096196949482)));

    constant weight_n1_55 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.00712354714050889)),(to_sfixed_a(-4.869938129559159e-05)),(to_sfixed_a(-4.280691427993588e-05)),(to_sfixed_a(-4.850503955822205e-06)),(to_sfixed_a(6.570303412445355e-06)),(to_sfixed_a(3.998699685325846e-05)),(to_sfixed_a(1.938427158165723e-05)),(to_sfixed_a(3.7052639527246356e-05)),(to_sfixed_a(-3.281294630141929e-05)),(to_sfixed_a(2.9780037948512472e-05)),(to_sfixed_a(2.3910410163807683e-05)),(to_sfixed_a(-5.047244485467672e-06)),(to_sfixed_a(2.9889797588111833e-05)),(to_sfixed_a(7.026300590950996e-05)),(to_sfixed_a(-6.631483847741038e-05)),(to_sfixed_a(5.4235839343164116e-05)),(to_sfixed_a(-5.271449845167808e-05)),(to_sfixed_a(5.200839223107323e-05)),(to_sfixed_a(2.8678674425464123e-05)),(to_sfixed_a(5.0790182285709307e-05)),(to_sfixed_a(1.0394325727247633e-05)),(to_sfixed_a(-6.320040483842604e-06)),(to_sfixed_a(-1.5741976312710904e-05)),(to_sfixed_a(-9.762735317053739e-06)),(to_sfixed_a(-2.757904258032795e-05)),(to_sfixed_a(4.316773629398085e-05)),(to_sfixed_a(5.7276582083432004e-05)),(to_sfixed_a(-3.5545228456612676e-05)),(to_sfixed_a(-8.909736607165541e-06)),(to_sfixed_a(-1.4095413689574343e-06)),(to_sfixed_a(4.5120214053895324e-05)),(to_sfixed_a(5.8194855228066444e-05)),(to_sfixed_a(-9.381403287989087e-06)),(to_sfixed_a(0.00011708301462931558)),(to_sfixed_a(-1.563924342917744e-05)),(to_sfixed_a(-5.5208067351486534e-05)),(to_sfixed_a(-7.002328402450075e-06)),(to_sfixed_a(-3.6909314076183364e-05)));

    constant weight_n1_56 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.032200492918491364)),(to_sfixed_a(0.006945925764739513)),(to_sfixed_a(-0.006539483088999987)),(to_sfixed_a(-0.000402995414333418)),(to_sfixed_a(0.00647975318133831)),(to_sfixed_a(-0.0016464883228763938)),(to_sfixed_a(0.004522024653851986)),(to_sfixed_a(-0.010588052682578564)),(to_sfixed_a(-0.023349862545728683)),(to_sfixed_a(0.0037821985315531492)),(to_sfixed_a(0.0058260043151676655)),(to_sfixed_a(-0.006236291490495205)),(to_sfixed_a(0.0058539854362607)),(to_sfixed_a(0.005502194631844759)),(to_sfixed_a(-0.020855581387877464)),(to_sfixed_a(-0.013357525691390038)),(to_sfixed_a(-0.00037734044599346817)),(to_sfixed_a(0.019293854013085365)),(to_sfixed_a(0.014606287702918053)),(to_sfixed_a(-0.025189585983753204)),(to_sfixed_a(-0.01563245616853237)),(to_sfixed_a(0.005294080823659897)),(to_sfixed_a(0.019130682572722435)),(to_sfixed_a(0.013585776090621948)),(to_sfixed_a(0.027056856080889702)),(to_sfixed_a(-0.0038683523889631033)),(to_sfixed_a(0.006013697944581509)),(to_sfixed_a(0.0005048805032856762)),(to_sfixed_a(0.0024632608983665705)),(to_sfixed_a(0.017412835732102394)),(to_sfixed_a(-0.007895641028881073)),(to_sfixed_a(0.0017205768963322043)),(to_sfixed_a(0.005356529727578163)),(to_sfixed_a(0.03547334298491478)),(to_sfixed_a(0.010235656052827835)),(to_sfixed_a(-0.009663945995271206)),(to_sfixed_a(0.0309356227517128)),(to_sfixed_a(-0.0061368634924292564)));

    constant weight_n1_57 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.04481665790081024)),(to_sfixed_a(1.6156020137714222e-05)),(to_sfixed_a(-8.095757948467508e-06)),(to_sfixed_a(6.702893642795971e-06)),(to_sfixed_a(3.980064138886519e-05)),(to_sfixed_a(-5.97320067754481e-05)),(to_sfixed_a(7.882335921749473e-05)),(to_sfixed_a(-2.6908714062301442e-05)),(to_sfixed_a(5.401002454163972e-06)),(to_sfixed_a(-6.429512268368853e-06)),(to_sfixed_a(-1.3463573850458488e-05)),(to_sfixed_a(-6.206007674336433e-05)),(to_sfixed_a(9.937405593518633e-06)),(to_sfixed_a(4.5961554860696197e-05)),(to_sfixed_a(5.872657857253216e-05)),(to_sfixed_a(-4.829472163692117e-05)),(to_sfixed_a(5.0550102059787605e-06)),(to_sfixed_a(-1.4014503904036246e-05)),(to_sfixed_a(6.172358553158119e-05)),(to_sfixed_a(-7.21284159226343e-05)),(to_sfixed_a(5.561840680456953e-06)),(to_sfixed_a(5.284658527671127e-06)),(to_sfixed_a(-6.478914292529225e-05)),(to_sfixed_a(-1.4049494438950205e-06)),(to_sfixed_a(2.3112618237064453e-06)),(to_sfixed_a(-2.525136551412288e-05)),(to_sfixed_a(-0.00010601292888168246)),(to_sfixed_a(8.243345291703008e-06)),(to_sfixed_a(-5.6541502999607474e-05)),(to_sfixed_a(-4.391768925415818e-06)),(to_sfixed_a(-6.423465674743056e-05)),(to_sfixed_a(0.0001159644962172024)),(to_sfixed_a(-4.707074913312681e-05)),(to_sfixed_a(2.8633850888581946e-05)),(to_sfixed_a(-9.708331344882026e-05)),(to_sfixed_a(5.8632133004721254e-05)),(to_sfixed_a(-2.5065546651603654e-05)),(to_sfixed_a(-7.48054007999599e-05)));

    constant weight_n1_58 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.00914741400629282)),(to_sfixed_a(-3.8891976146260276e-05)),(to_sfixed_a(-9.717681678012013e-06)),(to_sfixed_a(-4.0164431993616745e-05)),(to_sfixed_a(9.811470590648241e-06)),(to_sfixed_a(-1.261121633433504e-05)),(to_sfixed_a(-1.6104222311241756e-07)),(to_sfixed_a(3.850113716907799e-05)),(to_sfixed_a(2.0189767383271828e-05)),(to_sfixed_a(-1.2310478268773295e-05)),(to_sfixed_a(-3.547271262505092e-05)),(to_sfixed_a(-3.863491656375118e-06)),(to_sfixed_a(2.2557927877642214e-05)),(to_sfixed_a(1.4818063391430769e-05)),(to_sfixed_a(3.0657673050882295e-05)),(to_sfixed_a(1.1771858225984033e-05)),(to_sfixed_a(-6.5112399170175195e-06)),(to_sfixed_a(-2.102952203131281e-05)),(to_sfixed_a(4.097297278349288e-05)),(to_sfixed_a(4.8705471272114664e-05)),(to_sfixed_a(-8.638269355287775e-05)),(to_sfixed_a(3.3296673791483045e-05)),(to_sfixed_a(9.692674211692065e-05)),(to_sfixed_a(-4.653309588320553e-05)),(to_sfixed_a(-1.4533874491462484e-05)),(to_sfixed_a(-1.2050055374857038e-05)),(to_sfixed_a(2.4017221221583895e-05)),(to_sfixed_a(-1.672224243520759e-05)),(to_sfixed_a(5.166917253518477e-05)),(to_sfixed_a(5.277426680549979e-05)),(to_sfixed_a(-3.497413490549661e-05)),(to_sfixed_a(3.918374602562835e-08)),(to_sfixed_a(-4.6332472265930846e-05)),(to_sfixed_a(-7.133757662813878e-06)),(to_sfixed_a(7.518810889450833e-05)),(to_sfixed_a(-9.840492566581815e-05)),(to_sfixed_a(-7.686902245040983e-05)),(to_sfixed_a(5.004037666367367e-05)));

    constant weight_n1_59 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.5060866475105286)),(to_sfixed_a(-0.0019544532988220453)),(to_sfixed_a(0.021789399906992912)),(to_sfixed_a(0.019111456349492073)),(to_sfixed_a(0.033631831407547)),(to_sfixed_a(-0.004337341524660587)),(to_sfixed_a(-0.007810165174305439)),(to_sfixed_a(0.0031548975966870785)),(to_sfixed_a(-0.03471090644598007)),(to_sfixed_a(0.016196681186556816)),(to_sfixed_a(-0.03006800077855587)),(to_sfixed_a(-0.005883866921067238)),(to_sfixed_a(-0.0001940140500664711)),(to_sfixed_a(0.03591308370232582)),(to_sfixed_a(-0.02428504079580307)),(to_sfixed_a(0.0034526512026786804)),(to_sfixed_a(0.04638966545462608)),(to_sfixed_a(-0.03569979593157768)),(to_sfixed_a(0.04744739085435867)),(to_sfixed_a(-0.016803979873657227)),(to_sfixed_a(-0.018052732571959496)),(to_sfixed_a(-0.01708562858402729)),(to_sfixed_a(-0.0020447627175599337)),(to_sfixed_a(0.022899147123098373)),(to_sfixed_a(-0.05070533975958824)),(to_sfixed_a(0.009956936351954937)),(to_sfixed_a(-0.0004329135699663311)),(to_sfixed_a(0.02270352840423584)),(to_sfixed_a(0.026137687265872955)),(to_sfixed_a(-0.03169337660074234)),(to_sfixed_a(-0.011437827721238136)),(to_sfixed_a(0.044496629387140274)),(to_sfixed_a(-0.02464406006038189)),(to_sfixed_a(0.044839322566986084)),(to_sfixed_a(0.009054440073668957)),(to_sfixed_a(-0.0018465355969965458)),(to_sfixed_a(-0.0612424872815609)),(to_sfixed_a(-0.026476362720131874)));

    constant weight_n1_60 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.0321747325360775)),(to_sfixed_a(-0.003733262652531266)),(to_sfixed_a(-0.015194285660982132)),(to_sfixed_a(0.00594418914988637)),(to_sfixed_a(0.003489517141133547)),(to_sfixed_a(0.002778134774416685)),(to_sfixed_a(0.019029589369893074)),(to_sfixed_a(-0.02414056472480297)),(to_sfixed_a(0.0034002012107521296)),(to_sfixed_a(-0.016536174342036247)),(to_sfixed_a(-0.02759813703596592)),(to_sfixed_a(0.014535084366798401)),(to_sfixed_a(-0.022062284871935844)),(to_sfixed_a(-0.00024542456958442926)),(to_sfixed_a(0.005329374689608812)),(to_sfixed_a(0.007322376128286123)),(to_sfixed_a(-0.00236529135145247)),(to_sfixed_a(-0.014966894872486591)),(to_sfixed_a(8.398099453188479e-05)),(to_sfixed_a(-0.019460514187812805)),(to_sfixed_a(0.00786572229117155)),(to_sfixed_a(0.017095297574996948)),(to_sfixed_a(0.0049500479362905025)),(to_sfixed_a(-0.0036605794448405504)),(to_sfixed_a(0.003818678203970194)),(to_sfixed_a(0.0013406043872237206)),(to_sfixed_a(-0.015766266733407974)),(to_sfixed_a(-0.03285796940326691)),(to_sfixed_a(-0.033475346863269806)),(to_sfixed_a(-0.011830965988337994)),(to_sfixed_a(0.014150195755064487)),(to_sfixed_a(-0.024003639817237854)),(to_sfixed_a(-0.007098471280187368)),(to_sfixed_a(-0.01650046929717064)),(to_sfixed_a(0.012304050847887993)),(to_sfixed_a(-0.006644665263593197)),(to_sfixed_a(-0.005666332319378853)),(to_sfixed_a(0.012276223860681057)));

    constant weight_n1_61 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.02538255788385868)),(to_sfixed_a(0.019274622201919556)),(to_sfixed_a(-0.03503689914941788)),(to_sfixed_a(-0.01851755939424038)),(to_sfixed_a(0.022462299093604088)),(to_sfixed_a(-0.026641787961125374)),(to_sfixed_a(-0.026338716968894005)),(to_sfixed_a(-0.0007377025322057307)),(to_sfixed_a(0.03490261361002922)),(to_sfixed_a(-0.009724228642880917)),(to_sfixed_a(0.012207352556288242)),(to_sfixed_a(0.025164157152175903)),(to_sfixed_a(0.023730356246232986)),(to_sfixed_a(0.018907828256487846)),(to_sfixed_a(-0.04063567891716957)),(to_sfixed_a(0.015052316710352898)),(to_sfixed_a(-0.010927059687674046)),(to_sfixed_a(0.06291192770004272)),(to_sfixed_a(0.008296837098896503)),(to_sfixed_a(-0.0841807872056961)),(to_sfixed_a(-0.03419530764222145)),(to_sfixed_a(0.0004915576428174973)),(to_sfixed_a(0.011923067271709442)),(to_sfixed_a(0.05045298486948013)),(to_sfixed_a(0.032324325293302536)),(to_sfixed_a(0.0048428792506456375)),(to_sfixed_a(0.04513264074921608)),(to_sfixed_a(0.07498759776353836)),(to_sfixed_a(-0.008731693029403687)),(to_sfixed_a(-0.0479276180267334)),(to_sfixed_a(-0.07613252848386765)),(to_sfixed_a(0.07156310230493546)),(to_sfixed_a(-0.03879766911268234)),(to_sfixed_a(-0.015040382742881775)),(to_sfixed_a(0.025587091222405434)),(to_sfixed_a(0.06413526087999344)),(to_sfixed_a(-0.033124200999736786)),(to_sfixed_a(-0.003233914729207754)));

    constant weight_n1_62 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.04552634805440903)),(to_sfixed_a(-0.05576751008629799)),(to_sfixed_a(-0.027609866112470627)),(to_sfixed_a(0.017500272020697594)),(to_sfixed_a(0.05393300950527191)),(to_sfixed_a(-0.06452161073684692)),(to_sfixed_a(-0.12278691679239273)),(to_sfixed_a(0.06879982352256775)),(to_sfixed_a(0.05261589214205742)),(to_sfixed_a(-0.028608011081814766)),(to_sfixed_a(-0.01842605322599411)),(to_sfixed_a(-0.0009006980108097196)),(to_sfixed_a(0.07262331992387772)),(to_sfixed_a(-0.2126181721687317)),(to_sfixed_a(0.22920438647270203)),(to_sfixed_a(0.12710632383823395)),(to_sfixed_a(-0.0960664302110672)),(to_sfixed_a(-0.26916494965553284)),(to_sfixed_a(-0.0734485611319542)),(to_sfixed_a(0.13585583865642548)),(to_sfixed_a(0.20212788879871368)),(to_sfixed_a(5.866104402230121e-05)),(to_sfixed_a(-0.09961867332458496)),(to_sfixed_a(-0.0951654464006424)),(to_sfixed_a(-0.10517533123493195)),(to_sfixed_a(0.018836449831724167)),(to_sfixed_a(-0.010633595287799835)),(to_sfixed_a(-0.13445565104484558)),(to_sfixed_a(0.004085928667336702)),(to_sfixed_a(0.015323925763368607)),(to_sfixed_a(-0.06195066496729851)),(to_sfixed_a(-0.020040230825543404)),(to_sfixed_a(-0.10709786415100098)),(to_sfixed_a(-0.07407420873641968)),(to_sfixed_a(-0.010598286055028439)),(to_sfixed_a(-0.031408462673425674)),(to_sfixed_a(-0.26361083984375)),(to_sfixed_a(0.07337364554405212)));

    constant weight_n1_63 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.011922924779355526)),(to_sfixed_a(1.2673034689214546e-05)),(to_sfixed_a(-2.768872946035117e-05)),(to_sfixed_a(7.81378366809804e-06)),(to_sfixed_a(-3.6765672120964155e-05)),(to_sfixed_a(5.540591882891022e-05)),(to_sfixed_a(-1.7357968317810446e-05)),(to_sfixed_a(2.1316791389836e-05)),(to_sfixed_a(1.6012383639463224e-05)),(to_sfixed_a(-7.701554568484426e-05)),(to_sfixed_a(-3.4137767215725034e-05)),(to_sfixed_a(-2.8288020985201e-05)),(to_sfixed_a(9.01626845006831e-06)),(to_sfixed_a(-4.90884376631584e-05)),(to_sfixed_a(3.29402246279642e-05)),(to_sfixed_a(-2.6126743250642903e-05)),(to_sfixed_a(2.815519110299647e-05)),(to_sfixed_a(-8.915207581594586e-05)),(to_sfixed_a(5.4963027650956064e-05)),(to_sfixed_a(-1.4901394251864986e-06)),(to_sfixed_a(-4.4894637539982796e-05)),(to_sfixed_a(-8.654462817503372e-07)),(to_sfixed_a(-6.424757884815335e-05)),(to_sfixed_a(4.686828833655454e-05)),(to_sfixed_a(-7.587832897115732e-06)),(to_sfixed_a(5.179553045309149e-05)),(to_sfixed_a(-1.3755053259956185e-05)),(to_sfixed_a(2.6266612621839158e-05)),(to_sfixed_a(4.996057759854011e-05)),(to_sfixed_a(-5.5691674788249657e-05)),(to_sfixed_a(4.323139364714734e-06)),(to_sfixed_a(5.626348502119072e-05)),(to_sfixed_a(7.935443591122748e-07)),(to_sfixed_a(2.074806616292335e-05)),(to_sfixed_a(-6.4998930611182e-05)),(to_sfixed_a(3.2249118930849363e-07)),(to_sfixed_a(-9.550613867759239e-06)),(to_sfixed_a(4.4720189180225134e-05)));

    constant weight_n1_64 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.15831415355205536)),(to_sfixed_a(0.026853682473301888)),(to_sfixed_a(-0.10210394859313965)),(to_sfixed_a(-0.011193507350981236)),(to_sfixed_a(0.04258609563112259)),(to_sfixed_a(-0.16631044447422028)),(to_sfixed_a(0.10492265969514847)),(to_sfixed_a(0.22867360711097717)),(to_sfixed_a(0.12461443245410919)),(to_sfixed_a(0.17283882200717926)),(to_sfixed_a(0.07706400752067566)),(to_sfixed_a(0.2780294418334961)),(to_sfixed_a(-0.027570441365242004)),(to_sfixed_a(-0.05245685949921608)),(to_sfixed_a(-0.09405095130205154)),(to_sfixed_a(0.25483572483062744)),(to_sfixed_a(-0.15900662541389465)),(to_sfixed_a(0.13731029629707336)),(to_sfixed_a(-0.23710525035858154)),(to_sfixed_a(0.06508168578147888)),(to_sfixed_a(-0.24753963947296143)),(to_sfixed_a(-0.011836019344627857)),(to_sfixed_a(0.024066515266895294)),(to_sfixed_a(0.12652428448200226)),(to_sfixed_a(-0.07728955149650574)),(to_sfixed_a(0.00788357574492693)),(to_sfixed_a(-0.10558706521987915)),(to_sfixed_a(0.1666400134563446)),(to_sfixed_a(-0.09132913500070572)),(to_sfixed_a(0.0009165406227111816)),(to_sfixed_a(-0.2579912841320038)),(to_sfixed_a(0.12887048721313477)),(to_sfixed_a(-0.23376153409481049)),(to_sfixed_a(0.07227407395839691)),(to_sfixed_a(-0.017324751242995262)),(to_sfixed_a(0.05346110090613365)),(to_sfixed_a(0.057590682059526443)),(to_sfixed_a(-0.11153779178857803)));

    constant weight_n1_65 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.04273220896720886)),(to_sfixed_a(4.313618774176575e-05)),(to_sfixed_a(1.2261082702025305e-05)),(to_sfixed_a(-3.817126707872376e-05)),(to_sfixed_a(-5.6525565014453605e-05)),(to_sfixed_a(2.1446458049467765e-05)),(to_sfixed_a(-3.9874244066595566e-06)),(to_sfixed_a(-5.676785804098472e-06)),(to_sfixed_a(4.525435360847041e-05)),(to_sfixed_a(3.13379023282323e-05)),(to_sfixed_a(1.2333841368672438e-05)),(to_sfixed_a(-3.9073795051081106e-05)),(to_sfixed_a(-7.363365148194134e-05)),(to_sfixed_a(-2.5005403585964814e-05)),(to_sfixed_a(-6.565682997461408e-05)),(to_sfixed_a(1.2590651749633253e-05)),(to_sfixed_a(8.484045974910259e-05)),(to_sfixed_a(3.924991324311122e-05)),(to_sfixed_a(6.654411845374852e-05)),(to_sfixed_a(-9.579230209055822e-06)),(to_sfixed_a(8.909086318453774e-06)),(to_sfixed_a(-9.278279321733862e-05)),(to_sfixed_a(-2.186183337471448e-05)),(to_sfixed_a(-5.758234692621045e-05)),(to_sfixed_a(-7.774327968945727e-05)),(to_sfixed_a(-4.469548002816737e-05)),(to_sfixed_a(5.061834235675633e-05)),(to_sfixed_a(-3.5579003451857716e-05)),(to_sfixed_a(-3.848653068416752e-05)),(to_sfixed_a(-6.572336860699579e-05)),(to_sfixed_a(-1.957308313649264e-06)),(to_sfixed_a(-9.661842341301963e-05)),(to_sfixed_a(5.0169986934633926e-05)),(to_sfixed_a(6.218007183633745e-05)),(to_sfixed_a(1.1538775652297772e-05)),(to_sfixed_a(2.509033720343723e-06)),(to_sfixed_a(8.726574014872313e-05)),(to_sfixed_a(-5.674580825143494e-05)));

    constant weight_n1_66 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.10854636877775192)),(to_sfixed_a(0.29283273220062256)),(to_sfixed_a(0.18984395265579224)),(to_sfixed_a(-0.1048344075679779)),(to_sfixed_a(0.0728050172328949)),(to_sfixed_a(-0.003976179286837578)),(to_sfixed_a(-0.16187426447868347)),(to_sfixed_a(0.007467066403478384)),(to_sfixed_a(0.029842771589756012)),(to_sfixed_a(0.19606950879096985)),(to_sfixed_a(-0.12249623984098434)),(to_sfixed_a(-0.00893156137317419)),(to_sfixed_a(-0.04171709716320038)),(to_sfixed_a(0.065533347427845)),(to_sfixed_a(0.33821213245391846)),(to_sfixed_a(0.11300500482320786)),(to_sfixed_a(0.10561921447515488)),(to_sfixed_a(0.10720629245042801)),(to_sfixed_a(-0.008471129462122917)),(to_sfixed_a(-0.194168820977211)),(to_sfixed_a(-0.039151765406131744)),(to_sfixed_a(0.13396094739437103)),(to_sfixed_a(0.19562269747257233)),(to_sfixed_a(0.0432339571416378)),(to_sfixed_a(-0.028360914438962936)),(to_sfixed_a(0.09232060611248016)),(to_sfixed_a(-0.06909216195344925)),(to_sfixed_a(-0.06349315494298935)),(to_sfixed_a(-0.2980492115020752)),(to_sfixed_a(-0.044000327587127686)),(to_sfixed_a(-0.025263087823987007)),(to_sfixed_a(0.009662636555731297)),(to_sfixed_a(-0.0363110676407814)),(to_sfixed_a(0.1217353492975235)),(to_sfixed_a(0.16675573587417603)),(to_sfixed_a(-0.06747063994407654)),(to_sfixed_a(-0.006672275252640247)),(to_sfixed_a(0.02965421974658966)));

    constant weight_n1_67 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.02687550149857998)),(to_sfixed_a(-0.011866766959428787)),(to_sfixed_a(0.010284941643476486)),(to_sfixed_a(0.0032457115594297647)),(to_sfixed_a(0.008435701951384544)),(to_sfixed_a(0.00480466615408659)),(to_sfixed_a(-0.012204006314277649)),(to_sfixed_a(0.002984800608828664)),(to_sfixed_a(-0.008430739864706993)),(to_sfixed_a(0.0007876676390878856)),(to_sfixed_a(0.014269242994487286)),(to_sfixed_a(-0.02689010091125965)),(to_sfixed_a(0.009692137129604816)),(to_sfixed_a(-0.0021962416358292103)),(to_sfixed_a(-0.005629129707813263)),(to_sfixed_a(-0.002502195304259658)),(to_sfixed_a(0.0230467077344656)),(to_sfixed_a(0.016339022666215897)),(to_sfixed_a(0.017150919884443283)),(to_sfixed_a(0.002340982435271144)),(to_sfixed_a(0.003002665238454938)),(to_sfixed_a(-0.01092303916811943)),(to_sfixed_a(0.00966974999755621)),(to_sfixed_a(-0.009678232483565807)),(to_sfixed_a(0.001535404589958489)),(to_sfixed_a(0.011448785662651062)),(to_sfixed_a(0.008861205540597439)),(to_sfixed_a(-0.002999694785103202)),(to_sfixed_a(-0.001427841023541987)),(to_sfixed_a(0.01514950767159462)),(to_sfixed_a(-0.043461527675390244)),(to_sfixed_a(-0.02585257589817047)),(to_sfixed_a(-0.004794673528522253)),(to_sfixed_a(0.04228867590427399)),(to_sfixed_a(0.021226778626441956)),(to_sfixed_a(0.014373094774782658)),(to_sfixed_a(0.033832985907793045)),(to_sfixed_a(-0.035749346017837524)));

    constant weight_n1_68 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.015932437032461166)),(to_sfixed_a(1.2485414117691107e-05)),(to_sfixed_a(-1.9020921172341332e-05)),(to_sfixed_a(1.8494270989322104e-05)),(to_sfixed_a(4.435686605575029e-06)),(to_sfixed_a(-1.7362686776323244e-05)),(to_sfixed_a(-3.6651777918450534e-05)),(to_sfixed_a(-6.0497386584756896e-05)),(to_sfixed_a(2.519105873943772e-05)),(to_sfixed_a(-4.4498592615127563e-05)),(to_sfixed_a(2.7113248506793752e-05)),(to_sfixed_a(-2.197149660787545e-05)),(to_sfixed_a(8.2058621046599e-05)),(to_sfixed_a(-1.8671715224627405e-05)),(to_sfixed_a(-5.34035450527881e-07)),(to_sfixed_a(5.1852286560460925e-05)),(to_sfixed_a(1.6392186807934195e-05)),(to_sfixed_a(-9.132030754699372e-06)),(to_sfixed_a(-3.5820252378471196e-05)),(to_sfixed_a(5.5468339269282296e-05)),(to_sfixed_a(-1.590764441061765e-05)),(to_sfixed_a(3.4845914342440665e-05)),(to_sfixed_a(-6.619008490815759e-05)),(to_sfixed_a(-5.6810658861650154e-05)),(to_sfixed_a(6.135708827059716e-05)),(to_sfixed_a(8.937533493735828e-06)),(to_sfixed_a(3.25004912156146e-05)),(to_sfixed_a(-1.5885132597759366e-05)),(to_sfixed_a(4.741017983178608e-05)),(to_sfixed_a(0.0002104886807501316)),(to_sfixed_a(1.1634866496024188e-05)),(to_sfixed_a(7.112717139534652e-05)),(to_sfixed_a(4.469078703550622e-05)),(to_sfixed_a(2.6136984160984866e-05)),(to_sfixed_a(1.3853922609996516e-05)),(to_sfixed_a(-8.370693831238896e-05)),(to_sfixed_a(-6.644523818977177e-05)),(to_sfixed_a(8.113593503367156e-05)));

    constant weight_n1_69 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.30059128999710083)),(to_sfixed_a(-0.19843292236328125)),(to_sfixed_a(-0.05941928178071976)),(to_sfixed_a(-0.023916130885481834)),(to_sfixed_a(-0.07758259028196335)),(to_sfixed_a(0.0064984280616045)),(to_sfixed_a(-0.06901973485946655)),(to_sfixed_a(0.07745522260665894)),(to_sfixed_a(-0.07477644830942154)),(to_sfixed_a(0.1479446291923523)),(to_sfixed_a(-0.11638858914375305)),(to_sfixed_a(-0.02568785659968853)),(to_sfixed_a(-0.07596594095230103)),(to_sfixed_a(0.10088993608951569)),(to_sfixed_a(0.2249988615512848)),(to_sfixed_a(-0.09808415919542313)),(to_sfixed_a(0.03141532093286514)),(to_sfixed_a(0.03822409734129906)),(to_sfixed_a(-0.10282151401042938)),(to_sfixed_a(-0.07628049701452255)),(to_sfixed_a(0.05069858953356743)),(to_sfixed_a(-0.10014250874519348)),(to_sfixed_a(-0.041979629546403885)),(to_sfixed_a(0.11943496018648148)),(to_sfixed_a(0.34159326553344727)),(to_sfixed_a(0.20397262275218964)),(to_sfixed_a(-0.04316170886158943)),(to_sfixed_a(-0.010508173145353794)),(to_sfixed_a(0.2425571233034134)),(to_sfixed_a(0.06414955854415894)),(to_sfixed_a(0.005912561900913715)),(to_sfixed_a(0.24140557646751404)),(to_sfixed_a(-0.01114345621317625)),(to_sfixed_a(-0.08018511533737183)),(to_sfixed_a(-0.20639286935329437)),(to_sfixed_a(0.06325377523899078)),(to_sfixed_a(0.005528866313397884)),(to_sfixed_a(0.12454087287187576)));

    constant weight_n1_70 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.08288822323083878)),(to_sfixed_a(-0.12429346889257431)),(to_sfixed_a(0.06631514430046082)),(to_sfixed_a(-0.14744818210601807)),(to_sfixed_a(0.04750068485736847)),(to_sfixed_a(-0.06312884390354156)),(to_sfixed_a(0.011615087278187275)),(to_sfixed_a(-0.029191426932811737)),(to_sfixed_a(0.02492695115506649)),(to_sfixed_a(0.06460559368133545)),(to_sfixed_a(0.0360814705491066)),(to_sfixed_a(0.16991780698299408)),(to_sfixed_a(0.061075590550899506)),(to_sfixed_a(-0.08413823693990707)),(to_sfixed_a(-0.03980319947004318)),(to_sfixed_a(-0.0277326051145792)),(to_sfixed_a(0.08351609855890274)),(to_sfixed_a(-0.11797885596752167)),(to_sfixed_a(0.09024809300899506)),(to_sfixed_a(-0.00932466983795166)),(to_sfixed_a(-0.044930096715688705)),(to_sfixed_a(0.06458944827318192)),(to_sfixed_a(0.0676322653889656)),(to_sfixed_a(0.03197857737541199)),(to_sfixed_a(-0.11178668588399887)),(to_sfixed_a(0.14510951936244965)),(to_sfixed_a(0.09489130228757858)),(to_sfixed_a(-0.06207898631691933)),(to_sfixed_a(0.02664927951991558)),(to_sfixed_a(0.1298900842666626)),(to_sfixed_a(0.14004477858543396)),(to_sfixed_a(0.047237999737262726)),(to_sfixed_a(-0.03954213857650757)),(to_sfixed_a(0.04603291675448418)),(to_sfixed_a(-0.19480000436306)),(to_sfixed_a(-0.030456438660621643)),(to_sfixed_a(-0.04821375384926796)),(to_sfixed_a(0.08914975076913834)));

    constant weight_n1_71 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.24838581681251526)),(to_sfixed_a(-0.0068165273405611515)),(to_sfixed_a(0.03079892136156559)),(to_sfixed_a(0.016234174370765686)),(to_sfixed_a(-0.051308900117874146)),(to_sfixed_a(-0.03754320368170738)),(to_sfixed_a(0.0066346232779324055)),(to_sfixed_a(0.057128120213747025)),(to_sfixed_a(0.07888364791870117)),(to_sfixed_a(-0.010259074158966541)),(to_sfixed_a(0.1303286850452423)),(to_sfixed_a(0.04224000871181488)),(to_sfixed_a(-0.00809289887547493)),(to_sfixed_a(-0.10947246104478836)),(to_sfixed_a(0.07734763622283936)),(to_sfixed_a(0.0610358789563179)),(to_sfixed_a(-0.05914352834224701)),(to_sfixed_a(-0.030749348923563957)),(to_sfixed_a(-0.011597291566431522)),(to_sfixed_a(0.011981556192040443)),(to_sfixed_a(0.06057879328727722)),(to_sfixed_a(-0.01776224747300148)),(to_sfixed_a(-0.060895051807165146)),(to_sfixed_a(-0.12279883772134781)),(to_sfixed_a(0.04385983571410179)),(to_sfixed_a(-0.01891908422112465)),(to_sfixed_a(-0.1383107453584671)),(to_sfixed_a(0.019743718206882477)),(to_sfixed_a(-0.03530341386795044)),(to_sfixed_a(0.0008956361562013626)),(to_sfixed_a(-0.12421351671218872)),(to_sfixed_a(0.05821182578802109)),(to_sfixed_a(0.12322036176919937)),(to_sfixed_a(0.029652340337634087)),(to_sfixed_a(-0.11609333008527756)),(to_sfixed_a(-0.025655891746282578)),(to_sfixed_a(-0.04720497131347656)),(to_sfixed_a(-0.043077003210783005)));

    constant weight_n1_72 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.0263239573687315)),(to_sfixed_a(-7.93112485553138e-05)),(to_sfixed_a(1.762208921718411e-05)),(to_sfixed_a(-2.798556670313701e-05)),(to_sfixed_a(-2.509966361685656e-05)),(to_sfixed_a(2.9362456189119257e-05)),(to_sfixed_a(1.081064601748949e-05)),(to_sfixed_a(-1.5400890333694406e-05)),(to_sfixed_a(1.091547619580524e-05)),(to_sfixed_a(-3.285118145868182e-05)),(to_sfixed_a(-2.8364484023768455e-05)),(to_sfixed_a(-2.33777300309157e-05)),(to_sfixed_a(-3.341410410939716e-05)),(to_sfixed_a(3.4780543501256034e-05)),(to_sfixed_a(4.719590288004838e-05)),(to_sfixed_a(-2.5550267309881747e-05)),(to_sfixed_a(-4.701018406194635e-05)),(to_sfixed_a(-6.67260110276402e-06)),(to_sfixed_a(7.259678386617452e-05)),(to_sfixed_a(1.692240039119497e-05)),(to_sfixed_a(-3.942270632251166e-05)),(to_sfixed_a(-5.5305885325651616e-05)),(to_sfixed_a(-3.453492922744772e-07)),(to_sfixed_a(7.91253933130065e-06)),(to_sfixed_a(8.54973986861296e-05)),(to_sfixed_a(8.754673763178289e-05)),(to_sfixed_a(4.4528464059112594e-05)),(to_sfixed_a(3.987771924585104e-05)),(to_sfixed_a(3.4950120607391e-05)),(to_sfixed_a(6.659440259682015e-05)),(to_sfixed_a(-5.4169831855688244e-05)),(to_sfixed_a(-5.877995863556862e-05)),(to_sfixed_a(-6.444860628107563e-05)),(to_sfixed_a(-3.977297092205845e-05)),(to_sfixed_a(7.387586811091751e-05)),(to_sfixed_a(3.1746807508170605e-05)),(to_sfixed_a(-2.2104701201897115e-05)),(to_sfixed_a(5.543629595194943e-05)));

    constant weight_n1_73 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.010054564103484154)),(to_sfixed_a(-2.8360153009998612e-05)),(to_sfixed_a(2.805801159411203e-05)),(to_sfixed_a(7.912613000371493e-06)),(to_sfixed_a(-4.857964449911378e-05)),(to_sfixed_a(3.828441913356073e-05)),(to_sfixed_a(5.749508272856474e-05)),(to_sfixed_a(-5.518335092347115e-05)),(to_sfixed_a(-3.178750921506435e-05)),(to_sfixed_a(-1.101860198104987e-05)),(to_sfixed_a(-3.92728765064021e-07)),(to_sfixed_a(-1.2290111953916494e-05)),(to_sfixed_a(2.699421384022571e-05)),(to_sfixed_a(3.131885750917718e-05)),(to_sfixed_a(-0.00010256210953230038)),(to_sfixed_a(-3.435835969867185e-05)),(to_sfixed_a(1.6498648619744927e-05)),(to_sfixed_a(3.264402039349079e-05)),(to_sfixed_a(-2.3503573174821213e-05)),(to_sfixed_a(-3.397563432372408e-06)),(to_sfixed_a(-1.756916390149854e-05)),(to_sfixed_a(-8.899990461941343e-06)),(to_sfixed_a(7.00335658621043e-05)),(to_sfixed_a(-1.4872313158775796e-06)),(to_sfixed_a(-2.4006150852073915e-05)),(to_sfixed_a(6.409757043002173e-05)),(to_sfixed_a(-3.6392164474818856e-05)),(to_sfixed_a(-2.3519411115557887e-05)),(to_sfixed_a(-4.586591603583656e-05)),(to_sfixed_a(2.6967971280100755e-05)),(to_sfixed_a(-5.889995372854173e-05)),(to_sfixed_a(-2.9622156944242306e-05)),(to_sfixed_a(-4.156228169449605e-05)),(to_sfixed_a(4.213923239149153e-05)),(to_sfixed_a(1.2521317330538295e-05)),(to_sfixed_a(4.4868720578961074e-05)),(to_sfixed_a(7.832776645955164e-06)),(to_sfixed_a(-0.0001654562511248514)));

    constant weight_n1_74 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.018064986914396286)),(to_sfixed_a(-1.0985582775902003e-05)),(to_sfixed_a(4.3521875340957195e-05)),(to_sfixed_a(-1.3026373380853329e-05)),(to_sfixed_a(3.6919107515132055e-05)),(to_sfixed_a(2.5389501388417557e-05)),(to_sfixed_a(-2.2296026145340875e-05)),(to_sfixed_a(3.8770438550272956e-05)),(to_sfixed_a(-1.1063980309700128e-06)),(to_sfixed_a(9.826570021687075e-05)),(to_sfixed_a(-1.8924674805020913e-05)),(to_sfixed_a(5.917523958487436e-05)),(to_sfixed_a(-6.045269037713297e-05)),(to_sfixed_a(-3.9380454836646095e-05)),(to_sfixed_a(4.2957992263836786e-05)),(to_sfixed_a(9.97180450212909e-07)),(to_sfixed_a(-2.1386207663454115e-05)),(to_sfixed_a(5.761525244452059e-05)),(to_sfixed_a(-1.457490179745946e-05)),(to_sfixed_a(-3.7249945307848975e-05)),(to_sfixed_a(2.8130314149166225e-06)),(to_sfixed_a(-1.3826023860019632e-05)),(to_sfixed_a(5.722254718421027e-05)),(to_sfixed_a(2.7695305107044987e-05)),(to_sfixed_a(2.155700531147886e-05)),(to_sfixed_a(4.7338784497696906e-05)),(to_sfixed_a(4.0025925045483746e-06)),(to_sfixed_a(1.3722811672778334e-05)),(to_sfixed_a(4.6280660171760246e-05)),(to_sfixed_a(7.71569466451183e-06)),(to_sfixed_a(4.5177938545748475e-07)),(to_sfixed_a(4.638948666979559e-06)),(to_sfixed_a(-2.1815671061631292e-05)),(to_sfixed_a(6.096078141126782e-05)),(to_sfixed_a(-6.153310823719949e-05)),(to_sfixed_a(-6.65401530568488e-05)),(to_sfixed_a(6.742872938048095e-05)),(to_sfixed_a(-3.4353433875367045e-05)));

    constant weight_n1_75 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.3336969017982483)),(to_sfixed_a(0.055782873183488846)),(to_sfixed_a(0.02075355313718319)),(to_sfixed_a(0.04974014312028885)),(to_sfixed_a(-0.05762127786874771)),(to_sfixed_a(-0.048381634056568146)),(to_sfixed_a(-0.0983545184135437)),(to_sfixed_a(-0.07689255475997925)),(to_sfixed_a(0.30923327803611755)),(to_sfixed_a(-0.042600881308317184)),(to_sfixed_a(-0.09364135563373566)),(to_sfixed_a(0.11348334699869156)),(to_sfixed_a(-0.18180561065673828)),(to_sfixed_a(0.2443670630455017)),(to_sfixed_a(0.09050726890563965)),(to_sfixed_a(0.15245544910430908)),(to_sfixed_a(-0.08673351258039474)),(to_sfixed_a(-0.19461002945899963)),(to_sfixed_a(-0.04387940466403961)),(to_sfixed_a(-0.1846449077129364)),(to_sfixed_a(-0.04875333607196808)),(to_sfixed_a(-0.014586064033210278)),(to_sfixed_a(0.06950226426124573)),(to_sfixed_a(-0.07692615687847137)),(to_sfixed_a(0.11429334431886673)),(to_sfixed_a(-0.0580364428460598)),(to_sfixed_a(0.20986387133598328)),(to_sfixed_a(-0.10786264389753342)),(to_sfixed_a(0.11694255471229553)),(to_sfixed_a(0.04957651346921921)),(to_sfixed_a(-0.03139158710837364)),(to_sfixed_a(-0.08932279795408249)),(to_sfixed_a(-0.061484724283218384)),(to_sfixed_a(0.03441711515188217)),(to_sfixed_a(-0.006571502424776554)),(to_sfixed_a(0.01706230267882347)),(to_sfixed_a(-0.0027323684189468622)),(to_sfixed_a(-0.007874560542404652)));

    constant weight_n1_76 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.09432821720838547)),(to_sfixed_a(0.039074402302503586)),(to_sfixed_a(0.02550024539232254)),(to_sfixed_a(0.02198122628033161)),(to_sfixed_a(0.013352709822356701)),(to_sfixed_a(-0.01969103142619133)),(to_sfixed_a(-0.017378641292452812)),(to_sfixed_a(0.008484771475195885)),(to_sfixed_a(0.011263559572398663)),(to_sfixed_a(-0.024436069652438164)),(to_sfixed_a(0.017291367053985596)),(to_sfixed_a(-0.029454227536916733)),(to_sfixed_a(0.020933983847498894)),(to_sfixed_a(-0.051945872604846954)),(to_sfixed_a(0.01955539919435978)),(to_sfixed_a(-0.011532122269272804)),(to_sfixed_a(-0.003264766186475754)),(to_sfixed_a(-0.013838423416018486)),(to_sfixed_a(-0.03962979465723038)),(to_sfixed_a(0.034926217049360275)),(to_sfixed_a(-0.01263582706451416)),(to_sfixed_a(0.0016671806806698442)),(to_sfixed_a(0.01740437000989914)),(to_sfixed_a(-0.06305841356515884)),(to_sfixed_a(0.03996612876653671)),(to_sfixed_a(-0.022035649046301842)),(to_sfixed_a(-0.024223893880844116)),(to_sfixed_a(-0.0030795272905379534)),(to_sfixed_a(0.03306838870048523)),(to_sfixed_a(0.014041976071894169)),(to_sfixed_a(-0.007125793024897575)),(to_sfixed_a(-0.04725521057844162)),(to_sfixed_a(0.025846106931567192)),(to_sfixed_a(0.037007804960012436)),(to_sfixed_a(-0.05199568346142769)),(to_sfixed_a(0.014066777192056179)),(to_sfixed_a(-0.004561693873256445)),(to_sfixed_a(0.0036053035873919725)));

    constant weight_n1_77 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.014241009950637817)),(to_sfixed_a(-2.253475940960925e-05)),(to_sfixed_a(-2.527262768126093e-05)),(to_sfixed_a(6.821186980232596e-05)),(to_sfixed_a(1.5583858839818276e-05)),(to_sfixed_a(5.058405349700479e-06)),(to_sfixed_a(5.085697921458632e-05)),(to_sfixed_a(-3.29887043335475e-05)),(to_sfixed_a(-1.1913429261767305e-05)),(to_sfixed_a(3.848046253551729e-05)),(to_sfixed_a(4.142189573030919e-05)),(to_sfixed_a(-2.9990647817612626e-05)),(to_sfixed_a(-3.1724014206702122e-06)),(to_sfixed_a(-2.301045969943516e-05)),(to_sfixed_a(-4.5886852603871375e-05)),(to_sfixed_a(-4.823676135856658e-05)),(to_sfixed_a(3.0097684430074878e-05)),(to_sfixed_a(4.457420072867535e-05)),(to_sfixed_a(2.1608602764899842e-05)),(to_sfixed_a(3.940879105357453e-05)),(to_sfixed_a(-6.284979463089257e-05)),(to_sfixed_a(7.746441406197846e-05)),(to_sfixed_a(-2.9945025744382292e-05)),(to_sfixed_a(2.939319165307097e-05)),(to_sfixed_a(-3.781196937779896e-05)),(to_sfixed_a(5.112704457133077e-05)),(to_sfixed_a(-8.592804806539789e-05)),(to_sfixed_a(2.7870941266883165e-05)),(to_sfixed_a(3.5500704598234734e-06)),(to_sfixed_a(-1.9953611626988277e-05)),(to_sfixed_a(-5.816826887894422e-05)),(to_sfixed_a(5.159451757208444e-05)),(to_sfixed_a(7.033627480268478e-05)),(to_sfixed_a(0.00011299138714093715)),(to_sfixed_a(4.815321881324053e-05)),(to_sfixed_a(-4.325525515014306e-05)),(to_sfixed_a(3.782701605814509e-05)),(to_sfixed_a(3.6331432056613266e-05)));

    constant weight_n1_78 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.18302883207798004)),(to_sfixed_a(-0.10424985736608505)),(to_sfixed_a(0.2961113452911377)),(to_sfixed_a(0.14406709372997284)),(to_sfixed_a(-0.09612758457660675)),(to_sfixed_a(-0.25330862402915955)),(to_sfixed_a(-0.030055377632379532)),(to_sfixed_a(0.02246663346886635)),(to_sfixed_a(-0.012520184740424156)),(to_sfixed_a(-0.010443153791129589)),(to_sfixed_a(0.04309825226664543)),(to_sfixed_a(0.16211235523223877)),(to_sfixed_a(0.31473344564437866)),(to_sfixed_a(0.11583203822374344)),(to_sfixed_a(0.05188960209488869)),(to_sfixed_a(-0.012521804310381413)),(to_sfixed_a(-0.04751995578408241)),(to_sfixed_a(0.08401121944189072)),(to_sfixed_a(0.09116285294294357)),(to_sfixed_a(0.019986068829894066)),(to_sfixed_a(0.05008716508746147)),(to_sfixed_a(0.12647530436515808)),(to_sfixed_a(-0.03127451613545418)),(to_sfixed_a(0.024048740044236183)),(to_sfixed_a(-0.021299388259649277)),(to_sfixed_a(-0.22531667351722717)),(to_sfixed_a(-0.0451870858669281)),(to_sfixed_a(0.10360871255397797)),(to_sfixed_a(0.11715283989906311)),(to_sfixed_a(0.2787306010723114)),(to_sfixed_a(0.021968776360154152)),(to_sfixed_a(0.14582963287830353)),(to_sfixed_a(-0.06123623996973038)),(to_sfixed_a(0.12040628492832184)),(to_sfixed_a(0.09730522334575653)),(to_sfixed_a(0.14614270627498627)),(to_sfixed_a(-0.026425234973430634)),(to_sfixed_a(0.0916924923658371)));

    constant weight_n1_79 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.15201020240783691)),(to_sfixed_a(0.011255784891545773)),(to_sfixed_a(-0.014154440723359585)),(to_sfixed_a(-0.00631289416924119)),(to_sfixed_a(-0.00417175842449069)),(to_sfixed_a(0.025416914373636246)),(to_sfixed_a(0.003359974827617407)),(to_sfixed_a(0.0025030774995684624)),(to_sfixed_a(0.008829963393509388)),(to_sfixed_a(-0.0034676683135330677)),(to_sfixed_a(0.012273515574634075)),(to_sfixed_a(-0.015593121759593487)),(to_sfixed_a(-0.026817940175533295)),(to_sfixed_a(-0.007796221878379583)),(to_sfixed_a(0.0019522439688444138)),(to_sfixed_a(-0.012521602213382721)),(to_sfixed_a(-0.0011742357164621353)),(to_sfixed_a(0.0007448348915204406)),(to_sfixed_a(-0.006285522133111954)),(to_sfixed_a(-0.0031184705439954996)),(to_sfixed_a(0.007146394811570644)),(to_sfixed_a(-0.014036660082638264)),(to_sfixed_a(0.0021426372695714235)),(to_sfixed_a(-0.009662489406764507)),(to_sfixed_a(0.007406656630337238)),(to_sfixed_a(-0.010385435074567795)),(to_sfixed_a(-0.008228827267885208)),(to_sfixed_a(-0.004252637270838022)),(to_sfixed_a(0.002420805860310793)),(to_sfixed_a(-0.022688567638397217)),(to_sfixed_a(-0.01071985624730587)),(to_sfixed_a(-0.015885110944509506)),(to_sfixed_a(0.004519769921898842)),(to_sfixed_a(-0.01012544333934784)),(to_sfixed_a(0.025504522025585175)),(to_sfixed_a(0.00415379973128438)),(to_sfixed_a(-0.000262377638136968)),(to_sfixed_a(-0.013973761349916458)));

    constant weight_n1_80 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.10035869479179382)),(to_sfixed_a(3.780127735808492e-05)),(to_sfixed_a(-3.473725155345164e-05)),(to_sfixed_a(-7.892719622759614e-06)),(to_sfixed_a(3.856083276332356e-05)),(to_sfixed_a(1.1870905609612237e-06)),(to_sfixed_a(1.8876849935622886e-05)),(to_sfixed_a(6.164491992421972e-07)),(to_sfixed_a(4.024658119305968e-05)),(to_sfixed_a(-2.0453138859011233e-05)),(to_sfixed_a(-6.523432239191607e-05)),(to_sfixed_a(3.3351732326991623e-06)),(to_sfixed_a(-3.866711995215155e-05)),(to_sfixed_a(1.6109570424305275e-05)),(to_sfixed_a(7.348476356128231e-05)),(to_sfixed_a(-4.623668792191893e-05)),(to_sfixed_a(8.246724610216916e-05)),(to_sfixed_a(4.088501736987382e-05)),(to_sfixed_a(-6.90708384354366e-06)),(to_sfixed_a(1.0793450201163068e-05)),(to_sfixed_a(-1.4642621863458771e-05)),(to_sfixed_a(0.00012700256775133312)),(to_sfixed_a(7.866461237426847e-05)),(to_sfixed_a(-3.912859028787352e-05)),(to_sfixed_a(-4.290306969778612e-05)),(to_sfixed_a(9.471938028582372e-06)),(to_sfixed_a(4.2610805394360796e-05)),(to_sfixed_a(-2.551834040787071e-05)),(to_sfixed_a(-9.246122499462217e-05)),(to_sfixed_a(-7.623061537742615e-05)),(to_sfixed_a(4.057713158545084e-05)),(to_sfixed_a(3.627215119195171e-05)),(to_sfixed_a(-6.438461241486948e-06)),(to_sfixed_a(9.96910998196654e-09)),(to_sfixed_a(4.011119744973257e-05)),(to_sfixed_a(-1.2177624739706516e-05)),(to_sfixed_a(-3.629134880611673e-05)),(to_sfixed_a(3.0011264243512414e-05)));

    constant weight_n1_81 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.2509784996509552)),(to_sfixed_a(0.27725300192832947)),(to_sfixed_a(-0.08359826356172562)),(to_sfixed_a(0.07927782833576202)),(to_sfixed_a(-0.27644509077072144)),(to_sfixed_a(-0.06478491425514221)),(to_sfixed_a(-0.06683167070150375)),(to_sfixed_a(0.20329393446445465)),(to_sfixed_a(-0.11290600895881653)),(to_sfixed_a(-0.12874142825603485)),(to_sfixed_a(-0.05420779064297676)),(to_sfixed_a(0.05153267830610275)),(to_sfixed_a(0.13499857485294342)),(to_sfixed_a(0.1051950454711914)),(to_sfixed_a(0.025617578998208046)),(to_sfixed_a(0.0781463086605072)),(to_sfixed_a(0.030843017622828484)),(to_sfixed_a(0.029357561841607094)),(to_sfixed_a(0.17444278299808502)),(to_sfixed_a(0.047106459736824036)),(to_sfixed_a(-0.11934797465801239)),(to_sfixed_a(-0.1336418241262436)),(to_sfixed_a(-0.005289128050208092)),(to_sfixed_a(-0.2478068619966507)),(to_sfixed_a(0.19044002890586853)),(to_sfixed_a(-0.028634415939450264)),(to_sfixed_a(0.03319454938173294)),(to_sfixed_a(0.17684531211853027)),(to_sfixed_a(-0.030607091262936592)),(to_sfixed_a(-0.06979363411664963)),(to_sfixed_a(0.2204357236623764)),(to_sfixed_a(0.10182870924472809)),(to_sfixed_a(-0.1781836450099945)),(to_sfixed_a(0.11138378083705902)),(to_sfixed_a(-0.03435378149151802)),(to_sfixed_a(0.09302861988544464)),(to_sfixed_a(0.03208814188838005)),(to_sfixed_a(-0.07238547503948212)));

    constant weight_n1_82 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.07188867032527924)),(to_sfixed_a(0.030621174722909927)),(to_sfixed_a(0.0336703397333622)),(to_sfixed_a(0.0316285714507103)),(to_sfixed_a(-0.05079583451151848)),(to_sfixed_a(0.008595772087574005)),(to_sfixed_a(0.05091763660311699)),(to_sfixed_a(0.008216110989451408)),(to_sfixed_a(-0.02948288433253765)),(to_sfixed_a(-0.02585504949092865)),(to_sfixed_a(-0.020030563697218895)),(to_sfixed_a(0.054096635431051254)),(to_sfixed_a(-0.007678465452045202)),(to_sfixed_a(-0.02909964881837368)),(to_sfixed_a(0.017146021127700806)),(to_sfixed_a(-0.008992500603199005)),(to_sfixed_a(-0.017790446057915688)),(to_sfixed_a(-0.014581877738237381)),(to_sfixed_a(-0.09079005569219589)),(to_sfixed_a(-0.01160577591508627)),(to_sfixed_a(0.045786865055561066)),(to_sfixed_a(-0.01111601386219263)),(to_sfixed_a(0.03565646708011627)),(to_sfixed_a(0.020224163308739662)),(to_sfixed_a(0.022221826016902924)),(to_sfixed_a(-0.029682591557502747)),(to_sfixed_a(0.10099398344755173)),(to_sfixed_a(-0.04923476278781891)),(to_sfixed_a(0.02295028418302536)),(to_sfixed_a(0.011893647722899914)),(to_sfixed_a(-0.07968346774578094)),(to_sfixed_a(0.042099129408597946)),(to_sfixed_a(0.08194930106401443)),(to_sfixed_a(0.08703327924013138)),(to_sfixed_a(-0.009703213348984718)),(to_sfixed_a(0.09362587332725525)),(to_sfixed_a(0.0596235916018486)),(to_sfixed_a(-0.0374637134373188)));

    constant weight_n1_83 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.03390519693493843)),(to_sfixed_a(7.791625648678746e-06)),(to_sfixed_a(2.1774838387500495e-05)),(to_sfixed_a(3.671992089948617e-05)),(to_sfixed_a(-1.6502550352015533e-05)),(to_sfixed_a(-1.1410904335207306e-05)),(to_sfixed_a(2.6614552552928217e-06)),(to_sfixed_a(4.885668749921024e-05)),(to_sfixed_a(-3.185091190971434e-05)),(to_sfixed_a(-1.8505987100070342e-05)),(to_sfixed_a(3.0494922611978836e-05)),(to_sfixed_a(-1.1608466593315825e-05)),(to_sfixed_a(-3.792323332163505e-05)),(to_sfixed_a(-2.7300009151076665e-06)),(to_sfixed_a(-7.322012970689684e-05)),(to_sfixed_a(-2.4001888959901407e-05)),(to_sfixed_a(-1.3607826986117288e-05)),(to_sfixed_a(-5.512291318154894e-05)),(to_sfixed_a(-5.1617342251120135e-05)),(to_sfixed_a(-7.398921297863126e-05)),(to_sfixed_a(4.604981586453505e-05)),(to_sfixed_a(-3.366059536347166e-05)),(to_sfixed_a(-7.376731082331389e-05)),(to_sfixed_a(-3.47252243955154e-05)),(to_sfixed_a(1.1588012057472952e-05)),(to_sfixed_a(-4.207947858958505e-05)),(to_sfixed_a(1.6792992028058507e-05)),(to_sfixed_a(-9.208300070895348e-06)),(to_sfixed_a(1.7425067198928446e-05)),(to_sfixed_a(2.122803380188998e-05)),(to_sfixed_a(-3.451175143709406e-05)),(to_sfixed_a(6.14916134509258e-05)),(to_sfixed_a(8.334415724675637e-06)),(to_sfixed_a(-6.46893386146985e-05)),(to_sfixed_a(7.480188651243225e-05)),(to_sfixed_a(9.045621141012816e-07)),(to_sfixed_a(4.7355671995319426e-05)),(to_sfixed_a(-4.448660183697939e-05)));

    constant weight_n1_84 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.3384105861186981)),(to_sfixed_a(0.014084475114941597)),(to_sfixed_a(0.04407687485218048)),(to_sfixed_a(0.0991910770535469)),(to_sfixed_a(0.044490013271570206)),(to_sfixed_a(0.13045291602611542)),(to_sfixed_a(-0.03102361597120762)),(to_sfixed_a(0.009584181010723114)),(to_sfixed_a(0.009781359694898129)),(to_sfixed_a(-0.02566930651664734)),(to_sfixed_a(-0.011304670944809914)),(to_sfixed_a(-0.03731578588485718)),(to_sfixed_a(-0.006079232785850763)),(to_sfixed_a(0.02960256300866604)),(to_sfixed_a(0.0020792766008526087)),(to_sfixed_a(-0.01609220914542675)),(to_sfixed_a(-0.06325317174196243)),(to_sfixed_a(0.032132215797901154)),(to_sfixed_a(-0.022574134171009064)),(to_sfixed_a(-0.009333678521215916)),(to_sfixed_a(-0.010209983214735985)),(to_sfixed_a(-0.0072307707741856575)),(to_sfixed_a(0.02737307734787464)),(to_sfixed_a(0.0002816575870383531)),(to_sfixed_a(-0.011304432526230812)),(to_sfixed_a(0.02858590893447399)),(to_sfixed_a(-0.019521605223417282)),(to_sfixed_a(-0.02335743047297001)),(to_sfixed_a(0.04620889946818352)),(to_sfixed_a(0.04553570598363876)),(to_sfixed_a(-0.014293951913714409)),(to_sfixed_a(-0.08834795653820038)),(to_sfixed_a(-0.0396011658012867)),(to_sfixed_a(-0.023683372884988785)),(to_sfixed_a(-0.01704283617436886)),(to_sfixed_a(-0.010376404970884323)),(to_sfixed_a(-0.041825778782367706)),(to_sfixed_a(0.03918694704771042)));

    constant weight_n1_85 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.179833322763443)),(to_sfixed_a(-0.1257830709218979)),(to_sfixed_a(-0.08220607042312622)),(to_sfixed_a(0.07778328657150269)),(to_sfixed_a(-0.03598235920071602)),(to_sfixed_a(-0.03403109684586525)),(to_sfixed_a(0.030764136463403702)),(to_sfixed_a(0.005688684526830912)),(to_sfixed_a(0.09337769448757172)),(to_sfixed_a(0.016145825386047363)),(to_sfixed_a(-0.10158335417509079)),(to_sfixed_a(-0.0537961944937706)),(to_sfixed_a(0.03171314299106598)),(to_sfixed_a(0.014802265912294388)),(to_sfixed_a(0.09773781150579453)),(to_sfixed_a(0.0030098427087068558)),(to_sfixed_a(0.011095959693193436)),(to_sfixed_a(0.06906336545944214)),(to_sfixed_a(0.05380471795797348)),(to_sfixed_a(0.1371902972459793)),(to_sfixed_a(-0.02700357511639595)),(to_sfixed_a(0.0036024493165314198)),(to_sfixed_a(0.24951763451099396)),(to_sfixed_a(0.07679814100265503)),(to_sfixed_a(0.02469036914408207)),(to_sfixed_a(0.09672512114048004)),(to_sfixed_a(0.03685907647013664)),(to_sfixed_a(0.06741365045309067)),(to_sfixed_a(-0.17281940579414368)),(to_sfixed_a(-0.09958866238594055)),(to_sfixed_a(-0.07156626880168915)),(to_sfixed_a(0.1798466145992279)),(to_sfixed_a(0.17210231721401215)),(to_sfixed_a(-0.18187086284160614)),(to_sfixed_a(0.014844094403088093)),(to_sfixed_a(0.008786492981016636)),(to_sfixed_a(-0.04563109576702118)),(to_sfixed_a(-0.055336613208055496)));

    constant weight_n1_86 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.40086254477500916)),(to_sfixed_a(0.005186408758163452)),(to_sfixed_a(0.007991754449903965)),(to_sfixed_a(0.0275771114975214)),(to_sfixed_a(-0.015020010061562061)),(to_sfixed_a(-0.048346202820539474)),(to_sfixed_a(-0.045041490346193314)),(to_sfixed_a(0.013526994735002518)),(to_sfixed_a(0.09621106088161469)),(to_sfixed_a(-0.023891830816864967)),(to_sfixed_a(0.0031679319217801094)),(to_sfixed_a(-0.005817311350256205)),(to_sfixed_a(-0.0008789430721662939)),(to_sfixed_a(0.0722803920507431)),(to_sfixed_a(0.07015548646450043)),(to_sfixed_a(0.025605961680412292)),(to_sfixed_a(-0.029548337683081627)),(to_sfixed_a(-0.05781044065952301)),(to_sfixed_a(0.04034144803881645)),(to_sfixed_a(0.0203971229493618)),(to_sfixed_a(-0.03340433910489082)),(to_sfixed_a(-0.018671346828341484)),(to_sfixed_a(0.02680034190416336)),(to_sfixed_a(-0.008493627421557903)),(to_sfixed_a(-0.049977757036685944)),(to_sfixed_a(-0.04935380443930626)),(to_sfixed_a(0.048300616443157196)),(to_sfixed_a(-0.012257871218025684)),(to_sfixed_a(0.013195338658988476)),(to_sfixed_a(0.06256324797868729)),(to_sfixed_a(0.008068644441664219)),(to_sfixed_a(-0.014241809025406837)),(to_sfixed_a(-0.026095803827047348)),(to_sfixed_a(0.019618941470980644)),(to_sfixed_a(0.0719703882932663)),(to_sfixed_a(-0.004300993401557207)),(to_sfixed_a(-0.03368010371923447)),(to_sfixed_a(-0.020636219531297684)));

    constant weight_n1_87 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.14297477900981903)),(to_sfixed_a(2.441757715132553e-06)),(to_sfixed_a(-5.27388729096856e-05)),(to_sfixed_a(7.719941095274407e-06)),(to_sfixed_a(1.0297918379365001e-05)),(to_sfixed_a(2.6742542104329914e-05)),(to_sfixed_a(1.8980073946295306e-05)),(to_sfixed_a(2.33897335419897e-05)),(to_sfixed_a(6.0112146456958726e-05)),(to_sfixed_a(-9.027341548062395e-06)),(to_sfixed_a(3.1485376439377433e-06)),(to_sfixed_a(-8.968353540694807e-06)),(to_sfixed_a(7.184342848631786e-06)),(to_sfixed_a(-5.8001355682790745e-06)),(to_sfixed_a(1.3372876310313586e-05)),(to_sfixed_a(-8.669298404129222e-05)),(to_sfixed_a(2.637893339851871e-05)),(to_sfixed_a(4.344222543295473e-05)),(to_sfixed_a(-3.95190145354718e-05)),(to_sfixed_a(5.339904600987211e-05)),(to_sfixed_a(-1.9629851522040553e-05)),(to_sfixed_a(-3.1114803277887404e-05)),(to_sfixed_a(4.281218207324855e-05)),(to_sfixed_a(-7.077049758663634e-06)),(to_sfixed_a(-1.0655272490112111e-05)),(to_sfixed_a(-4.09851418226026e-05)),(to_sfixed_a(-5.6713914091233164e-05)),(to_sfixed_a(5.16033724125009e-05)),(to_sfixed_a(-0.00011902629194082692)),(to_sfixed_a(6.434482202166691e-05)),(to_sfixed_a(0.00013237344683147967)),(to_sfixed_a(6.9071252255525906e-06)),(to_sfixed_a(9.395218512509018e-05)),(to_sfixed_a(9.459762077312917e-05)),(to_sfixed_a(-2.5250488761230372e-05)),(to_sfixed_a(1.8728769646259025e-05)),(to_sfixed_a(7.55350265535526e-05)),(to_sfixed_a(-6.922057218616828e-05)));

    constant weight_n1_88 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.18598711490631104)),(to_sfixed_a(-5.050479376222938e-05)),(to_sfixed_a(3.522997576510534e-05)),(to_sfixed_a(-2.470292747602798e-05)),(to_sfixed_a(-3.590504275052808e-05)),(to_sfixed_a(9.57129850576166e-06)),(to_sfixed_a(1.2818527466151863e-05)),(to_sfixed_a(2.121715442626737e-05)),(to_sfixed_a(2.0462490283534862e-05)),(to_sfixed_a(2.0071089238626882e-05)),(to_sfixed_a(5.343676821212284e-05)),(to_sfixed_a(6.170755659695715e-05)),(to_sfixed_a(-6.468054925790057e-05)),(to_sfixed_a(-1.4228650798031595e-05)),(to_sfixed_a(5.6397943808406126e-06)),(to_sfixed_a(2.5243271011277102e-05)),(to_sfixed_a(1.0407724403194152e-05)),(to_sfixed_a(3.747004666365683e-05)),(to_sfixed_a(-1.0411884431960061e-05)),(to_sfixed_a(4.6321802074089646e-05)),(to_sfixed_a(-2.8983557058381848e-05)),(to_sfixed_a(-3.965282303397544e-05)),(to_sfixed_a(-4.1650688217487186e-05)),(to_sfixed_a(3.289306550868787e-05)),(to_sfixed_a(-6.532274710480124e-05)),(to_sfixed_a(-0.00010969312279485166)),(to_sfixed_a(-6.277955253608525e-05)),(to_sfixed_a(-2.587528433650732e-05)),(to_sfixed_a(-4.458893454284407e-05)),(to_sfixed_a(-3.107049997197464e-05)),(to_sfixed_a(-4.9116391892312095e-05)),(to_sfixed_a(-0.00012621242785826325)),(to_sfixed_a(7.232677307911217e-05)),(to_sfixed_a(1.4401866792468354e-06)),(to_sfixed_a(1.57683166435163e-06)),(to_sfixed_a(-2.578911153250374e-05)),(to_sfixed_a(5.883945050300099e-05)),(to_sfixed_a(-1.1215533049835358e-05)));

    constant weight_n1_89 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.2639009356498718)),(to_sfixed_a(-0.013977156020700932)),(to_sfixed_a(0.10137099027633667)),(to_sfixed_a(0.05199163779616356)),(to_sfixed_a(0.06945499032735825)),(to_sfixed_a(0.02429996058344841)),(to_sfixed_a(0.042274314910173416)),(to_sfixed_a(0.06300552189350128)),(to_sfixed_a(-0.03687789663672447)),(to_sfixed_a(-0.030579829588532448)),(to_sfixed_a(-0.17605651915073395)),(to_sfixed_a(-0.06408483535051346)),(to_sfixed_a(0.03533345088362694)),(to_sfixed_a(0.24608959257602692)),(to_sfixed_a(-0.3445795774459839)),(to_sfixed_a(-0.08556760102510452)),(to_sfixed_a(-0.021318236365914345)),(to_sfixed_a(0.07500114291906357)),(to_sfixed_a(-0.07949598133563995)),(to_sfixed_a(-0.17141962051391602)),(to_sfixed_a(-0.10539696365594864)),(to_sfixed_a(0.07237330079078674)),(to_sfixed_a(-0.02859978750348091)),(to_sfixed_a(0.20633968710899353)),(to_sfixed_a(-0.09654109179973602)),(to_sfixed_a(0.23975111544132233)),(to_sfixed_a(0.018729163333773613)),(to_sfixed_a(0.02237667888402939)),(to_sfixed_a(0.04985401779413223)),(to_sfixed_a(0.004093020223081112)),(to_sfixed_a(0.012492476962506771)),(to_sfixed_a(0.02835710346698761)),(to_sfixed_a(0.05931255966424942)),(to_sfixed_a(0.045157574117183685)),(to_sfixed_a(-0.023357879370450974)),(to_sfixed_a(-0.008664256893098354)),(to_sfixed_a(-0.2113082855939865)),(to_sfixed_a(-0.07689855247735977)));

    constant weight_n1_90 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.01397317461669445)),(to_sfixed_a(-5.763869467045879e-06)),(to_sfixed_a(5.4228421504376456e-05)),(to_sfixed_a(-7.958787136885803e-06)),(to_sfixed_a(-3.914824901585234e-06)),(to_sfixed_a(2.6453513783053495e-05)),(to_sfixed_a(1.8377295418758877e-05)),(to_sfixed_a(8.240245369961485e-05)),(to_sfixed_a(-3.42426574206911e-05)),(to_sfixed_a(-1.5047364286147058e-05)),(to_sfixed_a(-2.439318450342398e-05)),(to_sfixed_a(-3.401676440262236e-05)),(to_sfixed_a(-6.532689440064132e-05)),(to_sfixed_a(6.060115265427157e-05)),(to_sfixed_a(5.7240104069933295e-05)),(to_sfixed_a(5.418630098574795e-05)),(to_sfixed_a(4.226419696351513e-05)),(to_sfixed_a(-1.5657804397051223e-05)),(to_sfixed_a(0.00010628943709889427)),(to_sfixed_a(-3.28673304466065e-05)),(to_sfixed_a(8.460585377179086e-05)),(to_sfixed_a(-1.114586484618485e-05)),(to_sfixed_a(3.6080742574995384e-05)),(to_sfixed_a(6.868909258628264e-05)),(to_sfixed_a(-1.778713703970425e-05)),(to_sfixed_a(3.5631706850836053e-05)),(to_sfixed_a(2.919230973930098e-05)),(to_sfixed_a(-3.570337139535695e-05)),(to_sfixed_a(2.430095264571719e-06)),(to_sfixed_a(5.572058944380842e-05)),(to_sfixed_a(-2.4945644327090122e-05)),(to_sfixed_a(5.117378168506548e-05)),(to_sfixed_a(6.207801925484091e-05)),(to_sfixed_a(-6.241867959033698e-05)),(to_sfixed_a(-3.3094252103182953e-06)),(to_sfixed_a(1.3488877357303863e-06)),(to_sfixed_a(4.899083432974294e-05)),(to_sfixed_a(6.615971506107599e-05)));

    constant weight_n1_91 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.2417590618133545)),(to_sfixed_a(-0.010187830775976181)),(to_sfixed_a(-0.04451616853475571)),(to_sfixed_a(-0.004321523010730743)),(to_sfixed_a(0.04234263300895691)),(to_sfixed_a(0.0083008436486125)),(to_sfixed_a(-0.06163568049669266)),(to_sfixed_a(0.04177282005548477)),(to_sfixed_a(0.035386279225349426)),(to_sfixed_a(-0.015179627574980259)),(to_sfixed_a(0.007390317041426897)),(to_sfixed_a(-0.013968744315207005)),(to_sfixed_a(0.007384362630546093)),(to_sfixed_a(0.04287330061197281)),(to_sfixed_a(0.015726590529084206)),(to_sfixed_a(-0.09113836288452148)),(to_sfixed_a(0.0197521410882473)),(to_sfixed_a(-0.013800323940813541)),(to_sfixed_a(-0.02224653773009777)),(to_sfixed_a(0.011374100111424923)),(to_sfixed_a(-0.05968668684363365)),(to_sfixed_a(0.014362704008817673)),(to_sfixed_a(-0.06606251746416092)),(to_sfixed_a(-0.09855332225561142)),(to_sfixed_a(0.11138497292995453)),(to_sfixed_a(0.005910507403314114)),(to_sfixed_a(0.01630828157067299)),(to_sfixed_a(-0.11543598771095276)),(to_sfixed_a(-0.026047373190522194)),(to_sfixed_a(-0.006253812927752733)),(to_sfixed_a(-0.00984315387904644)),(to_sfixed_a(0.05135586857795715)),(to_sfixed_a(0.026926672086119652)),(to_sfixed_a(-0.019768238067626953)),(to_sfixed_a(0.08373171836137772)),(to_sfixed_a(-0.06920020282268524)),(to_sfixed_a(0.013754917308688164)),(to_sfixed_a(-0.03300435096025467)));

    constant weight_n1_92 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.0218121949583292)),(to_sfixed_a(2.0170989955659024e-05)),(to_sfixed_a(-3.280414966866374e-05)),(to_sfixed_a(-1.0243168617307674e-05)),(to_sfixed_a(1.9519386114552617e-05)),(to_sfixed_a(2.023242814175319e-05)),(to_sfixed_a(-1.3394748748396523e-05)),(to_sfixed_a(-4.3703032133635134e-05)),(to_sfixed_a(2.1154130081413314e-05)),(to_sfixed_a(4.4865981180919334e-05)),(to_sfixed_a(-5.213536041992484e-06)),(to_sfixed_a(4.052494477946311e-05)),(to_sfixed_a(3.1487459636991844e-05)),(to_sfixed_a(-4.019042171421461e-05)),(to_sfixed_a(-2.818745997501537e-06)),(to_sfixed_a(3.0941669137973804e-06)),(to_sfixed_a(-3.781053237617016e-06)),(to_sfixed_a(-4.1336312278872356e-05)),(to_sfixed_a(5.5150725529529154e-05)),(to_sfixed_a(-1.4907081094861496e-05)),(to_sfixed_a(-7.439322416757932e-06)),(to_sfixed_a(-3.9768045098753646e-05)),(to_sfixed_a(4.54694963991642e-05)),(to_sfixed_a(3.368063516973052e-07)),(to_sfixed_a(-7.930881838547066e-05)),(to_sfixed_a(4.364213964436203e-06)),(to_sfixed_a(6.933351414772915e-06)),(to_sfixed_a(-1.1030288987967651e-05)),(to_sfixed_a(-1.269897347810911e-05)),(to_sfixed_a(3.1342515285359696e-05)),(to_sfixed_a(7.804369488439988e-06)),(to_sfixed_a(-4.439019176061265e-05)),(to_sfixed_a(3.196535908500664e-05)),(to_sfixed_a(4.2412200855324045e-05)),(to_sfixed_a(4.206318044452928e-05)),(to_sfixed_a(-6.603623205592157e-06)),(to_sfixed_a(-2.08674136956688e-05)),(to_sfixed_a(5.751047410740284e-06)));

    constant weight_n1_93 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.29345107078552246)),(to_sfixed_a(-0.01027009915560484)),(to_sfixed_a(0.031460609287023544)),(to_sfixed_a(0.021131347864866257)),(to_sfixed_a(-0.06416763365268707)),(to_sfixed_a(-0.007310963235795498)),(to_sfixed_a(0.04067198187112808)),(to_sfixed_a(-0.026740161702036858)),(to_sfixed_a(-0.038330353796482086)),(to_sfixed_a(0.003717962419614196)),(to_sfixed_a(-0.06160745397210121)),(to_sfixed_a(0.00663868710398674)),(to_sfixed_a(-0.07456626743078232)),(to_sfixed_a(-0.041292402893304825)),(to_sfixed_a(0.04793568700551987)),(to_sfixed_a(0.03885607421398163)),(to_sfixed_a(-0.010796032845973969)),(to_sfixed_a(-0.033081624656915665)),(to_sfixed_a(0.030296145007014275)),(to_sfixed_a(0.06299217790365219)),(to_sfixed_a(-0.01891152746975422)),(to_sfixed_a(0.06946737319231033)),(to_sfixed_a(0.02629389427602291)),(to_sfixed_a(0.02618350088596344)),(to_sfixed_a(-0.03149513900279999)),(to_sfixed_a(0.05435282737016678)),(to_sfixed_a(-0.05682148039340973)),(to_sfixed_a(0.02885117381811142)),(to_sfixed_a(-0.05139870569109917)),(to_sfixed_a(0.11259973049163818)),(to_sfixed_a(-0.03535280004143715)),(to_sfixed_a(-0.13062156736850739)),(to_sfixed_a(-0.025047466158866882)),(to_sfixed_a(-0.04253844544291496)),(to_sfixed_a(0.032887618988752365)),(to_sfixed_a(0.017913948744535446)),(to_sfixed_a(-0.021529126912355423)),(to_sfixed_a(-0.022647950798273087)));

    constant weight_n1_94 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.16578339040279388)),(to_sfixed_a(0.003055874491110444)),(to_sfixed_a(-0.00045247634989209473)),(to_sfixed_a(-0.004258969333022833)),(to_sfixed_a(0.0075408658012747765)),(to_sfixed_a(-0.0015724677359685302)),(to_sfixed_a(0.001000222866423428)),(to_sfixed_a(0.00403329823166132)),(to_sfixed_a(-0.006261077243834734)),(to_sfixed_a(0.001555105671286583)),(to_sfixed_a(0.008873896673321724)),(to_sfixed_a(-0.00081034837057814)),(to_sfixed_a(0.004011866170912981)),(to_sfixed_a(0.00982827041298151)),(to_sfixed_a(0.002660309663042426)),(to_sfixed_a(0.003466569120064378)),(to_sfixed_a(0.001818910357542336)),(to_sfixed_a(-0.007546194829046726)),(to_sfixed_a(-0.0005611838423646986)),(to_sfixed_a(0.005861714947968721)),(to_sfixed_a(0.0006913284887559712)),(to_sfixed_a(-0.001751057105138898)),(to_sfixed_a(-0.004273240454494953)),(to_sfixed_a(0.003998854663223028)),(to_sfixed_a(-0.005966091528534889)),(to_sfixed_a(-0.00027722076629288495)),(to_sfixed_a(0.0036416940856724977)),(to_sfixed_a(-0.010775450617074966)),(to_sfixed_a(0.008052285760641098)),(to_sfixed_a(-0.002808439778164029)),(to_sfixed_a(0.00950173381716013)),(to_sfixed_a(-0.0016748878406360745)),(to_sfixed_a(0.008043731562793255)),(to_sfixed_a(0.0056413160637021065)),(to_sfixed_a(0.003298538736999035)),(to_sfixed_a(0.0025214296765625477)),(to_sfixed_a(0.004568107891827822)),(to_sfixed_a(-0.0019517544424161315)));

    constant weight_n1_95 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.0157876405864954)),(to_sfixed_a(1.228505152539583e-05)),(to_sfixed_a(2.1589858079096302e-05)),(to_sfixed_a(-6.248259160201997e-05)),(to_sfixed_a(-6.41718861515983e-06)),(to_sfixed_a(-3.7362804050644627e-07)),(to_sfixed_a(1.1723736861313228e-05)),(to_sfixed_a(3.505072891130112e-05)),(to_sfixed_a(-7.902237121015787e-05)),(to_sfixed_a(3.168599141645245e-05)),(to_sfixed_a(-5.42207999387756e-06)),(to_sfixed_a(-1.0526408686928335e-06)),(to_sfixed_a(2.707671228563413e-05)),(to_sfixed_a(6.762857810826972e-05)),(to_sfixed_a(3.6555582028086064e-06)),(to_sfixed_a(3.239434590796009e-05)),(to_sfixed_a(-7.49822793295607e-05)),(to_sfixed_a(0.00011637403804343194)),(to_sfixed_a(1.1864614862133749e-05)),(to_sfixed_a(8.306041127070785e-05)),(to_sfixed_a(2.890647556341719e-05)),(to_sfixed_a(8.835992957756389e-06)),(to_sfixed_a(8.866829739417881e-05)),(to_sfixed_a(6.571038829861209e-05)),(to_sfixed_a(-1.1189032989022962e-07)),(to_sfixed_a(8.49716379889287e-05)),(to_sfixed_a(4.6818924602121115e-05)),(to_sfixed_a(-5.116267493576743e-05)),(to_sfixed_a(7.337737042689696e-05)),(to_sfixed_a(8.627587703813333e-06)),(to_sfixed_a(-0.00011096313392044976)),(to_sfixed_a(6.243019015528262e-05)),(to_sfixed_a(7.900931814219803e-05)),(to_sfixed_a(-5.4558673582505435e-05)),(to_sfixed_a(-0.00011679487943183631)),(to_sfixed_a(-4.381437611300498e-05)),(to_sfixed_a(-1.1022168564522872e-06)),(to_sfixed_a(9.66690913628554e-06)));

    constant weight_n1_96 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.010441077873110771)),(to_sfixed_a(-8.679360803398595e-07)),(to_sfixed_a(-2.438689534756122e-06)),(to_sfixed_a(8.605237962910905e-05)),(to_sfixed_a(-3.610278872656636e-05)),(to_sfixed_a(-4.409810935612768e-05)),(to_sfixed_a(5.886978760827333e-05)),(to_sfixed_a(5.9610647440422326e-05)),(to_sfixed_a(4.314966645324603e-05)),(to_sfixed_a(1.5882247680565342e-05)),(to_sfixed_a(-4.767225618707016e-05)),(to_sfixed_a(-1.7279060557484627e-05)),(to_sfixed_a(-2.4412753191427328e-05)),(to_sfixed_a(-2.9668464776477776e-05)),(to_sfixed_a(7.014643779257312e-05)),(to_sfixed_a(1.0957677659462206e-05)),(to_sfixed_a(2.4513199605280533e-05)),(to_sfixed_a(8.424976840615273e-05)),(to_sfixed_a(-1.7889957462102757e-06)),(to_sfixed_a(1.5075977898959536e-05)),(to_sfixed_a(-1.135587808676064e-05)),(to_sfixed_a(-3.927315628970973e-05)),(to_sfixed_a(7.653198554180562e-05)),(to_sfixed_a(-3.4293541830265895e-05)),(to_sfixed_a(-3.807968460023403e-05)),(to_sfixed_a(2.8613811082323082e-05)),(to_sfixed_a(-9.192972356686369e-06)),(to_sfixed_a(-1.761336716299411e-05)),(to_sfixed_a(-2.819679139065556e-07)),(to_sfixed_a(1.575196256453637e-05)),(to_sfixed_a(-4.782411633641459e-05)),(to_sfixed_a(-2.5683686544653028e-05)),(to_sfixed_a(2.6245787012157962e-05)),(to_sfixed_a(-1.1135059139633086e-05)),(to_sfixed_a(-3.4268825402250513e-05)),(to_sfixed_a(3.932640902348794e-05)),(to_sfixed_a(4.2686384404078126e-05)),(to_sfixed_a(-1.412511664966587e-05)));

    constant weight_n1_97 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.02439234033226967)),(to_sfixed_a(-2.2198810256668366e-05)),(to_sfixed_a(-4.6300513645292085e-07)),(to_sfixed_a(1.9921868442906998e-05)),(to_sfixed_a(-5.776020771008916e-06)),(to_sfixed_a(-1.8182710846303962e-05)),(to_sfixed_a(1.1008894034603145e-05)),(to_sfixed_a(-1.5970613276294898e-06)),(to_sfixed_a(1.4460175407293718e-05)),(to_sfixed_a(2.2471011106972583e-05)),(to_sfixed_a(-1.0489207852515392e-05)),(to_sfixed_a(1.1202589121239726e-05)),(to_sfixed_a(3.429493517614901e-05)),(to_sfixed_a(-3.304038546048105e-05)),(to_sfixed_a(4.792128493136261e-06)),(to_sfixed_a(-1.0882621609198395e-05)),(to_sfixed_a(4.071595685672946e-05)),(to_sfixed_a(6.696467607980594e-06)),(to_sfixed_a(2.8209849915583618e-05)),(to_sfixed_a(-1.599736606294755e-05)),(to_sfixed_a(-2.582963315944653e-05)),(to_sfixed_a(1.3573018122770009e-06)),(to_sfixed_a(-3.4122767829103395e-05)),(to_sfixed_a(-8.61989155964693e-06)),(to_sfixed_a(2.9699813239858486e-05)),(to_sfixed_a(4.896526297670789e-05)),(to_sfixed_a(1.2306742291912087e-06)),(to_sfixed_a(6.829637277405709e-05)),(to_sfixed_a(-8.483509009238333e-05)),(to_sfixed_a(-3.147800816805102e-05)),(to_sfixed_a(7.79425899963826e-05)),(to_sfixed_a(3.250458757975139e-05)),(to_sfixed_a(-3.8254456740105525e-05)),(to_sfixed_a(-6.227912672329694e-05)),(to_sfixed_a(-1.5514131519012153e-05)),(to_sfixed_a(-6.21470348960429e-07)),(to_sfixed_a(8.400400838581845e-05)),(to_sfixed_a(4.135953531658743e-06)));

    constant weight_n1_98 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.0880594253540039)),(to_sfixed_a(-1.826176594477147e-05)),(to_sfixed_a(-3.178785391355632e-06)),(to_sfixed_a(2.8496331651695073e-05)),(to_sfixed_a(-1.686688483459875e-05)),(to_sfixed_a(-7.028061372693628e-05)),(to_sfixed_a(-1.1094344699813519e-05)),(to_sfixed_a(-2.71532353508519e-05)),(to_sfixed_a(3.26891677104868e-05)),(to_sfixed_a(-4.8019752284744754e-05)),(to_sfixed_a(7.952700798341539e-06)),(to_sfixed_a(2.47995340032503e-05)),(to_sfixed_a(2.661819053173531e-05)),(to_sfixed_a(5.229489761404693e-05)),(to_sfixed_a(-3.408478733035736e-05)),(to_sfixed_a(-3.815053787548095e-05)),(to_sfixed_a(1.5140745745156892e-05)),(to_sfixed_a(-3.691051824716851e-05)),(to_sfixed_a(5.702573980670422e-05)),(to_sfixed_a(2.9334254577406682e-05)),(to_sfixed_a(1.4999312043073587e-05)),(to_sfixed_a(4.6047181967878714e-05)),(to_sfixed_a(1.4547436876455322e-05)),(to_sfixed_a(2.9558310416177846e-05)),(to_sfixed_a(8.941731721279211e-06)),(to_sfixed_a(-1.6960713765001856e-05)),(to_sfixed_a(-8.955697558121756e-05)),(to_sfixed_a(3.9566202758578584e-05)),(to_sfixed_a(-3.700489105540328e-05)),(to_sfixed_a(1.0182978257944342e-05)),(to_sfixed_a(2.948874134744983e-05)),(to_sfixed_a(-5.39998545718845e-05)),(to_sfixed_a(4.946520857629366e-05)),(to_sfixed_a(-7.03791156411171e-05)),(to_sfixed_a(-2.6304553102818318e-05)),(to_sfixed_a(-5.559992860071361e-05)),(to_sfixed_a(-0.00011859378719236702)),(to_sfixed_a(1.0299731911800336e-05)));

    constant weight_n1_99 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.0770823210477829)),(to_sfixed_a(0.012878193520009518)),(to_sfixed_a(-0.02999105490744114)),(to_sfixed_a(-0.050864461809396744)),(to_sfixed_a(-0.014979931525886059)),(to_sfixed_a(-0.12074223905801773)),(to_sfixed_a(-0.01285032369196415)),(to_sfixed_a(-0.03131883591413498)),(to_sfixed_a(0.004316536709666252)),(to_sfixed_a(0.0046687438152730465)),(to_sfixed_a(0.0022393502295017242)),(to_sfixed_a(0.0705641508102417)),(to_sfixed_a(0.02146926335990429)),(to_sfixed_a(-0.02287346124649048)),(to_sfixed_a(0.035408973693847656)),(to_sfixed_a(-0.06146415323019028)),(to_sfixed_a(-0.0035621062852442265)),(to_sfixed_a(-0.026304597035050392)),(to_sfixed_a(0.04038284346461296)),(to_sfixed_a(0.009692908264696598)),(to_sfixed_a(-0.03818816691637039)),(to_sfixed_a(0.04021620750427246)),(to_sfixed_a(-0.08029469847679138)),(to_sfixed_a(0.0110880546271801)),(to_sfixed_a(-0.012400957755744457)),(to_sfixed_a(0.03040415048599243)),(to_sfixed_a(0.010199880227446556)),(to_sfixed_a(0.04589640349149704)),(to_sfixed_a(-0.009091569110751152)),(to_sfixed_a(-0.058465439826250076)),(to_sfixed_a(0.05334959924221039)),(to_sfixed_a(0.010954564437270164)),(to_sfixed_a(0.22397324442863464)),(to_sfixed_a(0.004812576808035374)),(to_sfixed_a(0.038104794919490814)),(to_sfixed_a(0.02154441736638546)),(to_sfixed_a(-0.01159703265875578)),(to_sfixed_a(0.06674802303314209)));

    constant weight_n1_100 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.2761847972869873)),(to_sfixed_a(0.0024357845541089773)),(to_sfixed_a(-0.02075275219976902)),(to_sfixed_a(0.008368476293981075)),(to_sfixed_a(0.018743883818387985)),(to_sfixed_a(0.010640906170010567)),(to_sfixed_a(0.010246221907436848)),(to_sfixed_a(0.012497379444539547)),(to_sfixed_a(0.011264602653682232)),(to_sfixed_a(-0.015564294531941414)),(to_sfixed_a(0.026641717180609703)),(to_sfixed_a(0.0390767902135849)),(to_sfixed_a(-0.011204284615814686)),(to_sfixed_a(0.0132606765255332)),(to_sfixed_a(0.019180983304977417)),(to_sfixed_a(-0.027603808790445328)),(to_sfixed_a(-0.017139393836259842)),(to_sfixed_a(0.02309880591928959)),(to_sfixed_a(-0.020223088562488556)),(to_sfixed_a(-0.04549451172351837)),(to_sfixed_a(-0.0018181886989623308)),(to_sfixed_a(0.07044017314910889)),(to_sfixed_a(0.0066137006506323814)),(to_sfixed_a(-0.033805351704359055)),(to_sfixed_a(-0.06222274526953697)),(to_sfixed_a(0.015111596323549747)),(to_sfixed_a(-0.022157950326800346)),(to_sfixed_a(0.024277782067656517)),(to_sfixed_a(-0.012677638791501522)),(to_sfixed_a(-0.005166096147149801)),(to_sfixed_a(0.007284353952854872)),(to_sfixed_a(0.035453423857688904)),(to_sfixed_a(-0.004058453720062971)),(to_sfixed_a(0.008482053875923157)),(to_sfixed_a(0.023294761776924133)),(to_sfixed_a(0.0035849011037498713)),(to_sfixed_a(0.0049766856245696545)),(to_sfixed_a(0.07417024672031403)));

    constant weight_n1_101 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.01821056194603443)),(to_sfixed_a(-3.0517858249368146e-06)),(to_sfixed_a(4.26784208684694e-05)),(to_sfixed_a(1.4229805856302846e-05)),(to_sfixed_a(3.9691454730927944e-05)),(to_sfixed_a(-4.678200639318675e-05)),(to_sfixed_a(5.677806711901212e-06)),(to_sfixed_a(-1.2377038729027845e-05)),(to_sfixed_a(2.6700954549596645e-05)),(to_sfixed_a(-6.337792729027569e-05)),(to_sfixed_a(-1.85869666893268e-05)),(to_sfixed_a(2.331710447833757e-06)),(to_sfixed_a(5.7631285017123446e-05)),(to_sfixed_a(1.551249260955956e-05)),(to_sfixed_a(-2.0246456188033335e-05)),(to_sfixed_a(-3.863593519781716e-05)),(to_sfixed_a(0.00010159921657759696)),(to_sfixed_a(8.988918852992356e-05)),(to_sfixed_a(4.671430724556558e-05)),(to_sfixed_a(9.79769083642168e-06)),(to_sfixed_a(4.690045170718804e-05)),(to_sfixed_a(-3.52746901626233e-05)),(to_sfixed_a(4.740710573969409e-05)),(to_sfixed_a(-1.8558956071501598e-05)),(to_sfixed_a(9.032450179802254e-05)),(to_sfixed_a(-2.3930095267132856e-05)),(to_sfixed_a(3.0798124498687685e-05)),(to_sfixed_a(-7.522392024839064e-06)),(to_sfixed_a(6.501773168565705e-05)),(to_sfixed_a(-8.571689249947667e-05)),(to_sfixed_a(-1.0219490832241718e-05)),(to_sfixed_a(2.8763153750333004e-05)),(to_sfixed_a(-6.036456034053117e-05)),(to_sfixed_a(-4.792965773958713e-05)),(to_sfixed_a(-3.018480583705241e-06)),(to_sfixed_a(7.504375844291644e-06)),(to_sfixed_a(-5.2954492275603116e-05)),(to_sfixed_a(-2.9997756428201683e-05)));

    constant weight_n1_102 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.3543364703655243)),(to_sfixed_a(0.07742490619421005)),(to_sfixed_a(-0.06221909448504448)),(to_sfixed_a(-0.009114387445151806)),(to_sfixed_a(0.12428738176822662)),(to_sfixed_a(0.0011045727878808975)),(to_sfixed_a(-0.07654326409101486)),(to_sfixed_a(0.08350339531898499)),(to_sfixed_a(-0.020929070189595222)),(to_sfixed_a(0.020419850945472717)),(to_sfixed_a(-0.0056418427266180515)),(to_sfixed_a(-0.08191962540149689)),(to_sfixed_a(0.06962624192237854)),(to_sfixed_a(-0.04708578437566757)),(to_sfixed_a(0.1518445461988449)),(to_sfixed_a(-0.004839859902858734)),(to_sfixed_a(0.016669323667883873)),(to_sfixed_a(-0.05713057518005371)),(to_sfixed_a(0.006537014152854681)),(to_sfixed_a(-0.08601433038711548)),(to_sfixed_a(-0.0461336225271225)),(to_sfixed_a(0.12073294818401337)),(to_sfixed_a(0.0698198601603508)),(to_sfixed_a(0.028272302821278572)),(to_sfixed_a(0.01733451895415783)),(to_sfixed_a(0.07715790718793869)),(to_sfixed_a(-0.009274374693632126)),(to_sfixed_a(0.012469240464270115)),(to_sfixed_a(0.05874727666378021)),(to_sfixed_a(-0.02764306217432022)),(to_sfixed_a(0.08342170715332031)),(to_sfixed_a(0.2097431868314743)),(to_sfixed_a(0.12513434886932373)),(to_sfixed_a(0.02346920222043991)),(to_sfixed_a(0.025466080754995346)),(to_sfixed_a(0.18610677123069763)),(to_sfixed_a(0.05252327397465706)),(to_sfixed_a(0.043155573308467865)));

    constant weight_n1_103 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.06728865206241608)),(to_sfixed_a(-0.0037387129850685596)),(to_sfixed_a(-0.06665140390396118)),(to_sfixed_a(-0.0030426110606640577)),(to_sfixed_a(-0.08172410726547241)),(to_sfixed_a(0.06428758800029755)),(to_sfixed_a(-0.09180614352226257)),(to_sfixed_a(0.19839295744895935)),(to_sfixed_a(-0.1468803733587265)),(to_sfixed_a(0.04140009358525276)),(to_sfixed_a(-0.1826845109462738)),(to_sfixed_a(0.025067780166864395)),(to_sfixed_a(0.02131779119372368)),(to_sfixed_a(0.046981289982795715)),(to_sfixed_a(0.1103004515171051)),(to_sfixed_a(-0.09206991642713547)),(to_sfixed_a(0.07853057980537415)),(to_sfixed_a(-0.08301099389791489)),(to_sfixed_a(0.04308497533202171)),(to_sfixed_a(0.03923855349421501)),(to_sfixed_a(0.09481780230998993)),(to_sfixed_a(0.06784530729055405)),(to_sfixed_a(-0.020542217418551445)),(to_sfixed_a(0.15972909331321716)),(to_sfixed_a(-0.07886172086000443)),(to_sfixed_a(0.08357483893632889)),(to_sfixed_a(0.05139817297458649)),(to_sfixed_a(0.0893167182803154)),(to_sfixed_a(0.07908512651920319)),(to_sfixed_a(0.1619855910539627)),(to_sfixed_a(0.001943659270182252)),(to_sfixed_a(-0.10012548416852951)),(to_sfixed_a(-0.07264187186956406)),(to_sfixed_a(-0.04774734750390053)),(to_sfixed_a(0.0042585995979607105)),(to_sfixed_a(-0.151402547955513)),(to_sfixed_a(0.0829809382557869)),(to_sfixed_a(0.05592551827430725)));

    constant weight_n1_104 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.4173811972141266)),(to_sfixed_a(0.0031150677241384983)),(to_sfixed_a(0.0011701994808390737)),(to_sfixed_a(-0.004110924433916807)),(to_sfixed_a(-0.03192473575472832)),(to_sfixed_a(6.987257802393287e-05)),(to_sfixed_a(-0.014697092585265636)),(to_sfixed_a(0.015844034031033516)),(to_sfixed_a(0.014072899706661701)),(to_sfixed_a(-0.05034314841032028)),(to_sfixed_a(0.05157193914055824)),(to_sfixed_a(-0.006704343482851982)),(to_sfixed_a(0.02932453341782093)),(to_sfixed_a(0.020610889419913292)),(to_sfixed_a(-0.0035089957527816296)),(to_sfixed_a(-0.03586605563759804)),(to_sfixed_a(-0.009047362022101879)),(to_sfixed_a(0.01856962777674198)),(to_sfixed_a(-0.020244566723704338)),(to_sfixed_a(-0.0012113854754716158)),(to_sfixed_a(-0.009971274062991142)),(to_sfixed_a(-0.010037138126790524)),(to_sfixed_a(0.0228856410831213)),(to_sfixed_a(-0.07356815785169601)),(to_sfixed_a(-0.018361184746026993)),(to_sfixed_a(-0.012369714677333832)),(to_sfixed_a(-0.03774894028902054)),(to_sfixed_a(-0.03820202499628067)),(to_sfixed_a(0.06959155201911926)),(to_sfixed_a(-0.019799476489424706)),(to_sfixed_a(0.004672922194004059)),(to_sfixed_a(0.07189473509788513)),(to_sfixed_a(-0.0025405173655599356)),(to_sfixed_a(0.05639045313000679)),(to_sfixed_a(-0.020724667236208916)),(to_sfixed_a(-0.023449420928955078)),(to_sfixed_a(0.0005386954289861023)),(to_sfixed_a(0.0029115905053913593)));

    constant weight_n1_105 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.01435128878802061)),(to_sfixed_a(-6.425131141440943e-05)),(to_sfixed_a(1.9526622054399922e-05)),(to_sfixed_a(1.1468458069430199e-05)),(to_sfixed_a(5.787859481642954e-05)),(to_sfixed_a(2.0006931663374417e-05)),(to_sfixed_a(5.858168879058212e-05)),(to_sfixed_a(-2.6210103897028603e-05)),(to_sfixed_a(3.21552470268216e-05)),(to_sfixed_a(4.4019958295393735e-05)),(to_sfixed_a(6.22759253019467e-05)),(to_sfixed_a(2.697222043934744e-05)),(to_sfixed_a(4.7567526053171605e-05)),(to_sfixed_a(4.3112606363138184e-05)),(to_sfixed_a(-7.0772516664874274e-06)),(to_sfixed_a(1.3480886991601437e-05)),(to_sfixed_a(3.481258318061009e-05)),(to_sfixed_a(2.249727549497038e-05)),(to_sfixed_a(-2.0014544134028256e-05)),(to_sfixed_a(-1.5231496945489198e-05)),(to_sfixed_a(-7.775842823321e-05)),(to_sfixed_a(-5.331095280780573e-07)),(to_sfixed_a(3.8526763091795146e-05)),(to_sfixed_a(-8.933777280617505e-06)),(to_sfixed_a(3.2133884815266356e-06)),(to_sfixed_a(6.473841494880617e-05)),(to_sfixed_a(-4.125884061068064e-06)),(to_sfixed_a(5.677992885466665e-05)),(to_sfixed_a(7.156580068112817e-06)),(to_sfixed_a(2.8775608370779082e-05)),(to_sfixed_a(1.2596767192007974e-05)),(to_sfixed_a(7.391061808448285e-05)),(to_sfixed_a(-3.8390404370147735e-05)),(to_sfixed_a(3.5498269426170737e-05)),(to_sfixed_a(-4.8487450840184465e-05)),(to_sfixed_a(-2.2009182430338115e-05)),(to_sfixed_a(6.0426460549933836e-05)),(to_sfixed_a(-3.0276502002379857e-05)));

    constant weight_n1_106 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.24410243332386017)),(to_sfixed_a(-0.0015007787151262164)),(to_sfixed_a(0.0024289945140480995)),(to_sfixed_a(0.0031379081774502993)),(to_sfixed_a(-0.00822539534419775)),(to_sfixed_a(-0.0029686246998608112)),(to_sfixed_a(-0.0023576710373163223)),(to_sfixed_a(0.0013324099127203226)),(to_sfixed_a(0.010666346177458763)),(to_sfixed_a(0.0005407774588093162)),(to_sfixed_a(0.006878227926790714)),(to_sfixed_a(-0.004903726279735565)),(to_sfixed_a(-0.0010960008949041367)),(to_sfixed_a(0.0022725139278918505)),(to_sfixed_a(0.0030715905595570803)),(to_sfixed_a(-1.0196355106018018e-05)),(to_sfixed_a(-9.369764302391559e-05)),(to_sfixed_a(0.0007508702110499144)),(to_sfixed_a(0.00023031760065350682)),(to_sfixed_a(-0.004074547905474901)),(to_sfixed_a(0.0018407877068966627)),(to_sfixed_a(0.0005287332460284233)),(to_sfixed_a(-0.0012241110671311617)),(to_sfixed_a(0.0025449004024267197)),(to_sfixed_a(-0.0053474255837500095)),(to_sfixed_a(-0.002519543981179595)),(to_sfixed_a(-0.0002696793817449361)),(to_sfixed_a(0.0006436375551857054)),(to_sfixed_a(-0.001075812499038875)),(to_sfixed_a(0.001619400572963059)),(to_sfixed_a(0.0014805304817855358)),(to_sfixed_a(0.005530699156224728)),(to_sfixed_a(0.0033963292371481657)),(to_sfixed_a(-0.002032396150752902)),(to_sfixed_a(-0.005339320283383131)),(to_sfixed_a(0.00249605905264616)),(to_sfixed_a(-0.00240531750023365)),(to_sfixed_a(-0.003033530432730913)));

    constant weight_n1_107 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.011954093351960182)),(to_sfixed_a(-4.178288236289518e-06)),(to_sfixed_a(-4.3217693018959835e-05)),(to_sfixed_a(-2.0036716250615427e-06)),(to_sfixed_a(5.1120397984050214e-05)),(to_sfixed_a(-1.386995063512586e-05)),(to_sfixed_a(3.2546522561460733e-05)),(to_sfixed_a(-2.5746592655195855e-05)),(to_sfixed_a(5.9125974075868726e-05)),(to_sfixed_a(4.2108869820367545e-05)),(to_sfixed_a(5.638194693347032e-07)),(to_sfixed_a(5.055367364548147e-05)),(to_sfixed_a(1.569491359987296e-05)),(to_sfixed_a(7.79920446802862e-05)),(to_sfixed_a(-5.763532044511521e-06)),(to_sfixed_a(1.7440593182982411e-06)),(to_sfixed_a(-1.7687380022834986e-05)),(to_sfixed_a(-3.7690158478653757e-06)),(to_sfixed_a(-4.355476994533092e-05)),(to_sfixed_a(-1.053516007232247e-05)),(to_sfixed_a(4.797924339072779e-05)),(to_sfixed_a(-1.1074799886046094e-06)),(to_sfixed_a(3.6658857425209135e-05)),(to_sfixed_a(2.342822335776873e-05)),(to_sfixed_a(2.183559990953654e-05)),(to_sfixed_a(-9.74545309873065e-06)),(to_sfixed_a(4.301106309867464e-05)),(to_sfixed_a(-6.84510450810194e-05)),(to_sfixed_a(-3.0000968763488345e-05)),(to_sfixed_a(-8.470425382256508e-05)),(to_sfixed_a(2.816604137478862e-05)),(to_sfixed_a(4.884830195805989e-05)),(to_sfixed_a(3.793146106545464e-06)),(to_sfixed_a(-2.2750555217498913e-05)),(to_sfixed_a(-2.6399035050417297e-05)),(to_sfixed_a(-9.19174199225381e-05)),(to_sfixed_a(-5.202354441280477e-05)),(to_sfixed_a(5.256627264316194e-05)));

    constant weight_n1_108 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.14963999390602112)),(to_sfixed_a(0.010941983200609684)),(to_sfixed_a(-0.008417832665145397)),(to_sfixed_a(0.07012486457824707)),(to_sfixed_a(0.02630290761590004)),(to_sfixed_a(0.0907537043094635)),(to_sfixed_a(-0.07667878270149231)),(to_sfixed_a(-0.04960418492555618)),(to_sfixed_a(0.014535712078213692)),(to_sfixed_a(-0.002635542768985033)),(to_sfixed_a(0.0359133705496788)),(to_sfixed_a(0.017604544758796692)),(to_sfixed_a(0.05771724134683609)),(to_sfixed_a(-0.019180288538336754)),(to_sfixed_a(-0.02679518237709999)),(to_sfixed_a(-0.08348783105611801)),(to_sfixed_a(0.004936676472425461)),(to_sfixed_a(-0.059659507125616074)),(to_sfixed_a(-0.027272524312138557)),(to_sfixed_a(-0.05317468196153641)),(to_sfixed_a(0.004874726757407188)),(to_sfixed_a(-0.060660623013973236)),(to_sfixed_a(0.006205914542078972)),(to_sfixed_a(0.010354837402701378)),(to_sfixed_a(0.028545530512928963)),(to_sfixed_a(-0.035910867154598236)),(to_sfixed_a(-0.04064109921455383)),(to_sfixed_a(0.037247758358716965)),(to_sfixed_a(0.009951299987733364)),(to_sfixed_a(0.11932899802923203)),(to_sfixed_a(0.010537725873291492)),(to_sfixed_a(0.006248867139220238)),(to_sfixed_a(-0.039350394159555435)),(to_sfixed_a(-0.019773749634623528)),(to_sfixed_a(0.013426903635263443)),(to_sfixed_a(0.02258153446018696)),(to_sfixed_a(-0.04848648980259895)),(to_sfixed_a(-0.006559513974934816)));

    constant weight_n1_109 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.3624887764453888)),(to_sfixed_a(0.048603687435388565)),(to_sfixed_a(-0.027156978845596313)),(to_sfixed_a(0.023873794823884964)),(to_sfixed_a(-0.011703195050358772)),(to_sfixed_a(-0.022846132516860962)),(to_sfixed_a(-0.004311526194214821)),(to_sfixed_a(-0.05593051761388779)),(to_sfixed_a(-0.014039479196071625)),(to_sfixed_a(0.11050569266080856)),(to_sfixed_a(-0.01662474311888218)),(to_sfixed_a(-0.11453390121459961)),(to_sfixed_a(0.11679467558860779)),(to_sfixed_a(-0.008506887592375278)),(to_sfixed_a(-0.16048268973827362)),(to_sfixed_a(-0.010287754237651825)),(to_sfixed_a(-0.06956516951322556)),(to_sfixed_a(0.106749027967453)),(to_sfixed_a(0.021576764062047005)),(to_sfixed_a(-0.2805052399635315)),(to_sfixed_a(-0.043455369770526886)),(to_sfixed_a(-0.04153444990515709)),(to_sfixed_a(0.10825547575950623)),(to_sfixed_a(0.01443424541503191)),(to_sfixed_a(0.20309914648532867)),(to_sfixed_a(-0.26528531312942505)),(to_sfixed_a(-0.04942312091588974)),(to_sfixed_a(-0.02440609596669674)),(to_sfixed_a(0.008368585258722305)),(to_sfixed_a(0.14910025894641876)),(to_sfixed_a(-0.08228755742311478)),(to_sfixed_a(0.09205524623394012)),(to_sfixed_a(0.21698226034641266)),(to_sfixed_a(0.16226856410503387)),(to_sfixed_a(-0.009216410107910633)),(to_sfixed_a(-0.33829042315483093)),(to_sfixed_a(0.14449506998062134)),(to_sfixed_a(0.025808576494455338)));

    constant weight_n1_110 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.03243264928460121)),(to_sfixed_a(4.841412737732753e-05)),(to_sfixed_a(-4.4326490751700476e-05)),(to_sfixed_a(2.3689872250542976e-05)),(to_sfixed_a(-1.7298461898462847e-05)),(to_sfixed_a(-4.473303124541417e-05)),(to_sfixed_a(1.8289378203917295e-05)),(to_sfixed_a(-3.541063779266551e-05)),(to_sfixed_a(-3.015018046426121e-05)),(to_sfixed_a(4.110737063456327e-05)),(to_sfixed_a(-1.6267576938844286e-05)),(to_sfixed_a(-5.243481427896768e-05)),(to_sfixed_a(3.4109409170923755e-05)),(to_sfixed_a(-4.675998570746742e-05)),(to_sfixed_a(6.519744056276977e-05)),(to_sfixed_a(1.6118798157549463e-05)),(to_sfixed_a(-6.34523166809231e-05)),(to_sfixed_a(2.184565892093815e-05)),(to_sfixed_a(-6.942728941794485e-05)),(to_sfixed_a(-3.640702925622463e-05)),(to_sfixed_a(-1.17611707537435e-05)),(to_sfixed_a(5.2537168812705204e-05)),(to_sfixed_a(9.80917684501037e-05)),(to_sfixed_a(1.4872075553284958e-05)),(to_sfixed_a(-1.2545709978439845e-05)),(to_sfixed_a(7.79413130658213e-06)),(to_sfixed_a(-1.5395922673633322e-05)),(to_sfixed_a(-5.3933548770146444e-05)),(to_sfixed_a(1.0089587476613815e-06)),(to_sfixed_a(1.5745305063319393e-05)),(to_sfixed_a(1.7823618691181764e-05)),(to_sfixed_a(-9.769250027602538e-06)),(to_sfixed_a(1.118171257985523e-05)),(to_sfixed_a(5.7213273976230994e-05)),(to_sfixed_a(3.477439531707205e-05)),(to_sfixed_a(4.039725172333419e-05)),(to_sfixed_a(2.4836845113895833e-05)),(to_sfixed_a(-1.1869853551615961e-05)));

    constant weight_n1_111 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.418648362159729)),(to_sfixed_a(-0.15873441100120544)),(to_sfixed_a(-0.102798692882061)),(to_sfixed_a(0.08782977610826492)),(to_sfixed_a(0.026807596907019615)),(to_sfixed_a(-0.08232899755239487)),(to_sfixed_a(0.09062501788139343)),(to_sfixed_a(-0.029563169926404953)),(to_sfixed_a(-0.07256454229354858)),(to_sfixed_a(-0.12849026918411255)),(to_sfixed_a(-0.012077338993549347)),(to_sfixed_a(0.07404050976037979)),(to_sfixed_a(-0.1107272133231163)),(to_sfixed_a(0.05516746640205383)),(to_sfixed_a(0.04740672931075096)),(to_sfixed_a(0.11933908611536026)),(to_sfixed_a(0.007086302153766155)),(to_sfixed_a(0.13690292835235596)),(to_sfixed_a(0.0013900600606575608)),(to_sfixed_a(0.0009578015888109803)),(to_sfixed_a(-0.15517181158065796)),(to_sfixed_a(-0.09407903254032135)),(to_sfixed_a(-0.07303530722856522)),(to_sfixed_a(-0.01134348101913929)),(to_sfixed_a(-0.07962729781866074)),(to_sfixed_a(0.031726427376270294)),(to_sfixed_a(0.030190398916602135)),(to_sfixed_a(0.08287981152534485)),(to_sfixed_a(0.00969650223851204)),(to_sfixed_a(0.06355025619268417)),(to_sfixed_a(0.028021786361932755)),(to_sfixed_a(0.12423817813396454)),(to_sfixed_a(0.19439338147640228)),(to_sfixed_a(-0.023701561614871025)),(to_sfixed_a(-0.03527094051241875)),(to_sfixed_a(-0.11112191528081894)),(to_sfixed_a(-0.1023220494389534)),(to_sfixed_a(-0.06196537986397743)));

    constant weight_n1_112 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.10766401886940002)),(to_sfixed_a(1.7308018868789077e-05)),(to_sfixed_a(-3.111406840616837e-05)),(to_sfixed_a(-2.056586708931718e-05)),(to_sfixed_a(2.887913433369249e-05)),(to_sfixed_a(-1.4960925909690559e-05)),(to_sfixed_a(1.8286475551576586e-06)),(to_sfixed_a(8.48401032271795e-06)),(to_sfixed_a(-8.94563527253922e-06)),(to_sfixed_a(6.111380935180932e-05)),(to_sfixed_a(2.8325281164143234e-05)),(to_sfixed_a(-6.361434498103335e-05)),(to_sfixed_a(3.5855151509167627e-05)),(to_sfixed_a(9.254626638721675e-05)),(to_sfixed_a(3.3619755868130596e-06)),(to_sfixed_a(2.01248076336924e-05)),(to_sfixed_a(6.589294935110956e-05)),(to_sfixed_a(2.5605611881474033e-05)),(to_sfixed_a(-4.915866156807169e-05)),(to_sfixed_a(-2.852821410215256e-07)),(to_sfixed_a(-1.078150307876058e-05)),(to_sfixed_a(-2.5243318305001594e-05)),(to_sfixed_a(-6.778033275622874e-05)),(to_sfixed_a(4.828982491744682e-05)),(to_sfixed_a(-4.542675014818087e-05)),(to_sfixed_a(7.53670246922411e-06)),(to_sfixed_a(-1.5787736629135907e-05)),(to_sfixed_a(-5.339542622095905e-05)),(to_sfixed_a(-8.268515375675634e-05)),(to_sfixed_a(0.00011388859275029972)),(to_sfixed_a(3.5882949305232614e-05)),(to_sfixed_a(-4.7853282012511045e-05)),(to_sfixed_a(-9.070067608263344e-05)),(to_sfixed_a(-1.0286911674484145e-05)),(to_sfixed_a(1.06968700492871e-05)),(to_sfixed_a(1.1121870556962676e-05)),(to_sfixed_a(-1.7134971130872145e-05)),(to_sfixed_a(5.0151262257713825e-05)));

    constant weight_n1_113 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.056508615612983704)),(to_sfixed_a(5.405093816079898e-06)),(to_sfixed_a(7.602135610795813e-06)),(to_sfixed_a(2.6887237254413776e-06)),(to_sfixed_a(-5.208828497416107e-06)),(to_sfixed_a(4.9213886086363345e-05)),(to_sfixed_a(-3.913186810677871e-05)),(to_sfixed_a(4.2343224777141586e-05)),(to_sfixed_a(-3.2042607926996425e-05)),(to_sfixed_a(1.3311143902683398e-06)),(to_sfixed_a(-1.8875196474255063e-05)),(to_sfixed_a(4.625585279427469e-05)),(to_sfixed_a(-1.3560559636971448e-05)),(to_sfixed_a(-9.80285676632775e-06)),(to_sfixed_a(2.8000738893751986e-05)),(to_sfixed_a(-8.47030823933892e-05)),(to_sfixed_a(4.745861951960251e-05)),(to_sfixed_a(-2.1324785848264582e-05)),(to_sfixed_a(-8.227872604038566e-05)),(to_sfixed_a(-2.3642141968593933e-05)),(to_sfixed_a(-6.107515946496278e-05)),(to_sfixed_a(1.638566936890129e-05)),(to_sfixed_a(3.65719897672534e-05)),(to_sfixed_a(3.3732725569279864e-05)),(to_sfixed_a(-1.5669551430619322e-05)),(to_sfixed_a(7.069518687785603e-06)),(to_sfixed_a(2.487619440216804e-06)),(to_sfixed_a(-1.3118720971760922e-06)),(to_sfixed_a(-3.4689324820647016e-05)),(to_sfixed_a(-5.163123205420561e-06)),(to_sfixed_a(-5.875769420526922e-05)),(to_sfixed_a(-5.966612297925167e-05)),(to_sfixed_a(2.176646921725478e-05)),(to_sfixed_a(-3.7608955608448014e-05)),(to_sfixed_a(9.25434724194929e-05)),(to_sfixed_a(-4.380469545139931e-05)),(to_sfixed_a(-6.816750101279467e-05)),(to_sfixed_a(8.665405175634078e-07)));

    constant weight_n1_114 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.33469027280807495)),(to_sfixed_a(0.0017114310758188367)),(to_sfixed_a(0.031418513506650925)),(to_sfixed_a(-0.03790511190891266)),(to_sfixed_a(-0.06650892645120621)),(to_sfixed_a(-0.0007063924567773938)),(to_sfixed_a(-0.009510669857263565)),(to_sfixed_a(-0.02092282846570015)),(to_sfixed_a(-0.06825421005487442)),(to_sfixed_a(-0.04759868234395981)),(to_sfixed_a(-0.02880851738154888)),(to_sfixed_a(-0.018138794228434563)),(to_sfixed_a(-0.12121125310659409)),(to_sfixed_a(0.024093197658658028)),(to_sfixed_a(0.013785992749035358)),(to_sfixed_a(-0.033787161111831665)),(to_sfixed_a(-0.051566366106271744)),(to_sfixed_a(-0.07756486535072327)),(to_sfixed_a(-0.05897410959005356)),(to_sfixed_a(0.019816812127828598)),(to_sfixed_a(-0.12441115081310272)),(to_sfixed_a(-0.058433886617422104)),(to_sfixed_a(-0.005087866447865963)),(to_sfixed_a(-0.0998155027627945)),(to_sfixed_a(-0.06055902689695358)),(to_sfixed_a(0.07923920452594757)),(to_sfixed_a(-0.07572480291128159)),(to_sfixed_a(0.04178917035460472)),(to_sfixed_a(-0.06818437576293945)),(to_sfixed_a(-0.06991156935691833)),(to_sfixed_a(0.015669576823711395)),(to_sfixed_a(0.0731709897518158)),(to_sfixed_a(0.002752767177298665)),(to_sfixed_a(-0.028482330963015556)),(to_sfixed_a(0.08613571524620056)),(to_sfixed_a(0.05062182992696762)),(to_sfixed_a(-0.10289423167705536)),(to_sfixed_a(0.032398466020822525)));

    constant weight_n1_115 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.10805870592594147)),(to_sfixed_a(0.030872300267219543)),(to_sfixed_a(0.032097816467285156)),(to_sfixed_a(0.012663248926401138)),(to_sfixed_a(0.0014462820254266262)),(to_sfixed_a(-0.01290671993046999)),(to_sfixed_a(0.03267591446638107)),(to_sfixed_a(0.004814714193344116)),(to_sfixed_a(-0.06302531808614731)),(to_sfixed_a(-0.005626995116472244)),(to_sfixed_a(0.09392733871936798)),(to_sfixed_a(-0.07769137620925903)),(to_sfixed_a(0.012501257471740246)),(to_sfixed_a(0.01038010511547327)),(to_sfixed_a(0.007483627647161484)),(to_sfixed_a(-0.04195577651262283)),(to_sfixed_a(-0.014299043454229832)),(to_sfixed_a(-0.014864935539662838)),(to_sfixed_a(0.05754738673567772)),(to_sfixed_a(-0.035125453025102615)),(to_sfixed_a(0.041212521493434906)),(to_sfixed_a(0.08110246807336807)),(to_sfixed_a(0.015130399726331234)),(to_sfixed_a(-0.028025353327393532)),(to_sfixed_a(-0.023316241800785065)),(to_sfixed_a(0.042817600071430206)),(to_sfixed_a(0.028585277497768402)),(to_sfixed_a(-0.011040437035262585)),(to_sfixed_a(0.019544964656233788)),(to_sfixed_a(0.020840810611844063)),(to_sfixed_a(-0.00808064453303814)),(to_sfixed_a(0.023579584434628487)),(to_sfixed_a(0.061009787023067474)),(to_sfixed_a(-0.012359168380498886)),(to_sfixed_a(0.07574861496686935)),(to_sfixed_a(-0.012823900207877159)),(to_sfixed_a(0.07332813739776611)),(to_sfixed_a(0.03757338970899582)));

    constant weight_n1_116 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.28173378109931946)),(to_sfixed_a(0.008770052343606949)),(to_sfixed_a(-0.01794291101396084)),(to_sfixed_a(-0.006126715801656246)),(to_sfixed_a(-0.020857417955994606)),(to_sfixed_a(0.025559764355421066)),(to_sfixed_a(0.015017210505902767)),(to_sfixed_a(-0.02111680991947651)),(to_sfixed_a(-0.009878628887236118)),(to_sfixed_a(-0.00931769423186779)),(to_sfixed_a(-0.012448769062757492)),(to_sfixed_a(-0.006867759861052036)),(to_sfixed_a(-0.004257471766322851)),(to_sfixed_a(-0.00046621516230516136)),(to_sfixed_a(-0.014257618226110935)),(to_sfixed_a(-0.0001696329127298668)),(to_sfixed_a(-0.0027965400367975235)),(to_sfixed_a(0.0009080010931938887)),(to_sfixed_a(0.007155527826398611)),(to_sfixed_a(-0.009245150722563267)),(to_sfixed_a(0.002799215028062463)),(to_sfixed_a(0.0026150071062147617)),(to_sfixed_a(-0.015404253266751766)),(to_sfixed_a(-0.005935049615800381)),(to_sfixed_a(-0.0005778252962045372)),(to_sfixed_a(0.002936406061053276)),(to_sfixed_a(0.003315393114462495)),(to_sfixed_a(-0.016278723254799843)),(to_sfixed_a(-0.02691805362701416)),(to_sfixed_a(-0.04772647097706795)),(to_sfixed_a(-0.004761512391269207)),(to_sfixed_a(-0.023821616545319557)),(to_sfixed_a(0.010203633457422256)),(to_sfixed_a(0.005878116935491562)),(to_sfixed_a(0.017435165122151375)),(to_sfixed_a(0.016265809535980225)),(to_sfixed_a(0.010484137572348118)),(to_sfixed_a(-0.008984025567770004)));

    constant weight_n1_117 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.009955125860869884)),(to_sfixed_a(-3.912572719855234e-05)),(to_sfixed_a(-2.8408985599526204e-05)),(to_sfixed_a(4.049644849146716e-05)),(to_sfixed_a(-9.143608622252941e-06)),(to_sfixed_a(3.885009573423304e-05)),(to_sfixed_a(4.273092054063454e-05)),(to_sfixed_a(7.973274591677182e-07)),(to_sfixed_a(8.887542207958177e-06)),(to_sfixed_a(7.839119643904269e-05)),(to_sfixed_a(-4.2172967368969694e-05)),(to_sfixed_a(2.573104211478494e-06)),(to_sfixed_a(-8.854800398694351e-06)),(to_sfixed_a(-4.036831887788139e-05)),(to_sfixed_a(-2.490179758751765e-05)),(to_sfixed_a(-2.830437006196007e-05)),(to_sfixed_a(2.9585642550955527e-05)),(to_sfixed_a(2.8597038181032985e-05)),(to_sfixed_a(-7.775060112180654e-06)),(to_sfixed_a(-4.6730398025829345e-05)),(to_sfixed_a(-5.8044595789397135e-05)),(to_sfixed_a(-5.037297887611203e-05)),(to_sfixed_a(-5.507988316821866e-05)),(to_sfixed_a(-1.9436745787970722e-05)),(to_sfixed_a(7.302882295334712e-05)),(to_sfixed_a(-1.962648411790724e-06)),(to_sfixed_a(-2.20800702663837e-05)),(to_sfixed_a(2.2447533410741016e-05)),(to_sfixed_a(-8.465816790703684e-05)),(to_sfixed_a(8.324659575009719e-05)),(to_sfixed_a(2.9505647489713738e-06)),(to_sfixed_a(2.5269559046137147e-05)),(to_sfixed_a(1.7956159354071133e-05)),(to_sfixed_a(-5.1865290515706874e-06)),(to_sfixed_a(7.06353530404158e-05)),(to_sfixed_a(-3.81936042685993e-05)),(to_sfixed_a(0.00011288648238405585)),(to_sfixed_a(-5.819256330141798e-05)));

    constant weight_n1_118 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.08028661459684372)),(to_sfixed_a(-0.039858292788267136)),(to_sfixed_a(0.01130594965070486)),(to_sfixed_a(0.002490229904651642)),(to_sfixed_a(-0.06057499349117279)),(to_sfixed_a(0.0048920470289886)),(to_sfixed_a(0.01994903013110161)),(to_sfixed_a(-0.055675629526376724)),(to_sfixed_a(-0.09073329716920853)),(to_sfixed_a(-0.0012340734247118235)),(to_sfixed_a(0.005831305868923664)),(to_sfixed_a(-0.042519837617874146)),(to_sfixed_a(-0.01940418966114521)),(to_sfixed_a(0.005294048227369785)),(to_sfixed_a(0.026975875720381737)),(to_sfixed_a(0.037452053278684616)),(to_sfixed_a(-0.04418900981545448)),(to_sfixed_a(0.1266031414270401)),(to_sfixed_a(-0.05934664234519005)),(to_sfixed_a(0.0762426033616066)),(to_sfixed_a(-0.05463737994432449)),(to_sfixed_a(-0.08413192629814148)),(to_sfixed_a(-0.050957802683115005)),(to_sfixed_a(0.010075910948216915)),(to_sfixed_a(0.06557325273752213)),(to_sfixed_a(0.08318259567022324)),(to_sfixed_a(-0.026315007358789444)),(to_sfixed_a(0.0866212472319603)),(to_sfixed_a(0.011994756758213043)),(to_sfixed_a(0.02052280865609646)),(to_sfixed_a(0.0011631682282313704)),(to_sfixed_a(0.03064299188554287)),(to_sfixed_a(-0.01996016316115856)),(to_sfixed_a(-0.014140068553388119)),(to_sfixed_a(0.048996761441230774)),(to_sfixed_a(0.12079425156116486)),(to_sfixed_a(0.004875475540757179)),(to_sfixed_a(-0.07210516929626465)));

    constant weight_n1_119 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.028810158371925354)),(to_sfixed_a(7.828422894817777e-06)),(to_sfixed_a(7.592173460579943e-06)),(to_sfixed_a(5.735917511628941e-05)),(to_sfixed_a(-4.7077723138500005e-05)),(to_sfixed_a(2.7506252081366256e-05)),(to_sfixed_a(2.216869870608207e-05)),(to_sfixed_a(-3.575503797037527e-05)),(to_sfixed_a(-1.081796654034406e-05)),(to_sfixed_a(8.603838978160638e-06)),(to_sfixed_a(-1.9364404579391703e-05)),(to_sfixed_a(-4.997290307073854e-05)),(to_sfixed_a(-4.632326090359129e-05)),(to_sfixed_a(3.981667759944685e-06)),(to_sfixed_a(2.1332185497158207e-05)),(to_sfixed_a(2.2244947103899904e-05)),(to_sfixed_a(-9.01875637282501e-07)),(to_sfixed_a(-1.0614444363454822e-05)),(to_sfixed_a(-3.5113993362756446e-05)),(to_sfixed_a(-5.256630902295001e-05)),(to_sfixed_a(-1.5326721040764824e-05)),(to_sfixed_a(2.3779992261552252e-05)),(to_sfixed_a(1.0724986168497708e-05)),(to_sfixed_a(2.1913609089097008e-05)),(to_sfixed_a(6.288835720624775e-05)),(to_sfixed_a(-8.5256906459108e-05)),(to_sfixed_a(-6.697799835819751e-05)),(to_sfixed_a(7.143841503420845e-05)),(to_sfixed_a(-2.5549543352099136e-05)),(to_sfixed_a(-4.926792826154269e-06)),(to_sfixed_a(-3.514010313665494e-05)),(to_sfixed_a(2.5730905690579675e-05)),(to_sfixed_a(-2.2611500753555447e-05)),(to_sfixed_a(8.901673027139623e-06)),(to_sfixed_a(-3.210398062947206e-05)),(to_sfixed_a(-4.882018765783869e-05)),(to_sfixed_a(-1.4792749425396323e-05)),(to_sfixed_a(-3.9452745113521814e-05)));

    constant weight_n1_120 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.15009868144989014)),(to_sfixed_a(2.642917024786584e-05)),(to_sfixed_a(2.9652966986759566e-05)),(to_sfixed_a(-9.598590622772463e-06)),(to_sfixed_a(-1.599383176653646e-05)),(to_sfixed_a(4.520822130871238e-06)),(to_sfixed_a(3.165595990139991e-05)),(to_sfixed_a(9.890169167192653e-06)),(to_sfixed_a(-3.117560481769033e-05)),(to_sfixed_a(-1.1789695236075204e-05)),(to_sfixed_a(2.6701391107053496e-05)),(to_sfixed_a(1.7781565475161187e-05)),(to_sfixed_a(6.856311665615067e-05)),(to_sfixed_a(5.947264435235411e-05)),(to_sfixed_a(2.6938396331388503e-05)),(to_sfixed_a(-5.7338475016877055e-05)),(to_sfixed_a(-1.4239408301364165e-05)),(to_sfixed_a(-8.484347745252308e-06)),(to_sfixed_a(2.374721589148976e-05)),(to_sfixed_a(9.535087883705273e-06)),(to_sfixed_a(-4.4607782911043614e-05)),(to_sfixed_a(-5.518754187505692e-05)),(to_sfixed_a(1.0129660040547606e-05)),(to_sfixed_a(-0.00014579670096281916)),(to_sfixed_a(-1.7850627045845613e-05)),(to_sfixed_a(-0.00010377240687375888)),(to_sfixed_a(1.1292663657513913e-05)),(to_sfixed_a(6.84588958392851e-05)),(to_sfixed_a(6.0678419686155394e-05)),(to_sfixed_a(8.550152415409684e-06)),(to_sfixed_a(6.1031798395561054e-05)),(to_sfixed_a(3.9479749830206856e-05)),(to_sfixed_a(4.4158459786558524e-05)),(to_sfixed_a(-3.050910891033709e-05)),(to_sfixed_a(4.4762193283531815e-05)),(to_sfixed_a(0.00010376008867751807)),(to_sfixed_a(-3.7557856558123603e-05)),(to_sfixed_a(-9.52945338212885e-05)));

    constant weight_n1_121 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.05272994562983513)),(to_sfixed_a(0.03747056424617767)),(to_sfixed_a(0.02152589149773121)),(to_sfixed_a(-0.03015931509435177)),(to_sfixed_a(0.03915870189666748)),(to_sfixed_a(0.027590693905949593)),(to_sfixed_a(0.004566673655062914)),(to_sfixed_a(0.02282687835395336)),(to_sfixed_a(-0.014094121754169464)),(to_sfixed_a(0.02218201942741871)),(to_sfixed_a(0.055086083710193634)),(to_sfixed_a(0.026865368708968163)),(to_sfixed_a(-0.015008711256086826)),(to_sfixed_a(0.05004388093948364)),(to_sfixed_a(0.009824736975133419)),(to_sfixed_a(-0.008128771558403969)),(to_sfixed_a(-0.009203704074025154)),(to_sfixed_a(-0.015008022077381611)),(to_sfixed_a(-0.042762771248817444)),(to_sfixed_a(0.09351364523172379)),(to_sfixed_a(-0.007924847304821014)),(to_sfixed_a(-0.05778080224990845)),(to_sfixed_a(-0.08885905891656876)),(to_sfixed_a(0.008057544007897377)),(to_sfixed_a(-0.02887369506061077)),(to_sfixed_a(0.025438617914915085)),(to_sfixed_a(0.028529921546578407)),(to_sfixed_a(0.031740639358758926)),(to_sfixed_a(0.012340160086750984)),(to_sfixed_a(-0.021518515422940254)),(to_sfixed_a(0.02590908110141754)),(to_sfixed_a(0.03360016271471977)),(to_sfixed_a(0.054459989070892334)),(to_sfixed_a(-0.006543116644024849)),(to_sfixed_a(0.010950087569653988)),(to_sfixed_a(-0.03929968550801277)),(to_sfixed_a(0.016447048634290695)),(to_sfixed_a(-0.015735439956188202)));

    constant weight_n1_122 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.16695624589920044)),(to_sfixed_a(1.5553567209281027e-05)),(to_sfixed_a(-3.873397872666828e-06)),(to_sfixed_a(-1.6899230104172602e-05)),(to_sfixed_a(-2.9754119168501347e-06)),(to_sfixed_a(-1.8850385458790697e-05)),(to_sfixed_a(1.7332804418401793e-05)),(to_sfixed_a(4.447947139851749e-05)),(to_sfixed_a(-2.28119533858262e-05)),(to_sfixed_a(-4.683709630626254e-05)),(to_sfixed_a(9.522244909021538e-06)),(to_sfixed_a(1.1865831766044721e-05)),(to_sfixed_a(2.803653296723496e-05)),(to_sfixed_a(1.4518279385811184e-05)),(to_sfixed_a(-2.5829240257735364e-05)),(to_sfixed_a(9.969933671527542e-06)),(to_sfixed_a(2.3622562366654165e-05)),(to_sfixed_a(6.417939403036144e-06)),(to_sfixed_a(2.0786423192475922e-05)),(to_sfixed_a(1.3593597941508051e-05)),(to_sfixed_a(9.690455044619739e-05)),(to_sfixed_a(-1.6227564628934488e-05)),(to_sfixed_a(2.3701343252469087e-06)),(to_sfixed_a(3.739784733625129e-05)),(to_sfixed_a(2.6595704184728675e-05)),(to_sfixed_a(-3.627682599471882e-05)),(to_sfixed_a(4.3624262616503984e-05)),(to_sfixed_a(4.5700955524807796e-05)),(to_sfixed_a(5.4384559916798025e-05)),(to_sfixed_a(4.562773392535746e-05)),(to_sfixed_a(-0.0001077213601092808)),(to_sfixed_a(3.143773938063532e-05)),(to_sfixed_a(3.062585528823547e-05)),(to_sfixed_a(-4.56566849607043e-05)),(to_sfixed_a(5.757279268436832e-06)),(to_sfixed_a(-5.304784281179309e-05)),(to_sfixed_a(-5.998702908982523e-05)),(to_sfixed_a(-6.048683280823752e-05)));

    constant weight_n1_123 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.13446144759655)),(to_sfixed_a(-5.644053544529015e-06)),(to_sfixed_a(-3.427603587624617e-05)),(to_sfixed_a(-6.584495622519171e-06)),(to_sfixed_a(2.203407575507299e-06)),(to_sfixed_a(1.0998324796673842e-05)),(to_sfixed_a(-5.582108860835433e-05)),(to_sfixed_a(7.804504275554791e-05)),(to_sfixed_a(-3.3190557587658986e-05)),(to_sfixed_a(-6.979900354053825e-05)),(to_sfixed_a(-0.0001256796094821766)),(to_sfixed_a(4.7306151827797294e-05)),(to_sfixed_a(-2.420806049485691e-05)),(to_sfixed_a(-3.3663025533314794e-05)),(to_sfixed_a(-2.3113896531867795e-05)),(to_sfixed_a(2.397595380898565e-05)),(to_sfixed_a(7.100640686985571e-06)),(to_sfixed_a(7.504619503606591e-08)),(to_sfixed_a(5.3037776524433866e-05)),(to_sfixed_a(7.26672078599222e-06)),(to_sfixed_a(4.7828951210249215e-05)),(to_sfixed_a(-4.872605131822638e-05)),(to_sfixed_a(1.3685244084626902e-06)),(to_sfixed_a(-1.623889329493977e-05)),(to_sfixed_a(5.344083547242917e-05)),(to_sfixed_a(0.00011829080176539719)),(to_sfixed_a(4.4339540181681514e-05)),(to_sfixed_a(6.2796869315207e-05)),(to_sfixed_a(-4.24580393882934e-05)),(to_sfixed_a(0.0001163550914498046)),(to_sfixed_a(9.27782166399993e-05)),(to_sfixed_a(1.4860018382023554e-05)),(to_sfixed_a(5.1290146075189114e-05)),(to_sfixed_a(4.942483428749256e-05)),(to_sfixed_a(4.122790051042102e-05)),(to_sfixed_a(-2.567970113886986e-05)),(to_sfixed_a(4.9491736717754975e-05)),(to_sfixed_a(4.4487296690931544e-05)));

    constant weight_n1_124 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.1343601793050766)),(to_sfixed_a(0.019505146890878677)),(to_sfixed_a(-0.11888498067855835)),(to_sfixed_a(0.05648198351264)),(to_sfixed_a(0.05655874311923981)),(to_sfixed_a(-0.01252006459981203)),(to_sfixed_a(0.15608908236026764)),(to_sfixed_a(0.13456003367900848)),(to_sfixed_a(0.1548534333705902)),(to_sfixed_a(0.049548178911209106)),(to_sfixed_a(0.18564975261688232)),(to_sfixed_a(0.09815704822540283)),(to_sfixed_a(-0.02507610246539116)),(to_sfixed_a(-0.07972061634063721)),(to_sfixed_a(0.02225556969642639)),(to_sfixed_a(0.13844750821590424)),(to_sfixed_a(-0.05659560114145279)),(to_sfixed_a(0.13812567293643951)),(to_sfixed_a(-0.16083720326423645)),(to_sfixed_a(-0.05681103095412254)),(to_sfixed_a(-0.14593657851219177)),(to_sfixed_a(0.0887083187699318)),(to_sfixed_a(0.06821379065513611)),(to_sfixed_a(0.062106773257255554)),(to_sfixed_a(0.09742762893438339)),(to_sfixed_a(0.0833258256316185)),(to_sfixed_a(-0.11828507483005524)),(to_sfixed_a(0.1126294806599617)),(to_sfixed_a(0.1024806946516037)),(to_sfixed_a(0.10292933136224747)),(to_sfixed_a(0.026034919545054436)),(to_sfixed_a(-0.20038637518882751)),(to_sfixed_a(0.08716000616550446)),(to_sfixed_a(-0.11147350072860718)),(to_sfixed_a(0.0474943108856678)),(to_sfixed_a(0.1213710606098175)),(to_sfixed_a(0.006434962153434753)),(to_sfixed_a(0.31865042448043823)));

    constant weight_n1_125 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.055833812803030014)),(to_sfixed_a(-0.010753578506410122)),(to_sfixed_a(-0.0011998343979939818)),(to_sfixed_a(0.008910313248634338)),(to_sfixed_a(0.03475072607398033)),(to_sfixed_a(0.06613340228796005)),(to_sfixed_a(0.018555238842964172)),(to_sfixed_a(0.007034618407487869)),(to_sfixed_a(-0.06490159779787064)),(to_sfixed_a(0.050143685191869736)),(to_sfixed_a(0.0094922399148345)),(to_sfixed_a(0.02714528888463974)),(to_sfixed_a(0.08702730387449265)),(to_sfixed_a(-0.028955379500985146)),(to_sfixed_a(0.0016389053780585527)),(to_sfixed_a(-0.11543481051921844)),(to_sfixed_a(0.01701902598142624)),(to_sfixed_a(0.00015210642595775425)),(to_sfixed_a(0.034269895404577255)),(to_sfixed_a(0.011058501899242401)),(to_sfixed_a(0.030703086405992508)),(to_sfixed_a(0.10034392029047012)),(to_sfixed_a(-0.1022915244102478)),(to_sfixed_a(-0.04888521507382393)),(to_sfixed_a(0.09571424871683121)),(to_sfixed_a(-0.041910819709300995)),(to_sfixed_a(-0.17601227760314941)),(to_sfixed_a(-0.011153008788824081)),(to_sfixed_a(0.009181173518300056)),(to_sfixed_a(-0.16647860407829285)),(to_sfixed_a(0.1268107146024704)),(to_sfixed_a(0.022502921521663666)),(to_sfixed_a(-0.10374213755130768)),(to_sfixed_a(0.1017298698425293)),(to_sfixed_a(0.10032222419977188)),(to_sfixed_a(-0.031619857996702194)),(to_sfixed_a(0.050876740366220474)),(to_sfixed_a(0.14838539063930511)));

    constant weight_n1_126 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.028336836025118828)),(to_sfixed_a(-4.2925483285216615e-05)),(to_sfixed_a(3.644277967396192e-05)),(to_sfixed_a(1.4400979125639424e-05)),(to_sfixed_a(6.47034994472051e-06)),(to_sfixed_a(1.5306857676478103e-05)),(to_sfixed_a(-2.0403081180120353e-06)),(to_sfixed_a(-7.788850780343637e-05)),(to_sfixed_a(-2.2444073692895472e-05)),(to_sfixed_a(-1.258540760318283e-05)),(to_sfixed_a(-1.2290023221339652e-07)),(to_sfixed_a(1.2866246834164485e-05)),(to_sfixed_a(-1.908737249323167e-05)),(to_sfixed_a(-1.3049981134827249e-05)),(to_sfixed_a(-3.0265455279732123e-06)),(to_sfixed_a(1.8111544704879634e-05)),(to_sfixed_a(-2.0114657672820613e-05)),(to_sfixed_a(-2.2358977957992465e-07)),(to_sfixed_a(-9.147642231255304e-06)),(to_sfixed_a(-2.1207713871262968e-05)),(to_sfixed_a(-3.5827823012368754e-05)),(to_sfixed_a(5.6934459280455485e-05)),(to_sfixed_a(-1.4759186342416797e-05)),(to_sfixed_a(9.935821253748145e-06)),(to_sfixed_a(-2.0793002022401197e-06)),(to_sfixed_a(-1.7744223441695794e-05)),(to_sfixed_a(-1.454924131394364e-05)),(to_sfixed_a(1.1839406397484709e-05)),(to_sfixed_a(-0.00012261046504136175)),(to_sfixed_a(3.8252241211012006e-05)),(to_sfixed_a(8.093562428257428e-06)),(to_sfixed_a(-2.678458031368791e-06)),(to_sfixed_a(8.423782855970785e-05)),(to_sfixed_a(3.647633275249973e-05)),(to_sfixed_a(-1.4378366358869243e-05)),(to_sfixed_a(-4.04586608055979e-05)),(to_sfixed_a(-4.634847573470324e-05)),(to_sfixed_a(5.594594040303491e-05)));

    constant weight_n1_127 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.018237117677927017)),(to_sfixed_a(-4.1346720536239445e-05)),(to_sfixed_a(6.490169198514195e-06)),(to_sfixed_a(4.133605398237705e-05)),(to_sfixed_a(4.000411354354583e-05)),(to_sfixed_a(6.414040399249643e-05)),(to_sfixed_a(2.7638989195111208e-05)),(to_sfixed_a(-5.023195626563393e-06)),(to_sfixed_a(5.549343768507242e-06)),(to_sfixed_a(7.877841562731192e-05)),(to_sfixed_a(-2.9447253837133758e-05)),(to_sfixed_a(2.9265562261571176e-05)),(to_sfixed_a(1.868655272119213e-05)),(to_sfixed_a(4.5225464418763295e-05)),(to_sfixed_a(3.998677129857242e-05)),(to_sfixed_a(1.4322244169306941e-05)),(to_sfixed_a(3.8830185076221824e-05)),(to_sfixed_a(3.142200148431584e-05)),(to_sfixed_a(3.486965943011455e-05)),(to_sfixed_a(-7.097291927493643e-06)),(to_sfixed_a(6.00926396145951e-05)),(to_sfixed_a(5.177245839149691e-05)),(to_sfixed_a(-2.258468339277897e-05)),(to_sfixed_a(8.338554471265525e-05)),(to_sfixed_a(2.9074356007185997e-06)),(to_sfixed_a(-1.1947070561291184e-05)),(to_sfixed_a(6.430298526538536e-05)),(to_sfixed_a(-0.00011736017768271267)),(to_sfixed_a(-3.893378743669018e-05)),(to_sfixed_a(-0.00015848909970372915)),(to_sfixed_a(-0.00014110376650933176)),(to_sfixed_a(-2.9687740607187152e-05)),(to_sfixed_a(-2.743398363236338e-05)),(to_sfixed_a(-0.0001277423434657976)),(to_sfixed_a(2.714663787628524e-05)),(to_sfixed_a(3.1746443710289896e-05)),(to_sfixed_a(9.917255738400854e-06)),(to_sfixed_a(-4.4448130211094394e-05)));

    constant weight_n1_128 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.008943295106291771)),(to_sfixed_a(5.248621164355427e-05)),(to_sfixed_a(2.098761615343392e-05)),(to_sfixed_a(-1.6746920664445497e-05)),(to_sfixed_a(-5.3481759096030146e-05)),(to_sfixed_a(-2.059406688204035e-05)),(to_sfixed_a(1.2694986253336538e-05)),(to_sfixed_a(-3.768906753975898e-05)),(to_sfixed_a(1.3305361790116876e-06)),(to_sfixed_a(4.8750189307611436e-05)),(to_sfixed_a(-2.1335712517611682e-05)),(to_sfixed_a(-4.907459515379742e-05)),(to_sfixed_a(1.8894414097303525e-05)),(to_sfixed_a(7.288990309461951e-05)),(to_sfixed_a(-7.277182157849893e-05)),(to_sfixed_a(-3.863453821395524e-05)),(to_sfixed_a(3.9290614950004965e-05)),(to_sfixed_a(-0.00010897943866439164)),(to_sfixed_a(-4.7510235162917525e-05)),(to_sfixed_a(1.331087332800962e-05)),(to_sfixed_a(2.6911024178843945e-05)),(to_sfixed_a(9.837193829298485e-06)),(to_sfixed_a(2.357160883548204e-05)),(to_sfixed_a(-2.0124902221141383e-05)),(to_sfixed_a(-6.805566954426467e-05)),(to_sfixed_a(2.7020787456422113e-05)),(to_sfixed_a(-7.702161383349448e-06)),(to_sfixed_a(1.6187666915357113e-05)),(to_sfixed_a(-2.9595357773359865e-05)),(to_sfixed_a(5.802194573334418e-05)),(to_sfixed_a(-5.9859488828806207e-05)),(to_sfixed_a(-5.018330193706788e-05)),(to_sfixed_a(6.583955109817907e-05)),(to_sfixed_a(-0.0001184591164928861)),(to_sfixed_a(-7.863147038733587e-05)),(to_sfixed_a(-1.1502528650453314e-05)),(to_sfixed_a(1.2894113332606594e-08)),(to_sfixed_a(-1.6646157746436074e-05)));

    constant weight_n1_129 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.03649440035223961)),(to_sfixed_a(-4.283906673663296e-05)),(to_sfixed_a(2.827495882229414e-05)),(to_sfixed_a(-2.341063918720465e-06)),(to_sfixed_a(1.3950786524219438e-05)),(to_sfixed_a(-6.2961539697425906e-06)),(to_sfixed_a(-1.1440564776421525e-05)),(to_sfixed_a(1.4693134289700538e-05)),(to_sfixed_a(7.823733176337555e-05)),(to_sfixed_a(-2.0097515516681597e-05)),(to_sfixed_a(2.1464951714733616e-05)),(to_sfixed_a(2.8891525289509445e-05)),(to_sfixed_a(3.0224422516766936e-05)),(to_sfixed_a(9.748384400154464e-06)),(to_sfixed_a(-3.2553787605138496e-05)),(to_sfixed_a(6.471350934589282e-05)),(to_sfixed_a(-0.00011876912321895361)),(to_sfixed_a(-2.3627420887351036e-05)),(to_sfixed_a(-2.5456980438320898e-05)),(to_sfixed_a(5.67534843867179e-05)),(to_sfixed_a(-2.204428892582655e-05)),(to_sfixed_a(-1.6599049558863044e-05)),(to_sfixed_a(-3.9578109863214195e-05)),(to_sfixed_a(-1.3672352906723972e-05)),(to_sfixed_a(1.9130702639813535e-05)),(to_sfixed_a(7.544254913227633e-05)),(to_sfixed_a(-1.1744726180040743e-05)),(to_sfixed_a(-5.578810305451043e-05)),(to_sfixed_a(-1.819725730456412e-05)),(to_sfixed_a(2.5373265089001507e-05)),(to_sfixed_a(0.00012402467837091535)),(to_sfixed_a(-1.754738696035929e-05)),(to_sfixed_a(-1.6569618310313672e-05)),(to_sfixed_a(1.826463449106086e-05)),(to_sfixed_a(-2.180896080972161e-05)),(to_sfixed_a(1.7288753952016123e-05)),(to_sfixed_a(6.556983134942129e-05)),(to_sfixed_a(6.24188469373621e-05)));

    constant weight_n1_130 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.027752352878451347)),(to_sfixed_a(4.0655271732248366e-05)),(to_sfixed_a(-7.289640052476898e-06)),(to_sfixed_a(-1.6494548617629334e-05)),(to_sfixed_a(-2.4616054361104034e-05)),(to_sfixed_a(-1.0520097021071706e-05)),(to_sfixed_a(-3.0376246286323294e-05)),(to_sfixed_a(2.3740294636809267e-05)),(to_sfixed_a(-5.084735676064156e-05)),(to_sfixed_a(3.440367436269298e-05)),(to_sfixed_a(3.3372016332577914e-05)),(to_sfixed_a(-2.768437479971908e-05)),(to_sfixed_a(3.085489879595116e-05)),(to_sfixed_a(2.9925857234047726e-05)),(to_sfixed_a(4.734755930257961e-05)),(to_sfixed_a(-9.548487469146494e-06)),(to_sfixed_a(3.059059235965833e-05)),(to_sfixed_a(-7.99760346126277e-06)),(to_sfixed_a(-1.6401540051447228e-05)),(to_sfixed_a(-1.5349374734796584e-05)),(to_sfixed_a(2.1473722881637514e-05)),(to_sfixed_a(8.230315870605409e-06)),(to_sfixed_a(3.509762609610334e-05)),(to_sfixed_a(6.060382293071598e-05)),(to_sfixed_a(-2.926067463704385e-05)),(to_sfixed_a(-1.6782499869805179e-06)),(to_sfixed_a(2.2358892238116823e-05)),(to_sfixed_a(-1.2482928468671162e-05)),(to_sfixed_a(5.939043694525026e-05)),(to_sfixed_a(1.9857870938722044e-05)),(to_sfixed_a(4.51013220299501e-05)),(to_sfixed_a(-1.4842005668924685e-07)),(to_sfixed_a(-2.078706893371418e-05)),(to_sfixed_a(6.522842886624858e-05)),(to_sfixed_a(-3.078651207033545e-05)),(to_sfixed_a(5.199812221690081e-05)),(to_sfixed_a(-2.834168481058441e-05)),(to_sfixed_a(5.6731762015260756e-05)));

    constant weight_n1_131 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.02611762098968029)),(to_sfixed_a(-0.019945595413446426)),(to_sfixed_a(0.02237250842154026)),(to_sfixed_a(0.10418523848056793)),(to_sfixed_a(0.013690716587007046)),(to_sfixed_a(0.08843636512756348)),(to_sfixed_a(-0.0669390931725502)),(to_sfixed_a(-0.03366951644420624)),(to_sfixed_a(-0.010053656995296478)),(to_sfixed_a(0.011306509375572205)),(to_sfixed_a(0.02972210943698883)),(to_sfixed_a(0.06545953452587128)),(to_sfixed_a(-0.03944621980190277)),(to_sfixed_a(-0.053841594606637955)),(to_sfixed_a(-0.010481237433850765)),(to_sfixed_a(-0.06840676814317703)),(to_sfixed_a(-0.02007300965487957)),(to_sfixed_a(-0.05051075667142868)),(to_sfixed_a(0.027707746252417564)),(to_sfixed_a(-0.06952237337827682)),(to_sfixed_a(-0.03432672470808029)),(to_sfixed_a(-0.05604211613535881)),(to_sfixed_a(0.017978854477405548)),(to_sfixed_a(0.020382514223456383)),(to_sfixed_a(0.032351791858673096)),(to_sfixed_a(0.026582365855574608)),(to_sfixed_a(-0.0002151855587726459)),(to_sfixed_a(0.06226818636059761)),(to_sfixed_a(-0.06352125108242035)),(to_sfixed_a(-0.008467601612210274)),(to_sfixed_a(0.013717716559767723)),(to_sfixed_a(0.020186617970466614)),(to_sfixed_a(-0.028377162292599678)),(to_sfixed_a(0.02718493528664112)),(to_sfixed_a(-0.006275986786931753)),(to_sfixed_a(-0.006527319084852934)),(to_sfixed_a(0.02242112159729004)),(to_sfixed_a(0.013748979195952415)));

    constant weight_n1_132 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.09913846105337143)),(to_sfixed_a(0.02163960039615631)),(to_sfixed_a(0.006911656819283962)),(to_sfixed_a(-0.011599992401897907)),(to_sfixed_a(0.0039034411311149597)),(to_sfixed_a(0.06127605214715004)),(to_sfixed_a(0.07554592192173004)),(to_sfixed_a(0.03960753232240677)),(to_sfixed_a(0.046281859278678894)),(to_sfixed_a(-0.03824806958436966)),(to_sfixed_a(-0.04513763636350632)),(to_sfixed_a(-0.020783916115760803)),(to_sfixed_a(-0.14743180572986603)),(to_sfixed_a(0.019497642293572426)),(to_sfixed_a(-0.02606998011469841)),(to_sfixed_a(-0.07970762252807617)),(to_sfixed_a(0.009693681262433529)),(to_sfixed_a(0.009447993710637093)),(to_sfixed_a(-0.06997793167829514)),(to_sfixed_a(0.06596623361110687)),(to_sfixed_a(0.01331548485904932)),(to_sfixed_a(-0.017239058390259743)),(to_sfixed_a(-0.00802986603230238)),(to_sfixed_a(-0.05011705309152603)),(to_sfixed_a(0.016197286546230316)),(to_sfixed_a(0.10176729410886765)),(to_sfixed_a(-0.010601040907204151)),(to_sfixed_a(0.02199786715209484)),(to_sfixed_a(-0.07705617696046829)),(to_sfixed_a(0.031106695532798767)),(to_sfixed_a(-0.08889463543891907)),(to_sfixed_a(0.0329061858355999)),(to_sfixed_a(-0.02610362507402897)),(to_sfixed_a(0.051568977534770966)),(to_sfixed_a(-0.059656526893377304)),(to_sfixed_a(0.023241152986884117)),(to_sfixed_a(0.14121940732002258)),(to_sfixed_a(0.07477789372205734)));

    constant weight_n1_133 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.05763981491327286)),(to_sfixed_a(1.796327887859661e-05)),(to_sfixed_a(-1.1396058653190266e-05)),(to_sfixed_a(-2.3260148736881092e-05)),(to_sfixed_a(-2.5843496587185655e-06)),(to_sfixed_a(-4.3843033381563146e-06)),(to_sfixed_a(6.98991652825498e-06)),(to_sfixed_a(-1.1898609955096617e-05)),(to_sfixed_a(-3.9978935092221946e-05)),(to_sfixed_a(-1.1418032954679802e-05)),(to_sfixed_a(-3.455563637544401e-05)),(to_sfixed_a(-3.577509778551757e-05)),(to_sfixed_a(1.9694914954015985e-05)),(to_sfixed_a(-7.951679208417772e-07)),(to_sfixed_a(-5.590418732026592e-05)),(to_sfixed_a(3.6600264138542116e-05)),(to_sfixed_a(-5.093717481940985e-05)),(to_sfixed_a(1.195144432131201e-05)),(to_sfixed_a(6.3986062741605565e-06)),(to_sfixed_a(-2.676432131920592e-06)),(to_sfixed_a(-5.349885395844467e-05)),(to_sfixed_a(-6.285797553573502e-06)),(to_sfixed_a(-3.7607305785058998e-06)),(to_sfixed_a(1.926454388012644e-05)),(to_sfixed_a(-6.844119980087271e-06)),(to_sfixed_a(4.012829958810471e-05)),(to_sfixed_a(-2.176018460886553e-05)),(to_sfixed_a(-1.2097742683181423e-06)),(to_sfixed_a(-8.708949462743476e-05)),(to_sfixed_a(-1.3625055544252973e-05)),(to_sfixed_a(2.5096439912886126e-06)),(to_sfixed_a(-1.4653030575573212e-06)),(to_sfixed_a(2.1662919607479125e-05)),(to_sfixed_a(-6.820609996793792e-05)),(to_sfixed_a(5.1997001719428226e-05)),(to_sfixed_a(-1.5444171367562376e-05)),(to_sfixed_a(-4.3717165681300685e-05)),(to_sfixed_a(5.698460154235363e-05)));

    constant weight_n1_134 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.02653462253510952)),(to_sfixed_a(2.0016415874124505e-05)),(to_sfixed_a(3.840000135824084e-05)),(to_sfixed_a(-4.086501576239243e-05)),(to_sfixed_a(3.350188126205467e-05)),(to_sfixed_a(-1.4032822036824655e-05)),(to_sfixed_a(-3.9864517020760104e-05)),(to_sfixed_a(-1.517254986538319e-06)),(to_sfixed_a(4.645327408070443e-06)),(to_sfixed_a(-6.677353667328134e-05)),(to_sfixed_a(-7.061439100652933e-05)),(to_sfixed_a(3.8915033655939624e-05)),(to_sfixed_a(1.2836264431825839e-05)),(to_sfixed_a(-4.3674808694049716e-05)),(to_sfixed_a(3.445893889875151e-05)),(to_sfixed_a(-3.045131597900763e-05)),(to_sfixed_a(6.901996130181942e-06)),(to_sfixed_a(7.749635187792592e-06)),(to_sfixed_a(-5.349260754883289e-05)),(to_sfixed_a(2.956126627395861e-05)),(to_sfixed_a(-6.694172043353319e-05)),(to_sfixed_a(1.3170605598133989e-05)),(to_sfixed_a(-1.1712836567312479e-05)),(to_sfixed_a(4.701728539657779e-05)),(to_sfixed_a(-4.0343871660297737e-05)),(to_sfixed_a(-3.083882256760262e-05)),(to_sfixed_a(-5.89858136663679e-05)),(to_sfixed_a(-1.7301379557466134e-05)),(to_sfixed_a(-1.384045299346326e-05)),(to_sfixed_a(-0.00010847557859960943)),(to_sfixed_a(-5.58749388801516e-06)),(to_sfixed_a(3.0299848731374368e-05)),(to_sfixed_a(3.261325036874041e-05)),(to_sfixed_a(6.159894837765023e-05)),(to_sfixed_a(0.00010546355770202354)),(to_sfixed_a(-4.139772954658838e-06)),(to_sfixed_a(-8.731681009521708e-05)),(to_sfixed_a(6.547218799823895e-05)));

    constant weight_n1_135 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.3782559931278229)),(to_sfixed_a(-0.010820984840393066)),(to_sfixed_a(-0.005481692496687174)),(to_sfixed_a(-0.07555495947599411)),(to_sfixed_a(-0.051212094724178314)),(to_sfixed_a(-0.020018320530653)),(to_sfixed_a(-0.3670213520526886)),(to_sfixed_a(0.04551337659358978)),(to_sfixed_a(0.1252230405807495)),(to_sfixed_a(-0.370170533657074)),(to_sfixed_a(0.09759804606437683)),(to_sfixed_a(-0.06571047753095627)),(to_sfixed_a(0.05112423002719879)),(to_sfixed_a(-0.028090182691812515)),(to_sfixed_a(-0.03533392772078514)),(to_sfixed_a(0.023097746074199677)),(to_sfixed_a(0.23352012038230896)),(to_sfixed_a(0.2322947084903717)),(to_sfixed_a(-0.007653191685676575)),(to_sfixed_a(0.17505903542041779)),(to_sfixed_a(0.00241011637263)),(to_sfixed_a(0.0116199916228652)),(to_sfixed_a(0.2652675211429596)),(to_sfixed_a(0.028026597574353218)),(to_sfixed_a(-0.10341337323188782)),(to_sfixed_a(0.1721828132867813)),(to_sfixed_a(-0.07946952432394028)),(to_sfixed_a(-0.017386525869369507)),(to_sfixed_a(0.10593977570533752)),(to_sfixed_a(-0.011040672659873962)),(to_sfixed_a(-0.07491234689950943)),(to_sfixed_a(0.059513937681913376)),(to_sfixed_a(0.009161075577139854)),(to_sfixed_a(0.07924922555685043)),(to_sfixed_a(0.05515085160732269)),(to_sfixed_a(-0.22041477262973785)),(to_sfixed_a(0.07221709191799164)),(to_sfixed_a(-0.015877334401011467)));

    constant weight_n1_136 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.12008633464574814)),(to_sfixed_a(0.025132622569799423)),(to_sfixed_a(-0.006992674432694912)),(to_sfixed_a(-0.024155838415026665)),(to_sfixed_a(-0.002509573008865118)),(to_sfixed_a(-0.007620303425937891)),(to_sfixed_a(-0.039724450558423996)),(to_sfixed_a(-0.028476212173700333)),(to_sfixed_a(0.1086641401052475)),(to_sfixed_a(-0.0707964226603508)),(to_sfixed_a(-0.07777378708124161)),(to_sfixed_a(-0.009234311990439892)),(to_sfixed_a(0.002283670473843813)),(to_sfixed_a(-0.007543953601270914)),(to_sfixed_a(-0.0332268550992012)),(to_sfixed_a(0.056257233023643494)),(to_sfixed_a(0.023847512900829315)),(to_sfixed_a(0.053522586822509766)),(to_sfixed_a(-0.024110540747642517)),(to_sfixed_a(0.032449886202812195)),(to_sfixed_a(0.043468721210956573)),(to_sfixed_a(0.041819892823696136)),(to_sfixed_a(0.07001552730798721)),(to_sfixed_a(0.015792502090334892)),(to_sfixed_a(-0.04430507495999336)),(to_sfixed_a(-0.021146655082702637)),(to_sfixed_a(-0.05156116187572479)),(to_sfixed_a(0.11807307600975037)),(to_sfixed_a(0.004725482780486345)),(to_sfixed_a(-0.09089621901512146)),(to_sfixed_a(0.07069490104913712)),(to_sfixed_a(0.1188773587346077)),(to_sfixed_a(0.0032505756244063377)),(to_sfixed_a(-0.05983958765864372)),(to_sfixed_a(0.032098352909088135)),(to_sfixed_a(-0.0319388248026371)),(to_sfixed_a(0.027095047757029533)),(to_sfixed_a(0.09754573553800583)));

    constant weight_n1_137 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.013911872170865536)),(to_sfixed_a(-1.794328636606224e-05)),(to_sfixed_a(5.318855255609378e-05)),(to_sfixed_a(-3.724473208421841e-05)),(to_sfixed_a(4.2189338273601606e-05)),(to_sfixed_a(8.437311407760717e-06)),(to_sfixed_a(2.3779131879564375e-05)),(to_sfixed_a(2.1711526642320678e-05)),(to_sfixed_a(6.222918273124378e-06)),(to_sfixed_a(1.999001506192144e-05)),(to_sfixed_a(9.017379852593876e-06)),(to_sfixed_a(4.072738374816254e-05)),(to_sfixed_a(-3.6681860365206376e-05)),(to_sfixed_a(-3.125567309325561e-05)),(to_sfixed_a(3.658147988971905e-06)),(to_sfixed_a(-3.915968773071654e-05)),(to_sfixed_a(-8.8236356532434e-06)),(to_sfixed_a(-4.871643795922864e-06)),(to_sfixed_a(9.535115532344207e-05)),(to_sfixed_a(-8.367337431991473e-05)),(to_sfixed_a(6.049329022062011e-05)),(to_sfixed_a(4.733021796710091e-06)),(to_sfixed_a(-3.8524740375578403e-05)),(to_sfixed_a(7.045813254080713e-05)),(to_sfixed_a(2.6896261260844767e-05)),(to_sfixed_a(-3.780272891162895e-05)),(to_sfixed_a(4.633402932086028e-05)),(to_sfixed_a(5.636197965941392e-05)),(to_sfixed_a(5.821287049911916e-05)),(to_sfixed_a(-3.7311488995328546e-05)),(to_sfixed_a(-2.0487237634370103e-05)),(to_sfixed_a(5.0653274229262024e-05)),(to_sfixed_a(5.957090252195485e-05)),(to_sfixed_a(-5.646671706927009e-05)),(to_sfixed_a(-5.5387721658917144e-05)),(to_sfixed_a(1.5763456758577377e-05)),(to_sfixed_a(1.3846270121575799e-05)),(to_sfixed_a(-3.8119109376566485e-05)));

    constant weight_n1_138 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.013911333866417408)),(to_sfixed_a(2.544147355365567e-05)),(to_sfixed_a(1.8993589037563652e-05)),(to_sfixed_a(1.975706618395634e-05)),(to_sfixed_a(5.695049367204774e-06)),(to_sfixed_a(-1.8632783849170664e-06)),(to_sfixed_a(3.741715045180172e-05)),(to_sfixed_a(2.585365109553095e-06)),(to_sfixed_a(5.003275873605162e-06)),(to_sfixed_a(1.292770502914209e-05)),(to_sfixed_a(-1.677745058259461e-05)),(to_sfixed_a(-5.0691051001194865e-05)),(to_sfixed_a(-1.7161712094093673e-05)),(to_sfixed_a(1.250627337867627e-05)),(to_sfixed_a(1.983188667509239e-05)),(to_sfixed_a(-3.451916199992411e-05)),(to_sfixed_a(1.6996769772958942e-05)),(to_sfixed_a(5.127242184244096e-05)),(to_sfixed_a(-2.631639836181421e-05)),(to_sfixed_a(3.659033609437756e-05)),(to_sfixed_a(1.8101331079378724e-05)),(to_sfixed_a(-3.8343147025443614e-05)),(to_sfixed_a(-3.594781082938425e-05)),(to_sfixed_a(-5.209679511608556e-05)),(to_sfixed_a(-6.384170410456136e-05)),(to_sfixed_a(-7.766922863083892e-06)),(to_sfixed_a(-0.00011014891788363457)),(to_sfixed_a(-1.3240228327049408e-05)),(to_sfixed_a(6.401179416570812e-05)),(to_sfixed_a(-1.7710453903418966e-05)),(to_sfixed_a(-2.430040512990672e-05)),(to_sfixed_a(-6.012067387928255e-05)),(to_sfixed_a(-1.560396958666388e-05)),(to_sfixed_a(-3.918636139133014e-05)),(to_sfixed_a(-4.121741221752018e-05)),(to_sfixed_a(4.952591098117409e-06)),(to_sfixed_a(-4.639543476514518e-05)),(to_sfixed_a(-5.438311563921161e-05)));

    constant weight_n1_139 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.17417477071285248)),(to_sfixed_a(-0.014531712047755718)),(to_sfixed_a(-0.06288982182741165)),(to_sfixed_a(0.07369698584079742)),(to_sfixed_a(0.002301538595929742)),(to_sfixed_a(-0.012017467059195042)),(to_sfixed_a(0.021631713956594467)),(to_sfixed_a(-0.006983216851949692)),(to_sfixed_a(-0.02291932888329029)),(to_sfixed_a(-0.045596588402986526)),(to_sfixed_a(0.03653758764266968)),(to_sfixed_a(-0.04220059514045715)),(to_sfixed_a(0.07469089329242706)),(to_sfixed_a(0.01349562220275402)),(to_sfixed_a(-0.048460446298122406)),(to_sfixed_a(0.004232123028486967)),(to_sfixed_a(-0.09900457412004471)),(to_sfixed_a(-0.004580573178827763)),(to_sfixed_a(0.017820989713072777)),(to_sfixed_a(0.12437949329614639)),(to_sfixed_a(0.04955938458442688)),(to_sfixed_a(-0.003446777816861868)),(to_sfixed_a(-0.03530440852046013)),(to_sfixed_a(0.07439938932657242)),(to_sfixed_a(0.033369068056344986)),(to_sfixed_a(-0.001391239813528955)),(to_sfixed_a(0.0948280394077301)),(to_sfixed_a(0.025362249463796616)),(to_sfixed_a(-0.021325362846255302)),(to_sfixed_a(0.09455481916666031)),(to_sfixed_a(0.046142324805259705)),(to_sfixed_a(-0.020819751545786858)),(to_sfixed_a(-0.05253154784440994)),(to_sfixed_a(0.07329178601503372)),(to_sfixed_a(-0.028957270085811615)),(to_sfixed_a(-0.12494339048862457)),(to_sfixed_a(-0.08828795701265335)),(to_sfixed_a(0.05659636855125427)));

    constant weight_n1_140 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.07514464110136032)),(to_sfixed_a(3.4844961191993207e-06)),(to_sfixed_a(-5.6670556659810245e-05)),(to_sfixed_a(3.2583458960289136e-05)),(to_sfixed_a(2.5214765628334135e-05)),(to_sfixed_a(1.230100588145433e-05)),(to_sfixed_a(-1.5993588021956384e-05)),(to_sfixed_a(-6.202108488650993e-05)),(to_sfixed_a(-1.93908217624994e-05)),(to_sfixed_a(-7.361808002315229e-06)),(to_sfixed_a(2.724012483668048e-05)),(to_sfixed_a(1.3158599358575884e-05)),(to_sfixed_a(7.5033531174995005e-06)),(to_sfixed_a(3.72887916455511e-05)),(to_sfixed_a(2.7053256417275406e-05)),(to_sfixed_a(-2.1836042378708953e-06)),(to_sfixed_a(-6.286506686592475e-05)),(to_sfixed_a(-6.0252910770941526e-05)),(to_sfixed_a(-1.5238539162965026e-05)),(to_sfixed_a(4.588323281495832e-05)),(to_sfixed_a(6.263814429985359e-05)),(to_sfixed_a(-3.47465138474945e-05)),(to_sfixed_a(5.2374602091731504e-05)),(to_sfixed_a(-1.1899177479790524e-05)),(to_sfixed_a(4.16465409216471e-05)),(to_sfixed_a(0.00012538211012724787)),(to_sfixed_a(-5.328696715878323e-05)),(to_sfixed_a(-8.679964230395854e-05)),(to_sfixed_a(-3.0708259146194905e-05)),(to_sfixed_a(4.270055069355294e-05)),(to_sfixed_a(-3.0742259696125984e-05)),(to_sfixed_a(2.820533154590521e-05)),(to_sfixed_a(3.7036720641481224e-06)),(to_sfixed_a(7.939418537716847e-06)),(to_sfixed_a(2.1947314962744713e-05)),(to_sfixed_a(1.4603770978283137e-05)),(to_sfixed_a(1.5846200767555274e-05)),(to_sfixed_a(-2.1885234673391096e-05)));

    constant weight_n1_141 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.016766933724284172)),(to_sfixed_a(-7.0339897320081946e-06)),(to_sfixed_a(-4.46337835455779e-05)),(to_sfixed_a(1.1195151273568626e-05)),(to_sfixed_a(-1.9212262486689724e-05)),(to_sfixed_a(-3.3753738534869626e-05)),(to_sfixed_a(-2.2277409073012677e-07)),(to_sfixed_a(-7.193077635747613e-06)),(to_sfixed_a(-5.232613602856873e-06)),(to_sfixed_a(0.00010629450844135135)),(to_sfixed_a(-0.00010156930511584505)),(to_sfixed_a(-2.5725161322043277e-05)),(to_sfixed_a(-1.4662931789644063e-05)),(to_sfixed_a(-4.40479516328196e-06)),(to_sfixed_a(2.3999524273676798e-05)),(to_sfixed_a(3.0184022762114182e-05)),(to_sfixed_a(-5.261702426651027e-06)),(to_sfixed_a(-1.6025031072786078e-05)),(to_sfixed_a(-3.794092845055275e-05)),(to_sfixed_a(-8.527958925697021e-06)),(to_sfixed_a(4.838505628868006e-05)),(to_sfixed_a(-2.7525888071977533e-05)),(to_sfixed_a(2.0604767996701412e-05)),(to_sfixed_a(3.473670221865177e-05)),(to_sfixed_a(-1.4863905562378932e-05)),(to_sfixed_a(1.8413018551655114e-05)),(to_sfixed_a(-5.0576629291754216e-05)),(to_sfixed_a(-4.9567104724701494e-05)),(to_sfixed_a(-6.464010948548093e-05)),(to_sfixed_a(5.098832116345875e-05)),(to_sfixed_a(3.1088045943761244e-05)),(to_sfixed_a(3.832266520475969e-05)),(to_sfixed_a(0.00010764671606011689)),(to_sfixed_a(-3.286470382590778e-05)),(to_sfixed_a(5.0503953389124945e-05)),(to_sfixed_a(-1.5913419701973908e-05)),(to_sfixed_a(8.400912338402122e-05)),(to_sfixed_a(5.9587982832454145e-05)));

    constant weight_n1_142 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.042253684252500534)),(to_sfixed_a(0.0348665826022625)),(to_sfixed_a(0.00046071773977018893)),(to_sfixed_a(-0.01375356875360012)),(to_sfixed_a(-0.009479868225753307)),(to_sfixed_a(0.012392857111990452)),(to_sfixed_a(0.019450608640909195)),(to_sfixed_a(-0.014747558161616325)),(to_sfixed_a(-0.004131569527089596)),(to_sfixed_a(-0.027729801833629608)),(to_sfixed_a(0.030505109578371048)),(to_sfixed_a(-0.01312269177287817)),(to_sfixed_a(-0.00036043766885995865)),(to_sfixed_a(0.0061921533197164536)),(to_sfixed_a(-0.003983674570918083)),(to_sfixed_a(0.0009963507764041424)),(to_sfixed_a(-0.03191615268588066)),(to_sfixed_a(-0.016462204977869987)),(to_sfixed_a(-0.03610633313655853)),(to_sfixed_a(-0.017058832570910454)),(to_sfixed_a(0.020306119695305824)),(to_sfixed_a(-0.015107779763638973)),(to_sfixed_a(-0.03854137659072876)),(to_sfixed_a(0.02051551826298237)),(to_sfixed_a(0.0027399456594139338)),(to_sfixed_a(-0.000528494012542069)),(to_sfixed_a(0.009239147417247295)),(to_sfixed_a(0.003881228156387806)),(to_sfixed_a(0.01816236786544323)),(to_sfixed_a(0.028515422716736794)),(to_sfixed_a(0.02871749736368656)),(to_sfixed_a(-0.018834363669157028)),(to_sfixed_a(-0.04770636558532715)),(to_sfixed_a(0.05704246833920479)),(to_sfixed_a(-0.05350315943360329)),(to_sfixed_a(0.0048622558824718)),(to_sfixed_a(0.0012088087387382984)),(to_sfixed_a(0.006269448436796665)));

    constant weight_n1_143 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.2181849479675293)),(to_sfixed_a(0.0366247221827507)),(to_sfixed_a(-0.03964253515005112)),(to_sfixed_a(-0.022095901891589165)),(to_sfixed_a(-0.13249267637729645)),(to_sfixed_a(0.08404255658388138)),(to_sfixed_a(-0.04946186766028404)),(to_sfixed_a(0.13673433661460876)),(to_sfixed_a(-0.04496212303638458)),(to_sfixed_a(-0.012730554677546024)),(to_sfixed_a(0.0033724759705364704)),(to_sfixed_a(0.00981360673904419)),(to_sfixed_a(0.052202511578798294)),(to_sfixed_a(-0.0007191224140115082)),(to_sfixed_a(-0.06365621834993362)),(to_sfixed_a(0.036679357290267944)),(to_sfixed_a(-0.07098256796598434)),(to_sfixed_a(-0.019789721816778183)),(to_sfixed_a(-0.005943066440522671)),(to_sfixed_a(0.005747673101723194)),(to_sfixed_a(-0.032917752861976624)),(to_sfixed_a(0.02811400778591633)),(to_sfixed_a(0.0191610436886549)),(to_sfixed_a(-0.05270885303616524)),(to_sfixed_a(-0.0024141755420714617)),(to_sfixed_a(0.003785169217735529)),(to_sfixed_a(0.0006846071337349713)),(to_sfixed_a(-0.03457939624786377)),(to_sfixed_a(-0.04997306317090988)),(to_sfixed_a(-0.003180833300575614)),(to_sfixed_a(0.040113914757966995)),(to_sfixed_a(0.06358341127634048)),(to_sfixed_a(-0.007718877401202917)),(to_sfixed_a(0.002074779476970434)),(to_sfixed_a(-0.024580424651503563)),(to_sfixed_a(-0.0012249568244442344)),(to_sfixed_a(0.01460556872189045)),(to_sfixed_a(-0.03227733448147774)));

    constant weight_n1_144 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.256603479385376)),(to_sfixed_a(0.004468761850148439)),(to_sfixed_a(0.011922852136194706)),(to_sfixed_a(-0.006624870467931032)),(to_sfixed_a(-0.004938516765832901)),(to_sfixed_a(-0.005406387150287628)),(to_sfixed_a(0.002208344405516982)),(to_sfixed_a(0.015578865073621273)),(to_sfixed_a(0.0097372867166996)),(to_sfixed_a(-0.017673930153250694)),(to_sfixed_a(0.03613457456231117)),(to_sfixed_a(-0.011969530023634434)),(to_sfixed_a(0.006238219328224659)),(to_sfixed_a(0.011584876105189323)),(to_sfixed_a(0.013801969587802887)),(to_sfixed_a(-0.024019936099648476)),(to_sfixed_a(-0.006424016319215298)),(to_sfixed_a(-0.006566192489117384)),(to_sfixed_a(0.0026275033596903086)),(to_sfixed_a(0.01641838252544403)),(to_sfixed_a(-0.012632431462407112)),(to_sfixed_a(0.0354728177189827)),(to_sfixed_a(0.007373819127678871)),(to_sfixed_a(-0.006430699955672026)),(to_sfixed_a(-0.006684142630547285)),(to_sfixed_a(0.030299736186861992)),(to_sfixed_a(0.011561780236661434)),(to_sfixed_a(-0.019605424255132675)),(to_sfixed_a(0.020434463396668434)),(to_sfixed_a(-0.0092870919033885)),(to_sfixed_a(-0.015499248169362545)),(to_sfixed_a(0.02522130310535431)),(to_sfixed_a(-0.025324249640107155)),(to_sfixed_a(0.01333553995937109)),(to_sfixed_a(-0.006096933502703905)),(to_sfixed_a(-0.045402005314826965)),(to_sfixed_a(0.0026127323508262634)),(to_sfixed_a(0.020857805386185646)));

    constant weight_n1_145 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.1021270677447319)),(to_sfixed_a(0.009230534546077251)),(to_sfixed_a(-0.0036888497415930033)),(to_sfixed_a(-0.026684079319238663)),(to_sfixed_a(0.003884996520355344)),(to_sfixed_a(-0.016479598358273506)),(to_sfixed_a(0.007610514760017395)),(to_sfixed_a(-0.0013045659288764)),(to_sfixed_a(-0.01611669547855854)),(to_sfixed_a(0.00853702612221241)),(to_sfixed_a(0.020587433129549026)),(to_sfixed_a(-0.030991196632385254)),(to_sfixed_a(0.012337383814156055)),(to_sfixed_a(0.016102826222777367)),(to_sfixed_a(-0.003052510553970933)),(to_sfixed_a(0.005961908493191004)),(to_sfixed_a(0.022029675543308258)),(to_sfixed_a(-0.023719847202301025)),(to_sfixed_a(-0.02666493132710457)),(to_sfixed_a(0.0035939423833042383)),(to_sfixed_a(-0.008635851554572582)),(to_sfixed_a(-0.009977219626307487)),(to_sfixed_a(-0.041289106011390686)),(to_sfixed_a(-0.008578353561460972)),(to_sfixed_a(0.012073537334799767)),(to_sfixed_a(0.013284667395055294)),(to_sfixed_a(0.02728075161576271)),(to_sfixed_a(-0.01772427000105381)),(to_sfixed_a(-0.01742442511022091)),(to_sfixed_a(-0.006926360540091991)),(to_sfixed_a(-0.02084708958864212)),(to_sfixed_a(0.008863838389515877)),(to_sfixed_a(-0.001486056367866695)),(to_sfixed_a(0.01749531738460064)),(to_sfixed_a(0.0023764558136463165)),(to_sfixed_a(-0.000823625479824841)),(to_sfixed_a(0.020032810047268867)),(to_sfixed_a(0.004088723100721836)));

    constant weight_n1_146 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.1323409527540207)),(to_sfixed_a(1.2117251571908128e-05)),(to_sfixed_a(-1.0767853382276371e-05)),(to_sfixed_a(6.142073107184842e-05)),(to_sfixed_a(5.327443068381399e-05)),(to_sfixed_a(0.00012062719906680286)),(to_sfixed_a(-1.774628253770061e-05)),(to_sfixed_a(-4.485070894588716e-05)),(to_sfixed_a(-2.8272566851228476e-05)),(to_sfixed_a(3.0625047656940296e-05)),(to_sfixed_a(-3.391010068298783e-06)),(to_sfixed_a(4.218743197270669e-05)),(to_sfixed_a(7.415356958517805e-05)),(to_sfixed_a(-5.4865620768396184e-05)),(to_sfixed_a(2.882048875108012e-06)),(to_sfixed_a(1.7330123228020966e-05)),(to_sfixed_a(8.918171806726605e-05)),(to_sfixed_a(-0.00010362280590925366)),(to_sfixed_a(-3.142471541650593e-05)),(to_sfixed_a(4.1870123823173344e-05)),(to_sfixed_a(-1.6846986909513362e-05)),(to_sfixed_a(-1.9732446162379347e-05)),(to_sfixed_a(-5.608598803519271e-05)),(to_sfixed_a(1.2011097169306595e-05)),(to_sfixed_a(-0.00010996322089340538)),(to_sfixed_a(-2.992042755067814e-05)),(to_sfixed_a(-1.7245542039745487e-05)),(to_sfixed_a(-3.2768944947747514e-05)),(to_sfixed_a(5.362475349102169e-05)),(to_sfixed_a(1.5846646419959143e-05)),(to_sfixed_a(-2.9104106943123043e-05)),(to_sfixed_a(8.262874325737357e-05)),(to_sfixed_a(1.5646495739929378e-05)),(to_sfixed_a(1.9134960894007236e-05)),(to_sfixed_a(-6.251316517591476e-05)),(to_sfixed_a(2.938350553449709e-05)),(to_sfixed_a(-7.096830086084083e-05)),(to_sfixed_a(5.508857066160999e-05)));

    constant weight_n1_147 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.008516574278473854)),(to_sfixed_a(-1.765231900208164e-05)),(to_sfixed_a(1.6919388144742697e-05)),(to_sfixed_a(6.536982709803851e-06)),(to_sfixed_a(6.963952046135091e-07)),(to_sfixed_a(-3.392025246284902e-05)),(to_sfixed_a(-7.670826744288206e-05)),(to_sfixed_a(-2.1060031940578483e-05)),(to_sfixed_a(3.419782660785131e-05)),(to_sfixed_a(-2.0386723917908967e-05)),(to_sfixed_a(-4.650802111427765e-06)),(to_sfixed_a(6.408845365513116e-05)),(to_sfixed_a(3.302729601273313e-05)),(to_sfixed_a(8.083176908257883e-06)),(to_sfixed_a(4.302049637772143e-05)),(to_sfixed_a(-2.58753243542742e-06)),(to_sfixed_a(5.006803621654399e-05)),(to_sfixed_a(-6.680985097773373e-05)),(to_sfixed_a(-4.783809345099144e-05)),(to_sfixed_a(3.5655408282764256e-05)),(to_sfixed_a(-1.5456129403901286e-05)),(to_sfixed_a(0.00012678596249315888)),(to_sfixed_a(-3.7006852835475e-06)),(to_sfixed_a(2.1218689653323963e-05)),(to_sfixed_a(1.8852015273296274e-05)),(to_sfixed_a(1.6853194892973988e-06)),(to_sfixed_a(6.0220325394766405e-05)),(to_sfixed_a(5.6279575801454484e-05)),(to_sfixed_a(-7.604670099681243e-05)),(to_sfixed_a(-4.935239121550694e-05)),(to_sfixed_a(1.6723728549550287e-05)),(to_sfixed_a(7.24437995813787e-05)),(to_sfixed_a(2.353954869249719e-06)),(to_sfixed_a(2.9321072361199185e-05)),(to_sfixed_a(8.506362064508721e-05)),(to_sfixed_a(-6.320383545244113e-05)),(to_sfixed_a(-3.017754715983756e-05)),(to_sfixed_a(-1.0343575922888704e-05)));

    constant weight_n1_148 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.15792615711688995)),(to_sfixed_a(-0.030241651460528374)),(to_sfixed_a(-0.005653179716318846)),(to_sfixed_a(0.0015765372663736343)),(to_sfixed_a(-0.04332064837217331)),(to_sfixed_a(0.002184156794101)),(to_sfixed_a(-0.013807201758027077)),(to_sfixed_a(-0.004658882971853018)),(to_sfixed_a(0.0123574398458004)),(to_sfixed_a(0.018457313999533653)),(to_sfixed_a(-0.012093763798475266)),(to_sfixed_a(0.007000316865742207)),(to_sfixed_a(0.0070856898091733456)),(to_sfixed_a(-0.029721064493060112)),(to_sfixed_a(-0.006098837126046419)),(to_sfixed_a(0.00732357706874609)),(to_sfixed_a(-0.026735275983810425)),(to_sfixed_a(0.022055380046367645)),(to_sfixed_a(0.009512120857834816)),(to_sfixed_a(-0.02436414547264576)),(to_sfixed_a(-0.0022856651339679956)),(to_sfixed_a(0.04434313252568245)),(to_sfixed_a(0.0007462732610292733)),(to_sfixed_a(0.03979798033833504)),(to_sfixed_a(0.007617240305989981)),(to_sfixed_a(-0.006770688109099865)),(to_sfixed_a(-0.042943645268678665)),(to_sfixed_a(0.017675725743174553)),(to_sfixed_a(-0.04698615521192551)),(to_sfixed_a(-0.036606114357709885)),(to_sfixed_a(-0.026356706395745277)),(to_sfixed_a(-0.012271786108613014)),(to_sfixed_a(-0.0052139610052108765)),(to_sfixed_a(0.0011706399964168668)),(to_sfixed_a(-0.030902696773409843)),(to_sfixed_a(-0.008502047508955002)),(to_sfixed_a(-0.043346405029296875)),(to_sfixed_a(-0.033150386065244675)));

    constant weight_n1_149 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.058288924396038055)),(to_sfixed_a(-1.566915125295054e-05)),(to_sfixed_a(8.701647857378703e-06)),(to_sfixed_a(-7.664570875931531e-05)),(to_sfixed_a(2.3098556994227692e-05)),(to_sfixed_a(4.507620906224474e-05)),(to_sfixed_a(3.3340740628773347e-05)),(to_sfixed_a(3.107244265265763e-05)),(to_sfixed_a(3.8210611819522455e-05)),(to_sfixed_a(7.060518692014739e-05)),(to_sfixed_a(1.5521274690399878e-05)),(to_sfixed_a(-1.4527719940815587e-05)),(to_sfixed_a(-6.233578005776508e-06)),(to_sfixed_a(3.25419896398671e-05)),(to_sfixed_a(1.8770825818137382e-06)),(to_sfixed_a(-7.26106227375567e-05)),(to_sfixed_a(-1.6625170246697962e-05)),(to_sfixed_a(-1.7440337614971213e-05)),(to_sfixed_a(-4.09347157983575e-05)),(to_sfixed_a(-3.3558975701453164e-05)),(to_sfixed_a(-4.296982297091745e-05)),(to_sfixed_a(-5.870259883522522e-06)),(to_sfixed_a(-1.8104316040989943e-05)),(to_sfixed_a(-3.6818059015786275e-05)),(to_sfixed_a(-4.634713695850223e-05)),(to_sfixed_a(-4.148454900132492e-05)),(to_sfixed_a(-4.129028820898384e-05)),(to_sfixed_a(-4.0239123336505145e-05)),(to_sfixed_a(-9.38007087825099e-06)),(to_sfixed_a(4.088714922545478e-05)),(to_sfixed_a(-4.560635261441348e-06)),(to_sfixed_a(0.0001223394792759791)),(to_sfixed_a(-7.871738489484414e-05)),(to_sfixed_a(8.985408203443512e-05)),(to_sfixed_a(7.352027751039714e-05)),(to_sfixed_a(-1.5067323147377465e-05)),(to_sfixed_a(5.676256841979921e-05)),(to_sfixed_a(1.8323744370718487e-05)));

    constant weight_n1_150 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.07871279865503311)),(to_sfixed_a(-8.49286952870898e-05)),(to_sfixed_a(3.8827205571578816e-05)),(to_sfixed_a(-7.109256330295466e-06)),(to_sfixed_a(-7.53613785491325e-05)),(to_sfixed_a(-1.2162819075456355e-05)),(to_sfixed_a(3.212753654224798e-05)),(to_sfixed_a(4.67588979518041e-05)),(to_sfixed_a(-8.762489414948504e-06)),(to_sfixed_a(-2.7093759854324162e-05)),(to_sfixed_a(4.9970367399509996e-05)),(to_sfixed_a(1.7947771993931383e-05)),(to_sfixed_a(3.90585046261549e-05)),(to_sfixed_a(-8.248217636719346e-05)),(to_sfixed_a(-3.262700920458883e-05)),(to_sfixed_a(1.9533295926521532e-05)),(to_sfixed_a(-5.408745437307516e-06)),(to_sfixed_a(1.4195470612321515e-05)),(to_sfixed_a(-4.9270376621279866e-05)),(to_sfixed_a(8.868724398780614e-05)),(to_sfixed_a(-4.7465739044127986e-05)),(to_sfixed_a(-1.7542957721161656e-05)),(to_sfixed_a(-5.789738497696817e-05)),(to_sfixed_a(-4.817467925022356e-05)),(to_sfixed_a(2.9391932912403718e-05)),(to_sfixed_a(-0.00016100675566121936)),(to_sfixed_a(-1.717764462227933e-05)),(to_sfixed_a(-9.500311716692522e-05)),(to_sfixed_a(-4.4735497795045376e-05)),(to_sfixed_a(2.6654894099920057e-05)),(to_sfixed_a(7.577568612759933e-05)),(to_sfixed_a(3.602154538384639e-05)),(to_sfixed_a(6.0385344113456085e-05)),(to_sfixed_a(1.353754851152189e-05)),(to_sfixed_a(-1.4462648323387839e-06)),(to_sfixed_a(2.534375016693957e-05)),(to_sfixed_a(-4.079970676684752e-05)),(to_sfixed_a(2.144641985069029e-05)));

    constant weight_n1_151 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.20059509575366974)),(to_sfixed_a(0.005504227709025145)),(to_sfixed_a(-0.008036253973841667)),(to_sfixed_a(0.02371777966618538)),(to_sfixed_a(0.0074083637446165085)),(to_sfixed_a(0.006037344224750996)),(to_sfixed_a(-0.019040612503886223)),(to_sfixed_a(0.017760159447789192)),(to_sfixed_a(-0.0077433413825929165)),(to_sfixed_a(0.00010026908421423286)),(to_sfixed_a(0.003930114675313234)),(to_sfixed_a(0.036204881966114044)),(to_sfixed_a(-0.060586050152778625)),(to_sfixed_a(-0.03128727152943611)),(to_sfixed_a(0.0038310782983899117)),(to_sfixed_a(0.008657561615109444)),(to_sfixed_a(-0.011459809727966785)),(to_sfixed_a(-0.025002729147672653)),(to_sfixed_a(-0.009113076142966747)),(to_sfixed_a(-0.02278841659426689)),(to_sfixed_a(-0.038407761603593826)),(to_sfixed_a(-0.05047912523150444)),(to_sfixed_a(0.018057042732834816)),(to_sfixed_a(-0.026460211724042892)),(to_sfixed_a(-0.05178886279463768)),(to_sfixed_a(0.009601948782801628)),(to_sfixed_a(-0.040424056351184845)),(to_sfixed_a(0.026098843663930893)),(to_sfixed_a(-0.01573793590068817)),(to_sfixed_a(0.01838955283164978)),(to_sfixed_a(0.010938339866697788)),(to_sfixed_a(0.0029440654907375574)),(to_sfixed_a(0.04749801382422447)),(to_sfixed_a(0.04409101977944374)),(to_sfixed_a(-0.011766382493078709)),(to_sfixed_a(-0.02824484184384346)),(to_sfixed_a(-0.01555678527802229)),(to_sfixed_a(0.0014908788725733757)));

    constant weight_n1_152 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.010537113063037395)),(to_sfixed_a(1.553635775053408e-05)),(to_sfixed_a(-3.6028490285389125e-05)),(to_sfixed_a(-8.519805305695627e-06)),(to_sfixed_a(-1.0937430488411337e-05)),(to_sfixed_a(-6.0774738813051954e-05)),(to_sfixed_a(-4.986835483578034e-05)),(to_sfixed_a(-7.415882282657549e-05)),(to_sfixed_a(-3.768296301132068e-05)),(to_sfixed_a(2.0633613530662842e-05)),(to_sfixed_a(3.6125547921983525e-05)),(to_sfixed_a(-6.162567842693534e-07)),(to_sfixed_a(4.6475954150082543e-05)),(to_sfixed_a(3.5139462397637544e-06)),(to_sfixed_a(9.1578485807986e-06)),(to_sfixed_a(-2.7700365535565652e-05)),(to_sfixed_a(-6.70471417834051e-05)),(to_sfixed_a(-4.777872527483851e-05)),(to_sfixed_a(-3.1375675462186337e-05)),(to_sfixed_a(-1.2775842151313554e-05)),(to_sfixed_a(-9.68347421803628e-07)),(to_sfixed_a(6.980648777243914e-06)),(to_sfixed_a(-6.169820699142292e-05)),(to_sfixed_a(7.916291360743344e-05)),(to_sfixed_a(4.61513627669774e-05)),(to_sfixed_a(-4.8022753617260605e-05)),(to_sfixed_a(1.2609091754711699e-05)),(to_sfixed_a(-2.7074458557763137e-05)),(to_sfixed_a(-3.688330252771266e-05)),(to_sfixed_a(6.0994207160547376e-05)),(to_sfixed_a(-2.585642687336076e-05)),(to_sfixed_a(8.956283272709697e-05)),(to_sfixed_a(-3.677808490465395e-05)),(to_sfixed_a(4.8496243834961206e-05)),(to_sfixed_a(-0.00011673079279717058)),(to_sfixed_a(-7.259777248691535e-06)),(to_sfixed_a(-1.5515835912083276e-05)),(to_sfixed_a(5.0654110964387655e-05)));

    constant weight_n1_153 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.07030119001865387)),(to_sfixed_a(-1.7995644157053903e-05)),(to_sfixed_a(-9.960450370272156e-06)),(to_sfixed_a(3.4942977436003275e-06)),(to_sfixed_a(-2.140736069122795e-05)),(to_sfixed_a(4.0008329960983247e-05)),(to_sfixed_a(-8.498386159772053e-05)),(to_sfixed_a(-7.335999544011429e-05)),(to_sfixed_a(2.7909538857784355e-06)),(to_sfixed_a(2.1107711290824227e-05)),(to_sfixed_a(3.0260060157161206e-05)),(to_sfixed_a(-3.795472366618924e-05)),(to_sfixed_a(-3.991214543930255e-05)),(to_sfixed_a(2.437399780319538e-05)),(to_sfixed_a(-2.640469574544113e-05)),(to_sfixed_a(9.252932613890152e-06)),(to_sfixed_a(2.078412398986984e-05)),(to_sfixed_a(-2.6716073989518918e-05)),(to_sfixed_a(-4.0827584598446265e-05)),(to_sfixed_a(0.00011996676767012104)),(to_sfixed_a(-1.1005398846464232e-05)),(to_sfixed_a(-4.927423651679419e-05)),(to_sfixed_a(-3.1380306609207764e-05)),(to_sfixed_a(1.449835781386355e-05)),(to_sfixed_a(-4.1090861486736685e-05)),(to_sfixed_a(-7.945421384647489e-05)),(to_sfixed_a(2.1090387235744856e-05)),(to_sfixed_a(-4.0996979805640876e-05)),(to_sfixed_a(2.3555279767606407e-05)),(to_sfixed_a(2.1731219021603465e-05)),(to_sfixed_a(-3.727246803464368e-05)),(to_sfixed_a(3.631763320299797e-05)),(to_sfixed_a(9.560107719153166e-05)),(to_sfixed_a(-8.744405931793153e-06)),(to_sfixed_a(-0.0001122977482737042)),(to_sfixed_a(-5.538156256079674e-05)),(to_sfixed_a(-0.0001714862883090973)),(to_sfixed_a(-6.602470875805011e-06)));

    constant weight_n1_154 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.10943152010440826)),(to_sfixed_a(0.02170414850115776)),(to_sfixed_a(-0.048202626407146454)),(to_sfixed_a(0.006138631142675877)),(to_sfixed_a(0.06776678562164307)),(to_sfixed_a(0.010870047844946384)),(to_sfixed_a(-0.03349132463335991)),(to_sfixed_a(0.0796092227101326)),(to_sfixed_a(0.043302763253450394)),(to_sfixed_a(-0.000514152692630887)),(to_sfixed_a(0.01708688959479332)),(to_sfixed_a(0.06781326234340668)),(to_sfixed_a(0.00632956949993968)),(to_sfixed_a(0.03469875454902649)),(to_sfixed_a(0.059914205223321915)),(to_sfixed_a(-0.02313772402703762)),(to_sfixed_a(0.028635451570153236)),(to_sfixed_a(-0.08644301444292068)),(to_sfixed_a(-0.1241266280412674)),(to_sfixed_a(-0.03400692716240883)),(to_sfixed_a(0.04358074814081192)),(to_sfixed_a(0.16818808019161224)),(to_sfixed_a(0.0811149999499321)),(to_sfixed_a(0.07182314246892929)),(to_sfixed_a(-0.02620047703385353)),(to_sfixed_a(-0.11117000132799149)),(to_sfixed_a(0.09489612281322479)),(to_sfixed_a(0.08836589753627777)),(to_sfixed_a(0.13949213922023773)),(to_sfixed_a(0.06358760595321655)),(to_sfixed_a(0.024861901998519897)),(to_sfixed_a(-0.048283617943525314)),(to_sfixed_a(0.036816515028476715)),(to_sfixed_a(-0.08358761668205261)),(to_sfixed_a(-0.0009803182911127806)),(to_sfixed_a(0.032981764525175095)),(to_sfixed_a(0.10581798851490021)),(to_sfixed_a(-0.07992745190858841)));

    constant weight_n1_155 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.02035353146493435)),(to_sfixed_a(2.0620429950213293e-06)),(to_sfixed_a(-3.1723015126772225e-05)),(to_sfixed_a(3.843639569822699e-05)),(to_sfixed_a(-1.1348396583343856e-05)),(to_sfixed_a(-0.00011121816351078451)),(to_sfixed_a(1.6561123629799113e-05)),(to_sfixed_a(-8.266638906206936e-05)),(to_sfixed_a(-2.2567484847968444e-05)),(to_sfixed_a(1.0957651284115855e-05)),(to_sfixed_a(4.45768419012893e-05)),(to_sfixed_a(-7.599936907354277e-06)),(to_sfixed_a(1.3932261026639026e-05)),(to_sfixed_a(-8.187210914911702e-05)),(to_sfixed_a(6.135419243946671e-05)),(to_sfixed_a(-6.0475758800748736e-05)),(to_sfixed_a(-2.8984351956751198e-05)),(to_sfixed_a(3.9475045923609287e-05)),(to_sfixed_a(-5.680082267645048e-06)),(to_sfixed_a(3.1988929549697787e-05)),(to_sfixed_a(-3.826415559160523e-05)),(to_sfixed_a(-7.595287024741992e-05)),(to_sfixed_a(-5.1670456741703674e-05)),(to_sfixed_a(-6.055960852791031e-07)),(to_sfixed_a(5.4163763707038015e-05)),(to_sfixed_a(-5.723734284401871e-05)),(to_sfixed_a(-1.4330054909805767e-05)),(to_sfixed_a(3.328278035041876e-05)),(to_sfixed_a(9.654147288529202e-05)),(to_sfixed_a(7.858149911044165e-05)),(to_sfixed_a(-7.999585068318993e-05)),(to_sfixed_a(-2.179698640247807e-05)),(to_sfixed_a(-3.1875199056230485e-05)),(to_sfixed_a(0.00013336693518795073)),(to_sfixed_a(4.448807885637507e-06)),(to_sfixed_a(7.735942199360579e-05)),(to_sfixed_a(8.943631110014394e-05)),(to_sfixed_a(0.00011247988732066005)));

    constant weight_n1_156 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.0816572979092598)),(to_sfixed_a(-0.007848934270441532)),(to_sfixed_a(-0.009098157286643982)),(to_sfixed_a(0.037814911454916)),(to_sfixed_a(-0.019204216077923775)),(to_sfixed_a(0.028646275401115417)),(to_sfixed_a(0.016072362661361694)),(to_sfixed_a(-0.010580458678305149)),(to_sfixed_a(0.03929847851395607)),(to_sfixed_a(0.014557759277522564)),(to_sfixed_a(0.0069676791317760944)),(to_sfixed_a(-0.01294022984802723)),(to_sfixed_a(-0.0006755802314728498)),(to_sfixed_a(-0.03602130338549614)),(to_sfixed_a(0.046531885862350464)),(to_sfixed_a(-0.036495573818683624)),(to_sfixed_a(0.036840178072452545)),(to_sfixed_a(0.08809193223714828)),(to_sfixed_a(-0.04250149056315422)),(to_sfixed_a(-0.0077972556464374065)),(to_sfixed_a(-0.02926955558359623)),(to_sfixed_a(0.046384893357753754)),(to_sfixed_a(-0.07413043826818466)),(to_sfixed_a(-0.04942317306995392)),(to_sfixed_a(-0.058579396456480026)),(to_sfixed_a(0.0644073337316513)),(to_sfixed_a(0.03563942760229111)),(to_sfixed_a(0.04088003933429718)),(to_sfixed_a(-0.08498282730579376)),(to_sfixed_a(0.1259547919034958)),(to_sfixed_a(0.0669797956943512)),(to_sfixed_a(0.02935461699962616)),(to_sfixed_a(0.01644941046833992)),(to_sfixed_a(0.0792527124285698)),(to_sfixed_a(0.06334861367940903)),(to_sfixed_a(0.02032136544585228)),(to_sfixed_a(-0.04290066286921501)),(to_sfixed_a(0.1334448754787445)));

    constant weight_n1_157 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.4024174213409424)),(to_sfixed_a(0.011853497475385666)),(to_sfixed_a(-0.00996487122029066)),(to_sfixed_a(0.01083659939467907)),(to_sfixed_a(-0.00017987402679864317)),(to_sfixed_a(-0.019831113517284393)),(to_sfixed_a(-8.462751429760829e-05)),(to_sfixed_a(-0.009419555775821209)),(to_sfixed_a(-0.0072759417816996574)),(to_sfixed_a(0.005889745429158211)),(to_sfixed_a(0.0014021340757608414)),(to_sfixed_a(-0.0007649605977348983)),(to_sfixed_a(0.003974770661443472)),(to_sfixed_a(0.0094258151948452)),(to_sfixed_a(-0.008398771286010742)),(to_sfixed_a(-0.008831159211695194)),(to_sfixed_a(-0.010569502599537373)),(to_sfixed_a(-0.0007308524218387902)),(to_sfixed_a(-0.01352381519973278)),(to_sfixed_a(-0.0010776249691843987)),(to_sfixed_a(0.011070581153035164)),(to_sfixed_a(0.0004566027782857418)),(to_sfixed_a(0.0048909373581409454)),(to_sfixed_a(-0.008646538481116295)),(to_sfixed_a(0.004155341070145369)),(to_sfixed_a(0.0029828171245753765)),(to_sfixed_a(0.0005631532985717058)),(to_sfixed_a(0.005407506134361029)),(to_sfixed_a(-0.0082633625715971)),(to_sfixed_a(-0.0034992313012480736)),(to_sfixed_a(0.009416542015969753)),(to_sfixed_a(-0.029182912781834602)),(to_sfixed_a(-0.0011080274125561118)),(to_sfixed_a(0.010963422246277332)),(to_sfixed_a(-0.01071970909833908)),(to_sfixed_a(-0.011526858434081078)),(to_sfixed_a(-0.029947614297270775)),(to_sfixed_a(0.015756534412503242)));

    constant weight_n1_158 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.14296528697013855)),(to_sfixed_a(4.181375970802037e-06)),(to_sfixed_a(3.2294187803927343e-06)),(to_sfixed_a(-2.9318703127501067e-06)),(to_sfixed_a(-2.2853605514683295e-06)),(to_sfixed_a(-1.4563269360223785e-05)),(to_sfixed_a(-2.5704221116029657e-05)),(to_sfixed_a(1.5697496564825997e-05)),(to_sfixed_a(6.982249760767445e-05)),(to_sfixed_a(-3.056129571632482e-06)),(to_sfixed_a(1.056368773788563e-06)),(to_sfixed_a(-1.6137637430801988e-05)),(to_sfixed_a(-2.824982857418945e-06)),(to_sfixed_a(4.299493866710691e-06)),(to_sfixed_a(5.7675541029311717e-05)),(to_sfixed_a(6.089644011808559e-05)),(to_sfixed_a(8.988003537524492e-05)),(to_sfixed_a(-1.3015737749810796e-05)),(to_sfixed_a(-3.580969132599421e-05)),(to_sfixed_a(2.9546332370955497e-05)),(to_sfixed_a(8.519766561221331e-05)),(to_sfixed_a(0.00010375535202911124)),(to_sfixed_a(-2.7530930310604163e-05)),(to_sfixed_a(5.154254176886752e-05)),(to_sfixed_a(-8.886076102498919e-06)),(to_sfixed_a(1.6264812074950896e-05)),(to_sfixed_a(8.978340338217095e-05)),(to_sfixed_a(7.234367512864992e-05)),(to_sfixed_a(-7.905740062597033e-07)),(to_sfixed_a(4.801362956641242e-05)),(to_sfixed_a(-9.158530156128109e-05)),(to_sfixed_a(2.0319828763604164e-05)),(to_sfixed_a(4.650789560400881e-05)),(to_sfixed_a(-4.332626849645749e-05)),(to_sfixed_a(7.1453265263699e-05)),(to_sfixed_a(-0.00013787085481453687)),(to_sfixed_a(2.6936770154861733e-05)),(to_sfixed_a(-5.334515662980266e-05)));

    constant weight_n1_159 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.054050691425800323)),(to_sfixed_a(2.1417865355033427e-05)),(to_sfixed_a(-5.307446917868219e-05)),(to_sfixed_a(3.0690720450365916e-05)),(to_sfixed_a(-3.662484959932044e-05)),(to_sfixed_a(4.9621626203588676e-06)),(to_sfixed_a(6.344455414364347e-06)),(to_sfixed_a(3.186697722412646e-05)),(to_sfixed_a(1.425995651516132e-05)),(to_sfixed_a(-3.905974517692812e-05)),(to_sfixed_a(1.110325047193328e-05)),(to_sfixed_a(-7.170481694629416e-06)),(to_sfixed_a(-1.3040485100646038e-05)),(to_sfixed_a(-3.4802412756107515e-06)),(to_sfixed_a(-2.5091698262258433e-05)),(to_sfixed_a(-4.264950257493183e-05)),(to_sfixed_a(3.9427895899279974e-06)),(to_sfixed_a(-1.1546096175152343e-05)),(to_sfixed_a(-4.092683957424015e-05)),(to_sfixed_a(2.8088414183002897e-05)),(to_sfixed_a(-0.00011403441749280319)),(to_sfixed_a(-3.395819658180699e-05)),(to_sfixed_a(2.902685446315445e-05)),(to_sfixed_a(-3.0512544526573038e-06)),(to_sfixed_a(6.532116094604135e-05)),(to_sfixed_a(-2.1525169358938e-05)),(to_sfixed_a(-7.793152326485142e-05)),(to_sfixed_a(1.6477215467602946e-05)),(to_sfixed_a(-2.8702756026177667e-05)),(to_sfixed_a(2.009933268709574e-05)),(to_sfixed_a(4.2915238736895844e-05)),(to_sfixed_a(7.160455425037071e-05)),(to_sfixed_a(-3.340498005854897e-05)),(to_sfixed_a(1.818508462747559e-05)),(to_sfixed_a(1.533093018224463e-05)),(to_sfixed_a(-6.745626160409302e-05)),(to_sfixed_a(8.690652066434268e-06)),(to_sfixed_a(4.146718492847867e-05)));

    constant weight_n1_160 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.018485886976122856)),(to_sfixed_a(3.212952651665546e-05)),(to_sfixed_a(7.856338197598234e-05)),(to_sfixed_a(-6.109546666266397e-05)),(to_sfixed_a(5.736670209444128e-05)),(to_sfixed_a(-4.754660767503083e-05)),(to_sfixed_a(4.236793756717816e-05)),(to_sfixed_a(-6.28314955974929e-06)),(to_sfixed_a(1.1928059393540025e-05)),(to_sfixed_a(2.7458727345219813e-05)),(to_sfixed_a(-1.9010334654012695e-05)),(to_sfixed_a(-5.612888344330713e-06)),(to_sfixed_a(1.832105772336945e-05)),(to_sfixed_a(1.7695283531793393e-05)),(to_sfixed_a(-2.5971514787670458e-06)),(to_sfixed_a(-1.010602409223793e-05)),(to_sfixed_a(-1.393117599945981e-05)),(to_sfixed_a(2.200178278144449e-05)),(to_sfixed_a(2.027614573307801e-05)),(to_sfixed_a(7.463113433914259e-05)),(to_sfixed_a(7.145421477616765e-06)),(to_sfixed_a(3.35625336447265e-05)),(to_sfixed_a(1.771906863723416e-05)),(to_sfixed_a(-1.6622632756480016e-05)),(to_sfixed_a(-4.45931545982603e-05)),(to_sfixed_a(5.209792288951576e-05)),(to_sfixed_a(1.4315645785245579e-05)),(to_sfixed_a(-1.2724292901111767e-05)),(to_sfixed_a(1.983356924029067e-05)),(to_sfixed_a(7.754950274829753e-06)),(to_sfixed_a(2.023014531005174e-05)),(to_sfixed_a(4.22063158111996e-06)),(to_sfixed_a(-7.32183616491966e-05)),(to_sfixed_a(5.578788841376081e-05)),(to_sfixed_a(2.1589532479993068e-05)),(to_sfixed_a(3.09779861709103e-05)),(to_sfixed_a(-7.278659904841334e-05)),(to_sfixed_a(-5.439580127131194e-05)));

    constant weight_n1_161 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.3709258437156677)),(to_sfixed_a(-0.0035115855280309916)),(to_sfixed_a(-0.0006381840794347227)),(to_sfixed_a(0.14972271025180817)),(to_sfixed_a(0.10159093886613846)),(to_sfixed_a(0.05001641437411308)),(to_sfixed_a(-0.024922188371419907)),(to_sfixed_a(0.07663683593273163)),(to_sfixed_a(0.12641118466854095)),(to_sfixed_a(0.06168639287352562)),(to_sfixed_a(0.04275994747877121)),(to_sfixed_a(0.12200150638818741)),(to_sfixed_a(0.03766511753201485)),(to_sfixed_a(-0.009570606052875519)),(to_sfixed_a(0.04620296508073807)),(to_sfixed_a(0.024470379576086998)),(to_sfixed_a(0.13281716406345367)),(to_sfixed_a(-0.04974937066435814)),(to_sfixed_a(-0.0773322582244873)),(to_sfixed_a(0.006579420994967222)),(to_sfixed_a(0.012578255496919155)),(to_sfixed_a(-0.08567190170288086)),(to_sfixed_a(-0.08010619878768921)),(to_sfixed_a(-0.09473419934511185)),(to_sfixed_a(0.04297560080885887)),(to_sfixed_a(-0.03051382675766945)),(to_sfixed_a(-0.04836747795343399)),(to_sfixed_a(0.02085777372121811)),(to_sfixed_a(-0.05539873242378235)),(to_sfixed_a(-0.11104936897754669)),(to_sfixed_a(-0.03518424928188324)),(to_sfixed_a(-0.030931266024708748)),(to_sfixed_a(0.1456466168165207)),(to_sfixed_a(0.07678178697824478)),(to_sfixed_a(-0.15757009387016296)),(to_sfixed_a(-0.16514965891838074)),(to_sfixed_a(-0.0023653744719922543)),(to_sfixed_a(0.037348419427871704)));

    constant weight_n1_162 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.05762486904859543)),(to_sfixed_a(0.014329244382679462)),(to_sfixed_a(0.0316382460296154)),(to_sfixed_a(0.0390157625079155)),(to_sfixed_a(-0.0881311446428299)),(to_sfixed_a(0.020193932577967644)),(to_sfixed_a(-0.009218416176736355)),(to_sfixed_a(-0.002705369843170047)),(to_sfixed_a(-0.036268219351768494)),(to_sfixed_a(-1.2146073459007312e-05)),(to_sfixed_a(0.025402769446372986)),(to_sfixed_a(-0.010991998948156834)),(to_sfixed_a(-0.0036110791843384504)),(to_sfixed_a(-0.06053854525089264)),(to_sfixed_a(-0.009748036973178387)),(to_sfixed_a(-0.050689924508333206)),(to_sfixed_a(0.03913086652755737)),(to_sfixed_a(0.04509493708610535)),(to_sfixed_a(-0.05811351165175438)),(to_sfixed_a(0.04386916756629944)),(to_sfixed_a(0.041007425636053085)),(to_sfixed_a(-0.018567871302366257)),(to_sfixed_a(0.060724079608917236)),(to_sfixed_a(-0.032569997012615204)),(to_sfixed_a(-0.06127263605594635)),(to_sfixed_a(-0.017411429435014725)),(to_sfixed_a(0.08827157318592072)),(to_sfixed_a(-0.029572851955890656)),(to_sfixed_a(-0.013103689067065716)),(to_sfixed_a(0.12291013449430466)),(to_sfixed_a(-0.03565807268023491)),(to_sfixed_a(0.009905756451189518)),(to_sfixed_a(0.049215905368328094)),(to_sfixed_a(0.011350139044225216)),(to_sfixed_a(-0.03142590820789337)),(to_sfixed_a(-0.004079571459442377)),(to_sfixed_a(0.01633242517709732)),(to_sfixed_a(-0.015727683901786804)));

    constant weight_n1_163 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.11680964380502701)),(to_sfixed_a(0.010528992861509323)),(to_sfixed_a(-0.018448974937200546)),(to_sfixed_a(0.01829030178487301)),(to_sfixed_a(-0.010313681326806545)),(to_sfixed_a(0.07172633707523346)),(to_sfixed_a(-0.04791552200913429)),(to_sfixed_a(-0.037073854357004166)),(to_sfixed_a(-0.0054710181429982185)),(to_sfixed_a(0.01250874437391758)),(to_sfixed_a(0.035634949803352356)),(to_sfixed_a(0.037915296852588654)),(to_sfixed_a(0.04625238850712776)),(to_sfixed_a(-0.022263094782829285)),(to_sfixed_a(-0.020007621496915817)),(to_sfixed_a(-0.03322368487715721)),(to_sfixed_a(-0.020214969292283058)),(to_sfixed_a(-0.042902037501335144)),(to_sfixed_a(-0.02853880263864994)),(to_sfixed_a(-0.07687176018953323)),(to_sfixed_a(-0.012053705751895905)),(to_sfixed_a(-0.06318626552820206)),(to_sfixed_a(-0.001824835897423327)),(to_sfixed_a(0.05195287615060806)),(to_sfixed_a(0.004347536247223616)),(to_sfixed_a(-0.020840154960751534)),(to_sfixed_a(-0.03589699789881706)),(to_sfixed_a(0.040410660207271576)),(to_sfixed_a(0.0051796226762235165)),(to_sfixed_a(0.0394902266561985)),(to_sfixed_a(0.03368060290813446)),(to_sfixed_a(-0.0013646832667291164)),(to_sfixed_a(0.0012866959441453218)),(to_sfixed_a(0.012982596643269062)),(to_sfixed_a(0.05409674718976021)),(to_sfixed_a(-0.04194014519453049)),(to_sfixed_a(0.012455865740776062)),(to_sfixed_a(-0.02062489464879036)));

    constant weight_n1_164 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.1328238546848297)),(to_sfixed_a(-0.003271864727139473)),(to_sfixed_a(-0.0031583246309310198)),(to_sfixed_a(0.06315986812114716)),(to_sfixed_a(-0.03246592357754707)),(to_sfixed_a(0.05437590181827545)),(to_sfixed_a(-0.03825460746884346)),(to_sfixed_a(0.11091317236423492)),(to_sfixed_a(0.010476925410330296)),(to_sfixed_a(-0.041161008179187775)),(to_sfixed_a(0.030752032995224)),(to_sfixed_a(0.029102226719260216)),(to_sfixed_a(0.11245160549879074)),(to_sfixed_a(0.016023579984903336)),(to_sfixed_a(0.05060208961367607)),(to_sfixed_a(-0.042419206351041794)),(to_sfixed_a(-0.006051347125321627)),(to_sfixed_a(-0.012386678718030453)),(to_sfixed_a(-0.08645126223564148)),(to_sfixed_a(0.013949917629361153)),(to_sfixed_a(0.017967738211154938)),(to_sfixed_a(-0.11267479509115219)),(to_sfixed_a(0.033373117446899414)),(to_sfixed_a(-0.06502074003219604)),(to_sfixed_a(-0.11317192018032074)),(to_sfixed_a(-0.03859329596161842)),(to_sfixed_a(-0.16598372161388397)),(to_sfixed_a(0.07498849928379059)),(to_sfixed_a(0.07045786082744598)),(to_sfixed_a(-0.03215546905994415)),(to_sfixed_a(0.009465333074331284)),(to_sfixed_a(-0.0721953809261322)),(to_sfixed_a(0.0034159484785050154)),(to_sfixed_a(0.09941542148590088)),(to_sfixed_a(-0.03002983145415783)),(to_sfixed_a(-0.11368779093027115)),(to_sfixed_a(0.03824812173843384)),(to_sfixed_a(-0.026721034198999405)));

    constant weight_n1_165 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.01698649302124977)),(to_sfixed_a(8.100284503598232e-06)),(to_sfixed_a(1.856123526522424e-05)),(to_sfixed_a(-2.1961619722787873e-07)),(to_sfixed_a(-1.7610245777177624e-05)),(to_sfixed_a(1.6337651686626486e-05)),(to_sfixed_a(-1.9090981368208304e-05)),(to_sfixed_a(3.24084862768359e-06)),(to_sfixed_a(2.4720638975850306e-05)),(to_sfixed_a(6.395441596396267e-05)),(to_sfixed_a(1.3460243280860595e-05)),(to_sfixed_a(1.4265936442825478e-05)),(to_sfixed_a(3.0370561944437213e-05)),(to_sfixed_a(2.7401016268413514e-05)),(to_sfixed_a(6.898325955262408e-05)),(to_sfixed_a(-1.269152471650159e-05)),(to_sfixed_a(3.732446930371225e-05)),(to_sfixed_a(1.4546688362315763e-05)),(to_sfixed_a(9.706453420221806e-05)),(to_sfixed_a(-3.878022835124284e-05)),(to_sfixed_a(-1.9336477635079063e-05)),(to_sfixed_a(7.507007831009105e-05)),(to_sfixed_a(1.4427307178266346e-05)),(to_sfixed_a(1.4030842066858895e-05)),(to_sfixed_a(-3.7195444747339934e-05)),(to_sfixed_a(-1.0357616702094674e-06)),(to_sfixed_a(8.406398592342157e-06)),(to_sfixed_a(-2.6425408577779308e-05)),(to_sfixed_a(2.337355363124516e-05)),(to_sfixed_a(-1.7929147361428477e-05)),(to_sfixed_a(1.911509571073111e-05)),(to_sfixed_a(-3.934789856430143e-05)),(to_sfixed_a(-4.557257125270553e-05)),(to_sfixed_a(-2.9136373996152543e-05)),(to_sfixed_a(1.3001699699088931e-05)),(to_sfixed_a(3.818326513282955e-05)),(to_sfixed_a(-1.6985461115837097e-05)),(to_sfixed_a(3.212899173377082e-05)));

    constant weight_n1_166 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.16304916143417358)),(to_sfixed_a(0.34312954545021057)),(to_sfixed_a(0.2985685467720032)),(to_sfixed_a(-0.1506289392709732)),(to_sfixed_a(0.16909605264663696)),(to_sfixed_a(-0.006658194586634636)),(to_sfixed_a(-0.173239603638649)),(to_sfixed_a(-0.004410916473716497)),(to_sfixed_a(0.0417947955429554)),(to_sfixed_a(0.10573562234640121)),(to_sfixed_a(0.08601371198892593)),(to_sfixed_a(0.036302994936704636)),(to_sfixed_a(-0.028887109830975533)),(to_sfixed_a(0.027297835797071457)),(to_sfixed_a(-0.0029033066239207983)),(to_sfixed_a(0.026868175715208054)),(to_sfixed_a(-0.019512411206960678)),(to_sfixed_a(0.11710642278194427)),(to_sfixed_a(0.0017740227049216628)),(to_sfixed_a(0.167699933052063)),(to_sfixed_a(-0.08189912140369415)),(to_sfixed_a(-0.13110265135765076)),(to_sfixed_a(-0.021285617724061012)),(to_sfixed_a(0.04688668251037598)),(to_sfixed_a(0.022052926942706108)),(to_sfixed_a(0.08168090134859085)),(to_sfixed_a(0.1468443125486374)),(to_sfixed_a(0.049978308379650116)),(to_sfixed_a(0.07068101316690445)),(to_sfixed_a(0.1898059993982315)),(to_sfixed_a(0.02914155274629593)),(to_sfixed_a(-0.0025528878904879093)),(to_sfixed_a(0.054400816559791565)),(to_sfixed_a(-0.050710562616586685)),(to_sfixed_a(-0.14418154954910278)),(to_sfixed_a(0.004376957658678293)),(to_sfixed_a(-0.019840853288769722)),(to_sfixed_a(0.0830332413315773)));

    constant weight_n1_167 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.04765930771827698)),(to_sfixed_a(2.1110055968165398e-05)),(to_sfixed_a(-9.960269380826503e-06)),(to_sfixed_a(-7.122028910089284e-05)),(to_sfixed_a(-2.5037927116500214e-05)),(to_sfixed_a(1.5805100701982155e-05)),(to_sfixed_a(-1.6880229622984189e-06)),(to_sfixed_a(-1.5389567124657333e-05)),(to_sfixed_a(7.454698788933456e-06)),(to_sfixed_a(1.5160258044488728e-05)),(to_sfixed_a(-3.048046892217826e-05)),(to_sfixed_a(8.382326996070333e-06)),(to_sfixed_a(6.899130676174536e-05)),(to_sfixed_a(-5.8735393395181745e-05)),(to_sfixed_a(-1.1144567906740122e-05)),(to_sfixed_a(4.486178113438655e-06)),(to_sfixed_a(-2.5346174879814498e-05)),(to_sfixed_a(-7.153535261750221e-05)),(to_sfixed_a(9.302410035161301e-05)),(to_sfixed_a(4.4913176679983735e-05)),(to_sfixed_a(5.221784249442862e-06)),(to_sfixed_a(1.8591159459901974e-05)),(to_sfixed_a(1.0569102414592635e-05)),(to_sfixed_a(5.765890023212705e-07)),(to_sfixed_a(-2.460205723764375e-05)),(to_sfixed_a(-1.61372336151544e-05)),(to_sfixed_a(1.1799659660027828e-05)),(to_sfixed_a(-1.280718879570486e-05)),(to_sfixed_a(8.668856753502041e-05)),(to_sfixed_a(5.2684012189274654e-05)),(to_sfixed_a(-1.1710946637322195e-05)),(to_sfixed_a(-1.5241451365000103e-05)),(to_sfixed_a(-2.3979695470188744e-05)),(to_sfixed_a(-2.9517224902519956e-05)),(to_sfixed_a(-5.0194379582535475e-05)),(to_sfixed_a(3.504000778775662e-05)),(to_sfixed_a(2.4263434170279652e-05)),(to_sfixed_a(8.595187682658434e-05)));

    constant weight_n1_168 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.037962958216667175)),(to_sfixed_a(1.947663986356929e-05)),(to_sfixed_a(-3.2498446671525016e-05)),(to_sfixed_a(3.771125420826138e-06)),(to_sfixed_a(-3.83260558010079e-05)),(to_sfixed_a(-3.768816441152012e-06)),(to_sfixed_a(-3.0329983928822912e-05)),(to_sfixed_a(2.7322765163262375e-05)),(to_sfixed_a(2.2814891053712927e-05)),(to_sfixed_a(-4.7643141442677006e-05)),(to_sfixed_a(-2.1484151147888042e-05)),(to_sfixed_a(-3.5535973438527435e-05)),(to_sfixed_a(-2.074338226520922e-05)),(to_sfixed_a(4.451953282114118e-05)),(to_sfixed_a(3.9922120777191594e-05)),(to_sfixed_a(-2.174654400732834e-05)),(to_sfixed_a(8.153659291565418e-05)),(to_sfixed_a(4.676598109654151e-05)),(to_sfixed_a(6.924064655322582e-05)),(to_sfixed_a(3.854317401419394e-05)),(to_sfixed_a(-4.2519201087998226e-05)),(to_sfixed_a(2.9225162506918423e-05)),(to_sfixed_a(-7.843877028790303e-06)),(to_sfixed_a(0.00010531816951697692)),(to_sfixed_a(-6.192110595293343e-05)),(to_sfixed_a(-2.0038454749737866e-05)),(to_sfixed_a(-3.0331910238601267e-05)),(to_sfixed_a(5.667601362802088e-05)),(to_sfixed_a(-4.006842209491879e-05)),(to_sfixed_a(-4.435586015461013e-05)),(to_sfixed_a(0.00014728319365531206)),(to_sfixed_a(-7.17120710760355e-05)),(to_sfixed_a(2.204619158874266e-05)),(to_sfixed_a(3.420665962039493e-05)),(to_sfixed_a(-4.294601967558265e-05)),(to_sfixed_a(2.491180202923715e-05)),(to_sfixed_a(1.1453968909336254e-05)),(to_sfixed_a(-2.2328102204483002e-05)));

    constant weight_n1_169 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.11858556419610977)),(to_sfixed_a(-0.03095490112900734)),(to_sfixed_a(-0.07047928869724274)),(to_sfixed_a(0.0619155615568161)),(to_sfixed_a(-0.021816516295075417)),(to_sfixed_a(-0.18899337947368622)),(to_sfixed_a(0.04302503913640976)),(to_sfixed_a(0.01799835078418255)),(to_sfixed_a(-0.09797124564647675)),(to_sfixed_a(-0.07487233728170395)),(to_sfixed_a(0.036666154861450195)),(to_sfixed_a(-0.04458865523338318)),(to_sfixed_a(-0.11999921500682831)),(to_sfixed_a(-0.1389600932598114)),(to_sfixed_a(-0.0419771745800972)),(to_sfixed_a(0.07739631831645966)),(to_sfixed_a(-0.045976605266332626)),(to_sfixed_a(0.07420812547206879)),(to_sfixed_a(0.02893490344285965)),(to_sfixed_a(-0.008684122003614902)),(to_sfixed_a(0.006105369422584772)),(to_sfixed_a(-0.09988800436258316)),(to_sfixed_a(-0.0974331870675087)),(to_sfixed_a(-0.0961364284157753)),(to_sfixed_a(6.91105960868299e-05)),(to_sfixed_a(0.19735054671764374)),(to_sfixed_a(0.11931045353412628)),(to_sfixed_a(0.03258656710386276)),(to_sfixed_a(0.030279535800218582)),(to_sfixed_a(0.03546953946352005)),(to_sfixed_a(0.07800928503274918)),(to_sfixed_a(-0.042696621268987656)),(to_sfixed_a(-0.027460088953375816)),(to_sfixed_a(0.06129182502627373)),(to_sfixed_a(0.011451821774244308)),(to_sfixed_a(0.007442581932991743)),(to_sfixed_a(0.030155370011925697)),(to_sfixed_a(0.062183719128370285)));

    constant weight_n1_170 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.20872575044631958)),(to_sfixed_a(0.0013202654663473368)),(to_sfixed_a(-0.00010241679410682991)),(to_sfixed_a(-0.001969127217307687)),(to_sfixed_a(-0.03525076061487198)),(to_sfixed_a(0.02628999389708042)),(to_sfixed_a(0.012030184268951416)),(to_sfixed_a(0.025457624346017838)),(to_sfixed_a(0.010289648547768593)),(to_sfixed_a(-0.023670833557844162)),(to_sfixed_a(0.05352318659424782)),(to_sfixed_a(0.026692332699894905)),(to_sfixed_a(0.030813096091151237)),(to_sfixed_a(0.055777981877326965)),(to_sfixed_a(0.006597296334803104)),(to_sfixed_a(-0.026786552742123604)),(to_sfixed_a(-0.05962293967604637)),(to_sfixed_a(-0.03530004248023033)),(to_sfixed_a(-0.022403830662369728)),(to_sfixed_a(0.032075583934783936)),(to_sfixed_a(0.013351657427847385)),(to_sfixed_a(0.014141653664410114)),(to_sfixed_a(-0.012719199992716312)),(to_sfixed_a(0.0030708429403603077)),(to_sfixed_a(-0.04358649253845215)),(to_sfixed_a(0.01249639131128788)),(to_sfixed_a(-0.010304944589734077)),(to_sfixed_a(0.05024410039186478)),(to_sfixed_a(-0.03907281160354614)),(to_sfixed_a(-0.01848328858613968)),(to_sfixed_a(-0.002332672942429781)),(to_sfixed_a(0.017407355830073357)),(to_sfixed_a(0.06146921217441559)),(to_sfixed_a(0.012917102314531803)),(to_sfixed_a(0.06394456326961517)),(to_sfixed_a(-0.014423087239265442)),(to_sfixed_a(0.006352557800710201)),(to_sfixed_a(-0.004980956204235554)));

    constant weight_n1_171 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.10045835375785828)),(to_sfixed_a(-0.025317562744021416)),(to_sfixed_a(-0.0010845860233530402)),(to_sfixed_a(0.014054866507649422)),(to_sfixed_a(0.004464203026145697)),(to_sfixed_a(-0.04100031033158302)),(to_sfixed_a(-0.0380406454205513)),(to_sfixed_a(0.027292722836136818)),(to_sfixed_a(0.05294708535075188)),(to_sfixed_a(-0.00471598282456398)),(to_sfixed_a(0.008558311499655247)),(to_sfixed_a(-0.02276037447154522)),(to_sfixed_a(0.02399798110127449)),(to_sfixed_a(-0.041373737156391144)),(to_sfixed_a(0.06301748752593994)),(to_sfixed_a(0.01702425442636013)),(to_sfixed_a(0.005270734429359436)),(to_sfixed_a(0.015003126114606857)),(to_sfixed_a(-0.020672636106610298)),(to_sfixed_a(-0.019165415316820145)),(to_sfixed_a(0.030339164659380913)),(to_sfixed_a(0.031977325677871704)),(to_sfixed_a(-0.01092161238193512)),(to_sfixed_a(0.008824017830193043)),(to_sfixed_a(-0.0309896357357502)),(to_sfixed_a(0.017513995990157127)),(to_sfixed_a(0.01593797281384468)),(to_sfixed_a(-0.05213276296854019)),(to_sfixed_a(0.051712069660425186)),(to_sfixed_a(0.003519331803545356)),(to_sfixed_a(0.027606435120105743)),(to_sfixed_a(0.04574928805232048)),(to_sfixed_a(-0.006215947214514017)),(to_sfixed_a(-0.05726275220513344)),(to_sfixed_a(0.0051806289702653885)),(to_sfixed_a(-0.054044418036937714)),(to_sfixed_a(-0.04015761986374855)),(to_sfixed_a(-0.044862210750579834)));

    constant weight_n1_172 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.011701256036758423)),(to_sfixed_a(-6.320178363239393e-05)),(to_sfixed_a(-1.1557872312550899e-06)),(to_sfixed_a(8.091356903605629e-06)),(to_sfixed_a(-2.026188485615421e-05)),(to_sfixed_a(-4.8091253120219335e-05)),(to_sfixed_a(-5.007955405744724e-05)),(to_sfixed_a(5.235735443420708e-05)),(to_sfixed_a(1.713456913421396e-05)),(to_sfixed_a(4.220953996991739e-05)),(to_sfixed_a(-3.5182097235519905e-06)),(to_sfixed_a(1.1772820471378509e-05)),(to_sfixed_a(-5.577604315476492e-05)),(to_sfixed_a(-6.246689736144617e-05)),(to_sfixed_a(4.32870319855283e-06)),(to_sfixed_a(-4.700997578765964e-06)),(to_sfixed_a(-1.7335929442197084e-05)),(to_sfixed_a(3.210593786207028e-05)),(to_sfixed_a(2.6724510462372564e-05)),(to_sfixed_a(-1.8739043298410252e-05)),(to_sfixed_a(-2.563730231486261e-05)),(to_sfixed_a(1.2734460597130237e-06)),(to_sfixed_a(-8.033560879994184e-05)),(to_sfixed_a(5.69272851862479e-05)),(to_sfixed_a(7.46066725696437e-05)),(to_sfixed_a(-5.3241936257109046e-05)),(to_sfixed_a(-4.23705751018133e-06)),(to_sfixed_a(4.764502227772027e-05)),(to_sfixed_a(-3.9961534639587626e-05)),(to_sfixed_a(-2.7120948288938962e-05)),(to_sfixed_a(-1.4491178262687754e-05)),(to_sfixed_a(-3.1875111744739115e-05)),(to_sfixed_a(-5.178237915970385e-05)),(to_sfixed_a(-1.2629047887458e-05)),(to_sfixed_a(6.833836232544854e-05)),(to_sfixed_a(3.850300345220603e-06)),(to_sfixed_a(-7.237902900669724e-05)),(to_sfixed_a(-1.0259908776788507e-05)));

    constant weight_n1_173 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.08198961615562439)),(to_sfixed_a(-0.061287425458431244)),(to_sfixed_a(-0.07199416309595108)),(to_sfixed_a(0.07442893832921982)),(to_sfixed_a(-0.01563175767660141)),(to_sfixed_a(-0.03377625346183777)),(to_sfixed_a(0.34530699253082275)),(to_sfixed_a(0.08989999443292618)),(to_sfixed_a(-0.11395382881164551)),(to_sfixed_a(0.3001696765422821)),(to_sfixed_a(0.24191758036613464)),(to_sfixed_a(-0.1569381058216095)),(to_sfixed_a(0.09209815412759781)),(to_sfixed_a(0.14067290723323822)),(to_sfixed_a(0.11834599822759628)),(to_sfixed_a(-0.06634824723005295)),(to_sfixed_a(0.1556435078382492)),(to_sfixed_a(-0.1288193017244339)),(to_sfixed_a(-0.08828971534967422)),(to_sfixed_a(0.007676247041672468)),(to_sfixed_a(-0.11924856156110764)),(to_sfixed_a(-0.05997046083211899)),(to_sfixed_a(0.1766039878129959)),(to_sfixed_a(-0.11345063149929047)),(to_sfixed_a(-0.2193308025598526)),(to_sfixed_a(0.025995459407567978)),(to_sfixed_a(0.15421423316001892)),(to_sfixed_a(-0.17488636076450348)),(to_sfixed_a(0.08191347867250443)),(to_sfixed_a(-0.1231246143579483)),(to_sfixed_a(0.08083692938089371)),(to_sfixed_a(0.11029066890478134)),(to_sfixed_a(-0.04427211731672287)),(to_sfixed_a(0.08625710755586624)),(to_sfixed_a(-0.03589755669236183)),(to_sfixed_a(0.004072707146406174)),(to_sfixed_a(0.0931214913725853)),(to_sfixed_a(-0.0033822960685938597)));

    constant weight_n1_174 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.16843871772289276)),(to_sfixed_a(-0.006430174224078655)),(to_sfixed_a(0.004038264974951744)),(to_sfixed_a(0.014500347897410393)),(to_sfixed_a(0.024100447073578835)),(to_sfixed_a(-0.043665338307619095)),(to_sfixed_a(-0.01933201402425766)),(to_sfixed_a(0.022770395502448082)),(to_sfixed_a(0.02889053337275982)),(to_sfixed_a(0.005474022589623928)),(to_sfixed_a(0.007674490101635456)),(to_sfixed_a(-0.0012766615254804492)),(to_sfixed_a(0.029837099835276604)),(to_sfixed_a(-0.027791576460003853)),(to_sfixed_a(0.027042347937822342)),(to_sfixed_a(0.007005220744758844)),(to_sfixed_a(-0.0013404481578618288)),(to_sfixed_a(0.007836690172553062)),(to_sfixed_a(-0.0015810682671144605)),(to_sfixed_a(-0.02183966524899006)),(to_sfixed_a(0.021929794922471046)),(to_sfixed_a(-0.00284789502620697)),(to_sfixed_a(-0.00657425494864583)),(to_sfixed_a(0.00020729529205709696)),(to_sfixed_a(-0.03196122124791145)),(to_sfixed_a(-0.01929224655032158)),(to_sfixed_a(0.02269763872027397)),(to_sfixed_a(-0.03315768763422966)),(to_sfixed_a(0.035149529576301575)),(to_sfixed_a(0.0402337945997715)),(to_sfixed_a(0.04817016422748566)),(to_sfixed_a(-0.0007017049938440323)),(to_sfixed_a(-0.00490364758297801)),(to_sfixed_a(-0.04605712369084358)),(to_sfixed_a(0.010115785524249077)),(to_sfixed_a(0.009512709453701973)),(to_sfixed_a(-0.01280661579221487)),(to_sfixed_a(-0.04006802290678024)));

    constant weight_n1_175 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.19803805649280548)),(to_sfixed_a(0.08440804481506348)),(to_sfixed_a(-0.0395955853164196)),(to_sfixed_a(0.05104059353470802)),(to_sfixed_a(0.050972770899534225)),(to_sfixed_a(-0.0362347774207592)),(to_sfixed_a(0.08257200568914413)),(to_sfixed_a(-0.03468726575374603)),(to_sfixed_a(0.03200565651059151)),(to_sfixed_a(0.008694524876773357)),(to_sfixed_a(0.052298229187726974)),(to_sfixed_a(-0.0375179685652256)),(to_sfixed_a(-0.08897413313388824)),(to_sfixed_a(0.030737128108739853)),(to_sfixed_a(0.04938855767250061)),(to_sfixed_a(-0.03370792418718338)),(to_sfixed_a(0.027606921270489693)),(to_sfixed_a(-0.030610572546720505)),(to_sfixed_a(0.07264365255832672)),(to_sfixed_a(0.00371400429867208)),(to_sfixed_a(-0.03333541378378868)),(to_sfixed_a(0.025345053523778915)),(to_sfixed_a(0.10998409986495972)),(to_sfixed_a(-0.09338915348052979)),(to_sfixed_a(0.09664618968963623)),(to_sfixed_a(-0.03890350088477135)),(to_sfixed_a(-0.05271795392036438)),(to_sfixed_a(-0.009665376506745815)),(to_sfixed_a(0.060867805033922195)),(to_sfixed_a(-0.02497093193233013)),(to_sfixed_a(0.026999490335583687)),(to_sfixed_a(0.06557536870241165)),(to_sfixed_a(0.018216382712125778)),(to_sfixed_a(0.023595765233039856)),(to_sfixed_a(0.12374956160783768)),(to_sfixed_a(0.04141346365213394)),(to_sfixed_a(0.012401117011904716)),(to_sfixed_a(0.0027008752804249525)));

    constant weight_n1_176 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.22192659974098206)),(to_sfixed_a(-0.003919451497495174)),(to_sfixed_a(-0.03187808766961098)),(to_sfixed_a(-0.007560476660728455)),(to_sfixed_a(-0.025680670514702797)),(to_sfixed_a(0.16949187219142914)),(to_sfixed_a(0.10227233916521072)),(to_sfixed_a(-0.01242757122963667)),(to_sfixed_a(0.08510599285364151)),(to_sfixed_a(-0.033692508935928345)),(to_sfixed_a(-0.028809456154704094)),(to_sfixed_a(0.10404311865568161)),(to_sfixed_a(0.0657617449760437)),(to_sfixed_a(0.039630331099033356)),(to_sfixed_a(0.029724910855293274)),(to_sfixed_a(-0.17642742395401)),(to_sfixed_a(0.0310997124761343)),(to_sfixed_a(0.1990208923816681)),(to_sfixed_a(-0.12071093916893005)),(to_sfixed_a(-0.04043235257267952)),(to_sfixed_a(0.007730549667030573)),(to_sfixed_a(0.22217358648777008)),(to_sfixed_a(-0.1189093068242073)),(to_sfixed_a(-0.2987063527107239)),(to_sfixed_a(-0.04186461865901947)),(to_sfixed_a(0.03987245261669159)),(to_sfixed_a(0.1428428441286087)),(to_sfixed_a(-0.02836724743247032)),(to_sfixed_a(-0.13664178550243378)),(to_sfixed_a(0.15957047045230865)),(to_sfixed_a(-0.14850136637687683)),(to_sfixed_a(0.10374059528112411)),(to_sfixed_a(-0.13452881574630737)),(to_sfixed_a(0.05045844241976738)),(to_sfixed_a(0.09440191835165024)),(to_sfixed_a(-0.061785001307725906)),(to_sfixed_a(-0.06452864408493042)),(to_sfixed_a(0.15733268857002258)));

    constant weight_n1_177 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.1536906659603119)),(to_sfixed_a(-0.07899069786071777)),(to_sfixed_a(0.056414760649204254)),(to_sfixed_a(0.05704674497246742)),(to_sfixed_a(-0.043398384004831314)),(to_sfixed_a(-0.08461941033601761)),(to_sfixed_a(0.07357113808393478)),(to_sfixed_a(-0.03666282817721367)),(to_sfixed_a(-0.0768902376294136)),(to_sfixed_a(0.052384186536073685)),(to_sfixed_a(-0.09253094345331192)),(to_sfixed_a(0.018022453412413597)),(to_sfixed_a(-0.019558778032660484)),(to_sfixed_a(0.04394761472940445)),(to_sfixed_a(0.07659032195806503)),(to_sfixed_a(0.22631680965423584)),(to_sfixed_a(0.03538535162806511)),(to_sfixed_a(0.08326302468776703)),(to_sfixed_a(0.20059140026569366)),(to_sfixed_a(0.0260000079870224)),(to_sfixed_a(-0.02359796315431595)),(to_sfixed_a(0.1928461343050003)),(to_sfixed_a(0.0033517328556627035)),(to_sfixed_a(0.027665602043271065)),(to_sfixed_a(-0.03422803804278374)),(to_sfixed_a(-0.061918556690216064)),(to_sfixed_a(-0.024692518636584282)),(to_sfixed_a(-0.041265424340963364)),(to_sfixed_a(0.10516972094774246)),(to_sfixed_a(-0.05460311844944954)),(to_sfixed_a(-0.11178365349769592)),(to_sfixed_a(-0.15779860317707062)),(to_sfixed_a(0.03044150397181511)),(to_sfixed_a(-0.028200233355164528)),(to_sfixed_a(-0.10584648698568344)),(to_sfixed_a(-0.09962183982133865)),(to_sfixed_a(0.05702771618962288)),(to_sfixed_a(-0.06618119031190872)));

    constant weight_n1_178 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.058876316994428635)),(to_sfixed_a(-0.08437737822532654)),(to_sfixed_a(0.17075315117835999)),(to_sfixed_a(-0.29055964946746826)),(to_sfixed_a(0.016879195347428322)),(to_sfixed_a(-0.15434996783733368)),(to_sfixed_a(0.2276814877986908)),(to_sfixed_a(0.2766950726509094)),(to_sfixed_a(0.14668208360671997)),(to_sfixed_a(-0.10999543964862823)),(to_sfixed_a(-0.10754801332950592)),(to_sfixed_a(0.01266290619969368)),(to_sfixed_a(-0.17843595147132874)),(to_sfixed_a(-0.04515041038393974)),(to_sfixed_a(-0.0034134462475776672)),(to_sfixed_a(-0.22675099968910217)),(to_sfixed_a(0.07207733392715454)),(to_sfixed_a(-0.036242272704839706)),(to_sfixed_a(0.17117850482463837)),(to_sfixed_a(0.005759031046181917)),(to_sfixed_a(0.12321974337100983)),(to_sfixed_a(0.04256761074066162)),(to_sfixed_a(0.020586878061294556)),(to_sfixed_a(-0.024777822196483612)),(to_sfixed_a(0.11594308167695999)),(to_sfixed_a(0.06110246106982231)),(to_sfixed_a(0.10479681938886642)),(to_sfixed_a(0.11110363900661469)),(to_sfixed_a(-0.18157030642032623)),(to_sfixed_a(-0.010990545153617859)),(to_sfixed_a(-0.021313006058335304)),(to_sfixed_a(-0.05716969072818756)),(to_sfixed_a(0.03418618068099022)),(to_sfixed_a(0.14815399050712585)),(to_sfixed_a(-0.2060050666332245)),(to_sfixed_a(0.001970230834558606)),(to_sfixed_a(0.14831209182739258)),(to_sfixed_a(0.01580881141126156)));

    constant weight_n1_179 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.1370323747396469)),(to_sfixed_a(0.005456695798784494)),(to_sfixed_a(0.010801258496940136)),(to_sfixed_a(-0.005461516324430704)),(to_sfixed_a(-0.013796263374388218)),(to_sfixed_a(0.004088421817868948)),(to_sfixed_a(-0.0024183138739317656)),(to_sfixed_a(-0.015946777537465096)),(to_sfixed_a(-0.003731442615389824)),(to_sfixed_a(-0.014586811885237694)),(to_sfixed_a(-0.0005125999450683594)),(to_sfixed_a(0.014473832212388515)),(to_sfixed_a(-0.011274718679487705)),(to_sfixed_a(-0.008617405779659748)),(to_sfixed_a(-0.01473701000213623)),(to_sfixed_a(-0.008873621933162212)),(to_sfixed_a(-0.007932644337415695)),(to_sfixed_a(0.02016732096672058)),(to_sfixed_a(-0.014330395497381687)),(to_sfixed_a(0.003655402222648263)),(to_sfixed_a(-0.008019128814339638)),(to_sfixed_a(0.01106270495802164)),(to_sfixed_a(-0.005543311592191458)),(to_sfixed_a(-0.013600016944110394)),(to_sfixed_a(0.0023920428939163685)),(to_sfixed_a(-0.017550231888890266)),(to_sfixed_a(0.007238158490508795)),(to_sfixed_a(-0.0013362381141632795)),(to_sfixed_a(-0.020018460229039192)),(to_sfixed_a(0.019105669111013412)),(to_sfixed_a(-0.011031728237867355)),(to_sfixed_a(-0.024925313889980316)),(to_sfixed_a(-0.011153128929436207)),(to_sfixed_a(-0.012457898817956448)),(to_sfixed_a(0.0115129379555583)),(to_sfixed_a(-0.005655509419739246)),(to_sfixed_a(0.0057809059508144855)),(to_sfixed_a(-0.0032275959383696318)));

    constant weight_n1_180 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.210197314620018)),(to_sfixed_a(0.013246554881334305)),(to_sfixed_a(0.014076389372348785)),(to_sfixed_a(-0.0004101865633856505)),(to_sfixed_a(-0.062182214111089706)),(to_sfixed_a(0.004690009634941816)),(to_sfixed_a(-0.009500572457909584)),(to_sfixed_a(0.024665016680955887)),(to_sfixed_a(0.02049744501709938)),(to_sfixed_a(0.08926310390233994)),(to_sfixed_a(-0.03434916213154793)),(to_sfixed_a(-0.0025402267929166555)),(to_sfixed_a(0.0033558669965714216)),(to_sfixed_a(0.002412100089713931)),(to_sfixed_a(0.18025745451450348)),(to_sfixed_a(-0.036932144314050674)),(to_sfixed_a(-0.06887132674455643)),(to_sfixed_a(-0.002605749061331153)),(to_sfixed_a(-0.07837921380996704)),(to_sfixed_a(-0.04323713853955269)),(to_sfixed_a(0.1614294797182083)),(to_sfixed_a(-0.025668032467365265)),(to_sfixed_a(-0.0017128816107288003)),(to_sfixed_a(0.020517531782388687)),(to_sfixed_a(0.15582922101020813)),(to_sfixed_a(0.20269638299942017)),(to_sfixed_a(-0.042230162769556046)),(to_sfixed_a(0.09835842996835709)),(to_sfixed_a(0.16238439083099365)),(to_sfixed_a(0.045226868242025375)),(to_sfixed_a(-0.023841558024287224)),(to_sfixed_a(0.1414758265018463)),(to_sfixed_a(-0.004579075612127781)),(to_sfixed_a(0.023455824702978134)),(to_sfixed_a(0.002934001386165619)),(to_sfixed_a(-0.10504589229822159)),(to_sfixed_a(-0.025949086993932724)),(to_sfixed_a(-0.13226161897182465)));

    constant weight_n1_181 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.020379148423671722)),(to_sfixed_a(9.239105565939099e-06)),(to_sfixed_a(-4.4464290112955496e-05)),(to_sfixed_a(3.3066971809603274e-05)),(to_sfixed_a(-2.2075029846746475e-05)),(to_sfixed_a(3.014275171153713e-05)),(to_sfixed_a(2.073277391900774e-05)),(to_sfixed_a(3.513978299451992e-05)),(to_sfixed_a(-4.755108420795295e-06)),(to_sfixed_a(1.3724497875955421e-05)),(to_sfixed_a(3.966917938669212e-05)),(to_sfixed_a(-4.6593568185926415e-06)),(to_sfixed_a(1.6087633412098512e-05)),(to_sfixed_a(-4.664734296966344e-05)),(to_sfixed_a(2.830830453603994e-05)),(to_sfixed_a(-2.9873242965550162e-05)),(to_sfixed_a(-5.613631583401002e-05)),(to_sfixed_a(2.847601535904687e-05)),(to_sfixed_a(-1.7116877643275075e-05)),(to_sfixed_a(-3.494730844977312e-05)),(to_sfixed_a(2.6357411115895957e-05)),(to_sfixed_a(-3.2599396945443004e-05)),(to_sfixed_a(1.314920973527478e-05)),(to_sfixed_a(5.055596193415113e-05)),(to_sfixed_a(-8.457613148493692e-06)),(to_sfixed_a(3.6236589949112386e-05)),(to_sfixed_a(-4.497586633078754e-05)),(to_sfixed_a(1.022140531858895e-05)),(to_sfixed_a(6.53538154438138e-05)),(to_sfixed_a(-5.327345206751488e-05)),(to_sfixed_a(-8.438668010057881e-05)),(to_sfixed_a(4.489295679377392e-05)),(to_sfixed_a(-4.379166421131231e-05)),(to_sfixed_a(5.605424667010084e-05)),(to_sfixed_a(7.299096614588052e-05)),(to_sfixed_a(5.212475298321806e-05)),(to_sfixed_a(-1.6054112847996294e-06)),(to_sfixed_a(4.724030804936774e-05)));

    constant weight_n1_182 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.055194806307554245)),(to_sfixed_a(-1.2799320757039823e-05)),(to_sfixed_a(-2.6429645004100166e-05)),(to_sfixed_a(-6.752013177901972e-06)),(to_sfixed_a(8.685768079885747e-06)),(to_sfixed_a(1.6306452380376868e-05)),(to_sfixed_a(-5.733177204092499e-06)),(to_sfixed_a(-4.595016434905119e-05)),(to_sfixed_a(1.8301062709724647e-06)),(to_sfixed_a(1.59646404540581e-07)),(to_sfixed_a(2.010147682085517e-06)),(to_sfixed_a(7.863505743443966e-05)),(to_sfixed_a(-1.914290351123782e-06)),(to_sfixed_a(-2.8266005756449886e-05)),(to_sfixed_a(4.879625703324564e-05)),(to_sfixed_a(-4.717812407761812e-05)),(to_sfixed_a(-1.2123662600060925e-05)),(to_sfixed_a(-3.5439352359389886e-05)),(to_sfixed_a(5.531435090233572e-05)),(to_sfixed_a(-2.385630295975716e-06)),(to_sfixed_a(-2.266043702547904e-05)),(to_sfixed_a(-3.3587533835088834e-05)),(to_sfixed_a(1.3535966900235508e-05)),(to_sfixed_a(-3.212415685993619e-05)),(to_sfixed_a(-9.75746206677286e-06)),(to_sfixed_a(-3.9201611798489466e-05)),(to_sfixed_a(5.586048791883513e-05)),(to_sfixed_a(-7.031605491647497e-05)),(to_sfixed_a(-1.8804498722602148e-06)),(to_sfixed_a(6.341520020214375e-06)),(to_sfixed_a(2.7953830795013346e-05)),(to_sfixed_a(-1.913257801788859e-05)),(to_sfixed_a(3.2174164516618475e-05)),(to_sfixed_a(-8.020789209695067e-06)),(to_sfixed_a(-0.0001074471729225479)),(to_sfixed_a(-2.4598268282716163e-05)),(to_sfixed_a(-0.00010682800348149613)),(to_sfixed_a(4.372495095594786e-05)));

    constant weight_n1_183 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.013391956686973572)),(to_sfixed_a(-4.035878737340681e-05)),(to_sfixed_a(2.1659343474311754e-05)),(to_sfixed_a(1.5094778063939884e-05)),(to_sfixed_a(-4.840337197720146e-08)),(to_sfixed_a(1.4542022654495668e-05)),(to_sfixed_a(7.945602192194201e-06)),(to_sfixed_a(-5.9108948335051537e-05)),(to_sfixed_a(4.535191328614019e-05)),(to_sfixed_a(3.9665621443418786e-05)),(to_sfixed_a(-2.6529696697252803e-05)),(to_sfixed_a(2.5223669581464492e-05)),(to_sfixed_a(-5.2616611355915666e-05)),(to_sfixed_a(5.178319952392485e-06)),(to_sfixed_a(-1.4881570677971467e-05)),(to_sfixed_a(-1.0933241355814971e-05)),(to_sfixed_a(-1.5044705833133776e-05)),(to_sfixed_a(-2.311681237188168e-05)),(to_sfixed_a(3.4668009902816266e-05)),(to_sfixed_a(3.9557820855407044e-05)),(to_sfixed_a(-2.8757844120264053e-05)),(to_sfixed_a(3.577667666831985e-05)),(to_sfixed_a(4.3290121539030224e-05)),(to_sfixed_a(-8.461092875222676e-06)),(to_sfixed_a(-4.9785587179940194e-05)),(to_sfixed_a(-3.7547186366282403e-05)),(to_sfixed_a(1.7402819139533676e-05)),(to_sfixed_a(-5.439186134026386e-05)),(to_sfixed_a(6.642656899202848e-06)),(to_sfixed_a(-1.9136128685204312e-05)),(to_sfixed_a(-2.545979805290699e-05)),(to_sfixed_a(-7.389055826934054e-05)),(to_sfixed_a(6.837592081865296e-05)),(to_sfixed_a(2.163254248443991e-05)),(to_sfixed_a(-1.709342177491635e-05)),(to_sfixed_a(-9.38847369980067e-06)),(to_sfixed_a(-2.932295683422126e-05)),(to_sfixed_a(1.6083145965239964e-05)));

    constant weight_n1_184 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.10231905430555344)),(to_sfixed_a(0.006342879496514797)),(to_sfixed_a(-0.0144991809502244)),(to_sfixed_a(0.02889443188905716)),(to_sfixed_a(-0.034762799739837646)),(to_sfixed_a(0.009228738024830818)),(to_sfixed_a(0.056203704327344894)),(to_sfixed_a(0.025912204757332802)),(to_sfixed_a(-0.06138576194643974)),(to_sfixed_a(-0.009307898581027985)),(to_sfixed_a(-0.03688035160303116)),(to_sfixed_a(0.05134217068552971)),(to_sfixed_a(0.05715280771255493)),(to_sfixed_a(0.0005474988138303161)),(to_sfixed_a(0.0435311421751976)),(to_sfixed_a(0.004494098015129566)),(to_sfixed_a(-0.055695563554763794)),(to_sfixed_a(0.004090665839612484)),(to_sfixed_a(-0.0289910975843668)),(to_sfixed_a(-0.014638441614806652)),(to_sfixed_a(0.0041299727745354176)),(to_sfixed_a(0.011765244416892529)),(to_sfixed_a(-0.040520086884498596)),(to_sfixed_a(0.054502375423908234)),(to_sfixed_a(-0.06379148364067078)),(to_sfixed_a(-0.011622166261076927)),(to_sfixed_a(0.04804510995745659)),(to_sfixed_a(0.01757495105266571)),(to_sfixed_a(-0.0666469931602478)),(to_sfixed_a(0.0622202530503273)),(to_sfixed_a(0.04018400236964226)),(to_sfixed_a(0.1127902939915657)),(to_sfixed_a(0.04526036977767944)),(to_sfixed_a(0.09234883636236191)),(to_sfixed_a(-0.023527665063738823)),(to_sfixed_a(-0.04918963462114334)),(to_sfixed_a(0.013412870466709137)),(to_sfixed_a(0.049848880618810654)));

    constant weight_n1_185 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.2381138801574707)),(to_sfixed_a(-0.005715264473110437)),(to_sfixed_a(-0.11345090717077255)),(to_sfixed_a(0.04177676513791084)),(to_sfixed_a(0.06807658076286316)),(to_sfixed_a(0.06642290949821472)),(to_sfixed_a(0.08843965083360672)),(to_sfixed_a(0.05904323235154152)),(to_sfixed_a(0.22125782072544098)),(to_sfixed_a(0.042459968477487564)),(to_sfixed_a(0.05840365216135979)),(to_sfixed_a(0.11771103739738464)),(to_sfixed_a(0.2678054869174957)),(to_sfixed_a(-0.08293411135673523)),(to_sfixed_a(0.0434684082865715)),(to_sfixed_a(-0.024346714839339256)),(to_sfixed_a(-0.00890273042023182)),(to_sfixed_a(0.3178127706050873)),(to_sfixed_a(-0.03816971927881241)),(to_sfixed_a(-0.01816190592944622)),(to_sfixed_a(0.13359099626541138)),(to_sfixed_a(0.15707823634147644)),(to_sfixed_a(-0.009281862527132034)),(to_sfixed_a(-0.0012827806640416384)),(to_sfixed_a(0.15120473504066467)),(to_sfixed_a(0.060668524354696274)),(to_sfixed_a(0.15971685945987701)),(to_sfixed_a(-0.060739945620298386)),(to_sfixed_a(0.09927820414304733)),(to_sfixed_a(-0.13071602582931519)),(to_sfixed_a(0.2819238603115082)),(to_sfixed_a(-0.1942223310470581)),(to_sfixed_a(0.05167309194803238)),(to_sfixed_a(-0.2260318100452423)),(to_sfixed_a(0.034403979778289795)),(to_sfixed_a(-0.017842380329966545)),(to_sfixed_a(0.10288752615451813)),(to_sfixed_a(-0.26425981521606445)));

    constant weight_n1_186 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.17303220927715302)),(to_sfixed_a(-0.0003757316735573113)),(to_sfixed_a(0.012512659654021263)),(to_sfixed_a(-0.00024861443671397865)),(to_sfixed_a(-0.012833784334361553)),(to_sfixed_a(0.005199226085096598)),(to_sfixed_a(0.024793488904833794)),(to_sfixed_a(0.0040023960173130035)),(to_sfixed_a(0.006863601040095091)),(to_sfixed_a(-0.004831724334508181)),(to_sfixed_a(-0.0068817539140582085)),(to_sfixed_a(-0.007753239944577217)),(to_sfixed_a(-0.007920486852526665)),(to_sfixed_a(0.014121051877737045)),(to_sfixed_a(-0.004808101803064346)),(to_sfixed_a(0.04215976223349571)),(to_sfixed_a(-0.02345506101846695)),(to_sfixed_a(0.044978294521570206)),(to_sfixed_a(0.04582515358924866)),(to_sfixed_a(0.007225809618830681)),(to_sfixed_a(-0.00511950021609664)),(to_sfixed_a(0.004737758543342352)),(to_sfixed_a(0.0019566714763641357)),(to_sfixed_a(0.0073518306016922)),(to_sfixed_a(-0.021764321252703667)),(to_sfixed_a(0.07644125819206238)),(to_sfixed_a(-0.02394280582666397)),(to_sfixed_a(-0.015342199243605137)),(to_sfixed_a(0.0032851386349648237)),(to_sfixed_a(-0.015917491167783737)),(to_sfixed_a(-0.008602398447692394)),(to_sfixed_a(0.0012647634139284492)),(to_sfixed_a(0.04588755592703819)),(to_sfixed_a(0.0354095920920372)),(to_sfixed_a(-0.030923478305339813)),(to_sfixed_a(0.0022223631385713816)),(to_sfixed_a(-0.03437737002968788)),(to_sfixed_a(0.019395610317587852)));

    constant weight_n1_187 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.059281639754772186)),(to_sfixed_a(0.011077646166086197)),(to_sfixed_a(-0.011379018425941467)),(to_sfixed_a(-0.0053727999329566956)),(to_sfixed_a(-0.005487427115440369)),(to_sfixed_a(0.01424458995461464)),(to_sfixed_a(0.010562943294644356)),(to_sfixed_a(0.0026083518750965595)),(to_sfixed_a(0.013591025955975056)),(to_sfixed_a(-0.0026414445601403713)),(to_sfixed_a(-0.019365180283784866)),(to_sfixed_a(-0.0029982533305883408)),(to_sfixed_a(-0.00976898055523634)),(to_sfixed_a(0.003917952999472618)),(to_sfixed_a(0.004462895914912224)),(to_sfixed_a(0.00012925133341923356)),(to_sfixed_a(-0.017427148297429085)),(to_sfixed_a(0.0017645664047449827)),(to_sfixed_a(-0.015531593933701515)),(to_sfixed_a(-0.0067016915418207645)),(to_sfixed_a(-0.002929327543824911)),(to_sfixed_a(-0.007466404233127832)),(to_sfixed_a(0.007470109965652227)),(to_sfixed_a(-0.0018938705325126648)),(to_sfixed_a(0.03134170174598694)),(to_sfixed_a(0.022440165281295776)),(to_sfixed_a(0.007723646238446236)),(to_sfixed_a(0.01368300523608923)),(to_sfixed_a(-0.03152547404170036)),(to_sfixed_a(-0.0001204788131872192)),(to_sfixed_a(-0.01096198707818985)),(to_sfixed_a(0.031147075816988945)),(to_sfixed_a(0.004528792109340429)),(to_sfixed_a(0.006261779926717281)),(to_sfixed_a(-0.0023447766434401274)),(to_sfixed_a(-0.010200314223766327)),(to_sfixed_a(-0.0016984886024147272)),(to_sfixed_a(0.0037181267980486155)));

    constant weight_n1_188 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.38805946707725525)),(to_sfixed_a(0.010045185685157776)),(to_sfixed_a(0.01633141189813614)),(to_sfixed_a(-0.008668382652103901)),(to_sfixed_a(0.04146168380975723)),(to_sfixed_a(0.007082877680659294)),(to_sfixed_a(0.0427737683057785)),(to_sfixed_a(-0.0044386968947947025)),(to_sfixed_a(-0.10123955458402634)),(to_sfixed_a(0.10762001574039459)),(to_sfixed_a(-0.020386267453432083)),(to_sfixed_a(-0.02281266637146473)),(to_sfixed_a(0.03449513018131256)),(to_sfixed_a(0.009519961662590504)),(to_sfixed_a(-0.023464906960725784)),(to_sfixed_a(-0.026115600019693375)),(to_sfixed_a(-0.023216629400849342)),(to_sfixed_a(0.028833620250225067)),(to_sfixed_a(0.004639809485524893)),(to_sfixed_a(0.10580015927553177)),(to_sfixed_a(-0.029652941972017288)),(to_sfixed_a(0.0005937485839240253)),(to_sfixed_a(-0.10968200117349625)),(to_sfixed_a(0.08303230255842209)),(to_sfixed_a(0.010591037571430206)),(to_sfixed_a(0.010057557374238968)),(to_sfixed_a(0.03700726479291916)),(to_sfixed_a(0.10645594447851181)),(to_sfixed_a(-0.01314384676516056)),(to_sfixed_a(-0.06647053360939026)),(to_sfixed_a(0.010742050595581532)),(to_sfixed_a(0.061502594500780106)),(to_sfixed_a(-0.012747466564178467)),(to_sfixed_a(0.023473558947443962)),(to_sfixed_a(0.031912896782159805)),(to_sfixed_a(-0.11644037812948227)),(to_sfixed_a(-0.02050809934735298)),(to_sfixed_a(0.04861881583929062)));

    constant weight_n1_189 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.18190154433250427)),(to_sfixed_a(0.006847519427537918)),(to_sfixed_a(0.019272079691290855)),(to_sfixed_a(0.008788537234067917)),(to_sfixed_a(-0.04238079860806465)),(to_sfixed_a(-0.020953845232725143)),(to_sfixed_a(0.013378402218222618)),(to_sfixed_a(-0.013128533028066158)),(to_sfixed_a(-0.03805921599268913)),(to_sfixed_a(0.019398268312215805)),(to_sfixed_a(0.04374014958739281)),(to_sfixed_a(-0.06687670201063156)),(to_sfixed_a(0.013365698978304863)),(to_sfixed_a(-0.033921074122190475)),(to_sfixed_a(-0.012323031201958656)),(to_sfixed_a(-0.013728833757340908)),(to_sfixed_a(-0.04176237806677818)),(to_sfixed_a(0.05550533905625343)),(to_sfixed_a(0.031067656353116035)),(to_sfixed_a(-0.03570958971977234)),(to_sfixed_a(-4.6486466089845635e-06)),(to_sfixed_a(-0.008018199354410172)),(to_sfixed_a(0.03679399937391281)),(to_sfixed_a(-0.0405820868909359)),(to_sfixed_a(-0.005691920407116413)),(to_sfixed_a(0.06593506038188934)),(to_sfixed_a(0.0027240756899118423)),(to_sfixed_a(-0.01993895135819912)),(to_sfixed_a(-0.012097004801034927)),(to_sfixed_a(0.017101889476180077)),(to_sfixed_a(0.011858719401061535)),(to_sfixed_a(-0.0031635938212275505)),(to_sfixed_a(0.045155011117458344)),(to_sfixed_a(-0.014916840940713882)),(to_sfixed_a(0.02417110651731491)),(to_sfixed_a(0.03762554004788399)),(to_sfixed_a(0.09210380911827087)),(to_sfixed_a(-0.047491058707237244)));

    constant weight_n1_190 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.016298454254865646)),(to_sfixed_a(3.0962117307353765e-05)),(to_sfixed_a(-5.0630820624064654e-05)),(to_sfixed_a(-3.8331661926349625e-05)),(to_sfixed_a(5.7036682846955955e-05)),(to_sfixed_a(2.6524169243202778e-06)),(to_sfixed_a(1.7426211343263276e-05)),(to_sfixed_a(-4.710745997726917e-05)),(to_sfixed_a(-3.208335328963585e-05)),(to_sfixed_a(-4.4429554691305384e-05)),(to_sfixed_a(8.230936509789899e-05)),(to_sfixed_a(6.407259206753224e-05)),(to_sfixed_a(7.65113509260118e-05)),(to_sfixed_a(-5.802858140668832e-05)),(to_sfixed_a(3.20007347909268e-05)),(to_sfixed_a(3.4290813346160576e-05)),(to_sfixed_a(6.787021266063675e-05)),(to_sfixed_a(-2.236420550616458e-05)),(to_sfixed_a(-6.685044809273677e-06)),(to_sfixed_a(1.0273131920257583e-05)),(to_sfixed_a(7.190401811385527e-05)),(to_sfixed_a(-1.6938716726144776e-05)),(to_sfixed_a(3.541938713169657e-05)),(to_sfixed_a(7.750057557132095e-05)),(to_sfixed_a(-4.678185359807685e-05)),(to_sfixed_a(-0.00010166845459025353)),(to_sfixed_a(-1.0123949323315173e-05)),(to_sfixed_a(-7.012677087914199e-05)),(to_sfixed_a(0.00010565459524514154)),(to_sfixed_a(4.523224924923852e-05)),(to_sfixed_a(4.009278927696869e-05)),(to_sfixed_a(2.9115475626895204e-05)),(to_sfixed_a(-8.205858466681093e-05)),(to_sfixed_a(0.00012038164277328178)),(to_sfixed_a(4.8859594244277105e-05)),(to_sfixed_a(1.3837167898600455e-05)),(to_sfixed_a(-2.609015064081177e-05)),(to_sfixed_a(-0.00022215482022147626)));

    constant weight_n1_191 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.2011478841304779)),(to_sfixed_a(0.0781405046582222)),(to_sfixed_a(0.08392807841300964)),(to_sfixed_a(-0.08554165065288544)),(to_sfixed_a(0.07700423896312714)),(to_sfixed_a(-0.0020303053315728903)),(to_sfixed_a(-0.04011780023574829)),(to_sfixed_a(-0.009251109324395657)),(to_sfixed_a(-0.0976710394024849)),(to_sfixed_a(0.021699974313378334)),(to_sfixed_a(0.07547741383314133)),(to_sfixed_a(0.001976604340597987)),(to_sfixed_a(-0.0312880240380764)),(to_sfixed_a(0.1116296574473381)),(to_sfixed_a(0.0020419659558683634)),(to_sfixed_a(-0.013026492670178413)),(to_sfixed_a(-0.01925147883594036)),(to_sfixed_a(-0.08038250356912613)),(to_sfixed_a(-0.1085968017578125)),(to_sfixed_a(0.08017272502183914)),(to_sfixed_a(-0.009319823235273361)),(to_sfixed_a(-0.05533970147371292)),(to_sfixed_a(-0.05315861850976944)),(to_sfixed_a(0.03809123486280441)),(to_sfixed_a(-0.025597818195819855)),(to_sfixed_a(-0.12666592001914978)),(to_sfixed_a(0.12321306765079498)),(to_sfixed_a(0.038245365023612976)),(to_sfixed_a(0.03418253734707832)),(to_sfixed_a(-0.07257082313299179)),(to_sfixed_a(0.07451089471578598)),(to_sfixed_a(0.015106488950550556)),(to_sfixed_a(0.02129128947854042)),(to_sfixed_a(-0.20745155215263367)),(to_sfixed_a(0.05678556114435196)),(to_sfixed_a(0.07589292526245117)),(to_sfixed_a(0.18649129569530487)),(to_sfixed_a(0.009386129677295685)));

    constant weight_n1_192 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.15308284759521484)),(to_sfixed_a(-0.006265909876674414)),(to_sfixed_a(0.07083327323198318)),(to_sfixed_a(0.11072918027639389)),(to_sfixed_a(0.1097131073474884)),(to_sfixed_a(0.023565830662846565)),(to_sfixed_a(0.011963172815740108)),(to_sfixed_a(0.11933538317680359)),(to_sfixed_a(-0.005921636708080769)),(to_sfixed_a(-0.029424399137496948)),(to_sfixed_a(0.03854987770318985)),(to_sfixed_a(-0.061838243156671524)),(to_sfixed_a(-0.05636409670114517)),(to_sfixed_a(0.0486786849796772)),(to_sfixed_a(-0.05025991052389145)),(to_sfixed_a(0.042705800384283066)),(to_sfixed_a(0.01566811464726925)),(to_sfixed_a(-0.030680609866976738)),(to_sfixed_a(-0.12227161228656769)),(to_sfixed_a(0.004722920712083578)),(to_sfixed_a(0.0678272545337677)),(to_sfixed_a(-0.0346391461789608)),(to_sfixed_a(0.006055878475308418)),(to_sfixed_a(-0.06645387411117554)),(to_sfixed_a(-0.0023369896225631237)),(to_sfixed_a(0.004160245414823294)),(to_sfixed_a(-0.034041136503219604)),(to_sfixed_a(-0.09696560353040695)),(to_sfixed_a(-0.05168551951646805)),(to_sfixed_a(0.00843896996229887)),(to_sfixed_a(0.02056465856730938)),(to_sfixed_a(-0.10754009336233139)),(to_sfixed_a(0.0361676886677742)),(to_sfixed_a(0.06242568418383598)),(to_sfixed_a(0.05192100629210472)),(to_sfixed_a(0.006854651030153036)),(to_sfixed_a(0.1719488948583603)),(to_sfixed_a(0.03219631314277649)));

    constant weight_n1_193 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.07964950054883957)),(to_sfixed_a(1.384579149998899e-06)),(to_sfixed_a(1.861368218669668e-05)),(to_sfixed_a(9.394311928190291e-05)),(to_sfixed_a(-4.614249746737187e-07)),(to_sfixed_a(-4.862928471993655e-05)),(to_sfixed_a(-1.2695571058429778e-05)),(to_sfixed_a(9.309573215432465e-06)),(to_sfixed_a(4.149332653469173e-06)),(to_sfixed_a(8.767979306867346e-05)),(to_sfixed_a(1.7244545233552344e-05)),(to_sfixed_a(2.899331593653187e-05)),(to_sfixed_a(1.0514860150578897e-05)),(to_sfixed_a(-1.622000490897335e-05)),(to_sfixed_a(-2.6053714464069344e-05)),(to_sfixed_a(1.3626063264382537e-05)),(to_sfixed_a(7.994314364623278e-05)),(to_sfixed_a(8.0141880971496e-06)),(to_sfixed_a(2.4071601728792302e-05)),(to_sfixed_a(-3.544277205946855e-05)),(to_sfixed_a(3.957690569222905e-05)),(to_sfixed_a(-2.4015427698032e-05)),(to_sfixed_a(1.5420875570271164e-05)),(to_sfixed_a(-4.0757557144388556e-05)),(to_sfixed_a(-1.3438906535157003e-05)),(to_sfixed_a(-3.779110193136148e-05)),(to_sfixed_a(-6.989749181229854e-06)),(to_sfixed_a(4.0481496398570016e-05)),(to_sfixed_a(-0.00010301629663445055)),(to_sfixed_a(8.466216740998789e-07)),(to_sfixed_a(1.782213189471804e-06)),(to_sfixed_a(-3.905354969901964e-05)),(to_sfixed_a(5.723802314605564e-05)),(to_sfixed_a(6.276211024669465e-06)),(to_sfixed_a(2.7503917863214156e-06)),(to_sfixed_a(7.826363435015082e-05)),(to_sfixed_a(-2.7594592211244162e-06)),(to_sfixed_a(3.609434861573391e-05)));

    constant weight_n1_194 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.04810601845383644)),(to_sfixed_a(-0.11013729125261307)),(to_sfixed_a(0.27508774399757385)),(to_sfixed_a(0.218402698636055)),(to_sfixed_a(0.09013793617486954)),(to_sfixed_a(0.3599816858768463)),(to_sfixed_a(0.04180912300944328)),(to_sfixed_a(0.14123627543449402)),(to_sfixed_a(0.022652659565210342)),(to_sfixed_a(-0.020771630108356476)),(to_sfixed_a(-0.06496359407901764)),(to_sfixed_a(0.03878036141395569)),(to_sfixed_a(-0.1505296677350998)),(to_sfixed_a(-0.09820390492677689)),(to_sfixed_a(0.09453504532575607)),(to_sfixed_a(0.06571224331855774)),(to_sfixed_a(-0.08699453622102737)),(to_sfixed_a(0.004022065084427595)),(to_sfixed_a(0.1518716961145401)),(to_sfixed_a(-0.0017247096402570605)),(to_sfixed_a(-0.10965780913829803)),(to_sfixed_a(-0.007575450465083122)),(to_sfixed_a(0.004311169032007456)),(to_sfixed_a(-0.0058663999661803246)),(to_sfixed_a(-0.03237098455429077)),(to_sfixed_a(0.0006820198032073677)),(to_sfixed_a(-0.059820033609867096)),(to_sfixed_a(0.01670018397271633)),(to_sfixed_a(0.06079808995127678)),(to_sfixed_a(0.13175883889198303)),(to_sfixed_a(0.19996052980422974)),(to_sfixed_a(-0.02228798344731331)),(to_sfixed_a(-0.023953920230269432)),(to_sfixed_a(0.018467819318175316)),(to_sfixed_a(-0.010458261705935001)),(to_sfixed_a(-0.12663187086582184)),(to_sfixed_a(0.16469885408878326)),(to_sfixed_a(-0.027998512610793114)));

    constant weight_n1_195 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.011521149426698685)),(to_sfixed_a(2.8833013857365586e-05)),(to_sfixed_a(-2.302724533365108e-05)),(to_sfixed_a(4.255978637957014e-05)),(to_sfixed_a(1.5355234381786431e-06)),(to_sfixed_a(4.8793222958920524e-05)),(to_sfixed_a(8.964016160462052e-06)),(to_sfixed_a(-3.2103068861033535e-06)),(to_sfixed_a(3.099662717431784e-05)),(to_sfixed_a(3.4353208320681006e-05)),(to_sfixed_a(-1.859907752077561e-05)),(to_sfixed_a(-6.798559297749307e-07)),(to_sfixed_a(-4.1169307223754004e-05)),(to_sfixed_a(-5.119938214193098e-05)),(to_sfixed_a(-2.368268178543076e-05)),(to_sfixed_a(-1.3371510249271523e-05)),(to_sfixed_a(-1.5790459656273015e-05)),(to_sfixed_a(-2.5036508304765448e-05)),(to_sfixed_a(0.00011238519073231146)),(to_sfixed_a(2.517052234907169e-05)),(to_sfixed_a(7.62783020036295e-05)),(to_sfixed_a(1.1894632734765764e-05)),(to_sfixed_a(1.4269297025748529e-05)),(to_sfixed_a(-7.4015138125105295e-06)),(to_sfixed_a(1.103004706237698e-05)),(to_sfixed_a(7.57331463319133e-06)),(to_sfixed_a(5.093742856843164e-06)),(to_sfixed_a(8.438845543423668e-05)),(to_sfixed_a(-4.0152597648557276e-05)),(to_sfixed_a(-5.159832653589547e-05)),(to_sfixed_a(9.443017188459635e-05)),(to_sfixed_a(-1.2750064342981204e-05)),(to_sfixed_a(-3.817294418695383e-05)),(to_sfixed_a(6.959708116482943e-05)),(to_sfixed_a(7.279652345459908e-05)),(to_sfixed_a(7.894532609498128e-05)),(to_sfixed_a(9.498254257778171e-06)),(to_sfixed_a(-5.214521297602914e-05)));

    constant weight_n1_196 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.21457096934318542)),(to_sfixed_a(0.011183719150722027)),(to_sfixed_a(0.013632369227707386)),(to_sfixed_a(-0.0037305632140487432)),(to_sfixed_a(0.01748654805123806)),(to_sfixed_a(0.008450916968286037)),(to_sfixed_a(0.017026416957378387)),(to_sfixed_a(0.02199324406683445)),(to_sfixed_a(-0.0732535719871521)),(to_sfixed_a(0.0056115020997822285)),(to_sfixed_a(0.10569917410612106)),(to_sfixed_a(-0.0015371141489595175)),(to_sfixed_a(0.06024930998682976)),(to_sfixed_a(-0.032944679260253906)),(to_sfixed_a(-0.027566900476813316)),(to_sfixed_a(-0.04465002939105034)),(to_sfixed_a(0.03724593669176102)),(to_sfixed_a(-0.008221408352255821)),(to_sfixed_a(0.031125523149967194)),(to_sfixed_a(-0.04201294854283333)),(to_sfixed_a(0.07923292368650436)),(to_sfixed_a(0.07372363656759262)),(to_sfixed_a(-0.05580293387174606)),(to_sfixed_a(-0.032330989837646484)),(to_sfixed_a(0.025303425267338753)),(to_sfixed_a(-0.039722975343465805)),(to_sfixed_a(-0.1166066825389862)),(to_sfixed_a(0.13082101941108704)),(to_sfixed_a(-0.04856221005320549)),(to_sfixed_a(-0.055592428892850876)),(to_sfixed_a(-0.07043731957674026)),(to_sfixed_a(-0.011837990954518318)),(to_sfixed_a(0.001548843109048903)),(to_sfixed_a(-0.047033146023750305)),(to_sfixed_a(0.033515531569719315)),(to_sfixed_a(-0.05174102634191513)),(to_sfixed_a(0.08203503489494324)),(to_sfixed_a(0.009549552574753761)));

    constant weight_n1_197 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.19379641115665436)),(to_sfixed_a(0.014524806290864944)),(to_sfixed_a(-0.0532015860080719)),(to_sfixed_a(0.046379804611206055)),(to_sfixed_a(0.13593007624149323)),(to_sfixed_a(0.006859967950731516)),(to_sfixed_a(0.10767962038516998)),(to_sfixed_a(-0.007371631450951099)),(to_sfixed_a(-0.1341080218553543)),(to_sfixed_a(0.017445623874664307)),(to_sfixed_a(-0.27495077252388)),(to_sfixed_a(0.07171208411455154)),(to_sfixed_a(0.14589199423789978)),(to_sfixed_a(-0.0483265183866024)),(to_sfixed_a(-0.09782557189464569)),(to_sfixed_a(0.04442322626709938)),(to_sfixed_a(-0.13401924073696136)),(to_sfixed_a(-0.154543936252594)),(to_sfixed_a(0.010908563621342182)),(to_sfixed_a(0.16335007548332214)),(to_sfixed_a(-0.06434301286935806)),(to_sfixed_a(0.031977877020835876)),(to_sfixed_a(0.16463540494441986)),(to_sfixed_a(-0.10916214436292648)),(to_sfixed_a(0.06492872536182404)),(to_sfixed_a(0.07169310748577118)),(to_sfixed_a(0.15514838695526123)),(to_sfixed_a(0.1500604748725891)),(to_sfixed_a(0.004013292491436005)),(to_sfixed_a(-0.059470899403095245)),(to_sfixed_a(-0.19600090384483337)),(to_sfixed_a(0.04146390035748482)),(to_sfixed_a(0.0014722100459039211)),(to_sfixed_a(-0.05638859421014786)),(to_sfixed_a(0.07950077950954437)),(to_sfixed_a(-0.19865459203720093)),(to_sfixed_a(0.10833361744880676)),(to_sfixed_a(-0.03295941278338432)));

    constant weight_n1_198 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.2206420600414276)),(to_sfixed_a(1.0530276085773949e-05)),(to_sfixed_a(4.158766387263313e-05)),(to_sfixed_a(-8.677745427121408e-06)),(to_sfixed_a(-9.954833330994006e-06)),(to_sfixed_a(3.5826909879688174e-05)),(to_sfixed_a(9.708654943096917e-06)),(to_sfixed_a(-3.106418080278672e-05)),(to_sfixed_a(-9.590120498614851e-06)),(to_sfixed_a(-2.3133148715714924e-05)),(to_sfixed_a(3.1279894756153226e-05)),(to_sfixed_a(-7.469094998668879e-05)),(to_sfixed_a(-7.027162791928276e-05)),(to_sfixed_a(5.799022801511455e-06)),(to_sfixed_a(4.1225870518246666e-05)),(to_sfixed_a(-8.914363570511341e-05)),(to_sfixed_a(3.2129584724316373e-05)),(to_sfixed_a(3.845108221867122e-05)),(to_sfixed_a(7.05959610058926e-05)),(to_sfixed_a(4.823960262001492e-05)),(to_sfixed_a(6.120728812675225e-06)),(to_sfixed_a(4.336009078542702e-05)),(to_sfixed_a(-6.320526881609112e-05)),(to_sfixed_a(2.9409689886961132e-05)),(to_sfixed_a(-8.067127782851458e-05)),(to_sfixed_a(5.0369468226563185e-05)),(to_sfixed_a(4.337666177889332e-05)),(to_sfixed_a(1.6279086594295222e-06)),(to_sfixed_a(2.026643414865248e-05)),(to_sfixed_a(-0.00012162020721007138)),(to_sfixed_a(7.44345088605769e-05)),(to_sfixed_a(-5.480261825141497e-05)),(to_sfixed_a(-1.339748087048065e-05)),(to_sfixed_a(-7.194506179075688e-05)),(to_sfixed_a(-6.0893911722814664e-05)),(to_sfixed_a(6.314808706520125e-05)),(to_sfixed_a(-5.099431655253284e-05)),(to_sfixed_a(3.4651522582862526e-05)));

    constant weight_n1_199 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.02769593894481659)),(to_sfixed_a(6.0222828324185684e-06)),(to_sfixed_a(-5.9034071455243975e-05)),(to_sfixed_a(4.1661711293272674e-05)),(to_sfixed_a(-4.119750883546658e-05)),(to_sfixed_a(1.7353571820422076e-05)),(to_sfixed_a(-1.5255328435159754e-05)),(to_sfixed_a(4.5263743231771514e-05)),(to_sfixed_a(-6.47285851300694e-05)),(to_sfixed_a(-4.9461614253232256e-05)),(to_sfixed_a(2.4393695639446378e-05)),(to_sfixed_a(-2.7655260055325925e-05)),(to_sfixed_a(4.4835695007350296e-05)),(to_sfixed_a(1.0118948011950124e-05)),(to_sfixed_a(-4.568359872791916e-05)),(to_sfixed_a(-1.1795547834481113e-05)),(to_sfixed_a(-8.343037188751623e-05)),(to_sfixed_a(-2.950189809780568e-05)),(to_sfixed_a(0.00010192307672696188)),(to_sfixed_a(-1.2128683920309413e-05)),(to_sfixed_a(8.748308755457401e-05)),(to_sfixed_a(2.046089866780676e-05)),(to_sfixed_a(0.00010695951641537249)),(to_sfixed_a(-4.964762047166005e-05)),(to_sfixed_a(-2.697303716558963e-05)),(to_sfixed_a(2.5475337679381482e-05)),(to_sfixed_a(-5.1553270168369636e-05)),(to_sfixed_a(1.6225500075961463e-05)),(to_sfixed_a(4.835708296013763e-06)),(to_sfixed_a(6.078867590986192e-05)),(to_sfixed_a(1.028435963235097e-05)),(to_sfixed_a(2.739492447290104e-05)),(to_sfixed_a(2.022442640736699e-05)),(to_sfixed_a(5.2864426834275946e-05)),(to_sfixed_a(-1.1810174328275025e-05)),(to_sfixed_a(2.7929385396419093e-05)),(to_sfixed_a(3.3044092560885474e-05)),(to_sfixed_a(1.1453374099801295e-05)));

    constant weight_n1_200 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.038346707820892334)),(to_sfixed_a(-1.577644252392929e-05)),(to_sfixed_a(-3.079499947489239e-05)),(to_sfixed_a(-1.011627864500042e-05)),(to_sfixed_a(-3.811539863818325e-05)),(to_sfixed_a(7.4182721618853975e-06)),(to_sfixed_a(2.615258017613087e-05)),(to_sfixed_a(-0.00010034939623437822)),(to_sfixed_a(-2.159517134714406e-05)),(to_sfixed_a(-4.92506933369441e-06)),(to_sfixed_a(-1.3612422662845347e-05)),(to_sfixed_a(2.143699566659052e-05)),(to_sfixed_a(-2.0032866814290173e-05)),(to_sfixed_a(-4.095722397323698e-05)),(to_sfixed_a(1.2683372005994897e-05)),(to_sfixed_a(-8.232083928305656e-05)),(to_sfixed_a(3.2653821108397096e-05)),(to_sfixed_a(3.0420400435104966e-05)),(to_sfixed_a(-1.8756692952592857e-05)),(to_sfixed_a(1.1284657375654206e-05)),(to_sfixed_a(2.7002704882761464e-05)),(to_sfixed_a(-1.7729204046190716e-05)),(to_sfixed_a(-0.00011042261030524969)),(to_sfixed_a(8.967489702627063e-05)),(to_sfixed_a(-3.7502341001527384e-05)),(to_sfixed_a(-3.108487726422027e-05)),(to_sfixed_a(3.442259912844747e-05)),(to_sfixed_a(-5.7750236010178924e-05)),(to_sfixed_a(8.459446689812467e-06)),(to_sfixed_a(1.7829436274041655e-06)),(to_sfixed_a(2.8342923542368226e-05)),(to_sfixed_a(5.717492240364663e-05)),(to_sfixed_a(7.654472574358806e-05)),(to_sfixed_a(-5.112470535095781e-05)),(to_sfixed_a(-5.150052857061382e-06)),(to_sfixed_a(6.116361328167841e-05)),(to_sfixed_a(1.4185272448230535e-05)),(to_sfixed_a(4.212004569126293e-05)));

    constant weight_n1_201 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.008721090853214264)),(to_sfixed_a(-2.1410804038168862e-05)),(to_sfixed_a(2.0330682673375122e-05)),(to_sfixed_a(-4.628606984624639e-05)),(to_sfixed_a(2.1352687326725572e-05)),(to_sfixed_a(-3.564562211977318e-05)),(to_sfixed_a(2.2164799702295568e-06)),(to_sfixed_a(-3.596020906115882e-05)),(to_sfixed_a(-5.7906868278223556e-06)),(to_sfixed_a(9.963930097001139e-06)),(to_sfixed_a(7.5085399657837115e-06)),(to_sfixed_a(2.3105447326088324e-05)),(to_sfixed_a(8.253319538198411e-05)),(to_sfixed_a(3.139883847325109e-05)),(to_sfixed_a(3.0154356863931753e-05)),(to_sfixed_a(-1.0085325811814982e-05)),(to_sfixed_a(-1.0512412700336426e-05)),(to_sfixed_a(-3.137060775770806e-05)),(to_sfixed_a(4.4844846343039535e-06)),(to_sfixed_a(-6.614547601202503e-05)),(to_sfixed_a(1.856671406130772e-05)),(to_sfixed_a(-3.365042357472703e-05)),(to_sfixed_a(7.475964957848191e-05)),(to_sfixed_a(3.434727113926783e-05)),(to_sfixed_a(3.2417450711363927e-05)),(to_sfixed_a(-5.187502029002644e-05)),(to_sfixed_a(-9.983243944589049e-05)),(to_sfixed_a(3.66852073057089e-05)),(to_sfixed_a(-2.1088826542836614e-05)),(to_sfixed_a(2.5991905204136856e-05)),(to_sfixed_a(-4.547846765490249e-05)),(to_sfixed_a(2.8958971597603522e-05)),(to_sfixed_a(8.481930854031816e-05)),(to_sfixed_a(-9.934563422575593e-05)),(to_sfixed_a(-4.813854320673272e-05)),(to_sfixed_a(-7.179927342804149e-05)),(to_sfixed_a(-7.04226185916923e-05)),(to_sfixed_a(8.084192813839763e-05)));

    constant weight_n1_202 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.013494838960468769)),(to_sfixed_a(-1.833812530094292e-05)),(to_sfixed_a(-1.1581069884414319e-05)),(to_sfixed_a(-4.134741175221279e-06)),(to_sfixed_a(2.4879367629182525e-05)),(to_sfixed_a(8.466233339277096e-06)),(to_sfixed_a(-3.478460348560475e-05)),(to_sfixed_a(-3.601459684432484e-05)),(to_sfixed_a(1.2990247341804206e-05)),(to_sfixed_a(-5.2667586714960635e-05)),(to_sfixed_a(-1.6921076166909188e-06)),(to_sfixed_a(-2.116727046086453e-05)),(to_sfixed_a(2.775044231384527e-05)),(to_sfixed_a(9.429321607967722e-07)),(to_sfixed_a(-5.497056554304436e-05)),(to_sfixed_a(7.856349111534655e-05)),(to_sfixed_a(-3.0438468456850387e-06)),(to_sfixed_a(6.930331437615678e-05)),(to_sfixed_a(6.5718348196242e-05)),(to_sfixed_a(5.821180820930749e-05)),(to_sfixed_a(7.482136425096542e-06)),(to_sfixed_a(1.3608821973321028e-05)),(to_sfixed_a(0.00010738275886978954)),(to_sfixed_a(1.8947455828310922e-05)),(to_sfixed_a(-1.6237416275544092e-05)),(to_sfixed_a(-4.310806980356574e-05)),(to_sfixed_a(6.543709605466574e-05)),(to_sfixed_a(5.8973528211936355e-05)),(to_sfixed_a(-6.657005724264309e-05)),(to_sfixed_a(-3.7149209674680606e-05)),(to_sfixed_a(-8.540104317944497e-06)),(to_sfixed_a(3.8210488128243014e-05)),(to_sfixed_a(-6.028883217368275e-05)),(to_sfixed_a(-2.407461215625517e-05)),(to_sfixed_a(0.0001041982977767475)),(to_sfixed_a(4.7691090003354475e-05)),(to_sfixed_a(7.468505828001071e-06)),(to_sfixed_a(-2.9475815608748235e-05)));

    constant weight_n1_203 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.014930598437786102)),(to_sfixed_a(-2.6936524591292255e-05)),(to_sfixed_a(5.1759583584498614e-05)),(to_sfixed_a(4.249957783031277e-06)),(to_sfixed_a(-1.3897791177441832e-05)),(to_sfixed_a(2.586303889984265e-05)),(to_sfixed_a(3.403036680538207e-05)),(to_sfixed_a(-8.925877409637906e-06)),(to_sfixed_a(-1.780162529030349e-05)),(to_sfixed_a(-2.100456003972795e-05)),(to_sfixed_a(-1.760196391842328e-05)),(to_sfixed_a(-7.93837352830451e-06)),(to_sfixed_a(7.24462661310099e-05)),(to_sfixed_a(-1.1500663958941004e-06)),(to_sfixed_a(-2.8350765205686912e-05)),(to_sfixed_a(-3.976880543632433e-05)),(to_sfixed_a(-3.791590279433876e-05)),(to_sfixed_a(-2.469388891768176e-05)),(to_sfixed_a(-2.8460792691475945e-06)),(to_sfixed_a(3.3477374472568044e-06)),(to_sfixed_a(3.233809184166603e-05)),(to_sfixed_a(-9.256966222892515e-06)),(to_sfixed_a(9.397772373631597e-06)),(to_sfixed_a(-1.726528353174217e-05)),(to_sfixed_a(-1.1414116670493968e-05)),(to_sfixed_a(3.8065454077695904e-07)),(to_sfixed_a(5.880732715013437e-05)),(to_sfixed_a(-3.336276859045029e-05)),(to_sfixed_a(-2.455477078910917e-05)),(to_sfixed_a(4.285381510271691e-05)),(to_sfixed_a(6.774851499358192e-05)),(to_sfixed_a(-2.7757805582950823e-05)),(to_sfixed_a(-5.6836088333511725e-05)),(to_sfixed_a(5.812910239910707e-05)),(to_sfixed_a(3.844561433652416e-05)),(to_sfixed_a(-6.004537863191217e-05)),(to_sfixed_a(5.880484604858793e-05)),(to_sfixed_a(4.101674858247861e-05)));

    constant weight_n1_204 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.11022815108299255)),(to_sfixed_a(0.009105628356337547)),(to_sfixed_a(-0.045192018151283264)),(to_sfixed_a(-0.03140706196427345)),(to_sfixed_a(-0.027815010398626328)),(to_sfixed_a(0.08727619051933289)),(to_sfixed_a(-0.028526687994599342)),(to_sfixed_a(0.066260926425457)),(to_sfixed_a(0.0017698591109365225)),(to_sfixed_a(-0.014061657711863518)),(to_sfixed_a(-0.03609084337949753)),(to_sfixed_a(0.014975575730204582)),(to_sfixed_a(0.07193756103515625)),(to_sfixed_a(0.032285988330841064)),(to_sfixed_a(-0.03211985155940056)),(to_sfixed_a(0.060681745409965515)),(to_sfixed_a(-0.038015078753232956)),(to_sfixed_a(-0.026104923337697983)),(to_sfixed_a(0.013761257752776146)),(to_sfixed_a(0.006545437965542078)),(to_sfixed_a(-0.03459296375513077)),(to_sfixed_a(-0.019469689577817917)),(to_sfixed_a(0.052043113857507706)),(to_sfixed_a(-0.005727572366595268)),(to_sfixed_a(0.005260365083813667)),(to_sfixed_a(-0.0515422560274601)),(to_sfixed_a(0.07786767929792404)),(to_sfixed_a(-0.022138196974992752)),(to_sfixed_a(-0.02146172523498535)),(to_sfixed_a(-0.07644744217395782)),(to_sfixed_a(-0.006994947325438261)),(to_sfixed_a(-0.04594938084483147)),(to_sfixed_a(-0.05124069005250931)),(to_sfixed_a(0.004602791275829077)),(to_sfixed_a(-0.004525929689407349)),(to_sfixed_a(-0.01986095868051052)),(to_sfixed_a(-0.04284023866057396)),(to_sfixed_a(0.00917670875787735)));

    constant weight_n1_205 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.1438216269016266)),(to_sfixed_a(0.22852616012096405)),(to_sfixed_a(0.04464361444115639)),(to_sfixed_a(0.15599140524864197)),(to_sfixed_a(-0.02524249441921711)),(to_sfixed_a(-0.04309559613466263)),(to_sfixed_a(0.2792976498603821)),(to_sfixed_a(-0.07643464207649231)),(to_sfixed_a(0.0003144429065287113)),(to_sfixed_a(-0.16426195204257965)),(to_sfixed_a(-0.048804473131895065)),(to_sfixed_a(0.01795388199388981)),(to_sfixed_a(-0.005939483642578125)),(to_sfixed_a(-0.056866176426410675)),(to_sfixed_a(0.15088306367397308)),(to_sfixed_a(-0.07561343908309937)),(to_sfixed_a(0.03973279893398285)),(to_sfixed_a(-0.07600148022174835)),(to_sfixed_a(-0.04123421385884285)),(to_sfixed_a(0.010321712121367455)),(to_sfixed_a(0.0019941406790167093)),(to_sfixed_a(-0.02635667286813259)),(to_sfixed_a(0.006482867524027824)),(to_sfixed_a(0.1332933008670807)),(to_sfixed_a(0.08172816783189774)),(to_sfixed_a(0.0037361846771091223)),(to_sfixed_a(-0.11683441698551178)),(to_sfixed_a(0.008490212261676788)),(to_sfixed_a(-0.04276883229613304)),(to_sfixed_a(0.047003958374261856)),(to_sfixed_a(0.13347183167934418)),(to_sfixed_a(0.0703062117099762)),(to_sfixed_a(-0.019231270998716354)),(to_sfixed_a(-0.09534415602684021)),(to_sfixed_a(-0.10990116745233536)),(to_sfixed_a(0.02653450332581997)),(to_sfixed_a(-0.05371421203017235)),(to_sfixed_a(-0.1434391885995865)));

    constant weight_n1_206 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.05072036758065224)),(to_sfixed_a(0.0686199814081192)),(to_sfixed_a(-0.1081402599811554)),(to_sfixed_a(0.04623199626803398)),(to_sfixed_a(0.025818636640906334)),(to_sfixed_a(-0.013241074047982693)),(to_sfixed_a(-0.015693819150328636)),(to_sfixed_a(-0.01960272528231144)),(to_sfixed_a(-0.031300805509090424)),(to_sfixed_a(0.10917089879512787)),(to_sfixed_a(0.02941099740564823)),(to_sfixed_a(0.15112775564193726)),(to_sfixed_a(-0.24171268939971924)),(to_sfixed_a(-0.05371762812137604)),(to_sfixed_a(0.05018133297562599)),(to_sfixed_a(-0.20712168514728546)),(to_sfixed_a(-0.25197720527648926)),(to_sfixed_a(0.24597738683223724)),(to_sfixed_a(0.18013525009155273)),(to_sfixed_a(0.08233215659856796)),(to_sfixed_a(0.041462503373622894)),(to_sfixed_a(-0.06430928409099579)),(to_sfixed_a(0.2616332769393921)),(to_sfixed_a(-0.017292017117142677)),(to_sfixed_a(-0.16703063249588013)),(to_sfixed_a(-0.1902473419904709)),(to_sfixed_a(-0.0653783529996872)),(to_sfixed_a(-0.1469212770462036)),(to_sfixed_a(0.10171516984701157)),(to_sfixed_a(-0.061646830290555954)),(to_sfixed_a(0.17835070192813873)),(to_sfixed_a(0.1069486141204834)),(to_sfixed_a(0.06717546284198761)),(to_sfixed_a(0.10657145082950592)),(to_sfixed_a(-0.13309715688228607)),(to_sfixed_a(0.011557353660464287)),(to_sfixed_a(-0.14474627375602722)),(to_sfixed_a(0.04701182246208191)));

    constant weight_n1_207 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.0012979559833183885)),(to_sfixed_a(0.011879668571054935)),(to_sfixed_a(-0.056600846350193024)),(to_sfixed_a(-0.11235130578279495)),(to_sfixed_a(-0.048520009964704514)),(to_sfixed_a(0.023203223943710327)),(to_sfixed_a(0.011342394165694714)),(to_sfixed_a(-0.033724345266819)),(to_sfixed_a(-0.05106232315301895)),(to_sfixed_a(0.03158823400735855)),(to_sfixed_a(0.03353795409202576)),(to_sfixed_a(-0.021700752899050713)),(to_sfixed_a(0.00514902314171195)),(to_sfixed_a(-0.05197978764772415)),(to_sfixed_a(0.038922663778066635)),(to_sfixed_a(-0.04911862313747406)),(to_sfixed_a(0.01041687373071909)),(to_sfixed_a(-0.019658032804727554)),(to_sfixed_a(0.0822867676615715)),(to_sfixed_a(0.06960189342498779)),(to_sfixed_a(-0.04764287918806076)),(to_sfixed_a(0.01207976695150137)),(to_sfixed_a(0.01602071337401867)),(to_sfixed_a(0.004979231394827366)),(to_sfixed_a(-0.08379244804382324)),(to_sfixed_a(-0.06336676329374313)),(to_sfixed_a(0.005118648987263441)),(to_sfixed_a(-0.018032187595963478)),(to_sfixed_a(0.07117060571908951)),(to_sfixed_a(0.12314695119857788)),(to_sfixed_a(0.013309899717569351)),(to_sfixed_a(0.021875392645597458)),(to_sfixed_a(-0.06872754544019699)),(to_sfixed_a(-0.026040835306048393)),(to_sfixed_a(0.011896241456270218)),(to_sfixed_a(0.025357460603117943)),(to_sfixed_a(0.01673145405948162)),(to_sfixed_a(0.01955467276275158)));

    constant weight_n1_208 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.1522538959980011)),(to_sfixed_a(-0.03466123715043068)),(to_sfixed_a(0.02679366059601307)),(to_sfixed_a(-0.09675215184688568)),(to_sfixed_a(-0.02141229808330536)),(to_sfixed_a(0.08553396910429001)),(to_sfixed_a(0.05668463185429573)),(to_sfixed_a(0.03577178716659546)),(to_sfixed_a(0.009255881421267986)),(to_sfixed_a(-0.04747674614191055)),(to_sfixed_a(0.048887789249420166)),(to_sfixed_a(-0.09266746044158936)),(to_sfixed_a(0.053481776267290115)),(to_sfixed_a(-0.027525687590241432)),(to_sfixed_a(0.05067300796508789)),(to_sfixed_a(0.06499343365430832)),(to_sfixed_a(0.10434851795434952)),(to_sfixed_a(0.04299656301736832)),(to_sfixed_a(-0.04232749715447426)),(to_sfixed_a(0.041349004954099655)),(to_sfixed_a(-0.1549915075302124)),(to_sfixed_a(-0.03685867413878441)),(to_sfixed_a(-0.014479754492640495)),(to_sfixed_a(0.040555499494075775)),(to_sfixed_a(-0.03135906532406807)),(to_sfixed_a(-0.08394459635019302)),(to_sfixed_a(0.017046838998794556)),(to_sfixed_a(-0.0019481773488223553)),(to_sfixed_a(0.07701302319765091)),(to_sfixed_a(0.03278278931975365)),(to_sfixed_a(0.10587043315172195)),(to_sfixed_a(0.05251232534646988)),(to_sfixed_a(0.027935001999139786)),(to_sfixed_a(-0.01576226018369198)),(to_sfixed_a(-0.08865660429000854)),(to_sfixed_a(-0.0605052150785923)),(to_sfixed_a(-0.001452879747375846)),(to_sfixed_a(0.05547986179590225)));

    constant weight_n1_209 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.031527724117040634)),(to_sfixed_a(-0.0007836144068278372)),(to_sfixed_a(-0.029713157564401627)),(to_sfixed_a(-0.04050597548484802)),(to_sfixed_a(-0.023013344034552574)),(to_sfixed_a(-0.002215868793427944)),(to_sfixed_a(0.006344348657876253)),(to_sfixed_a(-0.06857292354106903)),(to_sfixed_a(0.0347907729446888)),(to_sfixed_a(0.08825651556253433)),(to_sfixed_a(0.10086033493280411)),(to_sfixed_a(0.035490792244672775)),(to_sfixed_a(0.058176133781671524)),(to_sfixed_a(0.07948235422372818)),(to_sfixed_a(0.021262217313051224)),(to_sfixed_a(0.06427406519651413)),(to_sfixed_a(-0.029886487871408463)),(to_sfixed_a(-0.033032938838005066)),(to_sfixed_a(0.07578334957361221)),(to_sfixed_a(0.030050938948988914)),(to_sfixed_a(0.1016412153840065)),(to_sfixed_a(0.00552000617608428)),(to_sfixed_a(0.12414468824863434)),(to_sfixed_a(0.0007996258791536093)),(to_sfixed_a(0.08847958594560623)),(to_sfixed_a(0.06341221928596497)),(to_sfixed_a(0.01459964457899332)),(to_sfixed_a(0.016246018931269646)),(to_sfixed_a(-0.049296364188194275)),(to_sfixed_a(-0.0036991655360907316)),(to_sfixed_a(0.013347143307328224)),(to_sfixed_a(0.1802169382572174)),(to_sfixed_a(-0.03047524392604828)),(to_sfixed_a(-0.1543918401002884)),(to_sfixed_a(-0.07601594179868698)),(to_sfixed_a(-0.09312011301517487)),(to_sfixed_a(0.19835343956947327)),(to_sfixed_a(0.0018465286120772362)));

    constant weight_n1_210 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.007964972406625748)),(to_sfixed_a(-4.817503213416785e-05)),(to_sfixed_a(-1.2453607268980704e-05)),(to_sfixed_a(9.110014502766717e-07)),(to_sfixed_a(-3.6982601159252226e-05)),(to_sfixed_a(5.140521898283623e-05)),(to_sfixed_a(-5.088310717837885e-05)),(to_sfixed_a(4.971989619662054e-05)),(to_sfixed_a(2.0304922145442106e-05)),(to_sfixed_a(-9.806452681004885e-07)),(to_sfixed_a(1.0269268386764452e-05)),(to_sfixed_a(-7.791045391059015e-07)),(to_sfixed_a(2.4266815671580844e-05)),(to_sfixed_a(-1.8718294086284004e-05)),(to_sfixed_a(4.6981655032141134e-05)),(to_sfixed_a(-4.6220680815167725e-05)),(to_sfixed_a(2.2555599571205676e-05)),(to_sfixed_a(-2.5285937226726674e-05)),(to_sfixed_a(2.700195409488515e-06)),(to_sfixed_a(3.574359288904816e-05)),(to_sfixed_a(-9.34558738663327e-06)),(to_sfixed_a(-1.1037568583560642e-05)),(to_sfixed_a(-2.0085044525330886e-05)),(to_sfixed_a(-1.1808927411038894e-05)),(to_sfixed_a(-1.0246309102512896e-05)),(to_sfixed_a(-3.747127720998833e-06)),(to_sfixed_a(-2.4493941964465193e-05)),(to_sfixed_a(7.700813875999302e-05)),(to_sfixed_a(-2.3234879336087033e-05)),(to_sfixed_a(-1.3162796676624566e-05)),(to_sfixed_a(-5.345609679352492e-06)),(to_sfixed_a(1.8061566152027808e-05)),(to_sfixed_a(1.7183996533276513e-05)),(to_sfixed_a(3.434472455410287e-05)),(to_sfixed_a(-7.147745054680854e-05)),(to_sfixed_a(-3.3435397199355066e-05)),(to_sfixed_a(-7.875408482505009e-05)),(to_sfixed_a(-7.353541150223464e-05)));

    constant weight_n1_211 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.01362223457545042)),(to_sfixed_a(-2.9281729439389892e-05)),(to_sfixed_a(-1.758708276611287e-05)),(to_sfixed_a(4.599680323735811e-05)),(to_sfixed_a(-2.4498078801116208e-06)),(to_sfixed_a(-7.854446266719606e-06)),(to_sfixed_a(-9.052661908981463e-08)),(to_sfixed_a(1.0093035598401912e-05)),(to_sfixed_a(2.2161006199894473e-05)),(to_sfixed_a(-1.4808771084062755e-05)),(to_sfixed_a(4.501229398101714e-07)),(to_sfixed_a(6.971219136175932e-06)),(to_sfixed_a(8.181042176147457e-06)),(to_sfixed_a(-1.1671060747175943e-05)),(to_sfixed_a(-7.959495269460604e-05)),(to_sfixed_a(-5.8215282479068264e-05)),(to_sfixed_a(-7.602365803904831e-05)),(to_sfixed_a(4.8170812078751624e-05)),(to_sfixed_a(-1.5404553778353147e-05)),(to_sfixed_a(3.1485844374401495e-05)),(to_sfixed_a(4.898455154034309e-05)),(to_sfixed_a(-2.9329023163882084e-05)),(to_sfixed_a(-3.2390122214565054e-05)),(to_sfixed_a(4.7470575736952014e-06)),(to_sfixed_a(-8.407768291363027e-06)),(to_sfixed_a(3.9773862226866186e-05)),(to_sfixed_a(-8.181657904060557e-06)),(to_sfixed_a(4.05885475629475e-05)),(to_sfixed_a(-5.442331894300878e-05)),(to_sfixed_a(-8.176529809134081e-05)),(to_sfixed_a(1.6664038184899255e-06)),(to_sfixed_a(1.592505032022018e-05)),(to_sfixed_a(4.822608389076777e-05)),(to_sfixed_a(-2.15228610613849e-05)),(to_sfixed_a(1.8552727851783857e-05)),(to_sfixed_a(2.274379221489653e-05)),(to_sfixed_a(0.0001152868353528902)),(to_sfixed_a(-2.5982795705203898e-05)));

    constant weight_n1_212 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.009712628088891506)),(to_sfixed_a(-1.6168585716513917e-05)),(to_sfixed_a(4.111391899641603e-05)),(to_sfixed_a(-1.5197811990219634e-05)),(to_sfixed_a(-2.6509856979828328e-05)),(to_sfixed_a(2.9933489713585004e-05)),(to_sfixed_a(-2.613945434859488e-05)),(to_sfixed_a(-2.5968272893805988e-05)),(to_sfixed_a(-1.7338288671453483e-05)),(to_sfixed_a(-1.9698951291502453e-05)),(to_sfixed_a(6.984972515056143e-06)),(to_sfixed_a(4.247646211297251e-05)),(to_sfixed_a(1.5780733519932255e-05)),(to_sfixed_a(-2.4885406674002297e-05)),(to_sfixed_a(-4.132893081987277e-05)),(to_sfixed_a(-7.120676309568807e-05)),(to_sfixed_a(-3.262732207076624e-06)),(to_sfixed_a(-7.700589048909023e-05)),(to_sfixed_a(3.174923040205613e-05)),(to_sfixed_a(-7.172826735768467e-05)),(to_sfixed_a(4.7381679905811325e-05)),(to_sfixed_a(-4.0746101149125025e-05)),(to_sfixed_a(2.2344025637721643e-05)),(to_sfixed_a(3.1729156034998596e-05)),(to_sfixed_a(-1.9033526768907905e-05)),(to_sfixed_a(-4.635851291823201e-05)),(to_sfixed_a(-8.515476110915188e-06)),(to_sfixed_a(-2.4759809093666263e-05)),(to_sfixed_a(3.705786730279215e-05)),(to_sfixed_a(-5.185025656828657e-06)),(to_sfixed_a(-2.0709117961814627e-05)),(to_sfixed_a(1.6784086255938746e-05)),(to_sfixed_a(-7.455280137946829e-05)),(to_sfixed_a(-2.701585071918089e-05)),(to_sfixed_a(7.586064020870253e-05)),(to_sfixed_a(-8.162779704434797e-05)),(to_sfixed_a(7.144287337723654e-06)),(to_sfixed_a(8.378833445021883e-05)));

    constant weight_n1_213 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.06799939274787903)),(to_sfixed_a(4.31770968134515e-05)),(to_sfixed_a(-7.984826879692264e-06)),(to_sfixed_a(-6.553561252076179e-05)),(to_sfixed_a(-9.256448720407207e-06)),(to_sfixed_a(-2.5214205379597843e-05)),(to_sfixed_a(1.1801708751590922e-05)),(to_sfixed_a(-3.968278178945184e-05)),(to_sfixed_a(2.507460885681212e-05)),(to_sfixed_a(-4.50535626441706e-05)),(to_sfixed_a(6.364547880366445e-05)),(to_sfixed_a(-2.635139026097022e-05)),(to_sfixed_a(1.0099552127940115e-05)),(to_sfixed_a(5.594473350356566e-06)),(to_sfixed_a(3.7029636587249115e-05)),(to_sfixed_a(-3.516108336043544e-05)),(to_sfixed_a(1.245692965312628e-05)),(to_sfixed_a(6.584564835065976e-05)),(to_sfixed_a(3.0523038731189445e-05)),(to_sfixed_a(8.477393566863611e-05)),(to_sfixed_a(3.781026680371724e-05)),(to_sfixed_a(-1.7404014215571806e-05)),(to_sfixed_a(-2.6494810299482197e-05)),(to_sfixed_a(-8.234155757236294e-06)),(to_sfixed_a(7.262563303811476e-05)),(to_sfixed_a(-2.5082455977099016e-05)),(to_sfixed_a(7.127815479179844e-05)),(to_sfixed_a(-2.140043579856865e-05)),(to_sfixed_a(-2.1305586415110156e-05)),(to_sfixed_a(-1.5974854250089265e-05)),(to_sfixed_a(-2.812517595884856e-05)),(to_sfixed_a(3.957810258725658e-05)),(to_sfixed_a(4.989178341929801e-05)),(to_sfixed_a(-3.7892422710683604e-07)),(to_sfixed_a(6.557808956131339e-05)),(to_sfixed_a(-5.300230623106472e-05)),(to_sfixed_a(-2.5358433504152345e-06)),(to_sfixed_a(-6.957650384720182e-06)));

    constant weight_n1_214 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.023451078683137894)),(to_sfixed_a(1.5233455087582115e-05)),(to_sfixed_a(-7.792425458319485e-05)),(to_sfixed_a(-3.448241113801487e-05)),(to_sfixed_a(5.976506508886814e-05)),(to_sfixed_a(4.816798900719732e-05)),(to_sfixed_a(2.9221486329333857e-05)),(to_sfixed_a(1.723964487609919e-05)),(to_sfixed_a(5.51893244846724e-05)),(to_sfixed_a(8.384851389564574e-05)),(to_sfixed_a(-0.00010090740397572517)),(to_sfixed_a(1.619185695744818e-06)),(to_sfixed_a(2.3418777345796116e-05)),(to_sfixed_a(1.8274733520229347e-05)),(to_sfixed_a(2.828739889082499e-05)),(to_sfixed_a(-5.545942622120492e-05)),(to_sfixed_a(1.0872989150811918e-05)),(to_sfixed_a(-4.8041616537375376e-05)),(to_sfixed_a(1.3547729395213537e-05)),(to_sfixed_a(-8.398180943913758e-05)),(to_sfixed_a(1.1121455827378668e-05)),(to_sfixed_a(-3.5316439607413486e-05)),(to_sfixed_a(-6.730821041855961e-05)),(to_sfixed_a(1.7323663996648975e-05)),(to_sfixed_a(-1.1864523912663572e-05)),(to_sfixed_a(7.202534470707178e-05)),(to_sfixed_a(-1.3562477761297487e-05)),(to_sfixed_a(-5.46670489711687e-05)),(to_sfixed_a(4.9008427595254034e-05)),(to_sfixed_a(5.428555959952064e-05)),(to_sfixed_a(-6.593627404072322e-06)),(to_sfixed_a(-0.000126450730022043)),(to_sfixed_a(5.883779522264376e-06)),(to_sfixed_a(2.105837302224245e-05)),(to_sfixed_a(2.2882331904838793e-05)),(to_sfixed_a(-8.125887688947842e-06)),(to_sfixed_a(-6.121245678514242e-05)),(to_sfixed_a(1.2875336324214004e-05)));

    constant weight_n1_215 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.17339305579662323)),(to_sfixed_a(-0.01857994869351387)),(to_sfixed_a(0.010145802982151508)),(to_sfixed_a(0.027469199150800705)),(to_sfixed_a(-0.02143871784210205)),(to_sfixed_a(-0.02668570727109909)),(to_sfixed_a(0.006957967299968004)),(to_sfixed_a(-0.00019275544036645442)),(to_sfixed_a(0.019589992240071297)),(to_sfixed_a(0.04858004301786423)),(to_sfixed_a(0.012760939076542854)),(to_sfixed_a(-0.058588478714227676)),(to_sfixed_a(0.03907286375761032)),(to_sfixed_a(-0.032162293791770935)),(to_sfixed_a(0.00627486826851964)),(to_sfixed_a(-0.007379953283816576)),(to_sfixed_a(0.026675721630454063)),(to_sfixed_a(0.02237767167389393)),(to_sfixed_a(0.02011062018573284)),(to_sfixed_a(0.031225908547639847)),(to_sfixed_a(-0.010779635980725288)),(to_sfixed_a(-0.014602511189877987)),(to_sfixed_a(0.030408577993512154)),(to_sfixed_a(0.00337641267105937)),(to_sfixed_a(-0.053889594972133636)),(to_sfixed_a(0.00766875222325325)),(to_sfixed_a(0.008992601186037064)),(to_sfixed_a(0.02440517395734787)),(to_sfixed_a(-0.02930198796093464)),(to_sfixed_a(-0.023026777431368828)),(to_sfixed_a(0.002836410654708743)),(to_sfixed_a(0.04509880021214485)),(to_sfixed_a(0.009245914407074451)),(to_sfixed_a(-0.058318208903074265)),(to_sfixed_a(0.028224801644682884)),(to_sfixed_a(0.01739727333188057)),(to_sfixed_a(-0.034995194524526596)),(to_sfixed_a(0.03278268128633499)));

    constant weight_n1_216 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.027849331498146057)),(to_sfixed_a(0.041541147977113724)),(to_sfixed_a(-0.047833576798439026)),(to_sfixed_a(0.014949711970984936)),(to_sfixed_a(0.024246908724308014)),(to_sfixed_a(0.046348635107278824)),(to_sfixed_a(0.03980468213558197)),(to_sfixed_a(0.11728359758853912)),(to_sfixed_a(0.06837787479162216)),(to_sfixed_a(0.043042633682489395)),(to_sfixed_a(0.069705531001091)),(to_sfixed_a(0.031029395759105682)),(to_sfixed_a(-0.03463508561253548)),(to_sfixed_a(-0.07554863393306732)),(to_sfixed_a(0.05481014773249626)),(to_sfixed_a(0.039185650646686554)),(to_sfixed_a(0.03810657933354378)),(to_sfixed_a(-0.0786927193403244)),(to_sfixed_a(0.02693050540983677)),(to_sfixed_a(0.10774223506450653)),(to_sfixed_a(0.07684880495071411)),(to_sfixed_a(-0.03490881621837616)),(to_sfixed_a(-0.043307140469551086)),(to_sfixed_a(-0.012101937085390091)),(to_sfixed_a(-0.039422258734703064)),(to_sfixed_a(-0.09009438008069992)),(to_sfixed_a(-0.08113371580839157)),(to_sfixed_a(0.0016966803232207894)),(to_sfixed_a(-0.015629485249519348)),(to_sfixed_a(0.0976094901561737)),(to_sfixed_a(-0.08896099776029587)),(to_sfixed_a(0.01915903016924858)),(to_sfixed_a(0.1318979412317276)),(to_sfixed_a(-0.009177871979773045)),(to_sfixed_a(-0.12839096784591675)),(to_sfixed_a(-0.15174539387226105)),(to_sfixed_a(0.04749132692813873)),(to_sfixed_a(0.07576978206634521)));

    constant weight_n1_217 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.12548571825027466)),(to_sfixed_a(-0.09461696445941925)),(to_sfixed_a(0.024620525538921356)),(to_sfixed_a(-0.07873321324586868)),(to_sfixed_a(-0.01964803971350193)),(to_sfixed_a(0.08826438337564468)),(to_sfixed_a(0.09023820608854294)),(to_sfixed_a(-0.08619877696037292)),(to_sfixed_a(0.027748815715312958)),(to_sfixed_a(0.038580745458602905)),(to_sfixed_a(-0.032533738762140274)),(to_sfixed_a(-0.12536582350730896)),(to_sfixed_a(0.17509396374225616)),(to_sfixed_a(-0.007871502079069614)),(to_sfixed_a(0.028604086488485336)),(to_sfixed_a(0.08105115592479706)),(to_sfixed_a(-0.06587103009223938)),(to_sfixed_a(0.1245507225394249)),(to_sfixed_a(0.0877179279923439)),(to_sfixed_a(0.026941001415252686)),(to_sfixed_a(0.05966639518737793)),(to_sfixed_a(-0.27184322476387024)),(to_sfixed_a(-0.000757141737267375)),(to_sfixed_a(0.05139642953872681)),(to_sfixed_a(-0.035206105560064316)),(to_sfixed_a(0.09256388992071152)),(to_sfixed_a(-0.02339892089366913)),(to_sfixed_a(-0.15574952960014343)),(to_sfixed_a(0.03189171105623245)),(to_sfixed_a(0.04855061322450638)),(to_sfixed_a(-0.0905323177576065)),(to_sfixed_a(0.08477601408958435)),(to_sfixed_a(0.10435938835144043)),(to_sfixed_a(0.02089480124413967)),(to_sfixed_a(0.23224370181560516)),(to_sfixed_a(0.04712607339024544)),(to_sfixed_a(0.00451234495267272)),(to_sfixed_a(0.16497978568077087)));

    constant weight_n1_218 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.02138575166463852)),(to_sfixed_a(-3.986187948612496e-06)),(to_sfixed_a(-1.0107194611919113e-05)),(to_sfixed_a(1.1851152521558106e-05)),(to_sfixed_a(-2.339085767744109e-05)),(to_sfixed_a(3.054016997339204e-05)),(to_sfixed_a(-1.5247806913976092e-05)),(to_sfixed_a(4.041306601720862e-05)),(to_sfixed_a(-6.128615495981649e-05)),(to_sfixed_a(-1.4827947779849637e-05)),(to_sfixed_a(7.828597154002637e-05)),(to_sfixed_a(-1.8340631868341006e-05)),(to_sfixed_a(-1.2415021956257988e-05)),(to_sfixed_a(2.1123765691299923e-05)),(to_sfixed_a(1.9496486856951378e-05)),(to_sfixed_a(-3.863119491143152e-05)),(to_sfixed_a(-2.2292982976068743e-05)),(to_sfixed_a(1.5944351616781205e-05)),(to_sfixed_a(4.6429329813690856e-05)),(to_sfixed_a(2.300835149071645e-05)),(to_sfixed_a(-8.947487913246732e-06)),(to_sfixed_a(4.214476575725712e-05)),(to_sfixed_a(8.295386942336336e-05)),(to_sfixed_a(2.3154962036642246e-05)),(to_sfixed_a(7.777359860483557e-05)),(to_sfixed_a(4.1979478737630416e-06)),(to_sfixed_a(-1.2363744872345706e-06)),(to_sfixed_a(-3.64883744623512e-05)),(to_sfixed_a(-4.666926179197617e-05)),(to_sfixed_a(0.00013261102139949799)),(to_sfixed_a(3.2541316613787785e-05)),(to_sfixed_a(-4.52130516350735e-05)),(to_sfixed_a(-1.6116259757836815e-06)),(to_sfixed_a(8.350131793122273e-06)),(to_sfixed_a(-5.1579641876742244e-05)),(to_sfixed_a(-2.1373161871451885e-05)),(to_sfixed_a(2.717648385441862e-05)),(to_sfixed_a(-2.5413068215129897e-05)));

    constant weight_n1_219 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.009812843054533005)),(to_sfixed_a(-1.9990118744317442e-05)),(to_sfixed_a(-3.301770630059764e-05)),(to_sfixed_a(1.9724334379134234e-06)),(to_sfixed_a(2.890056566684507e-05)),(to_sfixed_a(-3.1386447517434135e-05)),(to_sfixed_a(-1.7799302440835163e-05)),(to_sfixed_a(1.3287295587360859e-05)),(to_sfixed_a(-3.3698488550726324e-05)),(to_sfixed_a(5.38682206752128e-06)),(to_sfixed_a(2.1948639187030494e-05)),(to_sfixed_a(-3.867034683935344e-05)),(to_sfixed_a(1.9138602510793135e-05)),(to_sfixed_a(5.0503538659540936e-05)),(to_sfixed_a(-4.978380093234591e-05)),(to_sfixed_a(2.2472608179668896e-05)),(to_sfixed_a(2.12605173146585e-05)),(to_sfixed_a(-1.5057173186505679e-05)),(to_sfixed_a(-2.5541387003613636e-05)),(to_sfixed_a(1.6397838408011012e-05)),(to_sfixed_a(-2.3675906390963064e-07)),(to_sfixed_a(-9.148946992354468e-05)),(to_sfixed_a(-7.163920963648707e-05)),(to_sfixed_a(-5.186896487430204e-06)),(to_sfixed_a(-1.5491190424654633e-05)),(to_sfixed_a(-5.2264345868024975e-05)),(to_sfixed_a(7.936331530800089e-05)),(to_sfixed_a(-6.216223118826747e-05)),(to_sfixed_a(2.7380485335015692e-05)),(to_sfixed_a(4.335261837695725e-05)),(to_sfixed_a(3.392211510799825e-05)),(to_sfixed_a(3.366901000845246e-05)),(to_sfixed_a(-4.5979319111211225e-05)),(to_sfixed_a(7.57341695134528e-06)),(to_sfixed_a(5.0515413022367284e-05)),(to_sfixed_a(-7.319832366192713e-05)),(to_sfixed_a(3.3637130400165915e-05)),(to_sfixed_a(1.4755599295313004e-05)));

    constant weight_n1_220 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.028062470257282257)),(to_sfixed_a(3.0166920623742044e-06)),(to_sfixed_a(8.358803825103678e-06)),(to_sfixed_a(-1.4811350411036983e-05)),(to_sfixed_a(6.175738235469908e-05)),(to_sfixed_a(2.7972504540230148e-05)),(to_sfixed_a(-7.506391739298124e-06)),(to_sfixed_a(2.1312984245014377e-05)),(to_sfixed_a(1.0527014637773391e-05)),(to_sfixed_a(-4.627181988325901e-05)),(to_sfixed_a(7.341991931753e-06)),(to_sfixed_a(1.5665440514567308e-05)),(to_sfixed_a(-3.120108158327639e-05)),(to_sfixed_a(-1.9178416550857946e-05)),(to_sfixed_a(-3.820920755970292e-05)),(to_sfixed_a(7.205609290394932e-05)),(to_sfixed_a(2.3898264771560207e-05)),(to_sfixed_a(8.882284600986168e-05)),(to_sfixed_a(-3.0170322133926675e-05)),(to_sfixed_a(-6.82985319144791e-06)),(to_sfixed_a(-4.220429673296167e-06)),(to_sfixed_a(2.564770147728268e-05)),(to_sfixed_a(-4.009074928035261e-06)),(to_sfixed_a(3.548709719325416e-05)),(to_sfixed_a(-7.900749915279448e-05)),(to_sfixed_a(6.165781815070659e-05)),(to_sfixed_a(-1.806538966775406e-05)),(to_sfixed_a(2.6999246983905323e-05)),(to_sfixed_a(-4.1013332520378754e-05)),(to_sfixed_a(-4.236196036799811e-05)),(to_sfixed_a(5.781164873042144e-05)),(to_sfixed_a(4.282345616957173e-05)),(to_sfixed_a(2.8660100724664517e-05)),(to_sfixed_a(2.5422141334274784e-05)),(to_sfixed_a(-7.328540232265368e-05)),(to_sfixed_a(-2.5753775844350457e-05)),(to_sfixed_a(-2.3470993255614303e-06)),(to_sfixed_a(4.765833182318602e-06)));

    constant weight_n1_221 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.026207871735095978)),(to_sfixed_a(-1.588656050444115e-05)),(to_sfixed_a(-8.466401595796924e-06)),(to_sfixed_a(2.451571162964683e-05)),(to_sfixed_a(-5.394697836891282e-06)),(to_sfixed_a(-2.823213071678765e-05)),(to_sfixed_a(5.964648153167218e-05)),(to_sfixed_a(-3.302856157461065e-06)),(to_sfixed_a(-6.773062523279805e-06)),(to_sfixed_a(4.688898116000928e-05)),(to_sfixed_a(1.6871144907781854e-05)),(to_sfixed_a(-4.7489644202869385e-05)),(to_sfixed_a(2.3937445803312585e-05)),(to_sfixed_a(1.0329656106478069e-05)),(to_sfixed_a(7.387023651972413e-05)),(to_sfixed_a(-8.014117156562861e-06)),(to_sfixed_a(-5.39407592441421e-05)),(to_sfixed_a(-2.517276516300626e-05)),(to_sfixed_a(-1.0293509149050806e-05)),(to_sfixed_a(-3.3579162845853716e-05)),(to_sfixed_a(-3.2773408747743815e-05)),(to_sfixed_a(-4.397971679281909e-06)),(to_sfixed_a(-0.00012649293057620525)),(to_sfixed_a(-1.5160919701884268e-06)),(to_sfixed_a(7.877500138420146e-06)),(to_sfixed_a(-1.06231027530157e-05)),(to_sfixed_a(-4.4421126403904054e-06)),(to_sfixed_a(2.7145973945152946e-05)),(to_sfixed_a(-1.5157757843553554e-05)),(to_sfixed_a(-2.985658056786633e-06)),(to_sfixed_a(2.0010260413982905e-05)),(to_sfixed_a(-2.427583785902243e-05)),(to_sfixed_a(1.3559567378251813e-05)),(to_sfixed_a(2.9932209145044908e-05)),(to_sfixed_a(3.6245797673473135e-05)),(to_sfixed_a(7.119127258192748e-05)),(to_sfixed_a(-8.460082608507946e-05)),(to_sfixed_a(0.00012224358215462416)));

    constant weight_n1_222 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.0898909643292427)),(to_sfixed_a(0.006079173646867275)),(to_sfixed_a(-0.041632384061813354)),(to_sfixed_a(-0.007057743147015572)),(to_sfixed_a(0.05714161694049835)),(to_sfixed_a(-0.01940731331706047)),(to_sfixed_a(-0.020522816106677055)),(to_sfixed_a(0.04119192063808441)),(to_sfixed_a(0.049335069954395294)),(to_sfixed_a(-0.036277636885643005)),(to_sfixed_a(0.06359367072582245)),(to_sfixed_a(-0.032004717737436295)),(to_sfixed_a(0.022261925041675568)),(to_sfixed_a(-0.04619995877146721)),(to_sfixed_a(0.0039322166703641415)),(to_sfixed_a(0.03035571612417698)),(to_sfixed_a(-0.02453826181590557)),(to_sfixed_a(-0.01897125504910946)),(to_sfixed_a(0.016618477180600166)),(to_sfixed_a(0.03225528076291084)),(to_sfixed_a(-0.04263800010085106)),(to_sfixed_a(0.03165898472070694)),(to_sfixed_a(-0.0371684767305851)),(to_sfixed_a(-0.03997129574418068)),(to_sfixed_a(-0.014138147234916687)),(to_sfixed_a(-0.08945470303297043)),(to_sfixed_a(0.0215336661785841)),(to_sfixed_a(-0.07551132887601852)),(to_sfixed_a(-0.061977703124284744)),(to_sfixed_a(0.027087895199656487)),(to_sfixed_a(0.006638317834585905)),(to_sfixed_a(-0.025392405688762665)),(to_sfixed_a(0.01718437671661377)),(to_sfixed_a(-0.038265109062194824)),(to_sfixed_a(-0.11200244724750519)),(to_sfixed_a(-0.030399398878216743)),(to_sfixed_a(-0.08812343329191208)),(to_sfixed_a(0.07704717665910721)));

    constant weight_n1_223 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.103602834045887)),(to_sfixed_a(-0.19706110656261444)),(to_sfixed_a(-0.013762356713414192)),(to_sfixed_a(-0.16208462417125702)),(to_sfixed_a(0.1726546734571457)),(to_sfixed_a(0.005138798151165247)),(to_sfixed_a(-0.1320897936820984)),(to_sfixed_a(-0.12130006402730942)),(to_sfixed_a(0.13097020983695984)),(to_sfixed_a(0.06371960788965225)),(to_sfixed_a(0.009560937993228436)),(to_sfixed_a(0.03282599151134491)),(to_sfixed_a(-0.09648729860782623)),(to_sfixed_a(0.03300045430660248)),(to_sfixed_a(-0.2672998011112213)),(to_sfixed_a(0.19093090295791626)),(to_sfixed_a(-0.015574718825519085)),(to_sfixed_a(-0.08519301563501358)),(to_sfixed_a(0.10660691559314728)),(to_sfixed_a(0.1001584455370903)),(to_sfixed_a(-0.04437866806983948)),(to_sfixed_a(0.1190771609544754)),(to_sfixed_a(0.05534753203392029)),(to_sfixed_a(-0.25969037413597107)),(to_sfixed_a(0.0551285594701767)),(to_sfixed_a(-0.024084215983748436)),(to_sfixed_a(-0.0008502501295879483)),(to_sfixed_a(-0.0006826221360825002)),(to_sfixed_a(0.08575572073459625)),(to_sfixed_a(0.04160560294985771)),(to_sfixed_a(0.08599300682544708)),(to_sfixed_a(0.2927974760532379)),(to_sfixed_a(0.04333435371518135)),(to_sfixed_a(-0.11589153856039047)),(to_sfixed_a(-0.01892399601638317)),(to_sfixed_a(0.03498339280486107)),(to_sfixed_a(0.09746342152357101)),(to_sfixed_a(0.015513496473431587)));

    constant weight_n1_224 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.03196924552321434)),(to_sfixed_a(-4.4048665586160496e-05)),(to_sfixed_a(-1.4924888091627508e-05)),(to_sfixed_a(-7.207190355984494e-05)),(to_sfixed_a(7.331107917707413e-05)),(to_sfixed_a(1.2370477634249255e-05)),(to_sfixed_a(2.9773145797662437e-05)),(to_sfixed_a(-1.8969587472383864e-05)),(to_sfixed_a(-4.408513177622808e-06)),(to_sfixed_a(-3.563659993233159e-05)),(to_sfixed_a(-4.381238977657631e-05)),(to_sfixed_a(3.733791527338326e-05)),(to_sfixed_a(-3.819439007202163e-05)),(to_sfixed_a(-3.405845563975163e-05)),(to_sfixed_a(-7.602386631333502e-06)),(to_sfixed_a(-3.1300451155402698e-06)),(to_sfixed_a(-1.7680678183751297e-06)),(to_sfixed_a(-2.0787454559467733e-05)),(to_sfixed_a(-6.345506699290127e-05)),(to_sfixed_a(-1.1721902410499752e-05)),(to_sfixed_a(2.074557232845109e-05)),(to_sfixed_a(4.932787123834714e-05)),(to_sfixed_a(-7.649202598258853e-05)),(to_sfixed_a(-3.135894803563133e-05)),(to_sfixed_a(6.425139144994318e-05)),(to_sfixed_a(4.0574544982519e-05)),(to_sfixed_a(2.8816686608479358e-05)),(to_sfixed_a(4.881871518591652e-06)),(to_sfixed_a(-8.112195791909471e-05)),(to_sfixed_a(7.705318421358243e-05)),(to_sfixed_a(7.143997208913788e-06)),(to_sfixed_a(3.081176691921428e-05)),(to_sfixed_a(-5.676868750015274e-05)),(to_sfixed_a(-5.5467030506406445e-06)),(to_sfixed_a(-2.114116568918689e-06)),(to_sfixed_a(-4.974147668690421e-05)),(to_sfixed_a(1.3354865586734377e-05)),(to_sfixed_a(0.00011946614540647715)));

    constant weight_n1_225 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.037106502801179886)),(to_sfixed_a(3.746619404410012e-05)),(to_sfixed_a(4.179280040261801e-06)),(to_sfixed_a(-4.350330345914699e-05)),(to_sfixed_a(-5.6096443586284295e-05)),(to_sfixed_a(2.364521424169652e-05)),(to_sfixed_a(-4.7804358473513275e-05)),(to_sfixed_a(4.660147533286363e-05)),(to_sfixed_a(1.776062708813697e-05)),(to_sfixed_a(2.2883883502800018e-05)),(to_sfixed_a(3.279232623754069e-05)),(to_sfixed_a(-1.828366112022195e-05)),(to_sfixed_a(-8.35733299027197e-05)),(to_sfixed_a(-2.045305518549867e-05)),(to_sfixed_a(2.3310152755584568e-05)),(to_sfixed_a(5.578715354204178e-05)),(to_sfixed_a(7.171644392656162e-05)),(to_sfixed_a(3.2160816772375256e-05)),(to_sfixed_a(0.00010383447079220787)),(to_sfixed_a(-1.5467136108782142e-05)),(to_sfixed_a(-1.7901014871313237e-05)),(to_sfixed_a(4.5485026930691674e-05)),(to_sfixed_a(-8.546008029952645e-05)),(to_sfixed_a(-7.661680865567178e-05)),(to_sfixed_a(0.00012212000729050487)),(to_sfixed_a(1.3965292964712717e-05)),(to_sfixed_a(-8.300003173644654e-06)),(to_sfixed_a(5.108975074108457e-06)),(to_sfixed_a(-1.705096656223759e-05)),(to_sfixed_a(-3.373446088517085e-05)),(to_sfixed_a(3.575701703084633e-05)),(to_sfixed_a(-5.768705887021497e-05)),(to_sfixed_a(3.499853119137697e-05)),(to_sfixed_a(-0.00012148371752118692)),(to_sfixed_a(4.859269756707363e-05)),(to_sfixed_a(8.914497448131442e-05)),(to_sfixed_a(-2.6479923690203577e-05)),(to_sfixed_a(2.635436067066621e-05)));

    constant weight_n1_226 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.02545987069606781)),(to_sfixed_a(-8.789826097199693e-06)),(to_sfixed_a(6.387831672327593e-05)),(to_sfixed_a(3.4748733014566824e-05)),(to_sfixed_a(-8.355692443728913e-06)),(to_sfixed_a(-1.7014930563163944e-05)),(to_sfixed_a(-2.3498545488109812e-05)),(to_sfixed_a(-5.224844426265918e-05)),(to_sfixed_a(6.151181878522038e-05)),(to_sfixed_a(1.4905552234267816e-05)),(to_sfixed_a(3.8184549566722126e-07)),(to_sfixed_a(-4.400027319206856e-05)),(to_sfixed_a(9.164683433482423e-06)),(to_sfixed_a(-7.858811295591295e-05)),(to_sfixed_a(3.925599958165549e-05)),(to_sfixed_a(1.3180508176446892e-05)),(to_sfixed_a(-4.5020715333521366e-05)),(to_sfixed_a(-3.402964648557827e-05)),(to_sfixed_a(5.107419929117896e-05)),(to_sfixed_a(-2.1614047000184655e-05)),(to_sfixed_a(-7.092631858540699e-05)),(to_sfixed_a(2.1826194824825507e-06)),(to_sfixed_a(-5.748986495746067e-06)),(to_sfixed_a(-9.075376874534413e-05)),(to_sfixed_a(-5.410680751083419e-05)),(to_sfixed_a(-2.31558096857043e-05)),(to_sfixed_a(3.074496635235846e-05)),(to_sfixed_a(-2.7924226742470637e-05)),(to_sfixed_a(-4.20835058321245e-05)),(to_sfixed_a(8.301267371280119e-05)),(to_sfixed_a(-2.944715197372716e-05)),(to_sfixed_a(9.527218026050832e-06)),(to_sfixed_a(9.341352415503934e-05)),(to_sfixed_a(9.746757132234052e-05)),(to_sfixed_a(0.00011765342060243711)),(to_sfixed_a(1.77129859366687e-05)),(to_sfixed_a(-2.491007762728259e-05)),(to_sfixed_a(1.033903936331626e-05)));

    constant weight_n1_227 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.12756170332431793)),(to_sfixed_a(0.04503527283668518)),(to_sfixed_a(-0.02444954216480255)),(to_sfixed_a(-0.02333042398095131)),(to_sfixed_a(0.2063496857881546)),(to_sfixed_a(0.0510086864233017)),(to_sfixed_a(0.017861366271972656)),(to_sfixed_a(-0.11211147159337997)),(to_sfixed_a(-0.009978367947041988)),(to_sfixed_a(0.19347454607486725)),(to_sfixed_a(-0.38670673966407776)),(to_sfixed_a(0.1435510367155075)),(to_sfixed_a(0.09204362332820892)),(to_sfixed_a(-0.20622658729553223)),(to_sfixed_a(-0.0933343842625618)),(to_sfixed_a(-0.00647076265886426)),(to_sfixed_a(0.0935150757431984)),(to_sfixed_a(0.0568925216794014)),(to_sfixed_a(-0.02270865999162197)),(to_sfixed_a(0.14477823674678802)),(to_sfixed_a(-0.015777355059981346)),(to_sfixed_a(-0.17470301687717438)),(to_sfixed_a(0.12237659096717834)),(to_sfixed_a(-0.19410720467567444)),(to_sfixed_a(0.08742647618055344)),(to_sfixed_a(0.02344891056418419)),(to_sfixed_a(-0.06517455726861954)),(to_sfixed_a(-0.036777328699827194)),(to_sfixed_a(0.06887584179639816)),(to_sfixed_a(0.040104735642671585)),(to_sfixed_a(0.06600851565599442)),(to_sfixed_a(-0.1107664704322815)),(to_sfixed_a(-0.03603369742631912)),(to_sfixed_a(0.014007233083248138)),(to_sfixed_a(0.09027576446533203)),(to_sfixed_a(0.1328711211681366)),(to_sfixed_a(-0.08630160242319107)),(to_sfixed_a(-0.030606862157583237)));

    constant weight_n1_228 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.15497596561908722)),(to_sfixed_a(0.0805223286151886)),(to_sfixed_a(-0.17698733508586884)),(to_sfixed_a(0.0017904757987707853)),(to_sfixed_a(0.19533266127109528)),(to_sfixed_a(-0.09610606729984283)),(to_sfixed_a(0.022019673138856888)),(to_sfixed_a(0.06142152100801468)),(to_sfixed_a(0.14278936386108398)),(to_sfixed_a(-0.04956602677702904)),(to_sfixed_a(-0.07391666620969772)),(to_sfixed_a(-0.021463271230459213)),(to_sfixed_a(0.1849546581506729)),(to_sfixed_a(0.20323683321475983)),(to_sfixed_a(0.08569373190402985)),(to_sfixed_a(-0.11030051112174988)),(to_sfixed_a(-0.12586145102977753)),(to_sfixed_a(0.05784430354833603)),(to_sfixed_a(0.31332826614379883)),(to_sfixed_a(-0.20878718793392181)),(to_sfixed_a(0.007192156743258238)),(to_sfixed_a(-0.26293039321899414)),(to_sfixed_a(-0.18327458202838898)),(to_sfixed_a(-0.14328213036060333)),(to_sfixed_a(-0.29743367433547974)),(to_sfixed_a(0.1300666630268097)),(to_sfixed_a(-0.1597280353307724)),(to_sfixed_a(0.0037475537974387407)),(to_sfixed_a(-0.008535024709999561)),(to_sfixed_a(0.1939748078584671)),(to_sfixed_a(-0.10505213588476181)),(to_sfixed_a(-0.04281610623002052)),(to_sfixed_a(-0.05949409678578377)),(to_sfixed_a(-0.23253712058067322)),(to_sfixed_a(-0.10839288681745529)),(to_sfixed_a(0.00424337200820446)),(to_sfixed_a(0.16061997413635254)),(to_sfixed_a(-0.00932370126247406)));

    constant weight_n1_229 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.1564747393131256)),(to_sfixed_a(-0.13790889084339142)),(to_sfixed_a(0.013850480318069458)),(to_sfixed_a(-0.13322509825229645)),(to_sfixed_a(-0.07519382983446121)),(to_sfixed_a(0.05010409280657768)),(to_sfixed_a(-0.10323379933834076)),(to_sfixed_a(0.1105283573269844)),(to_sfixed_a(-0.03406529873609543)),(to_sfixed_a(0.16195930540561676)),(to_sfixed_a(0.014846795238554478)),(to_sfixed_a(0.16849710047245026)),(to_sfixed_a(0.014260157011449337)),(to_sfixed_a(-0.0897059366106987)),(to_sfixed_a(-0.08859267085790634)),(to_sfixed_a(-0.057675302028656006)),(to_sfixed_a(-0.08275410532951355)),(to_sfixed_a(-0.09139865636825562)),(to_sfixed_a(0.10180087387561798)),(to_sfixed_a(-0.04384687542915344)),(to_sfixed_a(-0.07809129357337952)),(to_sfixed_a(0.09679756313562393)),(to_sfixed_a(0.01374909095466137)),(to_sfixed_a(0.11257272213697433)),(to_sfixed_a(-0.04841756075620651)),(to_sfixed_a(-0.017370570451021194)),(to_sfixed_a(-0.08340500295162201)),(to_sfixed_a(-0.2516948878765106)),(to_sfixed_a(-0.10014557093381882)),(to_sfixed_a(0.12514656782150269)),(to_sfixed_a(0.08644992113113403)),(to_sfixed_a(0.0662066712975502)),(to_sfixed_a(-0.11848019063472748)),(to_sfixed_a(-0.039222147315740585)),(to_sfixed_a(0.036919306963682175)),(to_sfixed_a(-0.020935148000717163)),(to_sfixed_a(0.04865493252873421)),(to_sfixed_a(-0.1483730971813202)));

    constant weight_n1_230 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.011495199985802174)),(to_sfixed_a(-7.0899163802096155e-06)),(to_sfixed_a(-1.4926359654054977e-05)),(to_sfixed_a(4.192472988506779e-05)),(to_sfixed_a(-1.748716204019729e-05)),(to_sfixed_a(3.821834616246633e-05)),(to_sfixed_a(5.195868288865313e-05)),(to_sfixed_a(-1.75611912709428e-05)),(to_sfixed_a(-1.5925754269119352e-05)),(to_sfixed_a(6.919189763721079e-05)),(to_sfixed_a(-0.00010005735384766012)),(to_sfixed_a(2.7748546926886775e-05)),(to_sfixed_a(3.3939511922653764e-05)),(to_sfixed_a(-5.6862019846448675e-05)),(to_sfixed_a(1.339833761448972e-05)),(to_sfixed_a(-1.1569616617634892e-05)),(to_sfixed_a(-3.1031479011289775e-05)),(to_sfixed_a(6.306929572019726e-05)),(to_sfixed_a(2.021906584559474e-05)),(to_sfixed_a(3.804538573604077e-05)),(to_sfixed_a(-2.955248419311829e-05)),(to_sfixed_a(-6.844925337645691e-06)),(to_sfixed_a(1.530422923678998e-05)),(to_sfixed_a(2.9677641578018665e-05)),(to_sfixed_a(-3.909883616870502e-06)),(to_sfixed_a(-3.140568878734484e-05)),(to_sfixed_a(7.598442607559264e-05)),(to_sfixed_a(-5.057904672867153e-06)),(to_sfixed_a(0.00010416975419502705)),(to_sfixed_a(-8.078062819549814e-06)),(to_sfixed_a(3.667881901492365e-05)),(to_sfixed_a(3.7826524931006134e-05)),(to_sfixed_a(-1.8059565263683908e-05)),(to_sfixed_a(0.0001000144038698636)),(to_sfixed_a(5.096045424579643e-05)),(to_sfixed_a(-1.5433388398378156e-05)),(to_sfixed_a(-2.0323952412582003e-05)),(to_sfixed_a(-7.086365258146543e-06)));

    constant weight_n1_231 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.007511806208640337)),(to_sfixed_a(4.234423613524996e-05)),(to_sfixed_a(-1.8038346752291545e-05)),(to_sfixed_a(2.153600325982552e-05)),(to_sfixed_a(4.054842793266289e-05)),(to_sfixed_a(-4.884950612904504e-05)),(to_sfixed_a(1.6572446384088835e-06)),(to_sfixed_a(2.584340654721018e-05)),(to_sfixed_a(-1.8150592950405553e-05)),(to_sfixed_a(7.943285891087726e-05)),(to_sfixed_a(3.955979263992049e-05)),(to_sfixed_a(2.494294494681526e-05)),(to_sfixed_a(1.0841683433682192e-05)),(to_sfixed_a(-3.416031540837139e-05)),(to_sfixed_a(2.47258176386822e-05)),(to_sfixed_a(-3.1843424949329346e-05)),(to_sfixed_a(-8.660363528179005e-05)),(to_sfixed_a(3.826237661996856e-05)),(to_sfixed_a(8.401108971156646e-06)),(to_sfixed_a(-8.43518409965327e-06)),(to_sfixed_a(-4.129290118726203e-06)),(to_sfixed_a(0.00010677660611690953)),(to_sfixed_a(-1.9668825189000927e-05)),(to_sfixed_a(-3.328453749418259e-05)),(to_sfixed_a(-6.351849879138172e-05)),(to_sfixed_a(-1.0578671208349988e-05)),(to_sfixed_a(-1.053590403898852e-05)),(to_sfixed_a(-2.3860809960751794e-05)),(to_sfixed_a(-1.6368343494832516e-05)),(to_sfixed_a(-1.3800616216030903e-05)),(to_sfixed_a(-5.365170363802463e-05)),(to_sfixed_a(-0.00011596005060710013)),(to_sfixed_a(8.149805944412947e-05)),(to_sfixed_a(-7.874556467868388e-05)),(to_sfixed_a(3.707632276928052e-05)),(to_sfixed_a(-9.579880861565471e-05)),(to_sfixed_a(-1.786008579074405e-05)),(to_sfixed_a(3.995920269517228e-05)));

    constant weight_n1_232 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.0077761756256222725)),(to_sfixed_a(-1.2292275641812012e-06)),(to_sfixed_a(1.5035702745080926e-05)),(to_sfixed_a(-4.3379161070333794e-05)),(to_sfixed_a(3.655116870504571e-06)),(to_sfixed_a(3.5566521546570584e-05)),(to_sfixed_a(-3.796459395744023e-06)),(to_sfixed_a(-1.5695737602072768e-05)),(to_sfixed_a(-4.49803592346143e-05)),(to_sfixed_a(-4.946316403220408e-05)),(to_sfixed_a(-7.188328163465485e-05)),(to_sfixed_a(-1.705714203126263e-05)),(to_sfixed_a(3.333702989039011e-05)),(to_sfixed_a(1.6694670193828642e-05)),(to_sfixed_a(-3.1415867852047086e-05)),(to_sfixed_a(2.585179390734993e-05)),(to_sfixed_a(5.326737664290704e-05)),(to_sfixed_a(-3.9184364140965044e-05)),(to_sfixed_a(3.553260467015207e-05)),(to_sfixed_a(-5.7289926189696416e-05)),(to_sfixed_a(2.3913069526315667e-05)),(to_sfixed_a(5.3174200729699805e-05)),(to_sfixed_a(3.26365880027879e-05)),(to_sfixed_a(4.86184362671338e-05)),(to_sfixed_a(-1.4323458344733808e-05)),(to_sfixed_a(1.3270304407342337e-05)),(to_sfixed_a(5.527624671231024e-05)),(to_sfixed_a(-1.7924308849615045e-05)),(to_sfixed_a(-1.0660824955266435e-05)),(to_sfixed_a(-1.6286201571347192e-05)),(to_sfixed_a(1.1407722013245802e-05)),(to_sfixed_a(5.885333303012885e-05)),(to_sfixed_a(5.510020491783507e-05)),(to_sfixed_a(3.226676199119538e-05)),(to_sfixed_a(1.9403689293540083e-05)),(to_sfixed_a(2.92111453745747e-05)),(to_sfixed_a(1.0410670256533194e-05)),(to_sfixed_a(1.4721363186254166e-05)));

    constant weight_n1_233 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.2585902214050293)),(to_sfixed_a(-0.012578031048178673)),(to_sfixed_a(-0.0016970658907666802)),(to_sfixed_a(0.010410075075924397)),(to_sfixed_a(0.023923536762595177)),(to_sfixed_a(-0.0001253922819159925)),(to_sfixed_a(-0.05166248604655266)),(to_sfixed_a(0.027994941920042038)),(to_sfixed_a(0.014175480231642723)),(to_sfixed_a(-0.011671802029013634)),(to_sfixed_a(0.015500720590353012)),(to_sfixed_a(0.013982213102281094)),(to_sfixed_a(0.0028014553245157003)),(to_sfixed_a(-0.0384613461792469)),(to_sfixed_a(0.017939480021595955)),(to_sfixed_a(-0.046866524964571)),(to_sfixed_a(-0.06311587989330292)),(to_sfixed_a(-0.0481363981962204)),(to_sfixed_a(-0.0312483049929142)),(to_sfixed_a(-0.002163292607292533)),(to_sfixed_a(-0.010191353969275951)),(to_sfixed_a(-0.0338742695748806)),(to_sfixed_a(0.016995064914226532)),(to_sfixed_a(0.03172145038843155)),(to_sfixed_a(-0.031779561191797256)),(to_sfixed_a(0.011425058357417583)),(to_sfixed_a(0.011895165778696537)),(to_sfixed_a(0.02927924506366253)),(to_sfixed_a(-0.010817211121320724)),(to_sfixed_a(-0.007030049804598093)),(to_sfixed_a(0.021937552839517593)),(to_sfixed_a(-0.007384744007140398)),(to_sfixed_a(-0.0398406907916069)),(to_sfixed_a(-0.016779227182269096)),(to_sfixed_a(0.017455479130148888)),(to_sfixed_a(0.04808450862765312)),(to_sfixed_a(0.000131741413497366)),(to_sfixed_a(-0.045919258147478104)));

    constant weight_n1_234 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.08158189058303833)),(to_sfixed_a(0.019897419959306717)),(to_sfixed_a(-0.00672896346077323)),(to_sfixed_a(0.002924447413533926)),(to_sfixed_a(0.0025013552512973547)),(to_sfixed_a(-0.04331120476126671)),(to_sfixed_a(-0.0002618332509882748)),(to_sfixed_a(0.023029984906315804)),(to_sfixed_a(0.0058055161498487)),(to_sfixed_a(0.017391206696629524)),(to_sfixed_a(0.004209456499665976)),(to_sfixed_a(-0.03640243038535118)),(to_sfixed_a(0.01724069193005562)),(to_sfixed_a(-0.030605394393205643)),(to_sfixed_a(-0.017412351444363594)),(to_sfixed_a(-0.025532366707921028)),(to_sfixed_a(-0.004189825616776943)),(to_sfixed_a(-0.014187411405146122)),(to_sfixed_a(0.02265278249979019)),(to_sfixed_a(-0.02801445871591568)),(to_sfixed_a(0.0011499070096760988)),(to_sfixed_a(0.02070818655192852)),(to_sfixed_a(0.03107963502407074)),(to_sfixed_a(-0.01480037160217762)),(to_sfixed_a(-0.006028526928275824)),(to_sfixed_a(0.024873623624444008)),(to_sfixed_a(-0.011966238729655743)),(to_sfixed_a(-0.011961313895881176)),(to_sfixed_a(-0.019813962280750275)),(to_sfixed_a(0.03289907053112984)),(to_sfixed_a(-0.029337655752897263)),(to_sfixed_a(-0.032304514199495316)),(to_sfixed_a(-0.026889238506555557)),(to_sfixed_a(0.016602715477347374)),(to_sfixed_a(-0.010311477817595005)),(to_sfixed_a(-0.03633382171392441)),(to_sfixed_a(0.031210601329803467)),(to_sfixed_a(0.011488466523587704)));

    constant weight_n1_235 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.011567567475140095)),(to_sfixed_a(-0.05571258068084717)),(to_sfixed_a(0.1469251811504364)),(to_sfixed_a(0.0995166152715683)),(to_sfixed_a(0.14289061725139618)),(to_sfixed_a(-0.09365817159414291)),(to_sfixed_a(-0.03419561684131622)),(to_sfixed_a(0.2117720991373062)),(to_sfixed_a(-0.02998960390686989)),(to_sfixed_a(-0.0329408198595047)),(to_sfixed_a(-0.023444635793566704)),(to_sfixed_a(-0.05177977681159973)),(to_sfixed_a(0.13216446340084076)),(to_sfixed_a(0.06856481730937958)),(to_sfixed_a(-0.23960307240486145)),(to_sfixed_a(0.09685196727514267)),(to_sfixed_a(0.03981856629252434)),(to_sfixed_a(-0.17541931569576263)),(to_sfixed_a(-0.2615495026111603)),(to_sfixed_a(-0.13715192675590515)),(to_sfixed_a(0.12013702839612961)),(to_sfixed_a(-0.10767960548400879)),(to_sfixed_a(0.11418814957141876)),(to_sfixed_a(-0.017442651093006134)),(to_sfixed_a(0.03977219760417938)),(to_sfixed_a(0.04239775240421295)),(to_sfixed_a(-0.10610228776931763)),(to_sfixed_a(-0.1356007307767868)),(to_sfixed_a(-0.09990163892507553)),(to_sfixed_a(0.10378607362508774)),(to_sfixed_a(0.19468523561954498)),(to_sfixed_a(0.060922689735889435)),(to_sfixed_a(0.02131601795554161)),(to_sfixed_a(-0.08187419176101685)),(to_sfixed_a(-0.015160397626459599)),(to_sfixed_a(0.0438968725502491)),(to_sfixed_a(0.04827078431844711)),(to_sfixed_a(0.027235889807343483)));

    constant weight_n1_236 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.012585005722939968)),(to_sfixed_a(1.3653486348630395e-05)),(to_sfixed_a(-5.510961273103021e-05)),(to_sfixed_a(3.890438892995007e-05)),(to_sfixed_a(2.566908733570017e-05)),(to_sfixed_a(-9.665512152423616e-06)),(to_sfixed_a(1.0739964636741206e-05)),(to_sfixed_a(3.266903877374716e-05)),(to_sfixed_a(-8.173336391337216e-05)),(to_sfixed_a(-1.1983298463746905e-05)),(to_sfixed_a(-1.840794902818743e-05)),(to_sfixed_a(1.4413243661692832e-05)),(to_sfixed_a(-6.082192703615874e-05)),(to_sfixed_a(-5.289326509227976e-06)),(to_sfixed_a(2.2369218640960753e-05)),(to_sfixed_a(5.954680091235787e-06)),(to_sfixed_a(6.114984444138827e-06)),(to_sfixed_a(5.052018241258338e-05)),(to_sfixed_a(4.284414171706885e-05)),(to_sfixed_a(-5.5584237998118624e-05)),(to_sfixed_a(-4.074173193657771e-05)),(to_sfixed_a(5.6280919125129e-06)),(to_sfixed_a(-3.117821688647382e-05)),(to_sfixed_a(-2.3837252228986472e-05)),(to_sfixed_a(-7.848019595257938e-05)),(to_sfixed_a(4.041227157358662e-07)),(to_sfixed_a(-0.00010289309284416959)),(to_sfixed_a(-7.617688970640302e-05)),(to_sfixed_a(5.4756288591306657e-05)),(to_sfixed_a(1.0207464583800174e-05)),(to_sfixed_a(-5.194517143536359e-05)),(to_sfixed_a(1.8203483705292456e-05)),(to_sfixed_a(3.4691340260906145e-05)),(to_sfixed_a(2.6993491701432504e-05)),(to_sfixed_a(9.10243579710368e-06)),(to_sfixed_a(3.208921407349408e-05)),(to_sfixed_a(-6.976459553698078e-05)),(to_sfixed_a(6.826207936683204e-06)));

    constant weight_n1_237 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.10138296335935593)),(to_sfixed_a(-0.0012866833712905645)),(to_sfixed_a(0.005217888858169317)),(to_sfixed_a(-0.009996401146054268)),(to_sfixed_a(0.002555137500166893)),(to_sfixed_a(-0.0008278582827188075)),(to_sfixed_a(-0.0076315151527523994)),(to_sfixed_a(0.004353985656052828)),(to_sfixed_a(0.0042342632077634335)),(to_sfixed_a(0.012018951587378979)),(to_sfixed_a(-0.0030106031335890293)),(to_sfixed_a(-0.0026365937665104866)),(to_sfixed_a(-0.0010181530378758907)),(to_sfixed_a(0.001670438447035849)),(to_sfixed_a(-0.003890013787895441)),(to_sfixed_a(-0.000387421838240698)),(to_sfixed_a(0.004314846359193325)),(to_sfixed_a(0.0012788847088813782)),(to_sfixed_a(0.0065599288791418076)),(to_sfixed_a(0.004032290540635586)),(to_sfixed_a(-0.006682706531137228)),(to_sfixed_a(0.00527567695826292)),(to_sfixed_a(-0.0040045431815087795)),(to_sfixed_a(-0.01182397361844778)),(to_sfixed_a(0.005887610372155905)),(to_sfixed_a(0.0043663703836500645)),(to_sfixed_a(-0.002232647268101573)),(to_sfixed_a(-0.0005223649204708636)),(to_sfixed_a(-0.004195898771286011)),(to_sfixed_a(0.010919235646724701)),(to_sfixed_a(-0.00313609023578465)),(to_sfixed_a(-0.013984959572553635)),(to_sfixed_a(-0.008367303758859634)),(to_sfixed_a(0.005897517316043377)),(to_sfixed_a(-0.0034052215050905943)),(to_sfixed_a(-0.00457456661388278)),(to_sfixed_a(-0.01074096281081438)),(to_sfixed_a(-0.010121593251824379)));

    constant weight_n1_238 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.017466960474848747)),(to_sfixed_a(1.0966742593154777e-05)),(to_sfixed_a(-4.321645974414423e-06)),(to_sfixed_a(-1.9404640624998137e-05)),(to_sfixed_a(-3.10422656184528e-05)),(to_sfixed_a(-2.428947846055962e-05)),(to_sfixed_a(-1.1866371096402872e-05)),(to_sfixed_a(6.336021033348516e-05)),(to_sfixed_a(-5.431670433608815e-05)),(to_sfixed_a(-4.56880297861062e-05)),(to_sfixed_a(5.372200121200876e-06)),(to_sfixed_a(1.6764823158155195e-05)),(to_sfixed_a(-7.215835040597085e-08)),(to_sfixed_a(-6.365161198118585e-07)),(to_sfixed_a(-9.906813147608773e-07)),(to_sfixed_a(2.5430235837120563e-05)),(to_sfixed_a(0.00012755265925079584)),(to_sfixed_a(-6.837466912656964e-07)),(to_sfixed_a(8.270076250482816e-06)),(to_sfixed_a(1.0438187928230036e-05)),(to_sfixed_a(-9.965917706722394e-05)),(to_sfixed_a(-2.6220225208817283e-06)),(to_sfixed_a(5.511179188033566e-05)),(to_sfixed_a(9.774946374818683e-05)),(to_sfixed_a(-5.468365634442307e-05)),(to_sfixed_a(-1.2246465303178411e-05)),(to_sfixed_a(-5.8999680732085835e-06)),(to_sfixed_a(-2.061701707134489e-05)),(to_sfixed_a(8.051897748373449e-05)),(to_sfixed_a(4.746539343614131e-05)),(to_sfixed_a(-9.43573809308873e-07)),(to_sfixed_a(3.991109042544849e-05)),(to_sfixed_a(6.617471808567643e-05)),(to_sfixed_a(-0.0001504043029854074)),(to_sfixed_a(-0.00013716172543354332)),(to_sfixed_a(0.00015771201287861913)),(to_sfixed_a(-2.335487624804955e-05)),(to_sfixed_a(5.036702350480482e-05)));

    constant weight_n1_239 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.4185349643230438)),(to_sfixed_a(-0.06057576462626457)),(to_sfixed_a(-0.02011050097644329)),(to_sfixed_a(0.02491292543709278)),(to_sfixed_a(-0.029656855389475822)),(to_sfixed_a(0.009480771608650684)),(to_sfixed_a(-0.03465600311756134)),(to_sfixed_a(0.02596265822649002)),(to_sfixed_a(-0.004340344108641148)),(to_sfixed_a(-0.06214392930269241)),(to_sfixed_a(0.0512617826461792)),(to_sfixed_a(0.009621505625545979)),(to_sfixed_a(-0.0786266103386879)),(to_sfixed_a(-0.11148817837238312)),(to_sfixed_a(-0.01959512196481228)),(to_sfixed_a(0.0050658113323152065)),(to_sfixed_a(-0.0349789597094059)),(to_sfixed_a(-0.01013726182281971)),(to_sfixed_a(-0.04245580732822418)),(to_sfixed_a(0.046503741294145584)),(to_sfixed_a(0.04277224466204643)),(to_sfixed_a(0.13478368520736694)),(to_sfixed_a(-0.10821899771690369)),(to_sfixed_a(0.10572204738855362)),(to_sfixed_a(0.1208723932504654)),(to_sfixed_a(0.13626256585121155)),(to_sfixed_a(-0.04848616570234299)),(to_sfixed_a(0.013311312533915043)),(to_sfixed_a(0.19911223649978638)),(to_sfixed_a(-0.09144969284534454)),(to_sfixed_a(0.10237301141023636)),(to_sfixed_a(0.07572674006223679)),(to_sfixed_a(-0.23652230203151703)),(to_sfixed_a(0.06634872406721115)),(to_sfixed_a(0.03399768844246864)),(to_sfixed_a(-0.15206797420978546)),(to_sfixed_a(-0.03717448189854622)),(to_sfixed_a(0.08303698897361755)));

    constant weight_n1_240 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.021449536085128784)),(to_sfixed_a(-5.441805478767492e-05)),(to_sfixed_a(-3.050589657505043e-05)),(to_sfixed_a(-6.250392470974475e-05)),(to_sfixed_a(5.5992142733884975e-05)),(to_sfixed_a(-6.741791003150865e-05)),(to_sfixed_a(6.97110499459086e-06)),(to_sfixed_a(4.1726092604221776e-05)),(to_sfixed_a(-1.1585445463424549e-05)),(to_sfixed_a(8.933011122280732e-05)),(to_sfixed_a(6.45286199869588e-05)),(to_sfixed_a(-7.637042290298268e-05)),(to_sfixed_a(1.8681317669688724e-05)),(to_sfixed_a(2.8512424250948243e-05)),(to_sfixed_a(-7.68165773479268e-05)),(to_sfixed_a(-2.933614086941816e-05)),(to_sfixed_a(-3.461191226961091e-06)),(to_sfixed_a(-3.8057991332607344e-05)),(to_sfixed_a(5.226629218668677e-05)),(to_sfixed_a(6.727692380081862e-05)),(to_sfixed_a(-2.060167935269419e-05)),(to_sfixed_a(-5.199105362407863e-05)),(to_sfixed_a(2.017093038375606e-06)),(to_sfixed_a(-8.729570254217833e-06)),(to_sfixed_a(-6.516427674796432e-05)),(to_sfixed_a(4.403336060931906e-05)),(to_sfixed_a(-7.141254172893241e-05)),(to_sfixed_a(5.4904798162169755e-05)),(to_sfixed_a(-2.96571397484513e-05)),(to_sfixed_a(3.0184270144673064e-05)),(to_sfixed_a(-2.6920677555608563e-05)),(to_sfixed_a(3.6733072192873806e-06)),(to_sfixed_a(7.154476043069735e-05)),(to_sfixed_a(-7.159139204304665e-05)),(to_sfixed_a(-0.00012142791820224375)),(to_sfixed_a(2.380688783887308e-05)),(to_sfixed_a(-3.444226967985742e-05)),(to_sfixed_a(6.832185317762196e-05)));

    constant weight_n1_241 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.3456396162509918)),(to_sfixed_a(-0.07250429689884186)),(to_sfixed_a(0.15432465076446533)),(to_sfixed_a(-0.09336686134338379)),(to_sfixed_a(-0.2980820834636688)),(to_sfixed_a(0.06556405127048492)),(to_sfixed_a(0.06782630831003189)),(to_sfixed_a(-0.11763327568769455)),(to_sfixed_a(-0.10810911655426025)),(to_sfixed_a(0.033389415591955185)),(to_sfixed_a(-0.034412868320941925)),(to_sfixed_a(0.1368841528892517)),(to_sfixed_a(0.0610562302172184)),(to_sfixed_a(0.09138597548007965)),(to_sfixed_a(-0.0030685153324157)),(to_sfixed_a(0.04896972328424454)),(to_sfixed_a(-0.09323985129594803)),(to_sfixed_a(0.093390092253685)),(to_sfixed_a(-0.12115160375833511)),(to_sfixed_a(0.02040836215019226)),(to_sfixed_a(-0.0371287502348423)),(to_sfixed_a(-0.010940918698906898)),(to_sfixed_a(0.021609045565128326)),(to_sfixed_a(-0.1718764454126358)),(to_sfixed_a(0.04239104315638542)),(to_sfixed_a(0.08994308114051819)),(to_sfixed_a(-0.14153748750686646)),(to_sfixed_a(-0.14572545886039734)),(to_sfixed_a(-0.06381065398454666)),(to_sfixed_a(-0.08590502291917801)),(to_sfixed_a(-0.02140686847269535)),(to_sfixed_a(-0.1349271982908249)),(to_sfixed_a(-0.002568613039329648)),(to_sfixed_a(-0.20469780266284943)),(to_sfixed_a(-0.1118248701095581)),(to_sfixed_a(-0.06092549487948418)),(to_sfixed_a(0.03548315539956093)),(to_sfixed_a(0.15239010751247406)));

    constant weight_n1_242 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.01422665175050497)),(to_sfixed_a(-2.3045244233799167e-05)),(to_sfixed_a(-5.093804247735534e-06)),(to_sfixed_a(-6.019173451932147e-05)),(to_sfixed_a(8.745023478695657e-06)),(to_sfixed_a(4.920989886159077e-05)),(to_sfixed_a(9.920840966515243e-06)),(to_sfixed_a(-1.4061984984437004e-05)),(to_sfixed_a(6.683372339466587e-05)),(to_sfixed_a(1.6844784113345668e-05)),(to_sfixed_a(8.200723823392764e-05)),(to_sfixed_a(-2.8117088731960393e-05)),(to_sfixed_a(6.234708416741341e-05)),(to_sfixed_a(8.73029712238349e-05)),(to_sfixed_a(-4.2994219256797805e-05)),(to_sfixed_a(-1.5369119864772074e-05)),(to_sfixed_a(-6.878799467813224e-05)),(to_sfixed_a(-2.4303586542373523e-05)),(to_sfixed_a(9.864461026154459e-05)),(to_sfixed_a(2.9857355912099592e-05)),(to_sfixed_a(2.922806015703827e-05)),(to_sfixed_a(-1.8284270481672138e-05)),(to_sfixed_a(1.1800049833254889e-05)),(to_sfixed_a(-8.249135134974495e-05)),(to_sfixed_a(-3.356353772687726e-05)),(to_sfixed_a(-8.468786109006032e-05)),(to_sfixed_a(2.811651211231947e-05)),(to_sfixed_a(-1.580635944264941e-05)),(to_sfixed_a(-1.3916208445152733e-05)),(to_sfixed_a(4.537427957984619e-05)),(to_sfixed_a(1.9597333448473364e-05)),(to_sfixed_a(-6.043140820111148e-05)),(to_sfixed_a(-6.481598393293098e-05)),(to_sfixed_a(-1.1292901035631076e-05)),(to_sfixed_a(-4.921802246826701e-05)),(to_sfixed_a(-2.298247636645101e-05)),(to_sfixed_a(-7.896963506937027e-05)),(to_sfixed_a(-2.144485551980324e-05)));

    constant weight_n1_243 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.0017546748276799917)),(to_sfixed_a(-0.05215568095445633)),(to_sfixed_a(0.06783121824264526)),(to_sfixed_a(-0.044513486325740814)),(to_sfixed_a(-0.03219150751829147)),(to_sfixed_a(-0.0838824212551117)),(to_sfixed_a(-0.1369992047548294)),(to_sfixed_a(-0.17051862180233002)),(to_sfixed_a(-0.09912218898534775)),(to_sfixed_a(-0.0750703513622284)),(to_sfixed_a(-0.09259271621704102)),(to_sfixed_a(0.028274361044168472)),(to_sfixed_a(0.09466245770454407)),(to_sfixed_a(0.08903595805168152)),(to_sfixed_a(0.06943882256746292)),(to_sfixed_a(-0.03003312088549137)),(to_sfixed_a(-0.20818372070789337)),(to_sfixed_a(0.07061270624399185)),(to_sfixed_a(-0.18667520582675934)),(to_sfixed_a(0.015719098970294)),(to_sfixed_a(-0.006756388116627932)),(to_sfixed_a(-0.048010632395744324)),(to_sfixed_a(-0.012424606829881668)),(to_sfixed_a(-0.03364245593547821)),(to_sfixed_a(-0.1133282333612442)),(to_sfixed_a(0.06415529549121857)),(to_sfixed_a(0.03639136254787445)),(to_sfixed_a(-0.11488030105829239)),(to_sfixed_a(-0.08712903410196304)),(to_sfixed_a(-0.10038385540246964)),(to_sfixed_a(0.04068822041153908)),(to_sfixed_a(0.00027663158834911883)),(to_sfixed_a(-0.15110857784748077)),(to_sfixed_a(0.04312599077820778)),(to_sfixed_a(-0.20561262965202332)),(to_sfixed_a(0.014039256609976292)),(to_sfixed_a(0.20178598165512085)),(to_sfixed_a(-0.1684211939573288)));

    constant weight_n1_244 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.11834007501602173)),(to_sfixed_a(-0.0028027743101119995)),(to_sfixed_a(-0.036950550973415375)),(to_sfixed_a(-0.0450618751347065)),(to_sfixed_a(-0.0423567071557045)),(to_sfixed_a(0.08116867393255234)),(to_sfixed_a(0.011411327868700027)),(to_sfixed_a(-0.06370092183351517)),(to_sfixed_a(0.008684339001774788)),(to_sfixed_a(-0.01316589955240488)),(to_sfixed_a(0.02244352176785469)),(to_sfixed_a(-0.04532739520072937)),(to_sfixed_a(-0.012364190071821213)),(to_sfixed_a(-0.059261538088321686)),(to_sfixed_a(0.1793517768383026)),(to_sfixed_a(0.04376061260700226)),(to_sfixed_a(-0.03852101415395737)),(to_sfixed_a(0.009109343402087688)),(to_sfixed_a(0.12172253429889679)),(to_sfixed_a(0.022238465026021004)),(to_sfixed_a(-0.1250474601984024)),(to_sfixed_a(0.05694492161273956)),(to_sfixed_a(-0.06642653793096542)),(to_sfixed_a(-0.06792642176151276)),(to_sfixed_a(-0.0031944916117936373)),(to_sfixed_a(-0.036326225847005844)),(to_sfixed_a(0.047845035791397095)),(to_sfixed_a(0.05863644555211067)),(to_sfixed_a(-0.009012183174490929)),(to_sfixed_a(0.01062572468072176)),(to_sfixed_a(0.030195461586117744)),(to_sfixed_a(0.08298584073781967)),(to_sfixed_a(0.015552929602563381)),(to_sfixed_a(-0.055373698472976685)),(to_sfixed_a(0.020982282236218452)),(to_sfixed_a(-0.009527844376862049)),(to_sfixed_a(0.03971979767084122)),(to_sfixed_a(-0.062228526920080185)));

    constant weight_n1_245 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.14216196537017822)),(to_sfixed_a(-0.0666775032877922)),(to_sfixed_a(0.21783101558685303)),(to_sfixed_a(0.05558232218027115)),(to_sfixed_a(0.17416392266750336)),(to_sfixed_a(0.3003716766834259)),(to_sfixed_a(0.17639727890491486)),(to_sfixed_a(0.22704526782035828)),(to_sfixed_a(0.08982249349355698)),(to_sfixed_a(-0.1646445095539093)),(to_sfixed_a(-0.08307139575481415)),(to_sfixed_a(-0.2530965507030487)),(to_sfixed_a(-0.09399648010730743)),(to_sfixed_a(0.05072346329689026)),(to_sfixed_a(0.0425010584294796)),(to_sfixed_a(0.03366614878177643)),(to_sfixed_a(-0.12599076330661774)),(to_sfixed_a(0.1648399382829666)),(to_sfixed_a(0.0016102828085422516)),(to_sfixed_a(0.038398221135139465)),(to_sfixed_a(0.06990903615951538)),(to_sfixed_a(-0.03912322223186493)),(to_sfixed_a(0.05024236440658569)),(to_sfixed_a(-0.016770385205745697)),(to_sfixed_a(0.020018599927425385)),(to_sfixed_a(-0.19767601788043976)),(to_sfixed_a(0.021780991926789284)),(to_sfixed_a(-0.04585632309317589)),(to_sfixed_a(0.043217018246650696)),(to_sfixed_a(-0.06935960054397583)),(to_sfixed_a(-0.18401704728603363)),(to_sfixed_a(0.15479102730751038)),(to_sfixed_a(-0.20268404483795166)),(to_sfixed_a(-0.07222986221313477)),(to_sfixed_a(0.0022611019667237997)),(to_sfixed_a(0.08790259808301926)),(to_sfixed_a(-0.06703346222639084)),(to_sfixed_a(-0.07602924853563309)));

    constant weight_n1_246 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.3781183362007141)),(to_sfixed_a(0.06473655253648758)),(to_sfixed_a(-0.19298851490020752)),(to_sfixed_a(-0.11279162764549255)),(to_sfixed_a(0.20296567678451538)),(to_sfixed_a(0.04645824059844017)),(to_sfixed_a(0.020787809044122696)),(to_sfixed_a(0.05926864221692085)),(to_sfixed_a(-0.11040893942117691)),(to_sfixed_a(-0.24519453942775726)),(to_sfixed_a(-0.05638844519853592)),(to_sfixed_a(-0.032694991677999496)),(to_sfixed_a(0.1965387463569641)),(to_sfixed_a(0.04788270965218544)),(to_sfixed_a(0.061827320605516434)),(to_sfixed_a(-0.04315727576613426)),(to_sfixed_a(-0.20126862823963165)),(to_sfixed_a(-0.07136039435863495)),(to_sfixed_a(0.0454377681016922)),(to_sfixed_a(0.17704181373119354)),(to_sfixed_a(-0.24314969778060913)),(to_sfixed_a(0.19707055389881134)),(to_sfixed_a(-0.014695807360112667)),(to_sfixed_a(0.036966267973184586)),(to_sfixed_a(0.29569658637046814)),(to_sfixed_a(0.004461788572371006)),(to_sfixed_a(-0.14915089309215546)),(to_sfixed_a(-0.2882896065711975)),(to_sfixed_a(-0.07580222189426422)),(to_sfixed_a(0.06392835080623627)),(to_sfixed_a(-0.030965497717261314)),(to_sfixed_a(-0.017866726964712143)),(to_sfixed_a(0.11802976578474045)),(to_sfixed_a(0.1806412637233734)),(to_sfixed_a(-0.1130947396159172)),(to_sfixed_a(0.14597901701927185)),(to_sfixed_a(0.09828009456396103)),(to_sfixed_a(0.09354159981012344)));

    constant weight_n1_247 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.06451129168272018)),(to_sfixed_a(1.880680247268174e-05)),(to_sfixed_a(5.8216719480697066e-05)),(to_sfixed_a(-4.090323727723444e-06)),(to_sfixed_a(1.736521335260477e-05)),(to_sfixed_a(-3.898415889125317e-05)),(to_sfixed_a(3.211406510672532e-05)),(to_sfixed_a(2.9873492167098448e-05)),(to_sfixed_a(-4.354498742031865e-05)),(to_sfixed_a(-6.490492523880675e-05)),(to_sfixed_a(6.827590550528839e-05)),(to_sfixed_a(-2.6063155019073747e-05)),(to_sfixed_a(2.269725882797502e-05)),(to_sfixed_a(2.1069534341222607e-05)),(to_sfixed_a(-5.006591891287826e-05)),(to_sfixed_a(-2.6389518097857945e-05)),(to_sfixed_a(-2.402340942353476e-05)),(to_sfixed_a(-2.999442040163558e-05)),(to_sfixed_a(-3.049960832868237e-05)),(to_sfixed_a(-5.878696538275108e-05)),(to_sfixed_a(3.0888566016074037e-06)),(to_sfixed_a(0.00010537595517234877)),(to_sfixed_a(-3.606654718169011e-05)),(to_sfixed_a(-7.0807000156492e-05)),(to_sfixed_a(-4.80980052088853e-05)),(to_sfixed_a(-3.758721868507564e-05)),(to_sfixed_a(-5.6538385251769796e-05)),(to_sfixed_a(6.197974926180905e-06)),(to_sfixed_a(-3.805350934271701e-05)),(to_sfixed_a(3.099089008173905e-05)),(to_sfixed_a(3.898250724887475e-06)),(to_sfixed_a(-2.2994196115178056e-05)),(to_sfixed_a(-9.149056495516561e-06)),(to_sfixed_a(7.005708903307095e-05)),(to_sfixed_a(-3.7362515286076814e-05)),(to_sfixed_a(3.424005626584403e-05)),(to_sfixed_a(-2.266779847559519e-05)),(to_sfixed_a(4.2525083699729294e-05)));

    constant weight_n1_248 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.14909620583057404)),(to_sfixed_a(0.00833887793123722)),(to_sfixed_a(-0.02060248702764511)),(to_sfixed_a(0.0131844412535429)),(to_sfixed_a(0.06528106331825256)),(to_sfixed_a(-0.09022417664527893)),(to_sfixed_a(-0.06351406127214432)),(to_sfixed_a(0.046895597130060196)),(to_sfixed_a(0.024099519476294518)),(to_sfixed_a(-0.03758816048502922)),(to_sfixed_a(0.01889009401202202)),(to_sfixed_a(-0.04204057157039642)),(to_sfixed_a(-0.00934368371963501)),(to_sfixed_a(-0.022445615381002426)),(to_sfixed_a(-0.004105754196643829)),(to_sfixed_a(-0.021098973229527473)),(to_sfixed_a(0.027839845046401024)),(to_sfixed_a(-0.09970701485872269)),(to_sfixed_a(0.04382454976439476)),(to_sfixed_a(-0.034396976232528687)),(to_sfixed_a(-0.0188850499689579)),(to_sfixed_a(-0.00037319454713724554)),(to_sfixed_a(-0.019997894763946533)),(to_sfixed_a(0.024352148175239563)),(to_sfixed_a(-0.02412502095103264)),(to_sfixed_a(0.04809577390551567)),(to_sfixed_a(0.01479173731058836)),(to_sfixed_a(0.055059973150491714)),(to_sfixed_a(-0.0005280945915728807)),(to_sfixed_a(0.016736513003706932)),(to_sfixed_a(0.038012776523828506)),(to_sfixed_a(-0.003274130867794156)),(to_sfixed_a(0.1111956313252449)),(to_sfixed_a(-0.009596971794962883)),(to_sfixed_a(0.13423344492912292)),(to_sfixed_a(-0.04885338246822357)),(to_sfixed_a(0.023597750812768936)),(to_sfixed_a(-0.052532706409692764)));

    constant weight_n1_249 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.23758837580680847)),(to_sfixed_a(0.0016473239520564675)),(to_sfixed_a(0.0008094183285720646)),(to_sfixed_a(0.013868667185306549)),(to_sfixed_a(-0.0028960632625967264)),(to_sfixed_a(0.001829120796173811)),(to_sfixed_a(-0.002895219950005412)),(to_sfixed_a(-0.002243733499199152)),(to_sfixed_a(0.007832536473870277)),(to_sfixed_a(0.009284342639148235)),(to_sfixed_a(0.006789674051105976)),(to_sfixed_a(0.016874445602297783)),(to_sfixed_a(-0.00573553703725338)),(to_sfixed_a(-0.012512974441051483)),(to_sfixed_a(0.001693323371000588)),(to_sfixed_a(0.006808658130466938)),(to_sfixed_a(-0.011580226942896843)),(to_sfixed_a(0.0016066712560132146)),(to_sfixed_a(0.014963982626795769)),(to_sfixed_a(-0.013203155249357224)),(to_sfixed_a(0.009599681943655014)),(to_sfixed_a(0.0005576141411438584)),(to_sfixed_a(-0.010161478072404861)),(to_sfixed_a(-0.0032764447387307882)),(to_sfixed_a(0.011783384718000889)),(to_sfixed_a(0.00487313698977232)),(to_sfixed_a(0.006556130014359951)),(to_sfixed_a(-0.0029880960937589407)),(to_sfixed_a(-0.015815021470189095)),(to_sfixed_a(-0.004860589746385813)),(to_sfixed_a(0.019839175045490265)),(to_sfixed_a(-0.003707817057147622)),(to_sfixed_a(0.004368945024907589)),(to_sfixed_a(9.983725612983108e-05)),(to_sfixed_a(-0.013827026821672916)),(to_sfixed_a(-0.005049613770097494)),(to_sfixed_a(0.0032099036034196615)),(to_sfixed_a(0.006178541574627161)));

    constant weight_n1_250 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.011148190125823021)),(to_sfixed_a(5.431669251265703e-06)),(to_sfixed_a(-3.170316631440073e-05)),(to_sfixed_a(-1.5503719623666257e-05)),(to_sfixed_a(-4.079308928339742e-05)),(to_sfixed_a(2.3253307517734356e-05)),(to_sfixed_a(-5.974019131826935e-06)),(to_sfixed_a(-1.3925746316090226e-05)),(to_sfixed_a(-4.9957936425926164e-05)),(to_sfixed_a(-3.320462565170601e-05)),(to_sfixed_a(-4.377641744213179e-05)),(to_sfixed_a(-2.254352148156613e-05)),(to_sfixed_a(-4.621616244548932e-05)),(to_sfixed_a(-7.516821642639115e-05)),(to_sfixed_a(-5.2039373258594424e-05)),(to_sfixed_a(-5.287980457069352e-05)),(to_sfixed_a(-2.645827225933317e-05)),(to_sfixed_a(1.9946566681028344e-05)),(to_sfixed_a(2.3008144125924446e-05)),(to_sfixed_a(-7.460678898496553e-05)),(to_sfixed_a(-2.382749880780466e-05)),(to_sfixed_a(6.342976121231914e-05)),(to_sfixed_a(8.4053332102485e-05)),(to_sfixed_a(-7.734106475254521e-05)),(to_sfixed_a(1.8931688828160986e-05)),(to_sfixed_a(6.11812574788928e-05)),(to_sfixed_a(-1.6319510905304924e-05)),(to_sfixed_a(-7.012479909462854e-05)),(to_sfixed_a(7.368065416812897e-05)),(to_sfixed_a(-8.796738256933168e-05)),(to_sfixed_a(9.265146945836022e-05)),(to_sfixed_a(2.795630507534952e-06)),(to_sfixed_a(1.3650320397573523e-05)),(to_sfixed_a(9.138521818385925e-06)),(to_sfixed_a(-5.581954610534012e-05)),(to_sfixed_a(-4.6211174776544794e-05)),(to_sfixed_a(-5.816928023705259e-05)),(to_sfixed_a(-5.1685103244381025e-05)));

    constant weight_n1_251 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.4111463129520416)),(to_sfixed_a(-0.017550483345985413)),(to_sfixed_a(0.015372354537248611)),(to_sfixed_a(0.0035856422036886215)),(to_sfixed_a(-0.03343158960342407)),(to_sfixed_a(-0.0034839536529034376)),(to_sfixed_a(0.021802853792905807)),(to_sfixed_a(-0.023620491847395897)),(to_sfixed_a(0.025706974789500237)),(to_sfixed_a(-0.009884594939649105)),(to_sfixed_a(-0.03969685360789299)),(to_sfixed_a(-0.026480525732040405)),(to_sfixed_a(-0.03462688997387886)),(to_sfixed_a(-0.05328044295310974)),(to_sfixed_a(0.004536386579275131)),(to_sfixed_a(0.0014328783145174384)),(to_sfixed_a(-0.07484563440084457)),(to_sfixed_a(0.0850720927119255)),(to_sfixed_a(0.07141714543104172)),(to_sfixed_a(0.09166313707828522)),(to_sfixed_a(-0.007641668897122145)),(to_sfixed_a(-0.10217326879501343)),(to_sfixed_a(-0.011928051710128784)),(to_sfixed_a(-0.0402451828122139)),(to_sfixed_a(0.011018304154276848)),(to_sfixed_a(0.08665785193443298)),(to_sfixed_a(-0.02807304635643959)),(to_sfixed_a(-0.015096492134034634)),(to_sfixed_a(-0.01496098842471838)),(to_sfixed_a(0.061474088579416275)),(to_sfixed_a(0.0017500050598755479)),(to_sfixed_a(-0.00805654190480709)),(to_sfixed_a(-0.03204480558633804)),(to_sfixed_a(0.009140405803918839)),(to_sfixed_a(0.06082088127732277)),(to_sfixed_a(0.07510961592197418)),(to_sfixed_a(0.018466288223862648)),(to_sfixed_a(0.026610152795910835)));

    constant weight_n1_252 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.09640305489301682)),(to_sfixed_a(-4.047319453093223e-05)),(to_sfixed_a(-1.2828415492549539e-05)),(to_sfixed_a(2.1895628378842957e-05)),(to_sfixed_a(-2.7316677005728707e-05)),(to_sfixed_a(-3.155375816277228e-05)),(to_sfixed_a(-5.620555043606146e-07)),(to_sfixed_a(-4.119388177059591e-05)),(to_sfixed_a(-1.849690670496784e-05)),(to_sfixed_a(-6.04684064455796e-05)),(to_sfixed_a(-3.465142071945593e-05)),(to_sfixed_a(-3.1912026315694675e-05)),(to_sfixed_a(-8.503048593411222e-05)),(to_sfixed_a(-4.488077320274897e-05)),(to_sfixed_a(3.2204625313170254e-06)),(to_sfixed_a(3.5625787859316915e-05)),(to_sfixed_a(-2.9823489967384376e-05)),(to_sfixed_a(6.269891309784725e-05)),(to_sfixed_a(-6.279900117078796e-05)),(to_sfixed_a(2.221162139903754e-05)),(to_sfixed_a(1.845855513238348e-05)),(to_sfixed_a(1.0757927157101221e-05)),(to_sfixed_a(3.856771218124777e-05)),(to_sfixed_a(8.105995220830664e-05)),(to_sfixed_a(-2.215228414570447e-05)),(to_sfixed_a(-9.961213800124824e-05)),(to_sfixed_a(-5.130687713972293e-05)),(to_sfixed_a(1.7378753909724765e-05)),(to_sfixed_a(4.046914182254113e-05)),(to_sfixed_a(8.907976734917611e-06)),(to_sfixed_a(-3.282081161160022e-05)),(to_sfixed_a(7.544736945419572e-06)),(to_sfixed_a(-5.148244963493198e-05)),(to_sfixed_a(2.0996109014959075e-05)),(to_sfixed_a(1.735566183924675e-05)),(to_sfixed_a(1.565248385304585e-05)),(to_sfixed_a(-2.0964318537153304e-05)),(to_sfixed_a(2.8540902349050157e-05)));

    constant weight_n1_253 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.013821960426867008)),(to_sfixed_a(-0.018037350848317146)),(to_sfixed_a(-0.00017117972311098129)),(to_sfixed_a(-0.005287542007863522)),(to_sfixed_a(0.00655452162027359)),(to_sfixed_a(-0.001470257993787527)),(to_sfixed_a(0.0006691787857562304)),(to_sfixed_a(0.015910709276795387)),(to_sfixed_a(-0.027345813810825348)),(to_sfixed_a(0.0019589518196880817)),(to_sfixed_a(0.04393209144473076)),(to_sfixed_a(-0.016823336482048035)),(to_sfixed_a(0.0012505479389801621)),(to_sfixed_a(0.022263681516051292)),(to_sfixed_a(0.012187103740870953)),(to_sfixed_a(-0.021591132506728172)),(to_sfixed_a(0.021229302510619164)),(to_sfixed_a(0.0008859615190885961)),(to_sfixed_a(-0.0059671299532055855)),(to_sfixed_a(0.01572553813457489)),(to_sfixed_a(-0.0632915198802948)),(to_sfixed_a(-0.013690117746591568)),(to_sfixed_a(-0.007757639512419701)),(to_sfixed_a(-0.011335432529449463)),(to_sfixed_a(0.023377085104584694)),(to_sfixed_a(0.0052634975872933865)),(to_sfixed_a(0.016745485365390778)),(to_sfixed_a(-0.026492012664675713)),(to_sfixed_a(-0.0006873037200421095)),(to_sfixed_a(0.001862932462245226)),(to_sfixed_a(-0.015345372259616852)),(to_sfixed_a(0.014637899585068226)),(to_sfixed_a(-0.019864030182361603)),(to_sfixed_a(-0.02127041295170784)),(to_sfixed_a(-0.026609497144818306)),(to_sfixed_a(-0.04184893146157265)),(to_sfixed_a(-0.019745593890547752)),(to_sfixed_a(-0.009945741854608059)));

    constant weight_n1_254 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.10084685683250427)),(to_sfixed_a(-0.044784318655729294)),(to_sfixed_a(0.10916507989168167)),(to_sfixed_a(-0.003875304479151964)),(to_sfixed_a(0.0392325222492218)),(to_sfixed_a(-0.06721488386392593)),(to_sfixed_a(-0.03880859166383743)),(to_sfixed_a(0.06968317925930023)),(to_sfixed_a(-0.04986365884542465)),(to_sfixed_a(-0.028671756386756897)),(to_sfixed_a(0.19806444644927979)),(to_sfixed_a(-0.040136322379112244)),(to_sfixed_a(0.04001254960894585)),(to_sfixed_a(0.12328445911407471)),(to_sfixed_a(0.06747626513242722)),(to_sfixed_a(-0.12120787054300308)),(to_sfixed_a(0.1159219816327095)),(to_sfixed_a(0.034094735980033875)),(to_sfixed_a(-0.062460269778966904)),(to_sfixed_a(0.04044393450021744)),(to_sfixed_a(-0.28455406427383423)),(to_sfixed_a(-0.06566653400659561)),(to_sfixed_a(0.015631526708602905)),(to_sfixed_a(-0.26958754658699036)),(to_sfixed_a(0.1603538990020752)),(to_sfixed_a(0.07536707818508148)),(to_sfixed_a(0.040599703788757324)),(to_sfixed_a(-0.07458633184432983)),(to_sfixed_a(0.1280173659324646)),(to_sfixed_a(0.013960999436676502)),(to_sfixed_a(-0.1386909931898117)),(to_sfixed_a(-0.08869699388742447)),(to_sfixed_a(-0.0322686992585659)),(to_sfixed_a(-0.03155355527997017)),(to_sfixed_a(-0.034205079078674316)),(to_sfixed_a(-0.20876477658748627)),(to_sfixed_a(-0.2189236581325531)),(to_sfixed_a(-0.12340577691793442)));

    constant weight_n1_255 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.2437620759010315)),(to_sfixed_a(0.07813221216201782)),(to_sfixed_a(-0.037888653576374054)),(to_sfixed_a(0.0384349450469017)),(to_sfixed_a(0.024105211719870567)),(to_sfixed_a(-0.06781723350286484)),(to_sfixed_a(0.06272082030773163)),(to_sfixed_a(-0.047589946538209915)),(to_sfixed_a(-0.05354980751872063)),(to_sfixed_a(0.08265293389558792)),(to_sfixed_a(-0.07900810241699219)),(to_sfixed_a(-0.11568865925073624)),(to_sfixed_a(-0.038661181926727295)),(to_sfixed_a(0.02561396360397339)),(to_sfixed_a(0.013541429303586483)),(to_sfixed_a(0.10887721180915833)),(to_sfixed_a(-0.203040212392807)),(to_sfixed_a(-0.0231606625020504)),(to_sfixed_a(0.021940868347883224)),(to_sfixed_a(-0.10710374265909195)),(to_sfixed_a(-0.04999411106109619)),(to_sfixed_a(0.08569775521755219)),(to_sfixed_a(0.016768014058470726)),(to_sfixed_a(-0.08191045373678207)),(to_sfixed_a(0.09528712928295135)),(to_sfixed_a(-0.08902017772197723)),(to_sfixed_a(0.18396610021591187)),(to_sfixed_a(0.08144637197256088)),(to_sfixed_a(0.029615504667162895)),(to_sfixed_a(0.12137436121702194)),(to_sfixed_a(0.04666982218623161)),(to_sfixed_a(-0.01717352122068405)),(to_sfixed_a(0.023686029016971588)),(to_sfixed_a(-0.026806164532899857)),(to_sfixed_a(-0.02707388810813427)),(to_sfixed_a(-0.23315463960170746)),(to_sfixed_a(-0.1981523185968399)),(to_sfixed_a(0.044803354889154434)));

    constant weight_n1_256 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.1262165755033493)),(to_sfixed_a(-1.1623184946074616e-05)),(to_sfixed_a(-9.392118954565376e-06)),(to_sfixed_a(-3.419159838813357e-05)),(to_sfixed_a(1.0530236977501772e-05)),(to_sfixed_a(-4.075668766745366e-05)),(to_sfixed_a(1.1290185284451582e-05)),(to_sfixed_a(4.1052146116271615e-05)),(to_sfixed_a(2.5368974092998542e-05)),(to_sfixed_a(4.19517164118588e-05)),(to_sfixed_a(-2.1241119156911736e-06)),(to_sfixed_a(1.3181410395191051e-05)),(to_sfixed_a(1.8597922462504357e-05)),(to_sfixed_a(-3.519144229358062e-05)),(to_sfixed_a(-2.628214133437723e-05)),(to_sfixed_a(-4.466877362574451e-05)),(to_sfixed_a(-1.8278296920470893e-05)),(to_sfixed_a(-9.283461258746684e-05)),(to_sfixed_a(3.813018702203408e-05)),(to_sfixed_a(2.3784788936609402e-05)),(to_sfixed_a(3.190897041349672e-05)),(to_sfixed_a(-3.3935571991605684e-05)),(to_sfixed_a(-4.801210525329225e-05)),(to_sfixed_a(1.3260570085549261e-05)),(to_sfixed_a(5.3657626267522573e-05)),(to_sfixed_a(-1.0871531230804976e-05)),(to_sfixed_a(5.679640526068397e-05)),(to_sfixed_a(6.8750350692425855e-06)),(to_sfixed_a(1.7391585060977377e-05)),(to_sfixed_a(3.4565735404612496e-05)),(to_sfixed_a(-8.718201570445672e-05)),(to_sfixed_a(9.910442167893052e-05)),(to_sfixed_a(-2.804011819534935e-05)),(to_sfixed_a(1.0275873592036078e-06)),(to_sfixed_a(2.3317539671552368e-05)),(to_sfixed_a(4.1949053411372006e-05)),(to_sfixed_a(-2.4233790099970065e-05)),(to_sfixed_a(1.1349558093343148e-07)));

    constant weight_n1_257 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.027986373752355576)),(to_sfixed_a(2.590182157291565e-05)),(to_sfixed_a(1.6635360111649788e-07)),(to_sfixed_a(5.134930324857123e-05)),(to_sfixed_a(2.741788193816319e-06)),(to_sfixed_a(5.368249276216375e-07)),(to_sfixed_a(4.176998118055053e-05)),(to_sfixed_a(7.647771781194024e-06)),(to_sfixed_a(-1.686273026280105e-05)),(to_sfixed_a(5.625559060717933e-05)),(to_sfixed_a(4.1709707147674635e-05)),(to_sfixed_a(-2.5633744371589273e-05)),(to_sfixed_a(-3.270692832302302e-05)),(to_sfixed_a(-3.855975955957547e-05)),(to_sfixed_a(-2.2535095922648907e-05)),(to_sfixed_a(6.137809396022931e-05)),(to_sfixed_a(1.3969237443234306e-05)),(to_sfixed_a(-3.643628224381246e-05)),(to_sfixed_a(1.239462108060252e-05)),(to_sfixed_a(5.482721462612972e-06)),(to_sfixed_a(3.4358265565970214e-06)),(to_sfixed_a(9.991304978029802e-05)),(to_sfixed_a(-5.766067624790594e-05)),(to_sfixed_a(2.7032021534978412e-05)),(to_sfixed_a(-1.4632665624958463e-05)),(to_sfixed_a(0.00010854643915081397)),(to_sfixed_a(1.4006699530000333e-05)),(to_sfixed_a(-4.331845775595866e-05)),(to_sfixed_a(0.00010746549378382042)),(to_sfixed_a(1.3488787772075739e-05)),(to_sfixed_a(-1.7308137103100307e-05)),(to_sfixed_a(-3.465424379101023e-05)),(to_sfixed_a(3.145889422739856e-05)),(to_sfixed_a(6.0620795920840465e-06)),(to_sfixed_a(1.6807560314191505e-05)),(to_sfixed_a(3.524444400682114e-05)),(to_sfixed_a(-4.331956006353721e-05)),(to_sfixed_a(-2.7033578589907847e-05)));

    constant weight_n1_258 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.054689355194568634)),(to_sfixed_a(-0.027271559461951256)),(to_sfixed_a(0.03203978016972542)),(to_sfixed_a(-0.18231286108493805)),(to_sfixed_a(-0.024215437471866608)),(to_sfixed_a(-0.15196000039577484)),(to_sfixed_a(0.1131240501999855)),(to_sfixed_a(0.1685912013053894)),(to_sfixed_a(0.058598265051841736)),(to_sfixed_a(-0.03122248500585556)),(to_sfixed_a(-0.11625384539365768)),(to_sfixed_a(0.03098328411579132)),(to_sfixed_a(-0.08782144635915756)),(to_sfixed_a(-0.0009226123802363873)),(to_sfixed_a(-0.026666032150387764)),(to_sfixed_a(-0.04627545177936554)),(to_sfixed_a(0.008196712471544743)),(to_sfixed_a(-0.0035775487776845694)),(to_sfixed_a(-0.0035051023587584496)),(to_sfixed_a(0.010789060033857822)),(to_sfixed_a(-0.011808514595031738)),(to_sfixed_a(-0.02622126415371895)),(to_sfixed_a(0.05082029476761818)),(to_sfixed_a(-0.016055718064308167)),(to_sfixed_a(0.04222101718187332)),(to_sfixed_a(-0.04547806829214096)),(to_sfixed_a(-0.018394239246845245)),(to_sfixed_a(0.06236277148127556)),(to_sfixed_a(-0.01979655586183071)),(to_sfixed_a(-0.052947547286748886)),(to_sfixed_a(0.06842146068811417)),(to_sfixed_a(-0.046338554471731186)),(to_sfixed_a(0.07687831670045853)),(to_sfixed_a(0.04932396113872528)),(to_sfixed_a(0.02418668568134308)),(to_sfixed_a(0.019949959591031075)),(to_sfixed_a(-0.07426206767559052)),(to_sfixed_a(0.011331175453960896)));

    constant weight_n1_259 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.10357283800840378)),(to_sfixed_a(-1.5809342585271224e-05)),(to_sfixed_a(3.500224556773901e-05)),(to_sfixed_a(-1.0001125474445871e-06)),(to_sfixed_a(-4.104826075490564e-05)),(to_sfixed_a(4.527834607870318e-05)),(to_sfixed_a(-6.174063310027122e-05)),(to_sfixed_a(-9.195672646455932e-06)),(to_sfixed_a(-3.4312477055209456e-06)),(to_sfixed_a(-2.155034053430427e-05)),(to_sfixed_a(-1.4000376722833607e-05)),(to_sfixed_a(-2.553475678723771e-05)),(to_sfixed_a(4.404597348184325e-05)),(to_sfixed_a(-2.4579123419243842e-05)),(to_sfixed_a(-6.333828059723601e-05)),(to_sfixed_a(1.9089315173914656e-05)),(to_sfixed_a(-6.29435307928361e-05)),(to_sfixed_a(-0.00010514597670407966)),(to_sfixed_a(4.773389809997752e-05)),(to_sfixed_a(-2.54630867857486e-05)),(to_sfixed_a(9.813769429456443e-05)),(to_sfixed_a(3.844229468086269e-06)),(to_sfixed_a(3.083820774918422e-05)),(to_sfixed_a(-0.00011803807137766853)),(to_sfixed_a(-9.09976297407411e-05)),(to_sfixed_a(4.9700087402015924e-05)),(to_sfixed_a(3.950787868234329e-05)),(to_sfixed_a(-5.2405699534574524e-05)),(to_sfixed_a(-4.042496584588662e-05)),(to_sfixed_a(3.2973854104056954e-05)),(to_sfixed_a(-2.72896395472344e-05)),(to_sfixed_a(2.0907747966703027e-05)),(to_sfixed_a(-3.214574826415628e-05)),(to_sfixed_a(3.3482185699540423e-06)),(to_sfixed_a(-2.0651776139857247e-05)),(to_sfixed_a(3.394480881979689e-05)),(to_sfixed_a(-4.952896051690914e-05)),(to_sfixed_a(-5.738185063819401e-05)));

    constant weight_n1_260 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.17119969427585602)),(to_sfixed_a(-0.014418101869523525)),(to_sfixed_a(-0.04777907207608223)),(to_sfixed_a(-0.014273270033299923)),(to_sfixed_a(-0.056766606867313385)),(to_sfixed_a(0.052483510226011276)),(to_sfixed_a(-0.08139237761497498)),(to_sfixed_a(0.10289344191551208)),(to_sfixed_a(-0.13351070880889893)),(to_sfixed_a(-0.04275871440768242)),(to_sfixed_a(-0.05364249274134636)),(to_sfixed_a(0.05592094361782074)),(to_sfixed_a(0.09863688051700592)),(to_sfixed_a(0.0143066281452775)),(to_sfixed_a(0.02503201737999916)),(to_sfixed_a(0.02602136880159378)),(to_sfixed_a(-0.0882510393857956)),(to_sfixed_a(0.04379257932305336)),(to_sfixed_a(-0.10089477151632309)),(to_sfixed_a(0.07104548811912537)),(to_sfixed_a(-0.12611396610736847)),(to_sfixed_a(-0.009132741950452328)),(to_sfixed_a(0.06565357744693756)),(to_sfixed_a(0.09352879971265793)),(to_sfixed_a(-0.12846754491329193)),(to_sfixed_a(-0.09329350292682648)),(to_sfixed_a(0.14646629989147186)),(to_sfixed_a(-0.03846200183033943)),(to_sfixed_a(-0.11513868719339371)),(to_sfixed_a(-0.05366159975528717)),(to_sfixed_a(0.07966706156730652)),(to_sfixed_a(-0.016043122857809067)),(to_sfixed_a(0.0682206079363823)),(to_sfixed_a(-0.028479577973484993)),(to_sfixed_a(-0.1945170909166336)),(to_sfixed_a(-0.021787719801068306)),(to_sfixed_a(-0.024319717660546303)),(to_sfixed_a(0.040887922048568726)));

    constant weight_n1_261 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.1959402710199356)),(to_sfixed_a(4.228017496643588e-05)),(to_sfixed_a(1.550085835333448e-05)),(to_sfixed_a(-3.9817481592763215e-05)),(to_sfixed_a(2.6730453100753948e-05)),(to_sfixed_a(-1.7059401216101833e-05)),(to_sfixed_a(-2.3764732759445906e-06)),(to_sfixed_a(7.595792703796178e-05)),(to_sfixed_a(3.481982639641501e-05)),(to_sfixed_a(2.733586916292552e-05)),(to_sfixed_a(7.317950803553686e-05)),(to_sfixed_a(-2.042422602244187e-05)),(to_sfixed_a(-1.0528337043069769e-05)),(to_sfixed_a(-2.1123390979482792e-05)),(to_sfixed_a(-2.8909291359013878e-05)),(to_sfixed_a(9.975833563657943e-06)),(to_sfixed_a(-5.737176616094075e-05)),(to_sfixed_a(1.086073461920023e-05)),(to_sfixed_a(-6.39381178189069e-05)),(to_sfixed_a(5.1163930038455874e-05)),(to_sfixed_a(-2.6986537704942748e-05)),(to_sfixed_a(2.1205578377703205e-05)),(to_sfixed_a(-2.2643578631686978e-05)),(to_sfixed_a(-8.922917913878337e-06)),(to_sfixed_a(-5.3822266636416316e-05)),(to_sfixed_a(-1.1970779212333582e-07)),(to_sfixed_a(-4.6251290768850595e-05)),(to_sfixed_a(3.511772956699133e-05)),(to_sfixed_a(4.797803740075324e-06)),(to_sfixed_a(-3.3003663702402264e-05)),(to_sfixed_a(-8.234872802859172e-05)),(to_sfixed_a(3.4090131521224976e-05)),(to_sfixed_a(-4.822171831619926e-05)),(to_sfixed_a(9.460347791900858e-05)),(to_sfixed_a(-0.00010812304390128702)),(to_sfixed_a(-7.007503154454753e-05)),(to_sfixed_a(7.983673276612535e-05)),(to_sfixed_a(-6.699898949591443e-05)));

    constant weight_n1_262 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.2855232357978821)),(to_sfixed_a(-0.012009457685053349)),(to_sfixed_a(0.016382595524191856)),(to_sfixed_a(-0.0009494824334979057)),(to_sfixed_a(-0.007986960001289845)),(to_sfixed_a(-0.009345650672912598)),(to_sfixed_a(-0.0034894326236099005)),(to_sfixed_a(-0.00044316297862678766)),(to_sfixed_a(-0.007842720486223698)),(to_sfixed_a(-0.0008521570125594735)),(to_sfixed_a(0.0016284298617392778)),(to_sfixed_a(0.007438482251018286)),(to_sfixed_a(0.016758719459176064)),(to_sfixed_a(0.006071758456528187)),(to_sfixed_a(0.0017645403277128935)),(to_sfixed_a(0.013219266198575497)),(to_sfixed_a(-0.008933383971452713)),(to_sfixed_a(0.0012750308960676193)),(to_sfixed_a(0.009280052967369556)),(to_sfixed_a(0.003594561479985714)),(to_sfixed_a(-0.01018866803497076)),(to_sfixed_a(-0.004435082897543907)),(to_sfixed_a(0.0008012870675884187)),(to_sfixed_a(0.010353920981287956)),(to_sfixed_a(0.01473205629736185)),(to_sfixed_a(-0.00863362941890955)),(to_sfixed_a(-0.00750513281673193)),(to_sfixed_a(0.006397109478712082)),(to_sfixed_a(-0.0018538394942879677)),(to_sfixed_a(0.010464725084602833)),(to_sfixed_a(-0.007720169611275196)),(to_sfixed_a(-0.025492992252111435)),(to_sfixed_a(-0.0007506797555834055)),(to_sfixed_a(-0.015484187752008438)),(to_sfixed_a(0.01580202579498291)),(to_sfixed_a(0.0035705692134797573)),(to_sfixed_a(-0.01352235022932291)),(to_sfixed_a(-0.010793164372444153)));

    constant weight_n1_263 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.025118069723248482)),(to_sfixed_a(1.8373853890807368e-05)),(to_sfixed_a(-5.154281097929925e-05)),(to_sfixed_a(-1.4688044757349417e-05)),(to_sfixed_a(-2.6783252906170674e-05)),(to_sfixed_a(4.218938192934729e-05)),(to_sfixed_a(2.7104088076157495e-05)),(to_sfixed_a(3.994382859673351e-05)),(to_sfixed_a(3.194859527866356e-05)),(to_sfixed_a(-3.577345341909677e-05)),(to_sfixed_a(5.637717549689114e-05)),(to_sfixed_a(-3.7980094930389896e-05)),(to_sfixed_a(-1.215906650031684e-06)),(to_sfixed_a(1.3277875723360921e-06)),(to_sfixed_a(6.761467375326902e-05)),(to_sfixed_a(7.049487612675875e-05)),(to_sfixed_a(4.905657624476589e-05)),(to_sfixed_a(-5.153948950464837e-05)),(to_sfixed_a(-7.777363498462364e-05)),(to_sfixed_a(-8.062774577410892e-05)),(to_sfixed_a(-3.083496994804591e-05)),(to_sfixed_a(-4.194413122604601e-05)),(to_sfixed_a(-7.390392056549899e-06)),(to_sfixed_a(-0.00010723681771196425)),(to_sfixed_a(-5.1169768994441256e-05)),(to_sfixed_a(2.2373031242750585e-05)),(to_sfixed_a(-2.795911484554381e-07)),(to_sfixed_a(-5.070502811577171e-05)),(to_sfixed_a(3.998948523076251e-05)),(to_sfixed_a(1.205043099616887e-05)),(to_sfixed_a(3.8176785892574117e-05)),(to_sfixed_a(-1.9905886802007444e-05)),(to_sfixed_a(-3.4692909594014054e-06)),(to_sfixed_a(7.800539606250823e-05)),(to_sfixed_a(9.467056224821135e-05)),(to_sfixed_a(-3.631187428254634e-05)),(to_sfixed_a(-1.6668052467139205e-06)),(to_sfixed_a(6.183432105899556e-06)));

    constant weight_n1_264 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.02477908693253994)),(to_sfixed_a(-0.019288891926407814)),(to_sfixed_a(0.015506207942962646)),(to_sfixed_a(0.06015670299530029)),(to_sfixed_a(-0.0035741347819566727)),(to_sfixed_a(-0.06525825709104538)),(to_sfixed_a(-0.038911692798137665)),(to_sfixed_a(-0.05510510876774788)),(to_sfixed_a(-0.07765734940767288)),(to_sfixed_a(-0.042760785669088364)),(to_sfixed_a(-0.05515104532241821)),(to_sfixed_a(-0.06800830364227295)),(to_sfixed_a(0.07014545053243637)),(to_sfixed_a(-0.057940997183322906)),(to_sfixed_a(0.057305868715047836)),(to_sfixed_a(0.03393867239356041)),(to_sfixed_a(-0.08886325359344482)),(to_sfixed_a(0.04616526886820793)),(to_sfixed_a(-0.11075863987207413)),(to_sfixed_a(-0.05938500910997391)),(to_sfixed_a(-0.004765186458826065)),(to_sfixed_a(0.009159451350569725)),(to_sfixed_a(0.09378679096698761)),(to_sfixed_a(-0.04158434271812439)),(to_sfixed_a(-0.04118884354829788)),(to_sfixed_a(0.045794207602739334)),(to_sfixed_a(0.10814567655324936)),(to_sfixed_a(-0.010431919246912003)),(to_sfixed_a(0.053056590259075165)),(to_sfixed_a(-0.0074803829193115234)),(to_sfixed_a(-0.0694463774561882)),(to_sfixed_a(-0.09940781444311142)),(to_sfixed_a(-0.0698736235499382)),(to_sfixed_a(-0.03904370591044426)),(to_sfixed_a(-0.14918029308319092)),(to_sfixed_a(0.035890646278858185)),(to_sfixed_a(0.016594503074884415)),(to_sfixed_a(0.11174057424068451)));

    constant weight_n1_265 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.01140575297176838)),(to_sfixed_a(1.944912401086185e-05)),(to_sfixed_a(-4.383268969831988e-05)),(to_sfixed_a(-3.141682827845216e-05)),(to_sfixed_a(1.9750405044760555e-05)),(to_sfixed_a(1.4573405678675044e-05)),(to_sfixed_a(9.65540311881341e-06)),(to_sfixed_a(-4.993536640540697e-05)),(to_sfixed_a(3.595332964323461e-05)),(to_sfixed_a(2.2144524336908944e-05)),(to_sfixed_a(2.2474245270132087e-05)),(to_sfixed_a(3.546551306499168e-05)),(to_sfixed_a(4.497759437072091e-05)),(to_sfixed_a(5.711020094167907e-06)),(to_sfixed_a(1.9226092263124883e-05)),(to_sfixed_a(-1.9597799109760672e-05)),(to_sfixed_a(3.347761230543256e-05)),(to_sfixed_a(6.316413055174053e-05)),(to_sfixed_a(-1.980233719223179e-05)),(to_sfixed_a(-2.723716534092091e-05)),(to_sfixed_a(3.125509465462528e-05)),(to_sfixed_a(7.657751666556578e-06)),(to_sfixed_a(-5.263443381409161e-05)),(to_sfixed_a(3.9794438634999096e-05)),(to_sfixed_a(-6.833297084085643e-05)),(to_sfixed_a(4.45602199761197e-05)),(to_sfixed_a(6.223218224477023e-05)),(to_sfixed_a(-2.6631971650203923e-06)),(to_sfixed_a(-4.875367449130863e-05)),(to_sfixed_a(-7.014566654106602e-05)),(to_sfixed_a(5.6388216762570664e-05)),(to_sfixed_a(3.603103095883853e-07)),(to_sfixed_a(2.1386878870544024e-05)),(to_sfixed_a(-6.511816172860563e-05)),(to_sfixed_a(1.2938985491928179e-05)),(to_sfixed_a(-7.93680919741746e-06)),(to_sfixed_a(-8.550210623070598e-05)),(to_sfixed_a(7.108946010703221e-05)));

    constant weight_n1_266 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.08651618659496307)),(to_sfixed_a(-3.06892761727795e-05)),(to_sfixed_a(4.4921775952389e-06)),(to_sfixed_a(1.6207755834329873e-05)),(to_sfixed_a(5.595830225502141e-05)),(to_sfixed_a(2.774448694253806e-05)),(to_sfixed_a(-1.3261817912280094e-05)),(to_sfixed_a(-2.176067755499389e-05)),(to_sfixed_a(-4.018019353679847e-06)),(to_sfixed_a(8.485700527671725e-05)),(to_sfixed_a(-2.1224637748673558e-05)),(to_sfixed_a(1.1668184924928937e-06)),(to_sfixed_a(2.3854325263528153e-05)),(to_sfixed_a(-8.229355444200337e-06)),(to_sfixed_a(-4.179045936325565e-05)),(to_sfixed_a(-6.947666861378821e-06)),(to_sfixed_a(1.1014752999471966e-05)),(to_sfixed_a(-4.5416014472721145e-05)),(to_sfixed_a(2.0459787265281193e-05)),(to_sfixed_a(-4.362263553048251e-06)),(to_sfixed_a(-1.6637201042613015e-05)),(to_sfixed_a(-1.3210345059633255e-05)),(to_sfixed_a(-0.0001171777694253251)),(to_sfixed_a(7.108573481673375e-05)),(to_sfixed_a(-5.5123080528574064e-05)),(to_sfixed_a(-2.4474298697896302e-05)),(to_sfixed_a(6.12157309660688e-05)),(to_sfixed_a(6.891584052937105e-05)),(to_sfixed_a(-7.429910328937694e-05)),(to_sfixed_a(1.6211913589359028e-07)),(to_sfixed_a(-3.285453567514196e-05)),(to_sfixed_a(1.6917805623961613e-05)),(to_sfixed_a(-5.9441601479193196e-05)),(to_sfixed_a(-1.2863194569945335e-05)),(to_sfixed_a(9.418804984306917e-05)),(to_sfixed_a(-2.2478281607618555e-05)),(to_sfixed_a(-7.33711349312216e-05)),(to_sfixed_a(0.0001636622764635831)));

    constant weight_n1_267 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.0536295622587204)),(to_sfixed_a(2.0616198526113294e-05)),(to_sfixed_a(1.9860955944750458e-05)),(to_sfixed_a(1.8695636754273437e-05)),(to_sfixed_a(-7.021222700132057e-06)),(to_sfixed_a(2.5302468202426098e-05)),(to_sfixed_a(-6.447012310673017e-06)),(to_sfixed_a(5.712843994842842e-05)),(to_sfixed_a(1.1788110896304715e-05)),(to_sfixed_a(-1.067588436853839e-05)),(to_sfixed_a(1.4983495020715054e-05)),(to_sfixed_a(6.8991071202617604e-06)),(to_sfixed_a(3.6528374039335176e-05)),(to_sfixed_a(-6.957101140869781e-05)),(to_sfixed_a(5.303024863678729e-06)),(to_sfixed_a(4.313078534323722e-05)),(to_sfixed_a(5.270748806651682e-05)),(to_sfixed_a(1.827456071623601e-05)),(to_sfixed_a(-4.888212060905062e-06)),(to_sfixed_a(0.00010099142673425376)),(to_sfixed_a(3.68246364814695e-05)),(to_sfixed_a(-4.291091318009421e-05)),(to_sfixed_a(-1.415697352058487e-05)),(to_sfixed_a(4.091101072845049e-05)),(to_sfixed_a(-6.19621278019622e-06)),(to_sfixed_a(6.516747816931456e-05)),(to_sfixed_a(-3.300037496956065e-05)),(to_sfixed_a(1.808389788493514e-05)),(to_sfixed_a(-8.009405064512976e-06)),(to_sfixed_a(1.85936860361835e-05)),(to_sfixed_a(0.00011464607814559713)),(to_sfixed_a(-1.074159263225738e-05)),(to_sfixed_a(2.422256784484489e-06)),(to_sfixed_a(3.8263075111899525e-05)),(to_sfixed_a(-1.764733315212652e-05)),(to_sfixed_a(-6.287500582402572e-05)),(to_sfixed_a(1.3183714145270642e-05)),(to_sfixed_a(-5.888039595447481e-05)));

    constant weight_n1_268 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.2709108591079712)),(to_sfixed_a(0.012121829204261303)),(to_sfixed_a(-0.018617091700434685)),(to_sfixed_a(0.004276081454008818)),(to_sfixed_a(-0.05284930020570755)),(to_sfixed_a(0.09579461067914963)),(to_sfixed_a(0.029992638155817986)),(to_sfixed_a(0.05601712316274643)),(to_sfixed_a(0.03034723363816738)),(to_sfixed_a(-0.07129666954278946)),(to_sfixed_a(0.050430383533239365)),(to_sfixed_a(0.06969772279262543)),(to_sfixed_a(-0.0509401336312294)),(to_sfixed_a(0.18041351437568665)),(to_sfixed_a(-0.013327508233487606)),(to_sfixed_a(-0.10017768293619156)),(to_sfixed_a(-0.19254954159259796)),(to_sfixed_a(-0.04052216187119484)),(to_sfixed_a(-0.014177285134792328)),(to_sfixed_a(0.09160775691270828)),(to_sfixed_a(-0.027776973322033882)),(to_sfixed_a(0.15416525304317474)),(to_sfixed_a(-0.07940360903739929)),(to_sfixed_a(0.04033343866467476)),(to_sfixed_a(-0.13875271379947662)),(to_sfixed_a(0.12435255944728851)),(to_sfixed_a(-0.04222894087433815)),(to_sfixed_a(0.022696377709507942)),(to_sfixed_a(-0.07972045987844467)),(to_sfixed_a(-0.051129404455423355)),(to_sfixed_a(0.06267987936735153)),(to_sfixed_a(0.07652270048856735)),(to_sfixed_a(0.11778531223535538)),(to_sfixed_a(-0.05972478166222572)),(to_sfixed_a(0.13196760416030884)),(to_sfixed_a(-0.051602981984615326)),(to_sfixed_a(-0.0048223827034235)),(to_sfixed_a(-0.03670242428779602)));

    constant weight_n1_269 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.09090588241815567)),(to_sfixed_a(0.20653146505355835)),(to_sfixed_a(0.10667987167835236)),(to_sfixed_a(-0.11129613220691681)),(to_sfixed_a(0.04893578216433525)),(to_sfixed_a(0.06423842906951904)),(to_sfixed_a(0.03845630958676338)),(to_sfixed_a(0.03737052530050278)),(to_sfixed_a(-0.027814345434308052)),(to_sfixed_a(0.061810847371816635)),(to_sfixed_a(0.1479017436504364)),(to_sfixed_a(-0.01780482567846775)),(to_sfixed_a(0.047876302152872086)),(to_sfixed_a(-0.0026486157439649105)),(to_sfixed_a(-0.10833846777677536)),(to_sfixed_a(-0.0019855026621371508)),(to_sfixed_a(-0.14021660387516022)),(to_sfixed_a(0.006913444492965937)),(to_sfixed_a(-0.05039491504430771)),(to_sfixed_a(0.1237754300236702)),(to_sfixed_a(0.06743653118610382)),(to_sfixed_a(-0.02218794822692871)),(to_sfixed_a(-0.1938343495130539)),(to_sfixed_a(-0.03188083693385124)),(to_sfixed_a(-0.030039189383387566)),(to_sfixed_a(0.09682638198137283)),(to_sfixed_a(-0.010419818572700024)),(to_sfixed_a(0.06438092887401581)),(to_sfixed_a(0.01791643165051937)),(to_sfixed_a(-0.03815428912639618)),(to_sfixed_a(0.07664895802736282)),(to_sfixed_a(0.028519507497549057)),(to_sfixed_a(0.0993911400437355)),(to_sfixed_a(0.019009022042155266)),(to_sfixed_a(0.08207280188798904)),(to_sfixed_a(-0.06739941239356995)),(to_sfixed_a(0.001349694444797933)),(to_sfixed_a(-0.10654909163713455)));

    constant weight_n1_270 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.023934610188007355)),(to_sfixed_a(-1.4337909306050278e-05)),(to_sfixed_a(-1.4912799088051543e-05)),(to_sfixed_a(-1.4821928743913304e-05)),(to_sfixed_a(3.625648969318718e-05)),(to_sfixed_a(-4.289431308279745e-05)),(to_sfixed_a(-1.279200387216406e-05)),(to_sfixed_a(-1.4168358575261664e-05)),(to_sfixed_a(-3.6734872992383316e-05)),(to_sfixed_a(3.6512901715468615e-05)),(to_sfixed_a(-4.4645810703514144e-05)),(to_sfixed_a(-1.9144743419019505e-05)),(to_sfixed_a(1.9994762624264695e-05)),(to_sfixed_a(4.7874884330667555e-05)),(to_sfixed_a(5.2366143791005015e-05)),(to_sfixed_a(-5.9164703998249024e-05)),(to_sfixed_a(8.596941256655555e-07)),(to_sfixed_a(5.4673055274179205e-06)),(to_sfixed_a(-5.757161488872953e-06)),(to_sfixed_a(-6.920578471181216e-06)),(to_sfixed_a(5.072130079497583e-05)),(to_sfixed_a(-6.868939817650244e-05)),(to_sfixed_a(2.3999955374165438e-05)),(to_sfixed_a(-2.1696690964745358e-05)),(to_sfixed_a(2.787970515782945e-06)),(to_sfixed_a(4.581723715091357e-06)),(to_sfixed_a(-4.330208412284264e-06)),(to_sfixed_a(-7.023267585282156e-07)),(to_sfixed_a(9.498933650320396e-05)),(to_sfixed_a(-0.00014111607742961496)),(to_sfixed_a(-2.1867228497285396e-05)),(to_sfixed_a(-1.5573275959468447e-05)),(to_sfixed_a(3.281051613157615e-05)),(to_sfixed_a(3.618720802478492e-05)),(to_sfixed_a(8.941495616454631e-05)),(to_sfixed_a(2.711335946514737e-05)),(to_sfixed_a(4.124908082303591e-05)),(to_sfixed_a(-3.8088550354586914e-05)));

    constant weight_n1_271 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.021533330902457237)),(to_sfixed_a(-1.3989964031679847e-07)),(to_sfixed_a(-9.342192242911551e-06)),(to_sfixed_a(-3.193292286596261e-05)),(to_sfixed_a(7.82609058660455e-05)),(to_sfixed_a(-6.74023385727196e-06)),(to_sfixed_a(7.877572897996288e-06)),(to_sfixed_a(-3.735786594916135e-05)),(to_sfixed_a(-3.963839844800532e-05)),(to_sfixed_a(7.038813055260107e-05)),(to_sfixed_a(1.999824416998308e-05)),(to_sfixed_a(3.4175579344264406e-07)),(to_sfixed_a(-6.859772838652134e-06)),(to_sfixed_a(4.0690811147214845e-06)),(to_sfixed_a(-6.423564627766609e-05)),(to_sfixed_a(2.454050991218537e-05)),(to_sfixed_a(-1.9838989828713238e-05)),(to_sfixed_a(2.5646522772149183e-05)),(to_sfixed_a(-5.500436600414105e-05)),(to_sfixed_a(1.9973822418251075e-05)),(to_sfixed_a(5.2492385293589905e-05)),(to_sfixed_a(-2.344514723517932e-05)),(to_sfixed_a(-0.0001123018009820953)),(to_sfixed_a(-3.334606662974693e-05)),(to_sfixed_a(-5.326601240085438e-05)),(to_sfixed_a(2.4895130991353653e-05)),(to_sfixed_a(2.8936838134541176e-05)),(to_sfixed_a(4.493001688388176e-05)),(to_sfixed_a(-2.6579244149615988e-05)),(to_sfixed_a(1.7436757843825035e-05)),(to_sfixed_a(-7.352286775130779e-05)),(to_sfixed_a(-0.0001181367042590864)),(to_sfixed_a(-4.50369443569798e-05)),(to_sfixed_a(-5.6351200328208506e-05)),(to_sfixed_a(5.1685852668015286e-05)),(to_sfixed_a(5.807870184071362e-05)),(to_sfixed_a(4.879822154180147e-05)),(to_sfixed_a(-1.6646943095111055e-06)));

    constant weight_n1_272 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.0069679380394518375)),(to_sfixed_a(1.501254882896319e-05)),(to_sfixed_a(-2.33866048802156e-05)),(to_sfixed_a(2.412778849247843e-05)),(to_sfixed_a(3.511815521051176e-05)),(to_sfixed_a(-1.9117744159302674e-05)),(to_sfixed_a(4.6763521822867915e-05)),(to_sfixed_a(1.1668395927699748e-05)),(to_sfixed_a(5.386089105741121e-05)),(to_sfixed_a(2.6271647584508173e-05)),(to_sfixed_a(4.033197183161974e-05)),(to_sfixed_a(1.920833528856747e-05)),(to_sfixed_a(1.8493783500161953e-05)),(to_sfixed_a(-2.3823296942282468e-05)),(to_sfixed_a(2.616000347188674e-05)),(to_sfixed_a(1.863338729890529e-05)),(to_sfixed_a(-7.330666267080233e-05)),(to_sfixed_a(-4.3890366214327514e-05)),(to_sfixed_a(-2.6064312805829104e-06)),(to_sfixed_a(-5.384000178310089e-05)),(to_sfixed_a(5.636464720737422e-06)),(to_sfixed_a(-5.148644413566217e-05)),(to_sfixed_a(1.1265385182923637e-05)),(to_sfixed_a(1.2296697605052032e-05)),(to_sfixed_a(-3.465605550445616e-05)),(to_sfixed_a(3.518240919220261e-05)),(to_sfixed_a(3.560736877261661e-05)),(to_sfixed_a(-6.569582183146849e-05)),(to_sfixed_a(-4.104225445189513e-05)),(to_sfixed_a(-4.6842742449371144e-05)),(to_sfixed_a(-4.2296931496821344e-05)),(to_sfixed_a(2.1687321350327693e-05)),(to_sfixed_a(1.1825098226836417e-05)),(to_sfixed_a(-6.183009190863231e-06)),(to_sfixed_a(2.873106495826505e-05)),(to_sfixed_a(-1.8488330169930123e-05)),(to_sfixed_a(-1.2092904398741666e-05)),(to_sfixed_a(-4.842328962695319e-06)));

    constant weight_n1_273 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.1439363956451416)),(to_sfixed_a(4.473391072679078e-06)),(to_sfixed_a(1.6226171055677696e-06)),(to_sfixed_a(-1.1908790611414588e-06)),(to_sfixed_a(2.5786750484257936e-05)),(to_sfixed_a(-3.845997343887575e-05)),(to_sfixed_a(4.3297714000800624e-05)),(to_sfixed_a(-1.1816334335890133e-05)),(to_sfixed_a(-1.6187301298487e-05)),(to_sfixed_a(2.5411662136320956e-05)),(to_sfixed_a(9.742587280925363e-06)),(to_sfixed_a(-9.084025805350393e-06)),(to_sfixed_a(1.648384022701066e-05)),(to_sfixed_a(-6.36133918305859e-05)),(to_sfixed_a(-1.7234317056136206e-05)),(to_sfixed_a(-2.049361683020834e-05)),(to_sfixed_a(7.668868056498468e-05)),(to_sfixed_a(-6.91183959133923e-05)),(to_sfixed_a(-9.789010800886899e-05)),(to_sfixed_a(7.4167808634229e-05)),(to_sfixed_a(0.00010372488759458065)),(to_sfixed_a(5.929194230702706e-05)),(to_sfixed_a(1.359299972136796e-06)),(to_sfixed_a(-2.037375270447228e-05)),(to_sfixed_a(-4.162466666457476e-06)),(to_sfixed_a(1.1920904398721177e-05)),(to_sfixed_a(-4.8064059228636324e-05)),(to_sfixed_a(-6.059658971935278e-06)),(to_sfixed_a(2.059578946500551e-05)),(to_sfixed_a(-4.89624471811112e-05)),(to_sfixed_a(-1.723919740470592e-05)),(to_sfixed_a(2.863433473976329e-05)),(to_sfixed_a(-4.226470264256932e-05)),(to_sfixed_a(-9.79885517153889e-05)),(to_sfixed_a(-9.968663107429165e-06)),(to_sfixed_a(-7.02863690094091e-05)),(to_sfixed_a(-4.558203727356158e-05)),(to_sfixed_a(3.7821195292053744e-05)));

    constant weight_n1_274 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.2833682894706726)),(to_sfixed_a(0.06736364215612411)),(to_sfixed_a(0.0959412232041359)),(to_sfixed_a(0.07500507682561874)),(to_sfixed_a(-0.0988767147064209)),(to_sfixed_a(0.0324171744287014)),(to_sfixed_a(-0.031115569174289703)),(to_sfixed_a(-0.025349998846650124)),(to_sfixed_a(0.10469494014978409)),(to_sfixed_a(0.11955595016479492)),(to_sfixed_a(-0.019722536206245422)),(to_sfixed_a(-0.07392393797636032)),(to_sfixed_a(-0.004625133704394102)),(to_sfixed_a(0.0075782896019518375)),(to_sfixed_a(-0.005693924613296986)),(to_sfixed_a(-0.17966563999652863)),(to_sfixed_a(-0.1206820160150528)),(to_sfixed_a(-0.10778584331274033)),(to_sfixed_a(-0.061861760914325714)),(to_sfixed_a(0.19210869073867798)),(to_sfixed_a(-0.14910437166690826)),(to_sfixed_a(0.10087059438228607)),(to_sfixed_a(0.009110260754823685)),(to_sfixed_a(-0.026321951299905777)),(to_sfixed_a(-0.024014940485358238)),(to_sfixed_a(0.0932726114988327)),(to_sfixed_a(-0.10831409692764282)),(to_sfixed_a(0.011574984528124332)),(to_sfixed_a(0.08470675349235535)),(to_sfixed_a(0.05946888402104378)),(to_sfixed_a(-0.02343805693089962)),(to_sfixed_a(-0.05834094062447548)),(to_sfixed_a(0.054633740335702896)),(to_sfixed_a(-0.03874765709042549)),(to_sfixed_a(-0.08605566620826721)),(to_sfixed_a(-0.12165069580078125)),(to_sfixed_a(0.060257695615291595)),(to_sfixed_a(-0.08705649524927139)));

    constant weight_n1_275 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.012518658302724361)),(to_sfixed_a(0.07668561488389969)),(to_sfixed_a(-0.002614077413454652)),(to_sfixed_a(-0.051420532166957855)),(to_sfixed_a(0.16417591273784637)),(to_sfixed_a(-0.012688889168202877)),(to_sfixed_a(-0.011804520152509212)),(to_sfixed_a(0.02429986000061035)),(to_sfixed_a(-0.17311398684978485)),(to_sfixed_a(0.04127948731184006)),(to_sfixed_a(0.005104245152324438)),(to_sfixed_a(-0.016280440613627434)),(to_sfixed_a(0.07527031749486923)),(to_sfixed_a(-0.046688925474882126)),(to_sfixed_a(0.0009014926617965102)),(to_sfixed_a(0.04018792882561684)),(to_sfixed_a(-0.016379455104470253)),(to_sfixed_a(-0.024096079170703888)),(to_sfixed_a(0.0418783538043499)),(to_sfixed_a(0.11747155338525772)),(to_sfixed_a(0.03180200979113579)),(to_sfixed_a(-0.025663599371910095)),(to_sfixed_a(-0.059752222150564194)),(to_sfixed_a(0.09095970541238785)),(to_sfixed_a(0.009109459817409515)),(to_sfixed_a(-0.019468730315566063)),(to_sfixed_a(0.04281075298786163)),(to_sfixed_a(0.054452553391456604)),(to_sfixed_a(-0.018839983269572258)),(to_sfixed_a(-0.0001928956771735102)),(to_sfixed_a(0.020802440121769905)),(to_sfixed_a(0.03374042734503746)),(to_sfixed_a(-0.03245437890291214)),(to_sfixed_a(0.05684492737054825)),(to_sfixed_a(0.09716375917196274)),(to_sfixed_a(-0.10619772225618362)),(to_sfixed_a(-0.130728080868721)),(to_sfixed_a(0.05784977599978447)));

    constant weight_n1_276 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.031037215143442154)),(to_sfixed_a(-0.012601389549672604)),(to_sfixed_a(-0.06916660815477371)),(to_sfixed_a(-0.012377538718283176)),(to_sfixed_a(-0.09974764287471771)),(to_sfixed_a(0.0942426398396492)),(to_sfixed_a(0.0026178888510912657)),(to_sfixed_a(-0.03199877217411995)),(to_sfixed_a(0.07723136246204376)),(to_sfixed_a(-0.02200993336737156)),(to_sfixed_a(-0.1136399433016777)),(to_sfixed_a(0.08251422643661499)),(to_sfixed_a(-0.012257360853254795)),(to_sfixed_a(-0.016432438045740128)),(to_sfixed_a(0.026192255318164825)),(to_sfixed_a(0.00043173145968466997)),(to_sfixed_a(0.018182015046477318)),(to_sfixed_a(0.0757492333650589)),(to_sfixed_a(-0.17391183972358704)),(to_sfixed_a(-0.07236877828836441)),(to_sfixed_a(0.011520648375153542)),(to_sfixed_a(0.10178365558385849)),(to_sfixed_a(-0.02733445167541504)),(to_sfixed_a(-0.15718351304531097)),(to_sfixed_a(-0.11573349684476852)),(to_sfixed_a(-0.04250534251332283)),(to_sfixed_a(-0.09016011655330658)),(to_sfixed_a(0.03662019595503807)),(to_sfixed_a(-0.09928867965936661)),(to_sfixed_a(0.056586019694805145)),(to_sfixed_a(0.15722349286079407)),(to_sfixed_a(0.09120552241802216)),(to_sfixed_a(0.00841178186237812)),(to_sfixed_a(-0.06205100193619728)),(to_sfixed_a(0.07991141080856323)),(to_sfixed_a(-0.07387077063322067)),(to_sfixed_a(0.0834999606013298)),(to_sfixed_a(0.10943973064422607)));

    constant weight_n1_277 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.0038026452530175447)),(to_sfixed_a(-0.015320259146392345)),(to_sfixed_a(0.0018455164972692728)),(to_sfixed_a(-0.02217993512749672)),(to_sfixed_a(0.0048056431114673615)),(to_sfixed_a(0.164385586977005)),(to_sfixed_a(0.07525914907455444)),(to_sfixed_a(-0.05724463611841202)),(to_sfixed_a(-0.07254447788000107)),(to_sfixed_a(-0.02949102595448494)),(to_sfixed_a(0.19216522574424744)),(to_sfixed_a(0.09013894200325012)),(to_sfixed_a(0.09735455363988876)),(to_sfixed_a(0.19587424397468567)),(to_sfixed_a(-0.11418907344341278)),(to_sfixed_a(0.023067589849233627)),(to_sfixed_a(0.08368521183729172)),(to_sfixed_a(-0.07108958065509796)),(to_sfixed_a(0.11210711300373077)),(to_sfixed_a(0.09766226261854172)),(to_sfixed_a(0.20626406371593475)),(to_sfixed_a(-0.05412275344133377)),(to_sfixed_a(0.317815899848938)),(to_sfixed_a(-0.08360674232244492)),(to_sfixed_a(0.09123747050762177)),(to_sfixed_a(0.06425527483224869)),(to_sfixed_a(-0.1227593943476677)),(to_sfixed_a(0.17857281863689423)),(to_sfixed_a(-0.09729181230068207)),(to_sfixed_a(0.04768436402082443)),(to_sfixed_a(-0.031884755939245224)),(to_sfixed_a(-0.09230542927980423)),(to_sfixed_a(-0.001456397701986134)),(to_sfixed_a(-0.10731910914182663)),(to_sfixed_a(-0.12313403189182281)),(to_sfixed_a(0.07975507527589798)),(to_sfixed_a(-0.19205647706985474)),(to_sfixed_a(0.056471746414899826)));

    constant weight_n1_278 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.39097559452056885)),(to_sfixed_a(0.05424775183200836)),(to_sfixed_a(-0.058898862451314926)),(to_sfixed_a(0.0020234589464962482)),(to_sfixed_a(-0.13854125142097473)),(to_sfixed_a(0.06578216701745987)),(to_sfixed_a(-0.04032213240861893)),(to_sfixed_a(0.19279904663562775)),(to_sfixed_a(-0.08523891121149063)),(to_sfixed_a(0.04835046827793121)),(to_sfixed_a(-0.05244262143969536)),(to_sfixed_a(0.08317595720291138)),(to_sfixed_a(-0.046711139380931854)),(to_sfixed_a(-0.018684737384319305)),(to_sfixed_a(-0.043795786798000336)),(to_sfixed_a(-0.005930733866989613)),(to_sfixed_a(0.04522937908768654)),(to_sfixed_a(-0.009236405603587627)),(to_sfixed_a(0.058702003210783005)),(to_sfixed_a(-0.06069190427660942)),(to_sfixed_a(0.010640977881848812)),(to_sfixed_a(-0.06559885293245316)),(to_sfixed_a(-0.0198160782456398)),(to_sfixed_a(0.08188146352767944)),(to_sfixed_a(-0.04012465849518776)),(to_sfixed_a(0.012901300564408302)),(to_sfixed_a(0.050755590200424194)),(to_sfixed_a(-0.08697325736284256)),(to_sfixed_a(0.05415770038962364)),(to_sfixed_a(-0.06322742998600006)),(to_sfixed_a(-0.1935914307832718)),(to_sfixed_a(0.06906428188085556)),(to_sfixed_a(0.09909181296825409)),(to_sfixed_a(-0.18471314013004303)),(to_sfixed_a(0.03424737975001335)),(to_sfixed_a(-0.042096033692359924)),(to_sfixed_a(0.060556646436452866)),(to_sfixed_a(0.22733233869075775)));

    constant weight_n1_279 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.024118540808558464)),(to_sfixed_a(-2.43294289248297e-05)),(to_sfixed_a(2.8410315280780196e-05)),(to_sfixed_a(-1.1064283171435818e-05)),(to_sfixed_a(4.279064523871057e-05)),(to_sfixed_a(4.79993577755522e-05)),(to_sfixed_a(-2.0645478798542172e-05)),(to_sfixed_a(-2.8695254513877444e-05)),(to_sfixed_a(3.070007005590014e-05)),(to_sfixed_a(-1.6440617400803603e-05)),(to_sfixed_a(4.140168312005699e-05)),(to_sfixed_a(5.971762220724486e-06)),(to_sfixed_a(-1.0908035619650036e-05)),(to_sfixed_a(3.0091248845565133e-05)),(to_sfixed_a(3.7710040487581864e-05)),(to_sfixed_a(2.0148057956248522e-05)),(to_sfixed_a(9.69041957432637e-06)),(to_sfixed_a(-4.046810499858111e-05)),(to_sfixed_a(8.514214641763829e-06)),(to_sfixed_a(3.7755973608000204e-05)),(to_sfixed_a(3.5060282243648544e-05)),(to_sfixed_a(5.9922786022070795e-05)),(to_sfixed_a(7.328332139877602e-05)),(to_sfixed_a(1.1902328878932167e-05)),(to_sfixed_a(6.487184873549268e-05)),(to_sfixed_a(6.743760604877025e-05)),(to_sfixed_a(-6.877968644403154e-06)),(to_sfixed_a(-1.3176971151551697e-05)),(to_sfixed_a(8.131572394631803e-05)),(to_sfixed_a(2.397196840320248e-05)),(to_sfixed_a(2.03956151381135e-05)),(to_sfixed_a(4.428171450854279e-05)),(to_sfixed_a(-2.3221065930556506e-05)),(to_sfixed_a(5.9127345593879e-05)),(to_sfixed_a(-8.107868052320555e-05)),(to_sfixed_a(3.4605777727847453e-06)),(to_sfixed_a(6.215405846887734e-06)),(to_sfixed_a(-7.49293394619599e-05)));

    constant weight_n1_280 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.017370225861668587)),(to_sfixed_a(-3.114174978691153e-05)),(to_sfixed_a(1.1764085684262682e-05)),(to_sfixed_a(4.165758582530543e-05)),(to_sfixed_a(-2.3625168978469446e-05)),(to_sfixed_a(4.5936340029584244e-05)),(to_sfixed_a(-3.613672379287891e-05)),(to_sfixed_a(-4.184772114967927e-05)),(to_sfixed_a(4.8792258894536644e-05)),(to_sfixed_a(-2.4958708308986388e-05)),(to_sfixed_a(1.963113209058065e-05)),(to_sfixed_a(3.352992280269973e-05)),(to_sfixed_a(-4.276878826203756e-05)),(to_sfixed_a(7.999797162483446e-06)),(to_sfixed_a(5.072744534118101e-05)),(to_sfixed_a(1.3692980246560182e-05)),(to_sfixed_a(-3.9658112882534624e-07)),(to_sfixed_a(-3.377349639777094e-05)),(to_sfixed_a(-7.175921837188071e-06)),(to_sfixed_a(-3.070419325013063e-06)),(to_sfixed_a(-6.507297712232685e-06)),(to_sfixed_a(-5.443937880045269e-06)),(to_sfixed_a(-5.5811005950090475e-06)),(to_sfixed_a(8.631959644844756e-05)),(to_sfixed_a(-9.64725695666857e-05)),(to_sfixed_a(-2.7020507332053967e-05)),(to_sfixed_a(-3.842843943857588e-05)),(to_sfixed_a(-4.644989166990854e-05)),(to_sfixed_a(3.306670987512916e-05)),(to_sfixed_a(-5.281511676002992e-06)),(to_sfixed_a(4.728382555185817e-05)),(to_sfixed_a(0.00012172941205790266)),(to_sfixed_a(1.4551125104844687e-06)),(to_sfixed_a(-6.926593414391391e-06)),(to_sfixed_a(-5.305755621520802e-06)),(to_sfixed_a(3.0072173103690147e-05)),(to_sfixed_a(-1.7012976968544535e-05)),(to_sfixed_a(5.916662757954327e-06)));

    constant weight_n1_281 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.11963588744401932)),(to_sfixed_a(3.2918011129368097e-05)),(to_sfixed_a(1.9855440768878907e-05)),(to_sfixed_a(1.0868356184801087e-05)),(to_sfixed_a(-9.089612831303384e-06)),(to_sfixed_a(-1.714102108962834e-05)),(to_sfixed_a(-4.730841737909941e-06)),(to_sfixed_a(1.378785691485973e-05)),(to_sfixed_a(-8.441261343250517e-07)),(to_sfixed_a(-2.783844138321001e-05)),(to_sfixed_a(-2.0233686882420443e-05)),(to_sfixed_a(-3.9371199818560854e-05)),(to_sfixed_a(8.054079444264062e-06)),(to_sfixed_a(7.48153543099761e-05)),(to_sfixed_a(1.3235616279416718e-05)),(to_sfixed_a(-4.34052744822111e-05)),(to_sfixed_a(-2.503582663848647e-06)),(to_sfixed_a(2.7016680178348906e-05)),(to_sfixed_a(-5.375401451601647e-05)),(to_sfixed_a(-1.4297487723524682e-05)),(to_sfixed_a(-4.826927397516556e-05)),(to_sfixed_a(2.1134474081918597e-05)),(to_sfixed_a(-1.993323712667916e-05)),(to_sfixed_a(1.3164564734324813e-05)),(to_sfixed_a(9.60506804403849e-06)),(to_sfixed_a(8.202653407352045e-05)),(to_sfixed_a(-3.354315776959993e-05)),(to_sfixed_a(2.0041445168317296e-05)),(to_sfixed_a(-2.3870254608482355e-06)),(to_sfixed_a(3.9905244193505496e-05)),(to_sfixed_a(-0.00010268310143146664)),(to_sfixed_a(-1.8678779269976076e-06)),(to_sfixed_a(2.4158774976967834e-05)),(to_sfixed_a(1.2809964573534671e-05)),(to_sfixed_a(4.222743882564828e-05)),(to_sfixed_a(-5.856570351170376e-05)),(to_sfixed_a(3.306213329778984e-05)),(to_sfixed_a(7.697906403336674e-05)));

    constant weight_n1_282 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.03734554722905159)),(to_sfixed_a(-0.003720561508089304)),(to_sfixed_a(0.00927024520933628)),(to_sfixed_a(-0.004645774606615305)),(to_sfixed_a(-0.007849730551242828)),(to_sfixed_a(-0.00978316180408001)),(to_sfixed_a(0.01879132352769375)),(to_sfixed_a(-0.004887694492936134)),(to_sfixed_a(-0.02688533440232277)),(to_sfixed_a(0.011374833062291145)),(to_sfixed_a(-0.001728131901472807)),(to_sfixed_a(-0.03725761920213699)),(to_sfixed_a(-0.0017374756280332804)),(to_sfixed_a(-0.006888478994369507)),(to_sfixed_a(0.0034551999997347593)),(to_sfixed_a(0.026415333151817322)),(to_sfixed_a(-0.03537596017122269)),(to_sfixed_a(0.03381207212805748)),(to_sfixed_a(0.0192733034491539)),(to_sfixed_a(-0.031116601079702377)),(to_sfixed_a(0.0015781113179400563)),(to_sfixed_a(0.04122023656964302)),(to_sfixed_a(0.03349613398313522)),(to_sfixed_a(-0.00011070526670664549)),(to_sfixed_a(0.0015719730872660875)),(to_sfixed_a(-0.020016666501760483)),(to_sfixed_a(0.02270672284066677)),(to_sfixed_a(-0.013527026399970055)),(to_sfixed_a(0.025169309228658676)),(to_sfixed_a(0.04708501324057579)),(to_sfixed_a(0.005839229561388493)),(to_sfixed_a(-0.019894305616617203)),(to_sfixed_a(-0.002975344192236662)),(to_sfixed_a(-0.04359135031700134)),(to_sfixed_a(-0.0030210530385375023)),(to_sfixed_a(-0.018899880349636078)),(to_sfixed_a(-0.007671207655221224)),(to_sfixed_a(-0.013373549096286297)));

    constant weight_n1_283 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.07417985051870346)),(to_sfixed_a(-2.548160955484491e-05)),(to_sfixed_a(-2.4028026018640958e-05)),(to_sfixed_a(2.173646498704329e-05)),(to_sfixed_a(7.604380698467139e-06)),(to_sfixed_a(7.139649369491963e-06)),(to_sfixed_a(2.0323157514212653e-05)),(to_sfixed_a(-8.17949421616504e-06)),(to_sfixed_a(-3.712144825840369e-05)),(to_sfixed_a(7.086272489686962e-06)),(to_sfixed_a(3.82936877940665e-06)),(to_sfixed_a(4.8324996896553785e-05)),(to_sfixed_a(-4.68374855699949e-05)),(to_sfixed_a(1.975342456717044e-05)),(to_sfixed_a(6.493507953564404e-06)),(to_sfixed_a(3.987286618212238e-05)),(to_sfixed_a(-2.2795107724959962e-05)),(to_sfixed_a(1.3045499144936912e-05)),(to_sfixed_a(1.2050995792378671e-05)),(to_sfixed_a(-7.602531695738435e-05)),(to_sfixed_a(4.8551159125054255e-05)),(to_sfixed_a(6.625342939514667e-05)),(to_sfixed_a(-4.1172308556269854e-05)),(to_sfixed_a(3.4290212624910055e-06)),(to_sfixed_a(-7.482822638849029e-06)),(to_sfixed_a(-1.67142832196987e-06)),(to_sfixed_a(8.430337766185403e-05)),(to_sfixed_a(-3.096520958933979e-05)),(to_sfixed_a(-6.183550340210786e-06)),(to_sfixed_a(1.843282916524913e-05)),(to_sfixed_a(5.926555604673922e-05)),(to_sfixed_a(-2.4302160454681143e-05)),(to_sfixed_a(7.013176946202293e-05)),(to_sfixed_a(-0.00010675506928237155)),(to_sfixed_a(-2.1190810002735816e-05)),(to_sfixed_a(5.071119448984973e-05)),(to_sfixed_a(3.537140855769394e-06)),(to_sfixed_a(-6.0300382756395265e-05)));

    constant weight_n1_284 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.030505316331982613)),(to_sfixed_a(-2.194713943026727e-06)),(to_sfixed_a(-8.033699486986734e-06)),(to_sfixed_a(8.980817801784724e-05)),(to_sfixed_a(-2.9330531106097624e-05)),(to_sfixed_a(3.3107950002886355e-05)),(to_sfixed_a(1.6129510186146945e-05)),(to_sfixed_a(6.669499271083623e-05)),(to_sfixed_a(2.6572450224193744e-05)),(to_sfixed_a(-4.318009814596735e-05)),(to_sfixed_a(-6.6451934799260926e-06)),(to_sfixed_a(-1.159758903668262e-05)),(to_sfixed_a(-4.70392478746362e-05)),(to_sfixed_a(4.798845111508854e-05)),(to_sfixed_a(-2.2186333808349445e-05)),(to_sfixed_a(-1.4480522168014431e-06)),(to_sfixed_a(4.785710189025849e-05)),(to_sfixed_a(1.7245802155230194e-05)),(to_sfixed_a(2.248744567623362e-05)),(to_sfixed_a(-8.638852159492671e-05)),(to_sfixed_a(6.895841215737164e-05)),(to_sfixed_a(-1.8994272977579385e-05)),(to_sfixed_a(6.599930202355608e-05)),(to_sfixed_a(3.0261715437518433e-05)),(to_sfixed_a(-7.608273881487548e-05)),(to_sfixed_a(-6.859212135168491e-06)),(to_sfixed_a(2.7129159207106568e-05)),(to_sfixed_a(-3.861932418658398e-05)),(to_sfixed_a(2.2938809706829488e-05)),(to_sfixed_a(7.831639959476888e-05)),(to_sfixed_a(-7.958870992297307e-05)),(to_sfixed_a(3.6914567317580804e-05)),(to_sfixed_a(2.6483050532988273e-05)),(to_sfixed_a(-6.21989747742191e-05)),(to_sfixed_a(4.460697527974844e-05)),(to_sfixed_a(1.6526504623470828e-05)),(to_sfixed_a(0.00011976833047810942)),(to_sfixed_a(-0.00010823615593835711)));

    constant weight_n1_285 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.15498720109462738)),(to_sfixed_a(0.0026776872109621763)),(to_sfixed_a(-0.0037142070941627026)),(to_sfixed_a(-0.02623279020190239)),(to_sfixed_a(-0.057957492768764496)),(to_sfixed_a(0.007420468609780073)),(to_sfixed_a(0.011048815213143826)),(to_sfixed_a(-0.026111265644431114)),(to_sfixed_a(0.008720392361283302)),(to_sfixed_a(0.028582122176885605)),(to_sfixed_a(0.026014775037765503)),(to_sfixed_a(0.011211913079023361)),(to_sfixed_a(0.033770594745874405)),(to_sfixed_a(-0.0249758530408144)),(to_sfixed_a(0.019595155492424965)),(to_sfixed_a(-0.0005603743484243751)),(to_sfixed_a(0.007188413757830858)),(to_sfixed_a(-0.0026014482136815786)),(to_sfixed_a(0.04030638560652733)),(to_sfixed_a(0.037486862391233444)),(to_sfixed_a(0.0011642674217000604)),(to_sfixed_a(0.021708009764552116)),(to_sfixed_a(0.03059788979589939)),(to_sfixed_a(-0.006763129029422998)),(to_sfixed_a(-0.017936989665031433)),(to_sfixed_a(-0.009353981353342533)),(to_sfixed_a(-0.011396088637411594)),(to_sfixed_a(0.03019394911825657)),(to_sfixed_a(-0.03742123767733574)),(to_sfixed_a(0.04468046501278877)),(to_sfixed_a(0.007835040800273418)),(to_sfixed_a(-0.028103990480303764)),(to_sfixed_a(0.03177084028720856)),(to_sfixed_a(-0.018792664632201195)),(to_sfixed_a(-0.05066857114434242)),(to_sfixed_a(-0.019582074135541916)),(to_sfixed_a(0.06156671419739723)),(to_sfixed_a(-0.01557457260787487)));

    constant weight_n1_286 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.4774242043495178)),(to_sfixed_a(0.0313040092587471)),(to_sfixed_a(0.06028437986969948)),(to_sfixed_a(-0.04368896782398224)),(to_sfixed_a(-0.011376624926924706)),(to_sfixed_a(-0.016493113711476326)),(to_sfixed_a(-0.03174189105629921)),(to_sfixed_a(-0.01778964325785637)),(to_sfixed_a(-0.012033785693347454)),(to_sfixed_a(-0.03597448393702507)),(to_sfixed_a(0.24164451658725739)),(to_sfixed_a(-0.04926976561546326)),(to_sfixed_a(-0.08027686178684235)),(to_sfixed_a(-0.01577550545334816)),(to_sfixed_a(-0.12933962047100067)),(to_sfixed_a(0.021587979048490524)),(to_sfixed_a(-0.13801975548267365)),(to_sfixed_a(0.1231796070933342)),(to_sfixed_a(0.0859910398721695)),(to_sfixed_a(-0.09937898069620132)),(to_sfixed_a(0.06583526730537415)),(to_sfixed_a(0.03155076131224632)),(to_sfixed_a(-0.18695975840091705)),(to_sfixed_a(0.037483133375644684)),(to_sfixed_a(0.14090067148208618)),(to_sfixed_a(-0.07061755657196045)),(to_sfixed_a(0.11104550957679749)),(to_sfixed_a(-0.06806783378124237)),(to_sfixed_a(-0.16783185303211212)),(to_sfixed_a(-0.05271899327635765)),(to_sfixed_a(0.022155769169330597)),(to_sfixed_a(0.038325801491737366)),(to_sfixed_a(-0.05513029173016548)),(to_sfixed_a(-0.18295198678970337)),(to_sfixed_a(-0.11375264078378677)),(to_sfixed_a(-0.022913511842489243)),(to_sfixed_a(-0.08449794352054596)),(to_sfixed_a(0.07433003932237625)));

    constant weight_n1_287 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.07903406769037247)),(to_sfixed_a(1.0000918337027542e-05)),(to_sfixed_a(-1.0431376722408459e-05)),(to_sfixed_a(4.841389454668388e-05)),(to_sfixed_a(6.8328508859849535e-06)),(to_sfixed_a(2.5712726710480638e-05)),(to_sfixed_a(2.718995528994128e-05)),(to_sfixed_a(-4.2416577343828976e-05)),(to_sfixed_a(4.202114723739214e-05)),(to_sfixed_a(5.74168325329083e-06)),(to_sfixed_a(-3.698106957017444e-05)),(to_sfixed_a(0.00011325735249556601)),(to_sfixed_a(-8.355843419849407e-06)),(to_sfixed_a(5.339848030416761e-06)),(to_sfixed_a(9.519627201370895e-05)),(to_sfixed_a(4.12024455727078e-05)),(to_sfixed_a(-3.509269663481973e-05)),(to_sfixed_a(-3.214595926692709e-05)),(to_sfixed_a(-5.409809818957001e-05)),(to_sfixed_a(-1.5266217587850406e-06)),(to_sfixed_a(2.509302976250183e-05)),(to_sfixed_a(2.5142053345916793e-05)),(to_sfixed_a(0.00010359884618083015)),(to_sfixed_a(7.534269388997927e-05)),(to_sfixed_a(-2.32660772780946e-06)),(to_sfixed_a(-5.754423000325914e-07)),(to_sfixed_a(-5.699690882465802e-05)),(to_sfixed_a(-8.329792763106525e-05)),(to_sfixed_a(-7.729310163995251e-05)),(to_sfixed_a(4.074950993526727e-05)),(to_sfixed_a(2.4745686459937133e-05)),(to_sfixed_a(8.985323074739426e-05)),(to_sfixed_a(2.033707824011799e-05)),(to_sfixed_a(-2.7141330065205693e-05)),(to_sfixed_a(-9.217548358719796e-05)),(to_sfixed_a(-2.3296943254536018e-05)),(to_sfixed_a(-7.973297033458948e-05)),(to_sfixed_a(8.74640500114765e-06)));

    constant weight_n1_288 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.06121509149670601)),(to_sfixed_a(0.19932720065116882)),(to_sfixed_a(0.1500130146741867)),(to_sfixed_a(0.09636067599058151)),(to_sfixed_a(-0.0034637022763490677)),(to_sfixed_a(-0.11668885499238968)),(to_sfixed_a(0.2395269125699997)),(to_sfixed_a(-0.13065117597579956)),(to_sfixed_a(0.04798204451799393)),(to_sfixed_a(-0.2779380977153778)),(to_sfixed_a(-0.03249204531311989)),(to_sfixed_a(0.20944899320602417)),(to_sfixed_a(0.05795677378773689)),(to_sfixed_a(-0.18872274458408356)),(to_sfixed_a(-0.04252968728542328)),(to_sfixed_a(-0.1293579339981079)),(to_sfixed_a(0.19484809041023254)),(to_sfixed_a(-0.06694295257329941)),(to_sfixed_a(0.04085693880915642)),(to_sfixed_a(-0.011686389334499836)),(to_sfixed_a(-0.19996468722820282)),(to_sfixed_a(-0.04311759024858475)),(to_sfixed_a(0.04595401510596275)),(to_sfixed_a(0.20672637224197388)),(to_sfixed_a(0.015894759446382523)),(to_sfixed_a(-0.011572130024433136)),(to_sfixed_a(-0.0022579459473490715)),(to_sfixed_a(-0.2385449856519699)),(to_sfixed_a(0.019683049991726875)),(to_sfixed_a(-0.024459006264805794)),(to_sfixed_a(-0.04625462368130684)),(to_sfixed_a(0.13044676184654236)),(to_sfixed_a(-0.06574054807424545)),(to_sfixed_a(-0.2743338942527771)),(to_sfixed_a(0.0735626295208931)),(to_sfixed_a(-0.1434391885995865)),(to_sfixed_a(-0.02025800198316574)),(to_sfixed_a(0.05996929481625557)));

    constant weight_n1_289 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.2938148081302643)),(to_sfixed_a(0.03104518912732601)),(to_sfixed_a(0.020731188356876373)),(to_sfixed_a(-0.042215097695589066)),(to_sfixed_a(0.01708052307367325)),(to_sfixed_a(-0.005302919074892998)),(to_sfixed_a(-0.01766001246869564)),(to_sfixed_a(0.0062851314432919025)),(to_sfixed_a(-0.024422260001301765)),(to_sfixed_a(0.017496168613433838)),(to_sfixed_a(0.013597279787063599)),(to_sfixed_a(-0.021143432706594467)),(to_sfixed_a(-0.017025211825966835)),(to_sfixed_a(0.005103029310703278)),(to_sfixed_a(-0.021630320698022842)),(to_sfixed_a(-0.007341337855905294)),(to_sfixed_a(-0.005816321820020676)),(to_sfixed_a(0.03236174210906029)),(to_sfixed_a(-0.01969306170940399)),(to_sfixed_a(0.03526407107710838)),(to_sfixed_a(0.029204629361629486)),(to_sfixed_a(0.046967703849077225)),(to_sfixed_a(-0.009404802694916725)),(to_sfixed_a(-0.005699943285435438)),(to_sfixed_a(0.0014094315702095628)),(to_sfixed_a(-0.04794807359576225)),(to_sfixed_a(-0.0003679454093798995)),(to_sfixed_a(-0.002977211493998766)),(to_sfixed_a(0.002359741134569049)),(to_sfixed_a(-0.007666326593607664)),(to_sfixed_a(-0.009516444057226181)),(to_sfixed_a(-0.0004326037596911192)),(to_sfixed_a(-0.014039811678230762)),(to_sfixed_a(-0.04349510744214058)),(to_sfixed_a(0.05372173711657524)),(to_sfixed_a(-0.014428570866584778)),(to_sfixed_a(0.0057450332678854465)),(to_sfixed_a(0.014946979470551014)));

    constant weight_n1_290 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.32488906383514404)),(to_sfixed_a(-0.027594614773988724)),(to_sfixed_a(0.020222188904881477)),(to_sfixed_a(-0.026104893535375595)),(to_sfixed_a(0.02121083252131939)),(to_sfixed_a(0.04328034818172455)),(to_sfixed_a(-0.03345341980457306)),(to_sfixed_a(0.01668495498597622)),(to_sfixed_a(-0.015696367248892784)),(to_sfixed_a(-0.003826610976830125)),(to_sfixed_a(0.017894523218274117)),(to_sfixed_a(0.06593739241361618)),(to_sfixed_a(0.08635153621435165)),(to_sfixed_a(-0.008231207728385925)),(to_sfixed_a(0.005145838018506765)),(to_sfixed_a(-0.052777811884880066)),(to_sfixed_a(-0.02257741056382656)),(to_sfixed_a(-0.028088735416531563)),(to_sfixed_a(-0.010255828499794006)),(to_sfixed_a(-0.0478544682264328)),(to_sfixed_a(0.03548588976264)),(to_sfixed_a(0.017810817807912827)),(to_sfixed_a(0.027973471209406853)),(to_sfixed_a(-0.014425192959606647)),(to_sfixed_a(0.06795480102300644)),(to_sfixed_a(-0.08280441164970398)),(to_sfixed_a(-0.04078613966703415)),(to_sfixed_a(-0.019478900358080864)),(to_sfixed_a(-0.03438418358564377)),(to_sfixed_a(-0.026186298578977585)),(to_sfixed_a(-0.00923915021121502)),(to_sfixed_a(0.013624017126858234)),(to_sfixed_a(-0.0737922415137291)),(to_sfixed_a(-0.014340213499963284)),(to_sfixed_a(0.05512343719601631)),(to_sfixed_a(0.0033824099227786064)),(to_sfixed_a(-0.08558829128742218)),(to_sfixed_a(-0.05277303606271744)));

    constant weight_n1_291 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.01803692989051342)),(to_sfixed_a(-0.009921497665345669)),(to_sfixed_a(0.09124439209699631)),(to_sfixed_a(0.05773346871137619)),(to_sfixed_a(-0.09205165505409241)),(to_sfixed_a(0.10243500024080276)),(to_sfixed_a(0.05519368126988411)),(to_sfixed_a(-0.0926409587264061)),(to_sfixed_a(-0.05031909421086311)),(to_sfixed_a(0.017227649688720703)),(to_sfixed_a(0.013320357538759708)),(to_sfixed_a(0.05596039816737175)),(to_sfixed_a(-0.08609278500080109)),(to_sfixed_a(-0.0072749340906739235)),(to_sfixed_a(-0.127702996134758)),(to_sfixed_a(-0.09581997990608215)),(to_sfixed_a(0.0848262757062912)),(to_sfixed_a(0.024310296401381493)),(to_sfixed_a(0.025076089426875114)),(to_sfixed_a(0.031881678849458694)),(to_sfixed_a(-0.06024899706244469)),(to_sfixed_a(0.030907809734344482)),(to_sfixed_a(0.07188834995031357)),(to_sfixed_a(-0.09473633021116257)),(to_sfixed_a(-0.050541896373033524)),(to_sfixed_a(0.005929839797317982)),(to_sfixed_a(0.1274806559085846)),(to_sfixed_a(0.15856891870498657)),(to_sfixed_a(0.02717314474284649)),(to_sfixed_a(0.11944819986820221)),(to_sfixed_a(0.09885250777006149)),(to_sfixed_a(0.009281039237976074)),(to_sfixed_a(-0.04303499311208725)),(to_sfixed_a(0.029085474088788033)),(to_sfixed_a(0.024240737780928612)),(to_sfixed_a(0.01599057950079441)),(to_sfixed_a(0.07177859544754028)),(to_sfixed_a(-0.04910143092274666)));

    constant weight_n1_292 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.012634140439331532)),(to_sfixed_a(1.0903922884608619e-05)),(to_sfixed_a(-8.202876051655039e-05)),(to_sfixed_a(2.841207606252283e-05)),(to_sfixed_a(-4.51622145192232e-05)),(to_sfixed_a(2.0014935216750018e-05)),(to_sfixed_a(7.591440862597665e-06)),(to_sfixed_a(1.46027259688708e-05)),(to_sfixed_a(2.1081599697936326e-05)),(to_sfixed_a(2.622338433866389e-05)),(to_sfixed_a(1.1548045222298242e-05)),(to_sfixed_a(4.63185961052659e-06)),(to_sfixed_a(-5.208502625464462e-05)),(to_sfixed_a(-1.5343464838224463e-05)),(to_sfixed_a(8.410094778810162e-06)),(to_sfixed_a(6.21435719949659e-06)),(to_sfixed_a(-4.196857480565086e-05)),(to_sfixed_a(-5.1890750910388306e-05)),(to_sfixed_a(1.1020166539310594e-06)),(to_sfixed_a(-5.991164925944759e-06)),(to_sfixed_a(4.0714476199354976e-05)),(to_sfixed_a(2.4132417820510454e-05)),(to_sfixed_a(0.0001119669177569449)),(to_sfixed_a(-1.728297138470225e-05)),(to_sfixed_a(1.2246920050529297e-05)),(to_sfixed_a(-3.990400000475347e-05)),(to_sfixed_a(8.660113235237077e-05)),(to_sfixed_a(8.009823432075791e-06)),(to_sfixed_a(-1.787952714948915e-05)),(to_sfixed_a(2.4339018636965193e-05)),(to_sfixed_a(3.738880332093686e-05)),(to_sfixed_a(2.233336454082746e-05)),(to_sfixed_a(-1.1505591828608885e-05)),(to_sfixed_a(-5.364006938179955e-05)),(to_sfixed_a(1.8955586710944772e-05)),(to_sfixed_a(-3.761840844163089e-06)),(to_sfixed_a(3.2259751606034115e-05)),(to_sfixed_a(2.0541112462524325e-05)));

    constant weight_n1_293 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.09827660769224167)),(to_sfixed_a(0.007736126892268658)),(to_sfixed_a(-0.0002997641859110445)),(to_sfixed_a(-0.052696529775857925)),(to_sfixed_a(-0.004962403792887926)),(to_sfixed_a(-0.010757622309029102)),(to_sfixed_a(0.0595187172293663)),(to_sfixed_a(0.01628093048930168)),(to_sfixed_a(-0.066990926861763)),(to_sfixed_a(0.0008858173387125134)),(to_sfixed_a(0.031089195981621742)),(to_sfixed_a(-0.051501210778951645)),(to_sfixed_a(0.014546651393175125)),(to_sfixed_a(0.05306513234972954)),(to_sfixed_a(-0.022013740614056587)),(to_sfixed_a(0.03788668289780617)),(to_sfixed_a(0.018420618027448654)),(to_sfixed_a(-0.006084825377911329)),(to_sfixed_a(-0.05718584358692169)),(to_sfixed_a(-0.0004286082985345274)),(to_sfixed_a(-0.02769073098897934)),(to_sfixed_a(0.061188843101263046)),(to_sfixed_a(0.012191136367619038)),(to_sfixed_a(0.02705351635813713)),(to_sfixed_a(-0.056332070380449295)),(to_sfixed_a(-0.0008105384767986834)),(to_sfixed_a(0.017367485910654068)),(to_sfixed_a(-0.07128685712814331)),(to_sfixed_a(0.0690373107790947)),(to_sfixed_a(0.005285607185214758)),(to_sfixed_a(0.025700606405735016)),(to_sfixed_a(-0.03003002144396305)),(to_sfixed_a(-0.004754595924168825)),(to_sfixed_a(0.07346654683351517)),(to_sfixed_a(0.049416396766901016)),(to_sfixed_a(-0.038708921521902084)),(to_sfixed_a(-0.011762098409235477)),(to_sfixed_a(0.052949853241443634)));

    constant weight_n1_294 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.19826844334602356)),(to_sfixed_a(-0.09035050123929977)),(to_sfixed_a(0.1282401829957962)),(to_sfixed_a(0.09025761485099792)),(to_sfixed_a(0.0673547238111496)),(to_sfixed_a(-0.20945735275745392)),(to_sfixed_a(-0.009750285185873508)),(to_sfixed_a(0.03619725629687309)),(to_sfixed_a(-0.02452705428004265)),(to_sfixed_a(-0.011059805750846863)),(to_sfixed_a(-0.041193313896656036)),(to_sfixed_a(0.030928073450922966)),(to_sfixed_a(0.038970235735177994)),(to_sfixed_a(0.08860638737678528)),(to_sfixed_a(0.013258431106805801)),(to_sfixed_a(-0.12004359066486359)),(to_sfixed_a(-0.06359665840864182)),(to_sfixed_a(0.0578620620071888)),(to_sfixed_a(-0.04058003053069115)),(to_sfixed_a(0.04941212385892868)),(to_sfixed_a(0.09586207568645477)),(to_sfixed_a(0.04492750018835068)),(to_sfixed_a(0.03588729724287987)),(to_sfixed_a(-0.05540447309613228)),(to_sfixed_a(0.03746660053730011)),(to_sfixed_a(-0.028052588924765587)),(to_sfixed_a(-0.1046086773276329)),(to_sfixed_a(0.018610430881381035)),(to_sfixed_a(-0.14415115118026733)),(to_sfixed_a(0.022757384926080704)),(to_sfixed_a(0.10125041007995605)),(to_sfixed_a(0.02347586862742901)),(to_sfixed_a(-0.04086398705840111)),(to_sfixed_a(-0.07439862191677094)),(to_sfixed_a(-0.020679611712694168)),(to_sfixed_a(-0.05584114044904709)),(to_sfixed_a(-0.14754068851470947)),(to_sfixed_a(0.1370982527732849)));

    constant weight_n1_295 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.23485298454761505)),(to_sfixed_a(0.009493929333984852)),(to_sfixed_a(0.024101098999381065)),(to_sfixed_a(0.007933643646538258)),(to_sfixed_a(0.010045337490737438)),(to_sfixed_a(0.0034517254680395126)),(to_sfixed_a(0.01190279982984066)),(to_sfixed_a(0.020017456263303757)),(to_sfixed_a(-0.024131817743182182)),(to_sfixed_a(0.00363722606562078)),(to_sfixed_a(0.004098030738532543)),(to_sfixed_a(0.013148123398423195)),(to_sfixed_a(-0.014150701463222504)),(to_sfixed_a(0.015851818025112152)),(to_sfixed_a(0.02155553735792637)),(to_sfixed_a(-0.014753598719835281)),(to_sfixed_a(0.00583539716899395)),(to_sfixed_a(-0.011831631883978844)),(to_sfixed_a(-0.0032919396180659533)),(to_sfixed_a(-0.007702155038714409)),(to_sfixed_a(-0.0002806690754368901)),(to_sfixed_a(-0.019815901294350624)),(to_sfixed_a(0.005893378518521786)),(to_sfixed_a(0.01587975025177002)),(to_sfixed_a(-0.01113112922757864)),(to_sfixed_a(2.93983357551042e-05)),(to_sfixed_a(0.009357931092381477)),(to_sfixed_a(-0.04333416745066643)),(to_sfixed_a(0.0021608308888971806)),(to_sfixed_a(-0.007579769939184189)),(to_sfixed_a(0.0006420702557079494)),(to_sfixed_a(-0.0006378993857651949)),(to_sfixed_a(0.008465421386063099)),(to_sfixed_a(0.007472262717783451)),(to_sfixed_a(0.005885730963200331)),(to_sfixed_a(0.026147158816456795)),(to_sfixed_a(0.040842022746801376)),(to_sfixed_a(0.013310317881405354)));

    constant weight_n1_296 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.08936900645494461)),(to_sfixed_a(-9.80710956355324e-06)),(to_sfixed_a(-2.238420711364597e-05)),(to_sfixed_a(3.739519161172211e-05)),(to_sfixed_a(-1.3017835044593085e-05)),(to_sfixed_a(3.5212081002100604e-06)),(to_sfixed_a(-4.674654337577522e-05)),(to_sfixed_a(3.720305903698318e-05)),(to_sfixed_a(-3.6426852602744475e-05)),(to_sfixed_a(3.834484959952533e-05)),(to_sfixed_a(-4.6285877033369616e-05)),(to_sfixed_a(-6.121103069745004e-05)),(to_sfixed_a(-5.9636557125486434e-05)),(to_sfixed_a(6.764213321730494e-05)),(to_sfixed_a(-5.460558531922288e-05)),(to_sfixed_a(6.360112456604838e-05)),(to_sfixed_a(-3.8982667319942266e-05)),(to_sfixed_a(5.2164985390845686e-05)),(to_sfixed_a(6.91357854520902e-05)),(to_sfixed_a(3.625578756327741e-05)),(to_sfixed_a(2.489211328793317e-05)),(to_sfixed_a(-0.00011995725071756169)),(to_sfixed_a(-7.528544665547088e-05)),(to_sfixed_a(4.434119910001755e-05)),(to_sfixed_a(1.0969094546453562e-05)),(to_sfixed_a(5.075658191344701e-05)),(to_sfixed_a(-1.4264647688833065e-05)),(to_sfixed_a(-3.6638809888245305e-06)),(to_sfixed_a(-6.804671284044161e-05)),(to_sfixed_a(7.51084735384211e-05)),(to_sfixed_a(3.823257429758087e-06)),(to_sfixed_a(-1.0194644346483983e-05)),(to_sfixed_a(3.373981962795369e-05)),(to_sfixed_a(4.439958865987137e-05)),(to_sfixed_a(-4.546520358417183e-05)),(to_sfixed_a(-0.00010208223102381453)),(to_sfixed_a(0.00010379073501098901)),(to_sfixed_a(-3.7974492443026975e-05)));

    constant weight_n1_297 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(0.08117362856864929)),(to_sfixed_a(-0.009324437938630581)),(to_sfixed_a(0.02069826051592827)),(to_sfixed_a(-0.041831228882074356)),(to_sfixed_a(-0.03339267894625664)),(to_sfixed_a(0.06158992648124695)),(to_sfixed_a(0.04798981547355652)),(to_sfixed_a(-0.130371555685997)),(to_sfixed_a(0.20860162377357483)),(to_sfixed_a(0.08119814842939377)),(to_sfixed_a(-0.11929849535226822)),(to_sfixed_a(0.13878850638866425)),(to_sfixed_a(-0.0497627891600132)),(to_sfixed_a(0.4302876591682434)),(to_sfixed_a(0.02456236630678177)),(to_sfixed_a(-0.04852021113038063)),(to_sfixed_a(0.010943898931145668)),(to_sfixed_a(-0.05706595256924629)),(to_sfixed_a(0.011049454100430012)),(to_sfixed_a(0.21669605374336243)),(to_sfixed_a(-0.03292899206280708)),(to_sfixed_a(-0.019640104845166206)),(to_sfixed_a(-0.1297282725572586)),(to_sfixed_a(0.12077336758375168)),(to_sfixed_a(0.023946885019540787)),(to_sfixed_a(-0.08008360117673874)),(to_sfixed_a(-0.051189567893743515)),(to_sfixed_a(-0.07122529298067093)),(to_sfixed_a(0.1068405881524086)),(to_sfixed_a(-0.10922123491764069)),(to_sfixed_a(0.008974460884928703)),(to_sfixed_a(-0.08928751200437546)),(to_sfixed_a(0.021097412332892418)),(to_sfixed_a(0.08930671960115433)),(to_sfixed_a(0.08391685038805008)),(to_sfixed_a(-0.022806761786341667)),(to_sfixed_a(-0.013277649879455566)),(to_sfixed_a(0.1502266824245453)));

    constant weight_n1_298 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.07293184101581573)),(to_sfixed_a(0.06656462699174881)),(to_sfixed_a(0.10438009351491928)),(to_sfixed_a(0.12297865003347397)),(to_sfixed_a(-0.22916410863399506)),(to_sfixed_a(-0.08121245354413986)),(to_sfixed_a(-0.07219179719686508)),(to_sfixed_a(0.015674451366066933)),(to_sfixed_a(0.35819190740585327)),(to_sfixed_a(0.22358949482440948)),(to_sfixed_a(-0.11011212319135666)),(to_sfixed_a(-0.39042192697525024)),(to_sfixed_a(0.1622074842453003)),(to_sfixed_a(-0.17522840201854706)),(to_sfixed_a(-0.15222196280956268)),(to_sfixed_a(-0.14168865978717804)),(to_sfixed_a(-0.004906178917735815)),(to_sfixed_a(-0.06078791990876198)),(to_sfixed_a(0.0008034229977056384)),(to_sfixed_a(0.12777094542980194)),(to_sfixed_a(-0.15900589525699615)),(to_sfixed_a(0.09862235933542252)),(to_sfixed_a(-0.059369783848524094)),(to_sfixed_a(-0.02197953127324581)),(to_sfixed_a(-0.04988323524594307)),(to_sfixed_a(-0.01115721557289362)),(to_sfixed_a(-0.01996438577771187)),(to_sfixed_a(0.007027185056358576)),(to_sfixed_a(-0.019625648856163025)),(to_sfixed_a(-0.08595611155033112)),(to_sfixed_a(-0.027850838378071785)),(to_sfixed_a(0.06010810285806656)),(to_sfixed_a(0.0010973665630444884)),(to_sfixed_a(-0.03169693425297737)),(to_sfixed_a(-0.09990599751472473)),(to_sfixed_a(0.09413562715053558)),(to_sfixed_a(-0.023425452411174774)),(to_sfixed_a(0.0795816034078598)));

    constant weight_n1_299 : sfixed_bus_array(37 downto 0) := ((to_sfixed_a(-0.043471332639455795)),(to_sfixed_a(0.00462960172444582)),(to_sfixed_a(0.029447250068187714)),(to_sfixed_a(0.06329707056283951)),(to_sfixed_a(0.07477883249521255)),(to_sfixed_a(-0.04786970838904381)),(to_sfixed_a(-0.036666322499513626)),(to_sfixed_a(0.07957089692354202)),(to_sfixed_a(-0.0006638221675530076)),(to_sfixed_a(-0.03141332417726517)),(to_sfixed_a(0.0576675608754158)),(to_sfixed_a(-0.013717909343540668)),(to_sfixed_a(-0.02756504900753498)),(to_sfixed_a(-0.07459476590156555)),(to_sfixed_a(0.04570676386356354)),(to_sfixed_a(-0.10189735889434814)),(to_sfixed_a(-0.15209239721298218)),(to_sfixed_a(-0.06258902698755264)),(to_sfixed_a(-0.020503360778093338)),(to_sfixed_a(0.05407082289457321)),(to_sfixed_a(0.046411968767642975)),(to_sfixed_a(0.17444133758544922)),(to_sfixed_a(0.1494518220424652)),(to_sfixed_a(-0.12376590073108673)),(to_sfixed_a(-0.10220236331224442)),(to_sfixed_a(0.021867450326681137)),(to_sfixed_a(0.109153151512146)),(to_sfixed_a(0.02460452727973461)),(to_sfixed_a(0.09530172497034073)),(to_sfixed_a(-0.01893080584704876)),(to_sfixed_a(-0.07033306360244751)),(to_sfixed_a(-0.006563478149473667)),(to_sfixed_a(-0.04257404804229736)),(to_sfixed_a(-0.05759034305810928)),(to_sfixed_a(0.02337595261633396)),(to_sfixed_a(0.05614641681313515)),(to_sfixed_a(-0.02624959498643875)),(to_sfixed_a(0.08900977671146393)));


    constant weight_n2_0 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.06503242254257202)),(to_sfixed_a(-0.3201495409011841)),(to_sfixed_a(-0.18904531002044678)),(to_sfixed_a(-0.00017916080832947046)),(to_sfixed_a(-0.002226591343060136)),(to_sfixed_a(5.700455221813172e-05)),(to_sfixed_a(-0.0015307648573070765)),(to_sfixed_a(0.00022695072402711958)),(to_sfixed_a(-6.170864071464166e-05)),(to_sfixed_a(-7.078427006490529e-05)),(to_sfixed_a(-0.00044694452662952244)),(to_sfixed_a(-0.0016299778362736106)),(to_sfixed_a(0.00029290010570548475)),(to_sfixed_a(-0.001841430552303791)),(to_sfixed_a(0.00013617367949336767)),(to_sfixed_a(6.265976116992533e-05)),(to_sfixed_a(0.00029594707302749157)),(to_sfixed_a(-6.8223278503865e-05)),(to_sfixed_a(-0.2603231370449066)),(to_sfixed_a(1.8663195078261197e-05)),(to_sfixed_a(0.00022071716375648975)),(to_sfixed_a(-0.0001930675789481029)),(to_sfixed_a(0.0001008526814985089)),(to_sfixed_a(0.011801455169916153)),(to_sfixed_a(0.0008108555339276791)),(to_sfixed_a(0.0022276942618191242)),(to_sfixed_a(-0.0001581604010425508)),(to_sfixed_a(-5.332746877684258e-05)),(to_sfixed_a(-8.29250129754655e-05)),(to_sfixed_a(-6.406808097381145e-07)),(to_sfixed_a(0.0011845771223306656)),(to_sfixed_a(7.022379577392712e-05)),(to_sfixed_a(0.0003243652172386646)),(to_sfixed_a(6.504469638457522e-06)),(to_sfixed_a(3.1587565899826586e-05)),(to_sfixed_a(-0.0003213939780835062)),(to_sfixed_a(-0.003550008637830615)),(to_sfixed_a(0.0017064189305528998)),(to_sfixed_a(-0.14093966782093048)),(to_sfixed_a(-9.37792137847282e-05)),(to_sfixed_a(0.1274830847978592)),(to_sfixed_a(-0.0003897250280715525)),(to_sfixed_a(-6.079021841287613e-05)),(to_sfixed_a(-4.856927989749238e-05)),(to_sfixed_a(-0.002561888424679637)),(to_sfixed_a(-1.8005535821430385e-05)),(to_sfixed_a(0.0004485829849727452)),(to_sfixed_a(-0.005033815745264292)),(to_sfixed_a(-0.0001927866687765345)),(to_sfixed_a(-0.0010583116672933102)),(to_sfixed_a(0.0003169199335388839)),(to_sfixed_a(0.000492364983074367)),(to_sfixed_a(0.00022169780277181417)),(to_sfixed_a(-0.38978666067123413)),(to_sfixed_a(-0.0007830478716641665)),(to_sfixed_a(-0.4035998582839966)),(to_sfixed_a(8.329894626513124e-06)),(to_sfixed_a(-0.0005339281051419675)),(to_sfixed_a(5.6237495300592855e-05)),(to_sfixed_a(-0.0002407604333711788)),(to_sfixed_a(-1.6503079677931964e-05)),(to_sfixed_a(-0.0009740635869093239)),(to_sfixed_a(0.0001892895088531077)),(to_sfixed_a(0.394731342792511)),(to_sfixed_a(-0.00012897609849460423)),(to_sfixed_a(4.863832145929337e-07)),(to_sfixed_a(-5.68242758163251e-05)),(to_sfixed_a(-0.002051222138106823)),(to_sfixed_a(-2.0342915377113968e-05)),(to_sfixed_a(-2.119540295097977e-05)),(to_sfixed_a(0.005512809846550226)),(to_sfixed_a(0.00024603004567325115)),(to_sfixed_a(0.014924348331987858)),(to_sfixed_a(3.114533319603652e-05)),(to_sfixed_a(-0.00010537973867030814)),(to_sfixed_a(-9.052062523551285e-06)),(to_sfixed_a(0.00024897276307456195)),(to_sfixed_a(0.0001256043033208698)),(to_sfixed_a(2.236445652670227e-06)),(to_sfixed_a(0.0012558209709823132)),(to_sfixed_a(0.00033506553154438734)),(to_sfixed_a(-3.631558865890838e-05)),(to_sfixed_a(-0.27795910835266113)),(to_sfixed_a(-0.008146814070641994)),(to_sfixed_a(0.00015091212117113173)),(to_sfixed_a(0.315836101770401)),(to_sfixed_a(-0.0037179940845817327)),(to_sfixed_a(-0.00010965008550556377)),(to_sfixed_a(-0.0002199954615207389)),(to_sfixed_a(0.00016734670498408377)),(to_sfixed_a(-0.5778124332427979)),(to_sfixed_a(7.057709444779903e-05)),(to_sfixed_a(0.39076292514801025)),(to_sfixed_a(-0.00015176644956227392)),(to_sfixed_a(0.011692794971168041)),(to_sfixed_a(0.00011661733879009262)),(to_sfixed_a(-6.725575076416135e-06)),(to_sfixed_a(-0.00017031609604600817)),(to_sfixed_a(-0.0003010049695149064)),(to_sfixed_a(2.36471532844007e-05)),(to_sfixed_a(0.6418099999427795)),(to_sfixed_a(0.2883972227573395)),(to_sfixed_a(0.0003023860335815698)),(to_sfixed_a(0.2279343456029892)),(to_sfixed_a(0.25919172167778015)),(to_sfixed_a(0.3766377568244934)),(to_sfixed_a(8.077664824668318e-05)),(to_sfixed_a(3.353131978656165e-05)),(to_sfixed_a(-0.00038381462218239903)),(to_sfixed_a(0.0006399316480383277)),(to_sfixed_a(0.005729239899665117)),(to_sfixed_a(0.00024041686265263706)),(to_sfixed_a(0.5716568231582642)),(to_sfixed_a(-1.2888078344985843e-05)),(to_sfixed_a(-0.000154887733515352)),(to_sfixed_a(0.0010657019447535276)),(to_sfixed_a(0.00135921745095402)),(to_sfixed_a(-0.0002274345315527171)),(to_sfixed_a(0.000158592956722714)),(to_sfixed_a(-0.001445532077923417)),(to_sfixed_a(-0.00015535690181422979)),(to_sfixed_a(-0.00021306266717147082)),(to_sfixed_a(-0.00029068320873193443)),(to_sfixed_a(0.00012959852756466717)),(to_sfixed_a(6.395742821041495e-05)),(to_sfixed_a(-0.0004319649306125939)),(to_sfixed_a(0.32946497201919556)),(to_sfixed_a(-0.00023769852123223245)),(to_sfixed_a(-6.595259765163064e-05)),(to_sfixed_a(2.6973983040079474e-05)),(to_sfixed_a(-2.0718289306387305e-07)),(to_sfixed_a(-0.0001507667184341699)),(to_sfixed_a(0.0032800936605781317)),(to_sfixed_a(0.014977428130805492)),(to_sfixed_a(0.00012939739099238068)),(to_sfixed_a(8.312798308907077e-05)),(to_sfixed_a(0.0014089160831645131)),(to_sfixed_a(-0.0006694017793051898)),(to_sfixed_a(3.6718476621899754e-05)),(to_sfixed_a(-0.00014972552889958024)),(to_sfixed_a(0.002266927855089307)),(to_sfixed_a(-0.0002736650640144944)),(to_sfixed_a(-2.3646483896300197e-05)),(to_sfixed_a(-2.5415751224500127e-05)),(to_sfixed_a(-0.00013726578617934138)),(to_sfixed_a(-0.00040707190055400133)),(to_sfixed_a(-0.17555439472198486)),(to_sfixed_a(-9.175590093946084e-06)),(to_sfixed_a(-6.770365871489048e-05)),(to_sfixed_a(-0.454326331615448)),(to_sfixed_a(-0.00011560162238311023)),(to_sfixed_a(-6.712695176247507e-05)),(to_sfixed_a(0.2872745096683502)),(to_sfixed_a(-3.6050943890586495e-05)),(to_sfixed_a(-1.0134501280845143e-05)),(to_sfixed_a(0.3202918767929077)),(to_sfixed_a(-0.00020234269322827458)),(to_sfixed_a(0.00035764736821874976)),(to_sfixed_a(1.935019827215001e-05)),(to_sfixed_a(2.2810807422501966e-05)),(to_sfixed_a(-0.00018696661572903395)),(to_sfixed_a(0.000136915419716388)),(to_sfixed_a(0.37244561314582825)),(to_sfixed_a(-0.05836920067667961)),(to_sfixed_a(0.0022535747848451138)),(to_sfixed_a(0.24840675294399261)),(to_sfixed_a(0.00015766927390359342)),(to_sfixed_a(-0.00020361211500130594)),(to_sfixed_a(0.0001671132631599903)),(to_sfixed_a(-6.226157711353153e-05)),(to_sfixed_a(0.013034544885158539)),(to_sfixed_a(0.000518349464982748)),(to_sfixed_a(0.10177900642156601)),(to_sfixed_a(0.0001468636910431087)),(to_sfixed_a(0.008441628888249397)),(to_sfixed_a(0.31264618039131165)),(to_sfixed_a(0.24731990694999695)),(to_sfixed_a(0.38471880555152893)),(to_sfixed_a(0.04906412214040756)),(to_sfixed_a(0.009812244214117527)),(to_sfixed_a(-7.06327919033356e-05)),(to_sfixed_a(-0.0011282312916591763)),(to_sfixed_a(0.00024355662753805518)),(to_sfixed_a(-5.519257683772594e-06)),(to_sfixed_a(-0.00017270719399675727)),(to_sfixed_a(-0.0022468280512839556)),(to_sfixed_a(0.12111204117536545)),(to_sfixed_a(4.493811138672754e-05)),(to_sfixed_a(6.0257265431573614e-05)),(to_sfixed_a(9.308053995482624e-05)),(to_sfixed_a(-0.0001141763204941526)),(to_sfixed_a(-0.00011589728092076257)),(to_sfixed_a(-0.0005291671259328723)),(to_sfixed_a(0.005761157721281052)),(to_sfixed_a(-3.457134880591184e-06)),(to_sfixed_a(-0.0025306581519544125)),(to_sfixed_a(6.851688522147015e-05)),(to_sfixed_a(0.004758994095027447)),(to_sfixed_a(0.001261427765712142)),(to_sfixed_a(-0.00020457638311199844)),(to_sfixed_a(4.226851160638034e-06)),(to_sfixed_a(-7.038642797851935e-05)),(to_sfixed_a(-3.3507276384625584e-05)),(to_sfixed_a(-3.72800714103505e-05)),(to_sfixed_a(0.00014558000839315355)),(to_sfixed_a(-0.28772222995758057)),(to_sfixed_a(-0.14147736132144928)),(to_sfixed_a(-0.1839216649532318)),(to_sfixed_a(-0.10814628005027771)),(to_sfixed_a(-0.27554768323898315)),(to_sfixed_a(-8.946954039856791e-05)),(to_sfixed_a(-0.00011710949911503121)),(to_sfixed_a(2.6328056264901534e-05)),(to_sfixed_a(0.0001333274703938514)),(to_sfixed_a(5.771003634436056e-05)),(to_sfixed_a(0.0002007288858294487)),(to_sfixed_a(0.018377408385276794)),(to_sfixed_a(0.4304310977458954)),(to_sfixed_a(-0.5485594272613525)),(to_sfixed_a(-8.161310688592494e-06)),(to_sfixed_a(-0.0001212596835102886)),(to_sfixed_a(5.590347427641973e-06)),(to_sfixed_a(-0.00045194875565357506)),(to_sfixed_a(0.0011681747855618596)),(to_sfixed_a(0.002732318127527833)),(to_sfixed_a(-5.830606824019924e-05)),(to_sfixed_a(1.5959863958414644e-05)),(to_sfixed_a(9.081899770535529e-05)),(to_sfixed_a(-0.0038033598102629185)),(to_sfixed_a(0.006789632141590118)),(to_sfixed_a(-0.03738853335380554)),(to_sfixed_a(7.251168426591903e-05)),(to_sfixed_a(-0.00022108056873548776)),(to_sfixed_a(-3.778886457439512e-05)),(to_sfixed_a(0.07592804729938507)),(to_sfixed_a(0.00447411322966218)),(to_sfixed_a(-0.37940725684165955)),(to_sfixed_a(-5.857194628333673e-05)),(to_sfixed_a(-9.138860332313925e-05)),(to_sfixed_a(0.00022082834038883448)),(to_sfixed_a(0.021230770274996758)),(to_sfixed_a(-8.417955541517586e-07)),(to_sfixed_a(-0.001325061428360641)),(to_sfixed_a(-0.0002470861072652042)),(to_sfixed_a(-0.0018783016130328178)),(to_sfixed_a(2.5808232749113813e-05)),(to_sfixed_a(-0.00223674182780087)),(to_sfixed_a(-0.005416049621999264)),(to_sfixed_a(-2.7419693651609123e-05)),(to_sfixed_a(0.0008846897981129587)),(to_sfixed_a(-0.0014011336024850607)),(to_sfixed_a(0.00038053406751714647)),(to_sfixed_a(-5.9523823438212276e-05)),(to_sfixed_a(-5.615243571810424e-05)),(to_sfixed_a(-9.959653107216582e-05)),(to_sfixed_a(8.182008605217561e-05)),(to_sfixed_a(0.1653849482536316)),(to_sfixed_a(-0.00016466487431898713)),(to_sfixed_a(-0.00017667392967268825)),(to_sfixed_a(-0.00012016935215797275)),(to_sfixed_a(3.685264164232649e-05)),(to_sfixed_a(4.798695590579882e-05)),(to_sfixed_a(7.099469075910747e-05)),(to_sfixed_a(6.911940727150068e-05)),(to_sfixed_a(-0.0001015395246213302)),(to_sfixed_a(0.03328287973999977)),(to_sfixed_a(-0.00014630061923526227)),(to_sfixed_a(-0.0002175799454562366)),(to_sfixed_a(8.732023707125336e-05)),(to_sfixed_a(-0.03759659826755524)),(to_sfixed_a(-0.0006318983505479991)),(to_sfixed_a(-1.688230986474082e-05)),(to_sfixed_a(4.2060521082021296e-05)),(to_sfixed_a(4.057132173329592e-06)),(to_sfixed_a(7.032173743937165e-05)),(to_sfixed_a(6.629426934523508e-05)),(to_sfixed_a(-0.0029028127901256084)),(to_sfixed_a(-0.0019953015726059675)),(to_sfixed_a(-0.4214950203895569)),(to_sfixed_a(-0.02023419179022312)),(to_sfixed_a(-1.6152021999005228e-05)),(to_sfixed_a(-3.012650995515287e-05)),(to_sfixed_a(6.948698137421161e-05)),(to_sfixed_a(-0.00048273103311657906)),(to_sfixed_a(-5.183328903513029e-05)),(to_sfixed_a(-8.77290585776791e-06)),(to_sfixed_a(0.002406578976660967)),(to_sfixed_a(0.00821943674236536)),(to_sfixed_a(3.710926102939993e-05)),(to_sfixed_a(-0.264583021402359)),(to_sfixed_a(0.00023337775201071054)),(to_sfixed_a(-0.0014758470933884382)),(to_sfixed_a(-0.20695717632770538)),(to_sfixed_a(0.00020510805188678205)),(to_sfixed_a(-0.20307843387126923)),(to_sfixed_a(0.004996892996132374)),(to_sfixed_a(-0.0036548995412886143)),(to_sfixed_a(3.63848521374166e-05)),(to_sfixed_a(0.23973427712917328)),(to_sfixed_a(0.003447110066190362)),(to_sfixed_a(0.47628164291381836)));

    constant weight_n2_1 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.025124521926045418)),(to_sfixed_a(0.02612602338194847)),(to_sfixed_a(0.06111837550997734)),(to_sfixed_a(-3.26566951116547e-05)),(to_sfixed_a(0.008441493846476078)),(to_sfixed_a(-6.203309749253094e-05)),(to_sfixed_a(0.00756555050611496)),(to_sfixed_a(-1.1038358934456483e-05)),(to_sfixed_a(0.00015455044922418892)),(to_sfixed_a(-0.00015011463256087154)),(to_sfixed_a(0.000322435749694705)),(to_sfixed_a(0.0006272050086408854)),(to_sfixed_a(0.004622453358024359)),(to_sfixed_a(6.462182500399649e-05)),(to_sfixed_a(-6.870023935334757e-05)),(to_sfixed_a(-0.00016945682000368834)),(to_sfixed_a(0.003633642103523016)),(to_sfixed_a(-0.000169271050253883)),(to_sfixed_a(-0.0020599523559212685)),(to_sfixed_a(6.069967639632523e-05)),(to_sfixed_a(-7.890643610153347e-05)),(to_sfixed_a(-0.0003160831402055919)),(to_sfixed_a(0.000699488737154752)),(to_sfixed_a(0.1456850916147232)),(to_sfixed_a(0.009555445052683353)),(to_sfixed_a(0.002240905538201332)),(to_sfixed_a(-0.00011355167953297496)),(to_sfixed_a(0.0003323159471619874)),(to_sfixed_a(0.00916819367557764)),(to_sfixed_a(-0.00012893389794044197)),(to_sfixed_a(0.30418944358825684)),(to_sfixed_a(6.720506644342095e-05)),(to_sfixed_a(0.0030911320354789495)),(to_sfixed_a(-3.028490027645603e-07)),(to_sfixed_a(0.00011817565246019512)),(to_sfixed_a(-1.3086813851259649e-05)),(to_sfixed_a(0.0037526795640587807)),(to_sfixed_a(0.26355651021003723)),(to_sfixed_a(0.0773925632238388)),(to_sfixed_a(8.294394501717761e-05)),(to_sfixed_a(0.17012836039066315)),(to_sfixed_a(0.24592408537864685)),(to_sfixed_a(-0.00013347939238883555)),(to_sfixed_a(9.80351833277382e-05)),(to_sfixed_a(0.0059973932802677155)),(to_sfixed_a(0.012807441875338554)),(to_sfixed_a(0.45586395263671875)),(to_sfixed_a(0.012935051694512367)),(to_sfixed_a(5.763114313594997e-05)),(to_sfixed_a(0.0065710037015378475)),(to_sfixed_a(0.0011989125050604343)),(to_sfixed_a(0.0005771306459791958)),(to_sfixed_a(-5.059438990429044e-06)),(to_sfixed_a(0.0002857789513655007)),(to_sfixed_a(0.012191352434456348)),(to_sfixed_a(-0.29129233956336975)),(to_sfixed_a(-0.0002441944379825145)),(to_sfixed_a(0.2700541019439697)),(to_sfixed_a(0.00015009191702120006)),(to_sfixed_a(-0.00020299776224419475)),(to_sfixed_a(0.001994896214455366)),(to_sfixed_a(0.0017708403756842017)),(to_sfixed_a(0.0005649558734148741)),(to_sfixed_a(-0.3191283345222473)),(to_sfixed_a(1.427740789949894e-05)),(to_sfixed_a(-0.3586217164993286)),(to_sfixed_a(-9.774570935405791e-05)),(to_sfixed_a(0.004725146107375622)),(to_sfixed_a(0.23448438942432404)),(to_sfixed_a(-6.79802760714665e-05)),(to_sfixed_a(0.00015875359531491995)),(to_sfixed_a(0.4631418287754059)),(to_sfixed_a(0.0036566394846886396)),(to_sfixed_a(6.027499694027938e-05)),(to_sfixed_a(-0.0001367642544209957)),(to_sfixed_a(-6.963533814996481e-05)),(to_sfixed_a(0.3427424132823944)),(to_sfixed_a(0.003198821097612381)),(to_sfixed_a(-0.00015503539179917425)),(to_sfixed_a(0.3028101921081543)),(to_sfixed_a(0.002416921779513359)),(to_sfixed_a(8.880160748958588e-06)),(to_sfixed_a(0.22848504781723022)),(to_sfixed_a(0.001906804507598281)),(to_sfixed_a(-0.0003246183041483164)),(to_sfixed_a(0.2244049459695816)),(to_sfixed_a(-0.23277053236961365)),(to_sfixed_a(0.24309797585010529)),(to_sfixed_a(0.00017180068243760616)),(to_sfixed_a(0.00010586007556412369)),(to_sfixed_a(-0.0014270443934947252)),(to_sfixed_a(-2.1333773474907503e-05)),(to_sfixed_a(0.0026921641547232866)),(to_sfixed_a(7.066696707624942e-05)),(to_sfixed_a(-0.31268176436424255)),(to_sfixed_a(-9.30314781726338e-05)),(to_sfixed_a(-7.328403444262221e-05)),(to_sfixed_a(-5.7792014558799565e-05)),(to_sfixed_a(-0.00044929378782399)),(to_sfixed_a(-7.638478564331308e-05)),(to_sfixed_a(0.0013577985810115933)),(to_sfixed_a(-0.001023145392537117)),(to_sfixed_a(-6.463335012085736e-06)),(to_sfixed_a(-0.14300444722175598)),(to_sfixed_a(-0.00354191311635077)),(to_sfixed_a(0.003626211080700159)),(to_sfixed_a(-8.972948126029223e-05)),(to_sfixed_a(0.0001000184565782547)),(to_sfixed_a(0.00014040875248610973)),(to_sfixed_a(0.00596236065030098)),(to_sfixed_a(0.006759504787623882)),(to_sfixed_a(5.534977753995918e-05)),(to_sfixed_a(0.002806998323649168)),(to_sfixed_a(-3.6335848562885076e-05)),(to_sfixed_a(-5.947522367932834e-05)),(to_sfixed_a(0.002623820211738348)),(to_sfixed_a(0.2384946048259735)),(to_sfixed_a(0.00019925610104110092)),(to_sfixed_a(0.00028283961000852287)),(to_sfixed_a(0.004436850547790527)),(to_sfixed_a(-6.312571349553764e-05)),(to_sfixed_a(-2.5043951609404758e-05)),(to_sfixed_a(-0.0012310208985581994)),(to_sfixed_a(-0.00022179623192641884)),(to_sfixed_a(6.985455547692254e-05)),(to_sfixed_a(-0.24623718857765198)),(to_sfixed_a(-0.00976000726222992)),(to_sfixed_a(3.657559136627242e-05)),(to_sfixed_a(0.0002028385642915964)),(to_sfixed_a(0.00015715285553596914)),(to_sfixed_a(-4.5354030589805916e-05)),(to_sfixed_a(7.19568706699647e-05)),(to_sfixed_a(-0.00038157738163135946)),(to_sfixed_a(0.03417704626917839)),(to_sfixed_a(-0.00015982580953277647)),(to_sfixed_a(2.4393812054768205e-06)),(to_sfixed_a(0.008713877759873867)),(to_sfixed_a(-0.00019816831627395004)),(to_sfixed_a(-3.795777229242958e-05)),(to_sfixed_a(-0.00015345927386078984)),(to_sfixed_a(-0.027700942009687424)),(to_sfixed_a(-5.5854005040600896e-05)),(to_sfixed_a(0.0001882986689452082)),(to_sfixed_a(-8.46093644213397e-06)),(to_sfixed_a(0.00023193232482299209)),(to_sfixed_a(0.00012205559323774651)),(to_sfixed_a(0.0036953571252524853)),(to_sfixed_a(-0.00029608028125949204)),(to_sfixed_a(6.466658669523895e-05)),(to_sfixed_a(-0.002862091874703765)),(to_sfixed_a(-0.0001612673804629594)),(to_sfixed_a(-8.033021003939211e-05)),(to_sfixed_a(0.1880967915058136)),(to_sfixed_a(-3.1502568162977695e-06)),(to_sfixed_a(-0.00023751400294713676)),(to_sfixed_a(-0.0006616500904783607)),(to_sfixed_a(7.919831114122644e-05)),(to_sfixed_a(0.13009783625602722)),(to_sfixed_a(8.932289347285405e-06)),(to_sfixed_a(-0.00023595723905600607)),(to_sfixed_a(0.00019006036745849997)),(to_sfixed_a(-4.372899638838135e-05)),(to_sfixed_a(-0.0005224003689363599)),(to_sfixed_a(0.0004061743966303766)),(to_sfixed_a(0.32781335711479187)),(to_sfixed_a(-0.0017479790840297937)),(to_sfixed_a(-3.799630212597549e-05)),(to_sfixed_a(0.003188453847542405)),(to_sfixed_a(-0.00037959308247081935)),(to_sfixed_a(0.00023772762506268919)),(to_sfixed_a(0.0020965165458619595)),(to_sfixed_a(-0.003448721021413803)),(to_sfixed_a(0.0014548853505402803)),(to_sfixed_a(-3.69702756870538e-05)),(to_sfixed_a(0.2136567234992981)),(to_sfixed_a(0.0013183113187551498)),(to_sfixed_a(0.0038790751714259386)),(to_sfixed_a(-6.564867362612858e-06)),(to_sfixed_a(-0.013008194975554943)),(to_sfixed_a(0.3394918739795685)),(to_sfixed_a(0.0004442712524905801)),(to_sfixed_a(0.023386720567941666)),(to_sfixed_a(-5.630256055155769e-05)),(to_sfixed_a(-9.422345101484098e-06)),(to_sfixed_a(-0.00015121695469133556)),(to_sfixed_a(0.008229967206716537)),(to_sfixed_a(0.0010231329360976815)),(to_sfixed_a(0.0017106266459450126)),(to_sfixed_a(0.000699665630236268)),(to_sfixed_a(-0.00029182538855820894)),(to_sfixed_a(-0.0004443297511897981)),(to_sfixed_a(-0.0001898916088975966)),(to_sfixed_a(-0.00033150595845654607)),(to_sfixed_a(0.18285827338695526)),(to_sfixed_a(-0.00020572349603753537)),(to_sfixed_a(-0.00030418025562539697)),(to_sfixed_a(4.594010897562839e-05)),(to_sfixed_a(-0.002294735750183463)),(to_sfixed_a(0.004549336154013872)),(to_sfixed_a(0.0001994111225940287)),(to_sfixed_a(0.0001872516586445272)),(to_sfixed_a(-0.00013649227912537754)),(to_sfixed_a(-1.2763688573613763e-05)),(to_sfixed_a(-8.077782695181668e-06)),(to_sfixed_a(2.5530142011120915e-05)),(to_sfixed_a(0.0015410315245389938)),(to_sfixed_a(0.1709200143814087)),(to_sfixed_a(0.0004758437571581453)),(to_sfixed_a(0.3678654134273529)),(to_sfixed_a(0.43811410665512085)),(to_sfixed_a(-0.0011372151784598827)),(to_sfixed_a(-0.000215317661059089)),(to_sfixed_a(0.00018119451124221087)),(to_sfixed_a(0.00022850741515867412)),(to_sfixed_a(-0.00012735059135593474)),(to_sfixed_a(2.1573832782451063e-06)),(to_sfixed_a(0.20142991840839386)),(to_sfixed_a(0.0019926647655665874)),(to_sfixed_a(0.19933202862739563)),(to_sfixed_a(2.8476701118052006e-05)),(to_sfixed_a(-0.00045032482012175024)),(to_sfixed_a(6.728377047693357e-05)),(to_sfixed_a(-0.00019383514882065356)),(to_sfixed_a(-0.23609140515327454)),(to_sfixed_a(0.5096491575241089)),(to_sfixed_a(3.617876427597366e-05)),(to_sfixed_a(1.683486334513873e-05)),(to_sfixed_a(0.00020285829668864608)),(to_sfixed_a(0.10052905976772308)),(to_sfixed_a(0.14588843286037445)),(to_sfixed_a(0.4560834765434265)),(to_sfixed_a(1.8566388462204486e-06)),(to_sfixed_a(0.00010864657815545797)),(to_sfixed_a(9.11920506041497e-06)),(to_sfixed_a(0.0030055269598960876)),(to_sfixed_a(-0.0054434072226285934)),(to_sfixed_a(0.17422431707382202)),(to_sfixed_a(0.00013880160986445844)),(to_sfixed_a(0.00019092141883447766)),(to_sfixed_a(0.00019323054584674537)),(to_sfixed_a(-0.29454946517944336)),(to_sfixed_a(0.00017994194058701396)),(to_sfixed_a(0.001071360893547535)),(to_sfixed_a(-0.00020053442858625203)),(to_sfixed_a(0.005243090447038412)),(to_sfixed_a(0.0004703705199062824)),(to_sfixed_a(0.37727048993110657)),(to_sfixed_a(-0.0007767313509248197)),(to_sfixed_a(-0.00011351343709975481)),(to_sfixed_a(0.18905971944332123)),(to_sfixed_a(0.016310956329107285)),(to_sfixed_a(-6.434749229811132e-05)),(to_sfixed_a(0.0006120280013419688)),(to_sfixed_a(0.00024368701269850135)),(to_sfixed_a(-0.00012274584150873125)),(to_sfixed_a(0.008522524498403072)),(to_sfixed_a(0.10351379960775375)),(to_sfixed_a(-4.536641790764406e-05)),(to_sfixed_a(-0.0002476563968230039)),(to_sfixed_a(0.003230493515729904)),(to_sfixed_a(-6.410744390450418e-05)),(to_sfixed_a(-0.41830599308013916)),(to_sfixed_a(0.0001569744636071846)),(to_sfixed_a(-4.4802458432968706e-05)),(to_sfixed_a(-6.49509092909284e-05)),(to_sfixed_a(0.00865948386490345)),(to_sfixed_a(-2.3550903279101476e-05)),(to_sfixed_a(0.00015023040759842843)),(to_sfixed_a(6.3864499679766595e-06)),(to_sfixed_a(0.004588947631418705)),(to_sfixed_a(0.01199676189571619)),(to_sfixed_a(-2.0517654775176197e-07)),(to_sfixed_a(-0.00015339608944486827)),(to_sfixed_a(-0.00041151835466735065)),(to_sfixed_a(-0.00011277063458692282)),(to_sfixed_a(0.014341229572892189)),(to_sfixed_a(0.016074402257800102)),(to_sfixed_a(0.0001263285957975313)),(to_sfixed_a(0.19884994626045227)),(to_sfixed_a(0.39691922068595886)),(to_sfixed_a(2.3360695195151493e-05)),(to_sfixed_a(0.0001172332267742604)),(to_sfixed_a(-0.0001192543059005402)),(to_sfixed_a(0.0001586202997714281)),(to_sfixed_a(-0.00019169662846252322)),(to_sfixed_a(-0.0001807674707379192)),(to_sfixed_a(1.3442995623336174e-06)),(to_sfixed_a(-0.005068455822765827)),(to_sfixed_a(0.00014958511746954173)),(to_sfixed_a(0.17415939271450043)),(to_sfixed_a(0.0020976215600967407)),(to_sfixed_a(0.007876832969486713)),(to_sfixed_a(-0.2591366767883301)),(to_sfixed_a(0.00010354076221119612)),(to_sfixed_a(0.06631049513816833)),(to_sfixed_a(-0.0017184449825435877)),(to_sfixed_a(0.014205435290932655)),(to_sfixed_a(-6.066940113669261e-05)),(to_sfixed_a(0.0031564312521368265)),(to_sfixed_a(-0.18049365282058716)),(to_sfixed_a(0.01249791495501995)));

    constant weight_n2_2 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.03955231234431267)),(to_sfixed_a(-0.019148925319314003)),(to_sfixed_a(-0.0008696437580510974)),(to_sfixed_a(-2.044631946773734e-05)),(to_sfixed_a(-0.0009482651948928833)),(to_sfixed_a(-0.00010839772585313767)),(to_sfixed_a(0.0012042538728564978)),(to_sfixed_a(-4.6095316065475345e-05)),(to_sfixed_a(-0.00011401988740544766)),(to_sfixed_a(0.00013008658424951136)),(to_sfixed_a(-0.00015795303625054657)),(to_sfixed_a(-0.00817969162017107)),(to_sfixed_a(0.28155481815338135)),(to_sfixed_a(-0.01195706706494093)),(to_sfixed_a(-0.00017450717859901488)),(to_sfixed_a(-0.00017105694860219955)),(to_sfixed_a(9.681381925474852e-06)),(to_sfixed_a(0.00014310010010376573)),(to_sfixed_a(-0.001107152784243226)),(to_sfixed_a(-0.002370130270719528)),(to_sfixed_a(3.827457840088755e-05)),(to_sfixed_a(4.5091743231751025e-05)),(to_sfixed_a(8.335162419825792e-06)),(to_sfixed_a(0.03564468026161194)),(to_sfixed_a(0.0010000292677432299)),(to_sfixed_a(-0.005422338843345642)),(to_sfixed_a(7.963104872033e-05)),(to_sfixed_a(-2.5640962121542543e-05)),(to_sfixed_a(0.0009685565601103008)),(to_sfixed_a(-4.746828562929295e-05)),(to_sfixed_a(0.00445939414203167)),(to_sfixed_a(0.00015874324890319258)),(to_sfixed_a(0.004136458970606327)),(to_sfixed_a(-1.704401074675843e-05)),(to_sfixed_a(7.761911547277123e-06)),(to_sfixed_a(7.814462878741324e-05)),(to_sfixed_a(0.21395140886306763)),(to_sfixed_a(0.024027789011597633)),(to_sfixed_a(-2.3170981876319274e-05)),(to_sfixed_a(0.00014983987784944475)),(to_sfixed_a(-0.2838882803916931)),(to_sfixed_a(9.437998232897371e-05)),(to_sfixed_a(-0.0002063833671854809)),(to_sfixed_a(-2.8985936296521686e-05)),(to_sfixed_a(-8.54067548061721e-06)),(to_sfixed_a(0.0013077222974970937)),(to_sfixed_a(3.5633211155072786e-06)),(to_sfixed_a(-4.5433789637172595e-06)),(to_sfixed_a(-0.00021517359709832817)),(to_sfixed_a(0.002202116884291172)),(to_sfixed_a(0.0007799723534844816)),(to_sfixed_a(-0.00016643131675664335)),(to_sfixed_a(1.2457094271667302e-05)),(to_sfixed_a(0.3276408314704895)),(to_sfixed_a(0.033003371208906174)),(to_sfixed_a(-0.023445066064596176)),(to_sfixed_a(-0.00016433358541689813)),(to_sfixed_a(0.0012084156041964889)),(to_sfixed_a(0.00016818908625282347)),(to_sfixed_a(-0.00011342031211825088)),(to_sfixed_a(4.698001794167794e-05)),(to_sfixed_a(0.00024684006348252296)),(to_sfixed_a(0.00040495622670277953)),(to_sfixed_a(-0.4869523346424103)),(to_sfixed_a(-6.082453910494223e-05)),(to_sfixed_a(0.24423231184482574)),(to_sfixed_a(7.007679232629016e-05)),(to_sfixed_a(-0.28444066643714905)),(to_sfixed_a(5.126983887748793e-05)),(to_sfixed_a(0.0001294496760237962)),(to_sfixed_a(-0.3011953830718994)),(to_sfixed_a(-0.3908132016658783)),(to_sfixed_a(0.0012733150506392121)),(to_sfixed_a(4.589090895024128e-05)),(to_sfixed_a(0.0001834297872846946)),(to_sfixed_a(-0.00017582577129360288)),(to_sfixed_a(-0.13137170672416687)),(to_sfixed_a(0.0014215053524821997)),(to_sfixed_a(0.00010830532119143754)),(to_sfixed_a(-0.003994747065007687)),(to_sfixed_a(-2.937748831755016e-06)),(to_sfixed_a(-0.00015666181570850313)),(to_sfixed_a(0.0006310823955573142)),(to_sfixed_a(4.6928653318900615e-06)),(to_sfixed_a(-2.283624780829996e-05)),(to_sfixed_a(-7.261569408001378e-06)),(to_sfixed_a(0.007348333019763231)),(to_sfixed_a(-2.72952820523642e-06)),(to_sfixed_a(-5.994435923639685e-06)),(to_sfixed_a(-0.00015325352433137596)),(to_sfixed_a(-5.876962859474588e-06)),(to_sfixed_a(-0.00018990162061527371)),(to_sfixed_a(0.008824077434837818)),(to_sfixed_a(3.297356306575239e-05)),(to_sfixed_a(-0.0029703467153012753)),(to_sfixed_a(-2.282461900904309e-05)),(to_sfixed_a(2.397684147581458e-05)),(to_sfixed_a(-5.295134906191379e-05)),(to_sfixed_a(-9.97233873931691e-05)),(to_sfixed_a(6.837413820903748e-06)),(to_sfixed_a(0.013239029794931412)),(to_sfixed_a(0.00045428265002556145)),(to_sfixed_a(3.6565241316566244e-05)),(to_sfixed_a(0.00039234539144672453)),(to_sfixed_a(4.675760283134878e-05)),(to_sfixed_a(3.692466634674929e-05)),(to_sfixed_a(4.527828423306346e-06)),(to_sfixed_a(-3.426857074373402e-05)),(to_sfixed_a(-0.0001576028880663216)),(to_sfixed_a(-0.39729923009872437)),(to_sfixed_a(0.002329785842448473)),(to_sfixed_a(-0.00011967499449383467)),(to_sfixed_a(0.002399349818006158)),(to_sfixed_a(1.3034208677709103e-05)),(to_sfixed_a(-0.0001363446790492162)),(to_sfixed_a(0.0014159911079332232)),(to_sfixed_a(0.013555475510656834)),(to_sfixed_a(-0.23819833993911743)),(to_sfixed_a(0.0004457532486412674)),(to_sfixed_a(-0.0013414528220891953)),(to_sfixed_a(0.00010325519542675465)),(to_sfixed_a(-1.4991601346991956e-06)),(to_sfixed_a(-8.796419933787547e-06)),(to_sfixed_a(-0.00010866673255804926)),(to_sfixed_a(4.53740794910118e-05)),(to_sfixed_a(-0.011491496115922928)),(to_sfixed_a(0.007831002585589886)),(to_sfixed_a(-0.00010122155072167516)),(to_sfixed_a(4.485467434278689e-05)),(to_sfixed_a(0.00020556450181175023)),(to_sfixed_a(1.0711846698541194e-05)),(to_sfixed_a(0.00014273291162680835)),(to_sfixed_a(-0.00016252111527137458)),(to_sfixed_a(-0.44425272941589355)),(to_sfixed_a(6.329829193418846e-05)),(to_sfixed_a(1.758872895152308e-05)),(to_sfixed_a(-0.0006980245234444737)),(to_sfixed_a(9.375009540235624e-06)),(to_sfixed_a(0.0002429070882499218)),(to_sfixed_a(-0.00010598882363410667)),(to_sfixed_a(6.616348400712013e-06)),(to_sfixed_a(-0.00010624275455484167)),(to_sfixed_a(0.00011517891107359901)),(to_sfixed_a(-0.00290560070425272)),(to_sfixed_a(0.0010342712048441172)),(to_sfixed_a(-4.773299951921217e-05)),(to_sfixed_a(-9.798195242183283e-05)),(to_sfixed_a(-7.739436841802672e-05)),(to_sfixed_a(4.291197910788469e-05)),(to_sfixed_a(0.0004457096219994128)),(to_sfixed_a(-0.0001164216228062287)),(to_sfixed_a(-0.00015104393241927028)),(to_sfixed_a(5.93444419791922e-05)),(to_sfixed_a(0.0004523209354374558)),(to_sfixed_a(-6.524276977870613e-05)),(to_sfixed_a(-0.00893430132418871)),(to_sfixed_a(3.346924495417625e-05)),(to_sfixed_a(0.002726121572777629)),(to_sfixed_a(-0.00014927706797607243)),(to_sfixed_a(5.7862016547005624e-05)),(to_sfixed_a(7.084964454406872e-05)),(to_sfixed_a(4.487257683649659e-06)),(to_sfixed_a(3.275966446381062e-05)),(to_sfixed_a(2.7423957362771034e-06)),(to_sfixed_a(6.38243873254396e-05)),(to_sfixed_a(-0.00040669666486792266)),(to_sfixed_a(7.592077599838376e-05)),(to_sfixed_a(0.0010984578402712941)),(to_sfixed_a(0.00011788733536377549)),(to_sfixed_a(-5.7628909416962415e-05)),(to_sfixed_a(0.19379599392414093)),(to_sfixed_a(0.002135002752766013)),(to_sfixed_a(-6.181978096719831e-05)),(to_sfixed_a(2.0654992113122717e-05)),(to_sfixed_a(0.31831637024879456)),(to_sfixed_a(2.1467294573085383e-06)),(to_sfixed_a(0.0010304473107680678)),(to_sfixed_a(2.41646575886989e-05)),(to_sfixed_a(-0.003330441890284419)),(to_sfixed_a(-0.02675768733024597)),(to_sfixed_a(3.283055411884561e-05)),(to_sfixed_a(0.0002387102722423151)),(to_sfixed_a(-0.00011674303095787764)),(to_sfixed_a(7.107111741788685e-05)),(to_sfixed_a(1.6792771930340677e-05)),(to_sfixed_a(-1.015991347230738e-05)),(to_sfixed_a(0.005456205923110247)),(to_sfixed_a(-0.0021357100922614336)),(to_sfixed_a(0.00010874112194869667)),(to_sfixed_a(0.0010701960418373346)),(to_sfixed_a(0.4001601040363312)),(to_sfixed_a(7.146720599848777e-05)),(to_sfixed_a(0.0015337216900661588)),(to_sfixed_a(-0.4595102369785309)),(to_sfixed_a(6.865539762657136e-05)),(to_sfixed_a(-0.006119419354945421)),(to_sfixed_a(6.55420299153775e-05)),(to_sfixed_a(0.01006265077739954)),(to_sfixed_a(-0.09429086744785309)),(to_sfixed_a(-0.00024666174431331456)),(to_sfixed_a(6.651649891864508e-05)),(to_sfixed_a(-7.851229020161554e-05)),(to_sfixed_a(0.00024369738821405917)),(to_sfixed_a(0.00018271389126311988)),(to_sfixed_a(-0.00017765641678124666)),(to_sfixed_a(-0.00033963093301281333)),(to_sfixed_a(-0.03907923027873039)),(to_sfixed_a(-0.014986705034971237)),(to_sfixed_a(0.0008257119916379452)),(to_sfixed_a(0.002139095216989517)),(to_sfixed_a(-0.00031351298093795776)),(to_sfixed_a(-0.00015142481424845755)),(to_sfixed_a(0.00024000411212909967)),(to_sfixed_a(-2.5365545297972858e-05)),(to_sfixed_a(-0.00016060721827670932)),(to_sfixed_a(3.6565863410942256e-05)),(to_sfixed_a(0.0019671705085784197)),(to_sfixed_a(-0.04737890884280205)),(to_sfixed_a(0.0012371808988973498)),(to_sfixed_a(-0.00014987291069701314)),(to_sfixed_a(-1.1258103768341243e-05)),(to_sfixed_a(0.00028928296524100006)),(to_sfixed_a(1.0024647053796798e-05)),(to_sfixed_a(1.3370958185987547e-05)),(to_sfixed_a(-1.0637857485562563e-05)),(to_sfixed_a(-0.00023031304590404034)),(to_sfixed_a(0.00010059537453344092)),(to_sfixed_a(7.623159763170406e-05)),(to_sfixed_a(0.00034419671283103526)),(to_sfixed_a(0.400529146194458)),(to_sfixed_a(-0.33347275853157043)),(to_sfixed_a(5.758833140134811e-06)),(to_sfixed_a(0.0003015384718310088)),(to_sfixed_a(-0.0002212945546489209)),(to_sfixed_a(6.92315079504624e-05)),(to_sfixed_a(0.003458113642409444)),(to_sfixed_a(-0.5927390456199646)),(to_sfixed_a(-0.00037721285480074584)),(to_sfixed_a(0.0004280005523469299)),(to_sfixed_a(-0.00028711959021165967)),(to_sfixed_a(0.0004944583051837981)),(to_sfixed_a(5.81259373575449e-05)),(to_sfixed_a(0.3567376732826233)),(to_sfixed_a(-0.0002973996743094176)),(to_sfixed_a(0.00016398978186771274)),(to_sfixed_a(0.00023234722902998328)),(to_sfixed_a(-0.015813304111361504)),(to_sfixed_a(-0.05991513282060623)),(to_sfixed_a(-2.0724537534988485e-05)),(to_sfixed_a(-9.941533789969981e-05)),(to_sfixed_a(0.00017214633408002555)),(to_sfixed_a(-0.0001913029554998502)),(to_sfixed_a(0.17313121259212494)),(to_sfixed_a(-7.8373916039709e-05)),(to_sfixed_a(-2.2902491764398292e-05)),(to_sfixed_a(0.0012438171543180943)),(to_sfixed_a(-5.427118594525382e-06)),(to_sfixed_a(-0.00015336228534579277)),(to_sfixed_a(-0.00013762630987912416)),(to_sfixed_a(-0.00465245358645916)),(to_sfixed_a(0.00018544610065873712)),(to_sfixed_a(2.7418216632213444e-05)),(to_sfixed_a(0.00011673678818624467)),(to_sfixed_a(1.18673087854404e-05)),(to_sfixed_a(5.721200432162732e-05)),(to_sfixed_a(0.0016550999134778976)),(to_sfixed_a(-4.931637522531673e-05)),(to_sfixed_a(-0.0001475833123549819)),(to_sfixed_a(-0.00015318648365791887)),(to_sfixed_a(-0.2277638167142868)),(to_sfixed_a(-0.00327738793566823)),(to_sfixed_a(-0.00025065435329452157)),(to_sfixed_a(-0.0003063681651838124)),(to_sfixed_a(1.860088377725333e-05)),(to_sfixed_a(-9.961282921722159e-05)),(to_sfixed_a(0.0005425019189715385)),(to_sfixed_a(0.00213454756885767)),(to_sfixed_a(-1.6300591596518643e-06)),(to_sfixed_a(-0.41925203800201416)),(to_sfixed_a(0.005653387866914272)),(to_sfixed_a(3.022466626134701e-05)),(to_sfixed_a(8.472114859614521e-05)),(to_sfixed_a(0.00015220293425954878)),(to_sfixed_a(-0.00020937428053002805)),(to_sfixed_a(-3.772874697460793e-05)),(to_sfixed_a(6.0120466514490545e-05)),(to_sfixed_a(0.004131362773478031)),(to_sfixed_a(0.07336941361427307)),(to_sfixed_a(-1.4318364264909178e-05)),(to_sfixed_a(-7.135715713957325e-05)),(to_sfixed_a(0.0009086515055969357)),(to_sfixed_a(0.006533759646117687)),(to_sfixed_a(-0.001838530763052404)),(to_sfixed_a(0.00017421602387912571)),(to_sfixed_a(0.003151330631226301)),(to_sfixed_a(0.2863685190677643)),(to_sfixed_a(0.0001864525256678462)),(to_sfixed_a(-0.0001406717929057777)),(to_sfixed_a(5.1772829465335235e-05)),(to_sfixed_a(-0.003435153979808092)),(to_sfixed_a(-0.00030218128813430667)));

    constant weight_n2_3 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.007740584667772055)),(to_sfixed_a(-6.750931788701564e-05)),(to_sfixed_a(0.0001923435484059155)),(to_sfixed_a(0.0001522120728623122)),(to_sfixed_a(-0.00013622251572087407)),(to_sfixed_a(-9.593717550160363e-05)),(to_sfixed_a(-0.0001822981284931302)),(to_sfixed_a(-0.0001052239749697037)),(to_sfixed_a(0.0001533032045699656)),(to_sfixed_a(-0.000154206165461801)),(to_sfixed_a(-0.00015681525110267103)),(to_sfixed_a(-2.072980350931175e-06)),(to_sfixed_a(-0.00011391338193789124)),(to_sfixed_a(-0.00024328078143298626)),(to_sfixed_a(-2.962484722957015e-05)),(to_sfixed_a(-7.042684592306614e-05)),(to_sfixed_a(0.00024165875220205635)),(to_sfixed_a(1.1888805602211505e-05)),(to_sfixed_a(0.00011313244613120332)),(to_sfixed_a(-0.0002701851481106132)),(to_sfixed_a(7.12782348273322e-05)),(to_sfixed_a(0.00010759717406472191)),(to_sfixed_a(-1.9491028069751337e-05)),(to_sfixed_a(0.00018645450472831726)),(to_sfixed_a(0.0001985708368010819)),(to_sfixed_a(-0.00013424627832137048)),(to_sfixed_a(-1.8516191630624235e-05)),(to_sfixed_a(0.00027760976809076965)),(to_sfixed_a(4.406006701174192e-05)),(to_sfixed_a(-0.0002875840582419187)),(to_sfixed_a(-0.0003759747778531164)),(to_sfixed_a(-6.854824459878728e-05)),(to_sfixed_a(1.2167420209152624e-05)),(to_sfixed_a(-8.251470717368647e-05)),(to_sfixed_a(0.0001578905648784712)),(to_sfixed_a(-4.996170900994912e-06)),(to_sfixed_a(6.715530616929755e-05)),(to_sfixed_a(-1.665226591285318e-05)),(to_sfixed_a(0.00013014423893764615)),(to_sfixed_a(-0.00015367490414064378)),(to_sfixed_a(0.00016673983191139996)),(to_sfixed_a(6.165671220514923e-05)),(to_sfixed_a(4.506880941335112e-05)),(to_sfixed_a(-0.00010837590525625274)),(to_sfixed_a(-7.148667646106333e-05)),(to_sfixed_a(0.00016883076750673354)),(to_sfixed_a(0.00024059780116658658)),(to_sfixed_a(-1.1778211046475917e-06)),(to_sfixed_a(0.0001140205204137601)),(to_sfixed_a(-0.00010286309407092631)),(to_sfixed_a(0.00019591290038079023)),(to_sfixed_a(0.00010379010200267658)),(to_sfixed_a(0.0003000791766680777)),(to_sfixed_a(-2.422473335172981e-05)),(to_sfixed_a(-0.00024769376614131033)),(to_sfixed_a(0.00020541853155009449)),(to_sfixed_a(-0.00015663787780795246)),(to_sfixed_a(-0.00015734744374640286)),(to_sfixed_a(0.0002922594721894711)),(to_sfixed_a(-1.1296113370917737e-05)),(to_sfixed_a(-0.0002012351615121588)),(to_sfixed_a(3.7379140849225223e-06)),(to_sfixed_a(-7.852238195482641e-05)),(to_sfixed_a(-1.112715108320117e-05)),(to_sfixed_a(-5.782426887890324e-05)),(to_sfixed_a(-6.0481488617369905e-05)),(to_sfixed_a(0.00018371225451119244)),(to_sfixed_a(-0.00017530818877276033)),(to_sfixed_a(-0.00011982407158939168)),(to_sfixed_a(-0.0002480612602084875)),(to_sfixed_a(-0.00011680874740704894)),(to_sfixed_a(-0.0001267248298972845)),(to_sfixed_a(0.00020380601927172393)),(to_sfixed_a(0.0001803253253456205)),(to_sfixed_a(6.64312465232797e-05)),(to_sfixed_a(-0.00013874647265765816)),(to_sfixed_a(3.754073622985743e-05)),(to_sfixed_a(-2.1483712771441787e-05)),(to_sfixed_a(-6.914781988598406e-05)),(to_sfixed_a(-0.00011178625572938472)),(to_sfixed_a(-5.7358840422239155e-05)),(to_sfixed_a(-0.00022073024592828006)),(to_sfixed_a(3.8286816561594605e-05)),(to_sfixed_a(-1.5345911378972232e-05)),(to_sfixed_a(-7.494804594898596e-05)),(to_sfixed_a(-0.00015111554239410907)),(to_sfixed_a(-0.000246017356403172)),(to_sfixed_a(-4.4008775148540735e-06)),(to_sfixed_a(-4.36652080679778e-05)),(to_sfixed_a(-6.963872874621302e-05)),(to_sfixed_a(2.4644552468089387e-05)),(to_sfixed_a(-0.0003058114380110055)),(to_sfixed_a(0.0003138573665637523)),(to_sfixed_a(3.7358699046308175e-05)),(to_sfixed_a(-0.00025197939248755574)),(to_sfixed_a(0.0001142383407568559)),(to_sfixed_a(-0.00017508228484075516)),(to_sfixed_a(7.107650162652135e-05)),(to_sfixed_a(-7.007969543337822e-06)),(to_sfixed_a(-6.609030242543668e-05)),(to_sfixed_a(4.798539157491177e-05)),(to_sfixed_a(-0.00019480804621707648)),(to_sfixed_a(0.00025146128609776497)),(to_sfixed_a(-6.729837332386523e-05)),(to_sfixed_a(-8.68791903485544e-05)),(to_sfixed_a(0.00011453617480583489)),(to_sfixed_a(-5.757990584243089e-05)),(to_sfixed_a(-0.00016818390577100217)),(to_sfixed_a(8.476887160213664e-05)),(to_sfixed_a(-9.24163541640155e-05)),(to_sfixed_a(-7.830934919184074e-05)),(to_sfixed_a(-0.00010587837459752336)),(to_sfixed_a(3.896684211213142e-05)),(to_sfixed_a(-4.211997293168679e-06)),(to_sfixed_a(-1.4916106010787189e-05)),(to_sfixed_a(0.00017027737339958549)),(to_sfixed_a(-8.707409142516553e-05)),(to_sfixed_a(-4.3293548515066504e-06)),(to_sfixed_a(-0.00015592173440381885)),(to_sfixed_a(0.00025028848904184997)),(to_sfixed_a(3.9031379856169224e-05)),(to_sfixed_a(-4.0320155676454306e-06)),(to_sfixed_a(0.00014695347636006773)),(to_sfixed_a(6.402533472282812e-07)),(to_sfixed_a(2.223876799689606e-05)),(to_sfixed_a(-3.769466275116429e-05)),(to_sfixed_a(9.792722266865894e-05)),(to_sfixed_a(1.0364523404859938e-05)),(to_sfixed_a(-0.00028420687885954976)),(to_sfixed_a(0.00028920595650561154)),(to_sfixed_a(-0.00013618086813949049)),(to_sfixed_a(-7.102253584889695e-05)),(to_sfixed_a(1.0346469935029745e-05)),(to_sfixed_a(-1.0706951798056252e-05)),(to_sfixed_a(-0.0002229366364190355)),(to_sfixed_a(-3.2640098652336746e-05)),(to_sfixed_a(1.0210205800831318e-05)),(to_sfixed_a(3.526296859490685e-05)),(to_sfixed_a(-6.648282578680664e-05)),(to_sfixed_a(-7.038432522676885e-05)),(to_sfixed_a(3.092103361268528e-05)),(to_sfixed_a(3.680909867398441e-05)),(to_sfixed_a(6.51837108307518e-05)),(to_sfixed_a(7.393541454803199e-05)),(to_sfixed_a(-0.00014880436356179416)),(to_sfixed_a(-7.073853339534253e-05)),(to_sfixed_a(0.0002892753982450813)),(to_sfixed_a(0.00010079440107801929)),(to_sfixed_a(-5.296044400893152e-05)),(to_sfixed_a(0.00018339364032726735)),(to_sfixed_a(3.01731051877141e-06)),(to_sfixed_a(7.127369462978095e-05)),(to_sfixed_a(-0.00017482541443314403)),(to_sfixed_a(-0.0002096860553137958)),(to_sfixed_a(1.0584626579657197e-05)),(to_sfixed_a(-2.6707581127993762e-05)),(to_sfixed_a(6.873628444736823e-05)),(to_sfixed_a(0.0001291045336984098)),(to_sfixed_a(-0.00010471278801560402)),(to_sfixed_a(8.08590411907062e-05)),(to_sfixed_a(-0.0002501612761989236)),(to_sfixed_a(-7.821520557627082e-05)),(to_sfixed_a(0.00020853776368312538)),(to_sfixed_a(-8.238490408984944e-05)),(to_sfixed_a(5.703095666831359e-05)),(to_sfixed_a(-5.7684999774210155e-05)),(to_sfixed_a(-1.432881981600076e-05)),(to_sfixed_a(-0.00011653183901216835)),(to_sfixed_a(-5.200706436880864e-05)),(to_sfixed_a(-0.00011699590686475858)),(to_sfixed_a(0.00011649603402474895)),(to_sfixed_a(-4.501394505496137e-05)),(to_sfixed_a(6.128264794824645e-05)),(to_sfixed_a(0.00023879132641013712)),(to_sfixed_a(0.00027364518609829247)),(to_sfixed_a(-0.00024675909662619233)),(to_sfixed_a(6.108463276177645e-05)),(to_sfixed_a(4.088535206392407e-06)),(to_sfixed_a(7.162422116380185e-05)),(to_sfixed_a(-0.00028105449746362865)),(to_sfixed_a(-0.0003163228102494031)),(to_sfixed_a(-0.00011373585584806278)),(to_sfixed_a(7.273921073647216e-05)),(to_sfixed_a(-3.896978887496516e-05)),(to_sfixed_a(-0.00013670364569406956)),(to_sfixed_a(-0.000291316129732877)),(to_sfixed_a(-3.952307451982051e-05)),(to_sfixed_a(-0.00013729938655160367)),(to_sfixed_a(-1.35546360979788e-05)),(to_sfixed_a(8.863376569934189e-05)),(to_sfixed_a(-0.00010856725566554815)),(to_sfixed_a(-0.00019242143025621772)),(to_sfixed_a(6.819171539973468e-05)),(to_sfixed_a(5.295532901072875e-05)),(to_sfixed_a(-0.00014869449660182)),(to_sfixed_a(2.9033792088739574e-05)),(to_sfixed_a(4.0899423765949905e-05)),(to_sfixed_a(0.0001951012818608433)),(to_sfixed_a(-0.00012075643462594599)),(to_sfixed_a(-3.533059498295188e-06)),(to_sfixed_a(-4.6210399887058884e-05)),(to_sfixed_a(-0.00017315236618742347)),(to_sfixed_a(-0.00013124954421073198)),(to_sfixed_a(-0.00012973518460057676)),(to_sfixed_a(2.612131356727332e-05)),(to_sfixed_a(-0.000185277676791884)),(to_sfixed_a(-3.365686279721558e-05)),(to_sfixed_a(1.2717035133391619e-05)),(to_sfixed_a(7.201004336820915e-05)),(to_sfixed_a(-1.7680526070762426e-05)),(to_sfixed_a(6.774303619749844e-05)),(to_sfixed_a(-0.0001937738707056269)),(to_sfixed_a(1.5241421351674944e-05)),(to_sfixed_a(-0.0001050718710757792)),(to_sfixed_a(-1.0363321052864194e-05)),(to_sfixed_a(1.9642617189674638e-05)),(to_sfixed_a(-0.000112843161332421)),(to_sfixed_a(-7.278230623342097e-05)),(to_sfixed_a(0.00010652674973243847)),(to_sfixed_a(0.00029238127171993256)),(to_sfixed_a(-0.0001884014200186357)),(to_sfixed_a(-0.00010850593389477581)),(to_sfixed_a(-0.0001487669360358268)),(to_sfixed_a(-0.00010009243851527572)),(to_sfixed_a(-4.672867362387478e-06)),(to_sfixed_a(0.00038230782956816256)),(to_sfixed_a(5.773087468696758e-05)),(to_sfixed_a(2.8027716325595975e-05)),(to_sfixed_a(-7.340728188864887e-05)),(to_sfixed_a(0.00010685468441806734)),(to_sfixed_a(6.720286910422146e-05)),(to_sfixed_a(0.0002169489162042737)),(to_sfixed_a(-0.00012950002565048635)),(to_sfixed_a(0.00017900530656334013)),(to_sfixed_a(-0.00020130653865635395)),(to_sfixed_a(-2.1514977561309934e-05)),(to_sfixed_a(3.9062990254024044e-05)),(to_sfixed_a(0.0001048676494974643)),(to_sfixed_a(-7.125853153411299e-05)),(to_sfixed_a(-0.00015015866665635258)),(to_sfixed_a(-0.0001283346355194226)),(to_sfixed_a(6.769183528376743e-05)),(to_sfixed_a(0.00012049036013195291)),(to_sfixed_a(0.00011223065666854382)),(to_sfixed_a(-1.208136382047087e-05)),(to_sfixed_a(0.00014910835307091475)),(to_sfixed_a(-2.834852784872055e-05)),(to_sfixed_a(6.920233863638714e-05)),(to_sfixed_a(-3.6867480957880616e-05)),(to_sfixed_a(8.675386925460771e-05)),(to_sfixed_a(-0.0002488226455170661)),(to_sfixed_a(0.00011390974395908415)),(to_sfixed_a(-5.583875463344157e-06)),(to_sfixed_a(0.00010641725384630263)),(to_sfixed_a(0.00015666615217924118)),(to_sfixed_a(-0.000448350008809939)),(to_sfixed_a(-7.953307795105502e-05)),(to_sfixed_a(-5.891280306968838e-05)),(to_sfixed_a(8.952191274147481e-05)),(to_sfixed_a(0.0002975659444928169)),(to_sfixed_a(-7.138049113564193e-05)),(to_sfixed_a(5.906422666157596e-05)),(to_sfixed_a(-0.00010081368964165449)),(to_sfixed_a(5.719756882172078e-05)),(to_sfixed_a(-0.00011683156481012702)),(to_sfixed_a(4.548845026874915e-06)),(to_sfixed_a(-6.982730701565742e-05)),(to_sfixed_a(-7.808180816937238e-05)),(to_sfixed_a(0.000242738620727323)),(to_sfixed_a(-3.067791840294376e-05)),(to_sfixed_a(0.00011268164962530136)),(to_sfixed_a(6.784722791053355e-05)),(to_sfixed_a(0.00031390751246362925)),(to_sfixed_a(0.00015904138854239136)),(to_sfixed_a(-0.0001885162782855332)),(to_sfixed_a(-4.459933552425355e-05)),(to_sfixed_a(-0.00012746002175845206)),(to_sfixed_a(-0.00011544136941665784)),(to_sfixed_a(-0.00013581718667410314)),(to_sfixed_a(-0.00015682254161220044)),(to_sfixed_a(0.0002419882221147418)),(to_sfixed_a(-0.0002173446409869939)),(to_sfixed_a(3.21953630191274e-05)),(to_sfixed_a(-0.00014648148498963565)),(to_sfixed_a(-0.0001368733064737171)),(to_sfixed_a(-7.141949026845396e-05)),(to_sfixed_a(-1.5838566469028592e-05)),(to_sfixed_a(0.00018750438175629824)),(to_sfixed_a(-1.0121482773683965e-05)),(to_sfixed_a(6.611261051148176e-05)),(to_sfixed_a(7.264682790264487e-05)),(to_sfixed_a(-4.052351869177073e-06)),(to_sfixed_a(-5.920762487221509e-05)),(to_sfixed_a(-2.079268051602412e-05)),(to_sfixed_a(-0.00017494325584266335)),(to_sfixed_a(-8.483888814225793e-05)),(to_sfixed_a(1.7454229237046093e-05)),(to_sfixed_a(3.9275080780498683e-05)),(to_sfixed_a(-0.00022846889623906463)),(to_sfixed_a(2.3154665541369468e-05)),(to_sfixed_a(-1.5326804714277387e-06)));

    constant weight_n2_4 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.31671884655952454)),(to_sfixed_a(-7.79757319833152e-05)),(to_sfixed_a(-9.329075692221522e-05)),(to_sfixed_a(-0.00022229657042771578)),(to_sfixed_a(7.786128844600171e-05)),(to_sfixed_a(-0.00021766126155853271)),(to_sfixed_a(-0.00010749198554549366)),(to_sfixed_a(-7.227936293929815e-05)),(to_sfixed_a(4.4531450839713216e-05)),(to_sfixed_a(0.00014635580009780824)),(to_sfixed_a(-7.147369615267962e-05)),(to_sfixed_a(7.031046698102728e-05)),(to_sfixed_a(8.255762077169493e-05)),(to_sfixed_a(5.7926787121687084e-05)),(to_sfixed_a(-4.531759623205289e-05)),(to_sfixed_a(-0.00012836442328989506)),(to_sfixed_a(1.4143253793008626e-05)),(to_sfixed_a(-0.00011183533933945)),(to_sfixed_a(-7.753628597129136e-05)),(to_sfixed_a(-0.00014864225522615016)),(to_sfixed_a(-0.00016241907724179327)),(to_sfixed_a(-0.00015425003948621452)),(to_sfixed_a(0.00028239371022209525)),(to_sfixed_a(-0.000176361805642955)),(to_sfixed_a(-0.00010471419955138117)),(to_sfixed_a(0.00018095967243425548)),(to_sfixed_a(0.00018077896675094962)),(to_sfixed_a(0.00015475966210942715)),(to_sfixed_a(-5.423644324764609e-07)),(to_sfixed_a(-0.0002477885573171079)),(to_sfixed_a(-7.301154255401343e-06)),(to_sfixed_a(-0.00016171307652257383)),(to_sfixed_a(-2.213520201621577e-05)),(to_sfixed_a(-0.00030149545636959374)),(to_sfixed_a(3.2677566196070984e-05)),(to_sfixed_a(7.996040949365124e-05)),(to_sfixed_a(-0.00011219541192986071)),(to_sfixed_a(2.6405221433378756e-05)),(to_sfixed_a(0.00013062532525509596)),(to_sfixed_a(-4.584027919918299e-06)),(to_sfixed_a(-6.946077337488532e-05)),(to_sfixed_a(6.835134990978986e-05)),(to_sfixed_a(-6.163265788927674e-05)),(to_sfixed_a(1.2828255421482027e-05)),(to_sfixed_a(-5.8503414038568735e-05)),(to_sfixed_a(-0.00016792632231954485)),(to_sfixed_a(0.0001673837541602552)),(to_sfixed_a(6.884850154165179e-05)),(to_sfixed_a(0.00015437659749295563)),(to_sfixed_a(-1.6999809304252267e-05)),(to_sfixed_a(5.2536590374074876e-05)),(to_sfixed_a(0.00011286504013696685)),(to_sfixed_a(-0.00013824165216647089)),(to_sfixed_a(-1.6905614756979048e-06)),(to_sfixed_a(5.631803651340306e-05)),(to_sfixed_a(-9.108279482461512e-05)),(to_sfixed_a(-0.00015488281496800482)),(to_sfixed_a(5.469555617310107e-07)),(to_sfixed_a(-0.0001823448546929285)),(to_sfixed_a(-0.00013532614684663713)),(to_sfixed_a(6.909073272254318e-05)),(to_sfixed_a(0.0001547507563373074)),(to_sfixed_a(4.41471638623625e-06)),(to_sfixed_a(-6.057283826521598e-05)),(to_sfixed_a(4.751775122713298e-06)),(to_sfixed_a(-0.0002852577017620206)),(to_sfixed_a(-0.00028302485588938)),(to_sfixed_a(0.0001697848638286814)),(to_sfixed_a(0.00016890074766706675)),(to_sfixed_a(0.00010639776883181185)),(to_sfixed_a(0.00019618759688455611)),(to_sfixed_a(-9.502274042461067e-05)),(to_sfixed_a(0.000246977258939296)),(to_sfixed_a(-7.023103535175323e-05)),(to_sfixed_a(9.116799628827721e-05)),(to_sfixed_a(-3.372895298525691e-05)),(to_sfixed_a(-4.304938192944974e-05)),(to_sfixed_a(-0.0002646452630870044)),(to_sfixed_a(-0.0002673296257853508)),(to_sfixed_a(-5.416528438217938e-06)),(to_sfixed_a(-2.302782377228141e-06)),(to_sfixed_a(-8.167067426256835e-05)),(to_sfixed_a(-0.0002126839099219069)),(to_sfixed_a(0.00029234460089355707)),(to_sfixed_a(4.977748176315799e-06)),(to_sfixed_a(-0.00019535001774784178)),(to_sfixed_a(-0.00014934818318579346)),(to_sfixed_a(9.662935553933494e-06)),(to_sfixed_a(6.732322799507529e-05)),(to_sfixed_a(7.004116923781112e-05)),(to_sfixed_a(-0.00028528799884952605)),(to_sfixed_a(0.00037640391383320093)),(to_sfixed_a(0.0002547256590332836)),(to_sfixed_a(-2.2466101654572412e-05)),(to_sfixed_a(2.9514638299588114e-05)),(to_sfixed_a(0.00011401281517464668)),(to_sfixed_a(-7.217891106847674e-05)),(to_sfixed_a(5.897018127143383e-06)),(to_sfixed_a(-0.00017412498709745705)),(to_sfixed_a(-8.278760651592165e-05)),(to_sfixed_a(-0.00015600120241288096)),(to_sfixed_a(-4.876144157606177e-05)),(to_sfixed_a(8.937480743043125e-05)),(to_sfixed_a(0.00010829311213456094)),(to_sfixed_a(-0.0003741882974281907)),(to_sfixed_a(-0.00010644538269843906)),(to_sfixed_a(-7.037406612653285e-05)),(to_sfixed_a(-0.00044690375216305256)),(to_sfixed_a(4.3933585402555764e-05)),(to_sfixed_a(-9.096143185161054e-05)),(to_sfixed_a(-4.0504364733351395e-05)),(to_sfixed_a(0.00015443461597897112)),(to_sfixed_a(-1.612680352991447e-05)),(to_sfixed_a(-2.4649400074849837e-05)),(to_sfixed_a(7.468104740837589e-05)),(to_sfixed_a(-0.00021372086484916508)),(to_sfixed_a(0.00023868704738561064)),(to_sfixed_a(0.0001552923204144463)),(to_sfixed_a(0.0003098099841736257)),(to_sfixed_a(-1.654891821090132e-05)),(to_sfixed_a(1.0040785127785057e-06)),(to_sfixed_a(0.00017672794638201594)),(to_sfixed_a(-0.0001573598856339231)),(to_sfixed_a(-0.00011549566988833249)),(to_sfixed_a(1.772275209077634e-05)),(to_sfixed_a(6.865945033496246e-05)),(to_sfixed_a(-0.00016774970572441816)),(to_sfixed_a(3.862376615870744e-05)),(to_sfixed_a(-0.0002843707916326821)),(to_sfixed_a(0.00028602004749700427)),(to_sfixed_a(-7.004493090789765e-05)),(to_sfixed_a(-6.915735139045864e-05)),(to_sfixed_a(0.00038395042065531015)),(to_sfixed_a(0.00014973175711929798)),(to_sfixed_a(-0.0001350999518763274)),(to_sfixed_a(-0.0002120661229128018)),(to_sfixed_a(3.1757677788846195e-05)),(to_sfixed_a(0.0001695563696557656)),(to_sfixed_a(3.909341467078775e-05)),(to_sfixed_a(-5.07899749209173e-05)),(to_sfixed_a(0.00032204881426878273)),(to_sfixed_a(1.8808867025654763e-05)),(to_sfixed_a(-0.0001536842464702204)),(to_sfixed_a(1.1461601388873532e-05)),(to_sfixed_a(0.00014178288984112442)),(to_sfixed_a(5.163343666936271e-05)),(to_sfixed_a(2.8783513698726892e-05)),(to_sfixed_a(-0.0002997973351739347)),(to_sfixed_a(3.742272383533418e-06)),(to_sfixed_a(4.048612026963383e-06)),(to_sfixed_a(0.0001806912332540378)),(to_sfixed_a(2.025110188696999e-05)),(to_sfixed_a(-3.8868674892000854e-05)),(to_sfixed_a(0.00011330514098517597)),(to_sfixed_a(-0.00041773583507165313)),(to_sfixed_a(0.00014849210856482387)),(to_sfixed_a(2.595530531834811e-05)),(to_sfixed_a(-0.00011371754226274788)),(to_sfixed_a(-0.0001392961567034945)),(to_sfixed_a(-2.425644197501242e-05)),(to_sfixed_a(3.0208713724277914e-05)),(to_sfixed_a(4.2809548176592216e-05)),(to_sfixed_a(4.63727192254737e-05)),(to_sfixed_a(-2.1023333829361945e-05)),(to_sfixed_a(2.478725218679756e-05)),(to_sfixed_a(-0.00016790714289527386)),(to_sfixed_a(-0.00011868079309351742)),(to_sfixed_a(5.794676690129563e-05)),(to_sfixed_a(0.0003015809052158147)),(to_sfixed_a(-3.709223528858274e-05)),(to_sfixed_a(1.9104714738205075e-05)),(to_sfixed_a(-1.1331954738125205e-05)),(to_sfixed_a(-3.6868172173853964e-05)),(to_sfixed_a(6.386890891008079e-05)),(to_sfixed_a(-6.850301724625751e-05)),(to_sfixed_a(0.00014771393034607172)),(to_sfixed_a(5.330366548150778e-08)),(to_sfixed_a(0.00011534554505487904)),(to_sfixed_a(-0.00016858884191606194)),(to_sfixed_a(-2.3128512111725286e-05)),(to_sfixed_a(-0.00011353186710039154)),(to_sfixed_a(-7.344193727476522e-05)),(to_sfixed_a(-6.815539381932467e-05)),(to_sfixed_a(5.657603105646558e-05)),(to_sfixed_a(-6.695660704281181e-05)),(to_sfixed_a(9.146597585640848e-05)),(to_sfixed_a(0.00011544707376742736)),(to_sfixed_a(-1.5005163731984794e-05)),(to_sfixed_a(-1.2558841262944043e-05)),(to_sfixed_a(-1.1753581929951906e-07)),(to_sfixed_a(-0.00021929747890681028)),(to_sfixed_a(0.00023337677703239024)),(to_sfixed_a(1.0275107342749834e-07)),(to_sfixed_a(6.923734326846898e-05)),(to_sfixed_a(-5.039306415710598e-06)),(to_sfixed_a(5.132577280164696e-05)),(to_sfixed_a(1.1236839782213792e-05)),(to_sfixed_a(4.342052125139162e-05)),(to_sfixed_a(0.00031684033456258476)),(to_sfixed_a(8.435027848463506e-05)),(to_sfixed_a(7.758604624541476e-05)),(to_sfixed_a(-0.00017479629605077207)),(to_sfixed_a(0.00020074195344932377)),(to_sfixed_a(-1.8498540157452226e-05)),(to_sfixed_a(-5.791020521428436e-05)),(to_sfixed_a(-6.818593828938901e-05)),(to_sfixed_a(6.722086982335895e-05)),(to_sfixed_a(8.581798465456814e-05)),(to_sfixed_a(-6.564932118635625e-05)),(to_sfixed_a(0.00021846065646968782)),(to_sfixed_a(1.1964184523094445e-06)),(to_sfixed_a(0.00010570694576017559)),(to_sfixed_a(-6.142090569483116e-05)),(to_sfixed_a(-0.00018645788077265024)),(to_sfixed_a(-0.00018915743567049503)),(to_sfixed_a(0.00010264242882840335)),(to_sfixed_a(3.263277903897688e-05)),(to_sfixed_a(0.0002519081172067672)),(to_sfixed_a(0.00017434614710509777)),(to_sfixed_a(-0.00020595778187271208)),(to_sfixed_a(0.00012958937440998852)),(to_sfixed_a(-1.8899409042205662e-06)),(to_sfixed_a(0.0004497824120335281)),(to_sfixed_a(-0.000287855276837945)),(to_sfixed_a(3.883015597239137e-05)),(to_sfixed_a(-1.139060259447433e-05)),(to_sfixed_a(-0.00024665554519742727)),(to_sfixed_a(-4.1689054341986775e-06)),(to_sfixed_a(-2.493720967322588e-05)),(to_sfixed_a(0.00014033925253897905)),(to_sfixed_a(0.00017506693257018924)),(to_sfixed_a(-0.00015692412853240967)),(to_sfixed_a(-0.0004595473292283714)),(to_sfixed_a(5.554204108193517e-06)),(to_sfixed_a(0.00025532866129651666)),(to_sfixed_a(-5.6681819842197e-06)),(to_sfixed_a(-3.412738078623079e-05)),(to_sfixed_a(0.0002354732423555106)),(to_sfixed_a(0.00017545963055454195)),(to_sfixed_a(-6.130342080723494e-05)),(to_sfixed_a(2.418482836219482e-05)),(to_sfixed_a(-6.766474689356983e-05)),(to_sfixed_a(-0.00013987146667204797)),(to_sfixed_a(-0.00012843564036302269)),(to_sfixed_a(-2.0204955944791436e-05)),(to_sfixed_a(-6.846994801890105e-05)),(to_sfixed_a(-4.776735295308754e-06)),(to_sfixed_a(7.228187314467505e-05)),(to_sfixed_a(6.935586134204641e-05)),(to_sfixed_a(-0.0001465928362449631)),(to_sfixed_a(3.146280869259499e-05)),(to_sfixed_a(1.218635225086473e-05)),(to_sfixed_a(-8.799906936474144e-08)),(to_sfixed_a(4.065470420755446e-06)),(to_sfixed_a(1.692720252322033e-05)),(to_sfixed_a(-5.660560418618843e-05)),(to_sfixed_a(-1.5535060811089352e-05)),(to_sfixed_a(0.000291523669147864)),(to_sfixed_a(-2.2713767975801602e-05)),(to_sfixed_a(-0.00010014694998972118)),(to_sfixed_a(1.954444269358646e-05)),(to_sfixed_a(2.375194526393898e-05)),(to_sfixed_a(0.0002465518191456795)),(to_sfixed_a(1.0824951459653676e-05)),(to_sfixed_a(0.00023838115157559514)),(to_sfixed_a(-0.0001153796911239624)),(to_sfixed_a(-6.362760905176401e-05)),(to_sfixed_a(0.0004161513352300972)),(to_sfixed_a(5.365567631088197e-06)),(to_sfixed_a(2.730610140133649e-05)),(to_sfixed_a(3.840997669612989e-05)),(to_sfixed_a(-0.00021974592527840286)),(to_sfixed_a(-6.193957960931584e-05)),(to_sfixed_a(0.00028836337151005864)),(to_sfixed_a(-1.7069527530111372e-05)),(to_sfixed_a(-3.5336754081072286e-05)),(to_sfixed_a(-0.00018440319399815053)),(to_sfixed_a(4.11831570090726e-05)),(to_sfixed_a(-0.00018559416639618576)),(to_sfixed_a(-3.416000981815159e-05)),(to_sfixed_a(3.730606840690598e-05)),(to_sfixed_a(-3.921132883988321e-05)),(to_sfixed_a(1.7614154785405844e-05)),(to_sfixed_a(0.00019896100275218487)),(to_sfixed_a(-7.159925735322759e-05)),(to_sfixed_a(-0.0002230927930213511)),(to_sfixed_a(5.640977178700268e-07)),(to_sfixed_a(-0.0001334675180260092)),(to_sfixed_a(-2.980972931254655e-05)),(to_sfixed_a(0.00024154788115993142)),(to_sfixed_a(-4.64366894448176e-06)),(to_sfixed_a(1.215009979205206e-05)),(to_sfixed_a(9.795991354621947e-05)),(to_sfixed_a(5.689087265636772e-05)),(to_sfixed_a(-9.466832125326619e-05)),(to_sfixed_a(-1.3721379218623042e-05)),(to_sfixed_a(0.00021818104141857475)),(to_sfixed_a(-2.2351490770233795e-05)),(to_sfixed_a(-6.488793587777764e-06)),(to_sfixed_a(4.189911123830825e-05)),(to_sfixed_a(1.6842976037878543e-05)));

    constant weight_n2_5 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.700954020023346)),(to_sfixed_a(-0.6477277278900146)),(to_sfixed_a(-0.25253212451934814)),(to_sfixed_a(-8.731603156775236e-05)),(to_sfixed_a(-0.0043187313713133335)),(to_sfixed_a(-4.611094482243061e-06)),(to_sfixed_a(-0.005776464007794857)),(to_sfixed_a(-6.37936609564349e-05)),(to_sfixed_a(8.853364852257073e-05)),(to_sfixed_a(-8.366370457224548e-05)),(to_sfixed_a(-1.1678079317789525e-05)),(to_sfixed_a(-0.0033364277333021164)),(to_sfixed_a(-0.008530442602932453)),(to_sfixed_a(0.47187188267707825)),(to_sfixed_a(-1.846016130002681e-05)),(to_sfixed_a(-0.0001817064912756905)),(to_sfixed_a(-0.007165838964283466)),(to_sfixed_a(-2.203495205321815e-05)),(to_sfixed_a(-0.0033731055445969105)),(to_sfixed_a(0.004975240211933851)),(to_sfixed_a(-2.3533957573818043e-05)),(to_sfixed_a(0.00021595493308268487)),(to_sfixed_a(-0.005266883876174688)),(to_sfixed_a(0.0036569724325090647)),(to_sfixed_a(-0.0012658395571634173)),(to_sfixed_a(-1.9424998754402623e-05)),(to_sfixed_a(-0.00023220588627737015)),(to_sfixed_a(-0.00045418826630339026)),(to_sfixed_a(0.00028539536288008094)),(to_sfixed_a(6.302106339717284e-05)),(to_sfixed_a(-0.0060454318299889565)),(to_sfixed_a(0.00013784246402792633)),(to_sfixed_a(0.2744829058647156)),(to_sfixed_a(-0.00019326535402797163)),(to_sfixed_a(-0.00011288975656498224)),(to_sfixed_a(0.0002038082602666691)),(to_sfixed_a(0.05086689814925194)),(to_sfixed_a(0.0004936995101161301)),(to_sfixed_a(-0.0010340814478695393)),(to_sfixed_a(-2.33794235100504e-05)),(to_sfixed_a(0.05720444768667221)),(to_sfixed_a(0.0026771575212478638)),(to_sfixed_a(-1.1269512469880283e-05)),(to_sfixed_a(-8.095172233879566e-06)),(to_sfixed_a(-0.012703870423138142)),(to_sfixed_a(-0.022060785442590714)),(to_sfixed_a(-0.6001166105270386)),(to_sfixed_a(-0.004691419191658497)),(to_sfixed_a(0.00019991231965832412)),(to_sfixed_a(-0.005109334830194712)),(to_sfixed_a(-0.021912308409810066)),(to_sfixed_a(-0.0005589653155766428)),(to_sfixed_a(-2.217545988969505e-05)),(to_sfixed_a(0.0005417696665972471)),(to_sfixed_a(-0.010545008815824986)),(to_sfixed_a(-0.004896146710962057)),(to_sfixed_a(0.00044674810487776995)),(to_sfixed_a(-0.0077691879123449326)),(to_sfixed_a(0.0001880114432424307)),(to_sfixed_a(-0.00017479804228059947)),(to_sfixed_a(-0.0020310510881245136)),(to_sfixed_a(-0.00926925428211689)),(to_sfixed_a(0.00028928762185387313)),(to_sfixed_a(-0.013571728020906448)),(to_sfixed_a(0.00012171184062026441)),(to_sfixed_a(-0.004897357430309057)),(to_sfixed_a(-1.9098923075944185e-05)),(to_sfixed_a(0.002742570359259844)),(to_sfixed_a(-7.796719000907615e-05)),(to_sfixed_a(0.00018214505689684302)),(to_sfixed_a(0.2542944848537445)),(to_sfixed_a(-0.0005763749359175563)),(to_sfixed_a(0.3645573556423187)),(to_sfixed_a(0.00017466655117459595)),(to_sfixed_a(-4.339090082794428e-06)),(to_sfixed_a(3.182672298862599e-05)),(to_sfixed_a(-0.006642149295657873)),(to_sfixed_a(-0.0008664547931402922)),(to_sfixed_a(2.9183538572397083e-05)),(to_sfixed_a(-0.36927375197410583)),(to_sfixed_a(-0.013223210349678993)),(to_sfixed_a(3.3076503314077854e-06)),(to_sfixed_a(-0.3563694655895233)),(to_sfixed_a(0.31050053238868713)),(to_sfixed_a(-7.805726636433974e-05)),(to_sfixed_a(-0.005308516789227724)),(to_sfixed_a(-0.0016095878090709448)),(to_sfixed_a(-0.0008789516286924481)),(to_sfixed_a(-1.499722566222772e-05)),(to_sfixed_a(0.00015601166523993015)),(to_sfixed_a(0.058729879558086395)),(to_sfixed_a(7.890582492109388e-05)),(to_sfixed_a(-0.009743627160787582)),(to_sfixed_a(2.312719152541831e-05)),(to_sfixed_a(0.0038892123848199844)),(to_sfixed_a(8.34367165225558e-05)),(to_sfixed_a(6.123566708993167e-05)),(to_sfixed_a(2.3724878701614216e-05)),(to_sfixed_a(0.00011272229312453419)),(to_sfixed_a(-0.00019648642046377063)),(to_sfixed_a(-0.0007512305164709687)),(to_sfixed_a(-0.005976264365017414)),(to_sfixed_a(-1.2444928870536387e-05)),(to_sfixed_a(-0.008306861855089664)),(to_sfixed_a(0.20632627606391907)),(to_sfixed_a(-0.0034442904870957136)),(to_sfixed_a(-0.0003816395183093846)),(to_sfixed_a(-5.8774810895556584e-05)),(to_sfixed_a(0.00018091774836648256)),(to_sfixed_a(-0.00769005948677659)),(to_sfixed_a(0.0012698880163952708)),(to_sfixed_a(7.087415724527091e-05)),(to_sfixed_a(0.00017605014727450907)),(to_sfixed_a(0.0002161342417821288)),(to_sfixed_a(2.2739310225006193e-05)),(to_sfixed_a(0.0011278139427304268)),(to_sfixed_a(0.00347122666426003)),(to_sfixed_a(-0.0020684716291725636)),(to_sfixed_a(1.8980950699187815e-05)),(to_sfixed_a(0.0008636231650598347)),(to_sfixed_a(-5.0365979404887185e-05)),(to_sfixed_a(0.00011391715088393539)),(to_sfixed_a(-0.0051992726512253284)),(to_sfixed_a(-0.0002514274965506047)),(to_sfixed_a(-6.121417391113937e-05)),(to_sfixed_a(-0.003969674464315176)),(to_sfixed_a(-0.00025235736393369734)),(to_sfixed_a(7.820306200301275e-05)),(to_sfixed_a(-2.5031506083905697e-05)),(to_sfixed_a(4.096531483810395e-06)),(to_sfixed_a(0.0003766969603020698)),(to_sfixed_a(-0.00020405159739311785)),(to_sfixed_a(-0.00031002829200588167)),(to_sfixed_a(0.2833787798881531)),(to_sfixed_a(-1.0454623406985775e-06)),(to_sfixed_a(-0.00024717889027670026)),(to_sfixed_a(-0.04704274237155914)),(to_sfixed_a(-0.0012163070496171713)),(to_sfixed_a(-1.5023972082417458e-05)),(to_sfixed_a(0.00017971289344131947)),(to_sfixed_a(-0.0016583655960857868)),(to_sfixed_a(-0.00013598120131064206)),(to_sfixed_a(-0.00010127616405952722)),(to_sfixed_a(-2.5640285457484424e-05)),(to_sfixed_a(-0.23676061630249023)),(to_sfixed_a(-1.9781000446528196e-05)),(to_sfixed_a(-0.002058093436062336)),(to_sfixed_a(0.00017085784929804504)),(to_sfixed_a(-7.170972821768373e-06)),(to_sfixed_a(0.0020301886834204197)),(to_sfixed_a(8.552378858439624e-05)),(to_sfixed_a(9.347969898954034e-05)),(to_sfixed_a(0.004462988581508398)),(to_sfixed_a(6.4317267970182e-05)),(to_sfixed_a(-4.5053402573103085e-05)),(to_sfixed_a(-0.001352975727058947)),(to_sfixed_a(0.0001157131337095052)),(to_sfixed_a(-0.006638485938310623)),(to_sfixed_a(-0.0001201057675643824)),(to_sfixed_a(-9.77824383880943e-05)),(to_sfixed_a(-7.721601286903024e-05)),(to_sfixed_a(1.558651274535805e-05)),(to_sfixed_a(-0.013214483857154846)),(to_sfixed_a(0.0005857159267179668)),(to_sfixed_a(0.004387448541820049)),(to_sfixed_a(-0.0047773863188922405)),(to_sfixed_a(-2.1184259821893647e-05)),(to_sfixed_a(0.002888783812522888)),(to_sfixed_a(-3.0211074772523716e-05)),(to_sfixed_a(-0.00011411697050789371)),(to_sfixed_a(0.0012235401663929224)),(to_sfixed_a(0.0877097025513649)),(to_sfixed_a(-0.0029870900325477123)),(to_sfixed_a(0.00012812355998903513)),(to_sfixed_a(-0.4065960943698883)),(to_sfixed_a(-2.2457545128418133e-05)),(to_sfixed_a(-0.5293416380882263)),(to_sfixed_a(-0.002121871104463935)),(to_sfixed_a(0.3342016935348511)),(to_sfixed_a(0.0018279997166246176)),(to_sfixed_a(0.205741286277771)),(to_sfixed_a(-0.0009667804697528481)),(to_sfixed_a(0.00010398278391221538)),(to_sfixed_a(-1.2267024430911988e-05)),(to_sfixed_a(-8.992335642687976e-05)),(to_sfixed_a(0.1441502571105957)),(to_sfixed_a(-0.020471742376685143)),(to_sfixed_a(0.0013354696566239)),(to_sfixed_a(0.0039354185573756695)),(to_sfixed_a(0.009615691378712654)),(to_sfixed_a(0.012826049700379372)),(to_sfixed_a(0.00019090827845502645)),(to_sfixed_a(-0.0003457023703958839)),(to_sfixed_a(-0.008652135729789734)),(to_sfixed_a(8.003562834346667e-05)),(to_sfixed_a(-0.007229460868984461)),(to_sfixed_a(-8.554878877475858e-05)),(to_sfixed_a(-0.0031348150223493576)),(to_sfixed_a(-0.4381624460220337)),(to_sfixed_a(0.0002519504923839122)),(to_sfixed_a(5.9082707593915984e-05)),(to_sfixed_a(-0.00011629838991211727)),(to_sfixed_a(-3.572707646526396e-05)),(to_sfixed_a(3.134644794045016e-05)),(to_sfixed_a(-0.00027432868955656886)),(to_sfixed_a(0.003810875816270709)),(to_sfixed_a(-0.3902503550052643)),(to_sfixed_a(0.004171999171376228)),(to_sfixed_a(-0.0031028054654598236)),(to_sfixed_a(-0.15224596858024597)),(to_sfixed_a(0.004784678108990192)),(to_sfixed_a(5.161428271094337e-05)),(to_sfixed_a(7.387364166788757e-05)),(to_sfixed_a(-0.00022569907014258206)),(to_sfixed_a(-0.0001944322430063039)),(to_sfixed_a(-6.735860370099545e-05)),(to_sfixed_a(0.0017572480719536543)),(to_sfixed_a(-0.0017425977857783437)),(to_sfixed_a(0.00500792171806097)),(to_sfixed_a(3.862675293930806e-05)),(to_sfixed_a(9.827414032770321e-05)),(to_sfixed_a(0.00015627781976945698)),(to_sfixed_a(7.090994040481746e-05)),(to_sfixed_a(-0.0013487943215295672)),(to_sfixed_a(-0.586677074432373)),(to_sfixed_a(-0.00014280213508754969)),(to_sfixed_a(0.00015355566574726254)),(to_sfixed_a(-0.00016286007303278893)),(to_sfixed_a(-0.1528584361076355)),(to_sfixed_a(-0.12940829992294312)),(to_sfixed_a(-5.836141644977033e-05)),(to_sfixed_a(1.140782842412591e-05)),(to_sfixed_a(-0.00018701504450291395)),(to_sfixed_a(-0.00018144377099815756)),(to_sfixed_a(-0.002697853371500969)),(to_sfixed_a(0.00572947459295392)),(to_sfixed_a(-0.013258382678031921)),(to_sfixed_a(0.00015021814033389091)),(to_sfixed_a(0.0026333671994507313)),(to_sfixed_a(-0.00016026460798457265)),(to_sfixed_a(0.0013503477675840259)),(to_sfixed_a(-1.5564168279524893e-05)),(to_sfixed_a(-0.0013151869643479586)),(to_sfixed_a(-8.788974082563072e-05)),(to_sfixed_a(-0.2706072926521301)),(to_sfixed_a(-0.3259141445159912)),(to_sfixed_a(-0.011061154305934906)),(to_sfixed_a(-0.3744824230670929)),(to_sfixed_a(-0.00022678848472423851)),(to_sfixed_a(-0.008983529172837734)),(to_sfixed_a(-0.011688588187098503)),(to_sfixed_a(-6.669870344921947e-08)),(to_sfixed_a(-0.0023673190735280514)),(to_sfixed_a(-0.00015078589785844088)),(to_sfixed_a(-0.00034708098974078894)),(to_sfixed_a(-0.10606450587511063)),(to_sfixed_a(0.010782398283481598)),(to_sfixed_a(7.240484410431236e-05)),(to_sfixed_a(-6.603699875995517e-05)),(to_sfixed_a(0.00043634235044009984)),(to_sfixed_a(2.2514010197483003e-05)),(to_sfixed_a(0.0010085366666316986)),(to_sfixed_a(-0.0001596693036844954)),(to_sfixed_a(0.00020214369578752667)),(to_sfixed_a(9.397872054250911e-05)),(to_sfixed_a(-0.010903057642281055)),(to_sfixed_a(0.0001331998937530443)),(to_sfixed_a(-5.8499186707194895e-05)),(to_sfixed_a(0.00011370475112926215)),(to_sfixed_a(0.27260327339172363)),(to_sfixed_a(0.11536074429750443)),(to_sfixed_a(-0.0001836737064877525)),(to_sfixed_a(-0.00022238836390897632)),(to_sfixed_a(-0.000168848957400769)),(to_sfixed_a(-3.3540898584760725e-05)),(to_sfixed_a(3.0062143196118996e-05)),(to_sfixed_a(-0.0036703599616885185)),(to_sfixed_a(-0.004110449925065041)),(to_sfixed_a(-0.030884843319654465)),(to_sfixed_a(0.00041839730693027377)),(to_sfixed_a(-0.00015004882880020887)),(to_sfixed_a(-0.00032314975396730006)),(to_sfixed_a(-0.0001527456915937364)),(to_sfixed_a(0.006635336205363274)),(to_sfixed_a(0.00015492131933569908)),(to_sfixed_a(0.00011486388393677771)),(to_sfixed_a(0.007098870817571878)),(to_sfixed_a(-0.0023716643918305635)),(to_sfixed_a(-3.128854586975649e-05)),(to_sfixed_a(-0.5418061017990112)),(to_sfixed_a(0.0002148549392586574)),(to_sfixed_a(-0.009875073097646236)),(to_sfixed_a(0.007134686689823866)),(to_sfixed_a(0.00013492688594851643)),(to_sfixed_a(-0.0005696553853340447)),(to_sfixed_a(-0.0027816486544907093)),(to_sfixed_a(-0.02389814518392086)),(to_sfixed_a(-6.711929745506495e-05)),(to_sfixed_a(0.17592626810073853)),(to_sfixed_a(0.009233646094799042)),(to_sfixed_a(-0.01634218357503414)));

    constant weight_n2_6 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.26528412103652954)),(to_sfixed_a(0.0014265391509979963)),(to_sfixed_a(0.002606589812785387)),(to_sfixed_a(7.445782830473036e-05)),(to_sfixed_a(0.24364909529685974)),(to_sfixed_a(0.0001182802880066447)),(to_sfixed_a(0.3479289710521698)),(to_sfixed_a(-0.00031785893952474)),(to_sfixed_a(-0.00010588712757453322)),(to_sfixed_a(-8.413182513322681e-05)),(to_sfixed_a(-0.00012906687334179878)),(to_sfixed_a(0.0004308058996684849)),(to_sfixed_a(0.0020606531761586666)),(to_sfixed_a(0.0038607793394476175)),(to_sfixed_a(-9.774496720638126e-05)),(to_sfixed_a(-2.5554872991051525e-05)),(to_sfixed_a(0.00013643589045386761)),(to_sfixed_a(2.4042019504122436e-05)),(to_sfixed_a(0.20477096736431122)),(to_sfixed_a(0.00037406524643301964)),(to_sfixed_a(-0.0003021068114321679)),(to_sfixed_a(0.00027632975252345204)),(to_sfixed_a(-0.002954831812530756)),(to_sfixed_a(-0.0028769795317202806)),(to_sfixed_a(-0.0007308869971893728)),(to_sfixed_a(-0.0013273765798658133)),(to_sfixed_a(-0.00016759807476773858)),(to_sfixed_a(0.00045314340968616307)),(to_sfixed_a(-0.0005141554865986109)),(to_sfixed_a(-0.0001994503109017387)),(to_sfixed_a(0.07282678037881851)),(to_sfixed_a(0.00031907224911265075)),(to_sfixed_a(-0.00994816329330206)),(to_sfixed_a(-7.274359813891351e-05)),(to_sfixed_a(4.3005853513022885e-05)),(to_sfixed_a(-6.846436008345336e-05)),(to_sfixed_a(-0.004365262575447559)),(to_sfixed_a(-0.19301259517669678)),(to_sfixed_a(-0.0001528681314084679)),(to_sfixed_a(-0.00023765896912664175)),(to_sfixed_a(-0.011005240492522717)),(to_sfixed_a(0.0028217583894729614)),(to_sfixed_a(0.00016020177281461656)),(to_sfixed_a(-0.00011543277651071548)),(to_sfixed_a(-0.01099495030939579)),(to_sfixed_a(-0.009300275705754757)),(to_sfixed_a(0.0032487413845956326)),(to_sfixed_a(-0.011371574364602566)),(to_sfixed_a(-0.0002971880603581667)),(to_sfixed_a(-0.003625885583460331)),(to_sfixed_a(-0.0003032323147635907)),(to_sfixed_a(-5.6172386393882334e-05)),(to_sfixed_a(7.12992186890915e-05)),(to_sfixed_a(0.0020570072811096907)),(to_sfixed_a(-0.021855734288692474)),(to_sfixed_a(0.003378975670784712)),(to_sfixed_a(0.0001333160325884819)),(to_sfixed_a(0.029692750424146652)),(to_sfixed_a(9.981760740629397e-06)),(to_sfixed_a(-6.087042856961489e-05)),(to_sfixed_a(-0.006505315657705069)),(to_sfixed_a(-0.005963814910501242)),(to_sfixed_a(0.0004977361531928182)),(to_sfixed_a(-0.006422140635550022)),(to_sfixed_a(0.0003083771443925798)),(to_sfixed_a(0.20679359138011932)),(to_sfixed_a(0.00016827418585307896)),(to_sfixed_a(0.002691263798624277)),(to_sfixed_a(0.0011335957096889615)),(to_sfixed_a(-1.7541577108204365e-05)),(to_sfixed_a(0.39621251821517944)),(to_sfixed_a(-0.0009289473528042436)),(to_sfixed_a(-0.010215901769697666)),(to_sfixed_a(-0.0004501432995311916)),(to_sfixed_a(0.00010226861923001707)),(to_sfixed_a(-0.000315461540594697)),(to_sfixed_a(-0.014994718134403229)),(to_sfixed_a(-0.011814611963927746)),(to_sfixed_a(-6.20353821432218e-05)),(to_sfixed_a(-0.5636654496192932)),(to_sfixed_a(-0.00897954124957323)),(to_sfixed_a(7.918386836536229e-05)),(to_sfixed_a(-0.0004341812455095351)),(to_sfixed_a(0.16928844153881073)),(to_sfixed_a(-5.984743620501831e-05)),(to_sfixed_a(-0.0014739230973646045)),(to_sfixed_a(0.005177181679755449)),(to_sfixed_a(0.005219887942075729)),(to_sfixed_a(-7.107558485586196e-05)),(to_sfixed_a(-7.030511915218085e-05)),(to_sfixed_a(0.0006950952229090035)),(to_sfixed_a(-0.0001486516703153029)),(to_sfixed_a(-0.00020638984278775752)),(to_sfixed_a(-3.6476489185588434e-05)),(to_sfixed_a(0.004912494216114283)),(to_sfixed_a(-0.00019827979849651456)),(to_sfixed_a(0.00013532652519643307)),(to_sfixed_a(-0.0001158832892542705)),(to_sfixed_a(-3.9434657082892954e-05)),(to_sfixed_a(-0.0001544599508633837)),(to_sfixed_a(-0.008361770771443844)),(to_sfixed_a(-0.008737833239138126)),(to_sfixed_a(0.00011049819295294583)),(to_sfixed_a(-0.265403687953949)),(to_sfixed_a(-0.007214811630547047)),(to_sfixed_a(-0.009256280027329922)),(to_sfixed_a(1.6362173482775688e-07)),(to_sfixed_a(6.915187259437516e-05)),(to_sfixed_a(0.0002693244314286858)),(to_sfixed_a(-0.007874496281147003)),(to_sfixed_a(-0.0007767790229991078)),(to_sfixed_a(2.864454290829599e-05)),(to_sfixed_a(0.0002347485424252227)),(to_sfixed_a(-4.902247746940702e-05)),(to_sfixed_a(1.6235302609857172e-05)),(to_sfixed_a(0.2193213552236557)),(to_sfixed_a(-0.0034475703723728657)),(to_sfixed_a(-0.006133331451565027)),(to_sfixed_a(-9.902614692691714e-05)),(to_sfixed_a(0.0009389068582095206)),(to_sfixed_a(0.0002825075061991811)),(to_sfixed_a(-7.095769251463935e-05)),(to_sfixed_a(0.0008491366170346737)),(to_sfixed_a(-6.170316191855818e-05)),(to_sfixed_a(0.00029041600646451116)),(to_sfixed_a(-0.001344442367553711)),(to_sfixed_a(0.004649010952562094)),(to_sfixed_a(-1.457634789403528e-05)),(to_sfixed_a(-5.611769302049652e-05)),(to_sfixed_a(0.00015222970978356898)),(to_sfixed_a(4.987952706869692e-06)),(to_sfixed_a(-5.603214958682656e-06)),(to_sfixed_a(-0.00012548510858323425)),(to_sfixed_a(0.12140340358018875)),(to_sfixed_a(3.2107127481140196e-06)),(to_sfixed_a(-4.02333025704138e-05)),(to_sfixed_a(-0.001411468256264925)),(to_sfixed_a(-0.33164528012275696)),(to_sfixed_a(0.00024042368750087917)),(to_sfixed_a(-0.00011051780165871605)),(to_sfixed_a(0.005643330514431)),(to_sfixed_a(-9.698295616544783e-05)),(to_sfixed_a(0.00016552193847019225)),(to_sfixed_a(0.0003340370603837073)),(to_sfixed_a(0.21633251011371613)),(to_sfixed_a(0.0007269278867170215)),(to_sfixed_a(0.0008854061597958207)),(to_sfixed_a(0.00044797544251196086)),(to_sfixed_a(-7.003647624514997e-05)),(to_sfixed_a(0.0024894673842936754)),(to_sfixed_a(-1.941218761203345e-05)),(to_sfixed_a(-9.877415868686512e-05)),(to_sfixed_a(0.009645630605518818)),(to_sfixed_a(-8.576331310905516e-06)),(to_sfixed_a(3.892877430189401e-05)),(to_sfixed_a(-0.004191793035715818)),(to_sfixed_a(6.659291102550924e-05)),(to_sfixed_a(0.003305060788989067)),(to_sfixed_a(7.474372978322208e-05)),(to_sfixed_a(0.0001368807425023988)),(to_sfixed_a(-7.037125760689378e-05)),(to_sfixed_a(2.910957846324891e-06)),(to_sfixed_a(-0.0012087933719158173)),(to_sfixed_a(0.000572235556319356)),(to_sfixed_a(-0.001245353021658957)),(to_sfixed_a(0.0006325097638182342)),(to_sfixed_a(-0.0002836017229128629)),(to_sfixed_a(0.0013551705051213503)),(to_sfixed_a(-6.140695768408477e-05)),(to_sfixed_a(-0.00015986693324521184)),(to_sfixed_a(-0.29685649275779724)),(to_sfixed_a(0.0003167958930134773)),(to_sfixed_a(0.0020505802240222692)),(to_sfixed_a(7.254909723997116e-05)),(to_sfixed_a(-0.4699210822582245)),(to_sfixed_a(0.002867873990908265)),(to_sfixed_a(-0.026015231385827065)),(to_sfixed_a(-0.1415480524301529)),(to_sfixed_a(0.0037555929739028215)),(to_sfixed_a(-0.0056982035748660564)),(to_sfixed_a(-0.00038075121119618416)),(to_sfixed_a(0.0020147927571088076)),(to_sfixed_a(-0.00011684911441989243)),(to_sfixed_a(-0.00018256397743243724)),(to_sfixed_a(-4.7138018999248743e-07)),(to_sfixed_a(-0.0213484987616539)),(to_sfixed_a(0.004081740975379944)),(to_sfixed_a(0.0025690440088510513)),(to_sfixed_a(0.002422104123979807)),(to_sfixed_a(0.009102145209908485)),(to_sfixed_a(0.002638117875903845)),(to_sfixed_a(-0.0002884298446588218)),(to_sfixed_a(-0.019669130444526672)),(to_sfixed_a(-0.000939980847761035)),(to_sfixed_a(-4.3284191633574665e-05)),(to_sfixed_a(-0.009362920187413692)),(to_sfixed_a(-5.990015051793307e-05)),(to_sfixed_a(0.17157483100891113)),(to_sfixed_a(-0.3397224545478821)),(to_sfixed_a(-0.0001173438795376569)),(to_sfixed_a(9.871826478047296e-05)),(to_sfixed_a(0.00031600543297827244)),(to_sfixed_a(0.00016981427324935794)),(to_sfixed_a(0.00020407570991665125)),(to_sfixed_a(3.784777072723955e-05)),(to_sfixed_a(0.006806597579270601)),(to_sfixed_a(0.001293464214541018)),(to_sfixed_a(-0.006737754214555025)),(to_sfixed_a(0.0009659967618063092)),(to_sfixed_a(-0.19960737228393555)),(to_sfixed_a(0.004738093353807926)),(to_sfixed_a(-0.00023872285964898765)),(to_sfixed_a(0.0001470318966312334)),(to_sfixed_a(5.034380592405796e-06)),(to_sfixed_a(0.00011477078078314662)),(to_sfixed_a(-0.0001788583176676184)),(to_sfixed_a(0.01310998946428299)),(to_sfixed_a(0.00024773430777713656)),(to_sfixed_a(0.01891469396650791)),(to_sfixed_a(0.00011191458179382607)),(to_sfixed_a(-0.00013017850869800895)),(to_sfixed_a(-8.426416025031358e-05)),(to_sfixed_a(-0.00012078622239641845)),(to_sfixed_a(0.004369175061583519)),(to_sfixed_a(0.24968497455120087)),(to_sfixed_a(-4.5132161176297814e-05)),(to_sfixed_a(1.0179537639487535e-06)),(to_sfixed_a(1.2427804904291406e-05)),(to_sfixed_a(-0.0029965618159621954)),(to_sfixed_a(-0.003609391860663891)),(to_sfixed_a(0.30761855840682983)),(to_sfixed_a(0.0001622092822799459)),(to_sfixed_a(-8.790145511738956e-05)),(to_sfixed_a(-8.212296233978122e-05)),(to_sfixed_a(-0.0052141472697257996)),(to_sfixed_a(-0.010094915516674519)),(to_sfixed_a(-0.0012302044779062271)),(to_sfixed_a(-8.451072062598541e-05)),(to_sfixed_a(0.0028561302460730076)),(to_sfixed_a(-1.5521509340032935e-05)),(to_sfixed_a(0.002003098139539361)),(to_sfixed_a(0.00029478195938281715)),(to_sfixed_a(-0.44342663884162903)),(to_sfixed_a(-0.00023646051704417914)),(to_sfixed_a(-0.182326078414917)),(to_sfixed_a(-0.12958712875843048)),(to_sfixed_a(-0.00882173515856266)),(to_sfixed_a(-0.4897874593734741)),(to_sfixed_a(-0.00016848492668941617)),(to_sfixed_a(-0.008296843618154526)),(to_sfixed_a(0.2636699378490448)),(to_sfixed_a(0.00011597694538068026)),(to_sfixed_a(0.0014709413517266512)),(to_sfixed_a(0.00011364345846232027)),(to_sfixed_a(-0.00047351577086374164)),(to_sfixed_a(-0.0025801830925047398)),(to_sfixed_a(-0.5581392645835876)),(to_sfixed_a(-0.00029366122907958925)),(to_sfixed_a(-2.3600503482157364e-05)),(to_sfixed_a(-0.0017286977963522077)),(to_sfixed_a(2.407978172414005e-06)),(to_sfixed_a(1.5804340364411473e-05)),(to_sfixed_a(2.7196714654564857e-05)),(to_sfixed_a(-0.0004207080928608775)),(to_sfixed_a(-0.00010197124356636778)),(to_sfixed_a(-0.014681131578981876)),(to_sfixed_a(-9.836933895712718e-05)),(to_sfixed_a(2.178657814511098e-05)),(to_sfixed_a(1.8871360225602984e-05)),(to_sfixed_a(0.3612056076526642)),(to_sfixed_a(0.3126886188983917)),(to_sfixed_a(6.0713304264936596e-05)),(to_sfixed_a(0.0002523849834688008)),(to_sfixed_a(8.611082739662379e-05)),(to_sfixed_a(-2.8426729841157794e-06)),(to_sfixed_a(0.003764854511246085)),(to_sfixed_a(-0.004780816379934549)),(to_sfixed_a(-0.003662492148578167)),(to_sfixed_a(0.29845306277275085)),(to_sfixed_a(0.004131993744522333)),(to_sfixed_a(-0.00023797503672540188)),(to_sfixed_a(-0.0001576106733409688)),(to_sfixed_a(-5.009886444895528e-05)),(to_sfixed_a(-0.0007906057871878147)),(to_sfixed_a(5.858535587321967e-06)),(to_sfixed_a(0.0001481141080148518)),(to_sfixed_a(0.0022471975535154343)),(to_sfixed_a(0.20134490728378296)),(to_sfixed_a(-0.0002753533481154591)),(to_sfixed_a(0.0003101366455666721)),(to_sfixed_a(0.00037710031028836966)),(to_sfixed_a(-0.006549830082803965)),(to_sfixed_a(0.12935394048690796)),(to_sfixed_a(-2.5627803552197292e-05)),(to_sfixed_a(0.005019231699407101)),(to_sfixed_a(0.0020470088347792625)),(to_sfixed_a(-0.02570774033665657)),(to_sfixed_a(0.00011073026689700782)),(to_sfixed_a(-0.0036987094208598137)),(to_sfixed_a(0.009762370958924294)),(to_sfixed_a(-0.012978555634617805)));

    constant weight_n2_7 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.37494099140167236)),(to_sfixed_a(-0.0013854816788807511)),(to_sfixed_a(0.0015076019335538149)),(to_sfixed_a(0.0001321657036896795)),(to_sfixed_a(0.005800063721835613)),(to_sfixed_a(9.282575047109276e-05)),(to_sfixed_a(-0.008664250373840332)),(to_sfixed_a(4.965637708664872e-05)),(to_sfixed_a(-0.0002929912880063057)),(to_sfixed_a(-0.00041811494156718254)),(to_sfixed_a(5.917776434216648e-06)),(to_sfixed_a(-0.33173590898513794)),(to_sfixed_a(-0.0037969842087477446)),(to_sfixed_a(0.004098434001207352)),(to_sfixed_a(0.00010516795009607449)),(to_sfixed_a(-0.0002861304674297571)),(to_sfixed_a(-0.20432783663272858)),(to_sfixed_a(0.00014986497990321368)),(to_sfixed_a(-0.43244102597236633)),(to_sfixed_a(-0.0008784350357018411)),(to_sfixed_a(9.164144285023212e-05)),(to_sfixed_a(-3.72577051166445e-05)),(to_sfixed_a(-1.2545693607535213e-05)),(to_sfixed_a(-0.0046748011372983456)),(to_sfixed_a(-0.008202413097023964)),(to_sfixed_a(-0.34125515818595886)),(to_sfixed_a(-0.00013057823525741696)),(to_sfixed_a(-5.77559694647789e-05)),(to_sfixed_a(-0.0001465214736526832)),(to_sfixed_a(-9.080665040528402e-05)),(to_sfixed_a(-0.0022831421811133623)),(to_sfixed_a(-7.054384332150221e-05)),(to_sfixed_a(-0.006562685128301382)),(to_sfixed_a(8.503813296556473e-05)),(to_sfixed_a(-0.00022000136959832162)),(to_sfixed_a(-9.532097465125844e-05)),(to_sfixed_a(0.27953022718429565)),(to_sfixed_a(0.008276814594864845)),(to_sfixed_a(-0.0033779062796384096)),(to_sfixed_a(-1.7238380678463727e-06)),(to_sfixed_a(-0.001494887052103877)),(to_sfixed_a(0.0024509700015187263)),(to_sfixed_a(6.878076965222135e-05)),(to_sfixed_a(-4.651581548387185e-06)),(to_sfixed_a(-6.0350008425302804e-05)),(to_sfixed_a(0.3079454302787781)),(to_sfixed_a(-0.0003340825205668807)),(to_sfixed_a(-0.000657907803542912)),(to_sfixed_a(-9.126169607043266e-05)),(to_sfixed_a(-0.019824370741844177)),(to_sfixed_a(0.0001120478700613603)),(to_sfixed_a(0.0011504215653985739)),(to_sfixed_a(2.164051511499565e-05)),(to_sfixed_a(-0.00014798398478887975)),(to_sfixed_a(0.0010745920008048415)),(to_sfixed_a(-0.008446692489087582)),(to_sfixed_a(7.604320853715762e-05)),(to_sfixed_a(-0.009914983995258808)),(to_sfixed_a(-0.00016855962167028338)),(to_sfixed_a(6.32587616564706e-05)),(to_sfixed_a(-2.8711972845485434e-05)),(to_sfixed_a(0.002433893270790577)),(to_sfixed_a(9.00727536645718e-06)),(to_sfixed_a(-0.1365237683057785)),(to_sfixed_a(3.104133429587819e-05)),(to_sfixed_a(0.4108608365058899)),(to_sfixed_a(0.00025132534210570157)),(to_sfixed_a(-0.16941572725772858)),(to_sfixed_a(0.4414290189743042)),(to_sfixed_a(-2.538977059884928e-05)),(to_sfixed_a(0.15482540428638458)),(to_sfixed_a(-0.07674811035394669)),(to_sfixed_a(0.23395417630672455)),(to_sfixed_a(-3.725872375071049e-07)),(to_sfixed_a(-0.00016796511772554368)),(to_sfixed_a(0.0002789534046314657)),(to_sfixed_a(-0.029464654624462128)),(to_sfixed_a(-0.03304990008473396)),(to_sfixed_a(7.129653386073187e-05)),(to_sfixed_a(-0.20005974173545837)),(to_sfixed_a(0.0006216607289388776)),(to_sfixed_a(-9.468572534387931e-05)),(to_sfixed_a(-0.00028872699476778507)),(to_sfixed_a(0.43736156821250916)),(to_sfixed_a(0.00010616061626933515)),(to_sfixed_a(-0.005266993306577206)),(to_sfixed_a(-0.0014821043005213141)),(to_sfixed_a(-0.0009299051598645747)),(to_sfixed_a(-1.9234823412261903e-05)),(to_sfixed_a(4.662246647058055e-05)),(to_sfixed_a(-0.009202517569065094)),(to_sfixed_a(-0.0002911825431510806)),(to_sfixed_a(-0.0030578237492591143)),(to_sfixed_a(6.996742740739137e-05)),(to_sfixed_a(-0.009872139431536198)),(to_sfixed_a(-5.1182141760364175e-05)),(to_sfixed_a(-1.8837235984392464e-05)),(to_sfixed_a(0.000305001565720886)),(to_sfixed_a(3.5277189454063773e-06)),(to_sfixed_a(-0.00021811803162563592)),(to_sfixed_a(-0.022120194509625435)),(to_sfixed_a(-0.0019755028188228607)),(to_sfixed_a(0.00011926385923288763)),(to_sfixed_a(-0.21463078260421753)),(to_sfixed_a(0.25797733664512634)),(to_sfixed_a(-0.20692075788974762)),(to_sfixed_a(-0.00010017328168032691)),(to_sfixed_a(-3.800229751504958e-05)),(to_sfixed_a(-5.960100679658353e-08)),(to_sfixed_a(-0.0077036479488015175)),(to_sfixed_a(0.2201349139213562)),(to_sfixed_a(0.0001087540658772923)),(to_sfixed_a(-0.004114903509616852)),(to_sfixed_a(2.199807931901887e-05)),(to_sfixed_a(-6.952405965421349e-05)),(to_sfixed_a(-0.01121607981622219)),(to_sfixed_a(-0.0011163903400301933)),(to_sfixed_a(-0.010449678637087345)),(to_sfixed_a(0.0001425209775334224)),(to_sfixed_a(0.0003374338266439736)),(to_sfixed_a(3.042240859940648e-05)),(to_sfixed_a(-4.59989532828331e-05)),(to_sfixed_a(-0.0006113765994086862)),(to_sfixed_a(0.0001532544702058658)),(to_sfixed_a(1.2527394574135542e-05)),(to_sfixed_a(-0.46685710549354553)),(to_sfixed_a(-0.30836033821105957)),(to_sfixed_a(1.0563089745119214e-05)),(to_sfixed_a(-0.00015329662710428238)),(to_sfixed_a(-0.00012939280713908374)),(to_sfixed_a(-3.141622801194899e-05)),(to_sfixed_a(-5.791756484541111e-05)),(to_sfixed_a(-0.0003802456194534898)),(to_sfixed_a(0.01322912611067295)),(to_sfixed_a(0.00030535575933754444)),(to_sfixed_a(-7.778585859341547e-05)),(to_sfixed_a(-0.4315844476222992)),(to_sfixed_a(3.8821352063678205e-05)),(to_sfixed_a(-0.00010394143464509398)),(to_sfixed_a(6.27929694019258e-06)),(to_sfixed_a(0.0001598572125658393)),(to_sfixed_a(5.927881284151226e-05)),(to_sfixed_a(7.908446423243731e-05)),(to_sfixed_a(-0.0017821252113208175)),(to_sfixed_a(0.0003893183311447501)),(to_sfixed_a(8.83784523466602e-05)),(to_sfixed_a(0.0010511847212910652)),(to_sfixed_a(3.3367363357683644e-05)),(to_sfixed_a(-7.90720951044932e-05)),(to_sfixed_a(-0.017184458673000336)),(to_sfixed_a(-0.00013413617853075266)),(to_sfixed_a(4.20695505454205e-06)),(to_sfixed_a(0.00039349490543827415)),(to_sfixed_a(0.00014700222527608275)),(to_sfixed_a(4.174908099230379e-07)),(to_sfixed_a(-0.0007253959192894399)),(to_sfixed_a(-0.00029894683393649757)),(to_sfixed_a(0.16936691105365753)),(to_sfixed_a(-0.00013402361946646124)),(to_sfixed_a(3.917516733054072e-05)),(to_sfixed_a(0.00011321804049657658)),(to_sfixed_a(0.00012910942314192653)),(to_sfixed_a(-0.002458865288645029)),(to_sfixed_a(0.406732976436615)),(to_sfixed_a(-0.006193993147462606)),(to_sfixed_a(-0.4582895040512085)),(to_sfixed_a(0.00016954075545072556)),(to_sfixed_a(-0.006893766112625599)),(to_sfixed_a(-1.8035658285953104e-05)),(to_sfixed_a(0.00029409962007775903)),(to_sfixed_a(0.00023020146181806922)),(to_sfixed_a(-0.007036096416413784)),(to_sfixed_a(-1.4317425666376948e-05)),(to_sfixed_a(2.2568921849597245e-05)),(to_sfixed_a(0.010944902896881104)),(to_sfixed_a(0.00011680133320624009)),(to_sfixed_a(-0.3033207058906555)),(to_sfixed_a(-0.19033239781856537)),(to_sfixed_a(-0.005063421092927456)),(to_sfixed_a(0.0006538142333738506)),(to_sfixed_a(0.0007836225559003651)),(to_sfixed_a(0.012164684943854809)),(to_sfixed_a(-0.0001010111445793882)),(to_sfixed_a(0.00011365683167241514)),(to_sfixed_a(-6.131833652034402e-05)),(to_sfixed_a(-0.001306014135479927)),(to_sfixed_a(-0.3139943778514862)),(to_sfixed_a(-0.000669403001666069)),(to_sfixed_a(0.004054185003042221)),(to_sfixed_a(0.003939380403608084)),(to_sfixed_a(0.28238505125045776)),(to_sfixed_a(-9.962882177205756e-05)),(to_sfixed_a(-0.44919607043266296)),(to_sfixed_a(-0.00015618883480783552)),(to_sfixed_a(1.526341657154262e-05)),(to_sfixed_a(-0.00030542287277057767)),(to_sfixed_a(-0.0001825220388127491)),(to_sfixed_a(-0.006721279583871365)),(to_sfixed_a(0.0039009773172438145)),(to_sfixed_a(2.100565325235948e-05)),(to_sfixed_a(4.4237825932214037e-05)),(to_sfixed_a(-2.04566094907932e-05)),(to_sfixed_a(-3.4688637242652476e-06)),(to_sfixed_a(-0.00010541847586864606)),(to_sfixed_a(-3.6142198950983584e-05)),(to_sfixed_a(0.0013750821817666292)),(to_sfixed_a(0.018209436908364296)),(to_sfixed_a(0.42796826362609863)),(to_sfixed_a(0.35523557662963867)),(to_sfixed_a(0.2501193583011627)),(to_sfixed_a(0.22798483073711395)),(to_sfixed_a(-5.1856914069503546e-06)),(to_sfixed_a(8.002499089343473e-05)),(to_sfixed_a(2.857997787941713e-05)),(to_sfixed_a(0.0002875477075576782)),(to_sfixed_a(-0.00017512797785457224)),(to_sfixed_a(0.0014566672034561634)),(to_sfixed_a(0.005834379233419895)),(to_sfixed_a(0.24340850114822388)),(to_sfixed_a(-0.00029311139951460063)),(to_sfixed_a(0.00010531340376473963)),(to_sfixed_a(0.0001533980539534241)),(to_sfixed_a(6.803488940931857e-05)),(to_sfixed_a(-4.8073590733110905e-05)),(to_sfixed_a(0.0322091169655323)),(to_sfixed_a(7.089956488925964e-05)),(to_sfixed_a(-6.762355769751593e-05)),(to_sfixed_a(0.00022470889962278306)),(to_sfixed_a(-0.3262193500995636)),(to_sfixed_a(0.28067007660865784)),(to_sfixed_a(0.12674809992313385)),(to_sfixed_a(0.00011340751370880753)),(to_sfixed_a(-3.745917638298124e-05)),(to_sfixed_a(-1.154860365204513e-05)),(to_sfixed_a(0.0010979034705087543)),(to_sfixed_a(-0.004462232813239098)),(to_sfixed_a(-0.001119227847084403)),(to_sfixed_a(2.1873711375519633e-07)),(to_sfixed_a(0.0026337753515690565)),(to_sfixed_a(0.00011514886864461005)),(to_sfixed_a(-0.5324495434761047)),(to_sfixed_a(-0.0001033646403811872)),(to_sfixed_a(-0.3374772369861603)),(to_sfixed_a(-0.00011738685861928388)),(to_sfixed_a(-0.49616706371307373)),(to_sfixed_a(0.30775564908981323)),(to_sfixed_a(-0.4893435537815094)),(to_sfixed_a(0.33309465646743774)),(to_sfixed_a(3.92971487599425e-05)),(to_sfixed_a(-0.17172040045261383)),(to_sfixed_a(-0.013285069726407528)),(to_sfixed_a(0.00013026950182393193)),(to_sfixed_a(0.0016811762470752)),(to_sfixed_a(-0.00010417841258458793)),(to_sfixed_a(-5.9334339312044904e-05)),(to_sfixed_a(-0.5243262648582458)),(to_sfixed_a(-0.002537125488743186)),(to_sfixed_a(-0.00018935555999632925)),(to_sfixed_a(5.991200669086538e-05)),(to_sfixed_a(-0.4100492596626282)),(to_sfixed_a(-5.809332651551813e-05)),(to_sfixed_a(0.0010282306466251612)),(to_sfixed_a(-2.970072819152847e-05)),(to_sfixed_a(0.00013452455459628254)),(to_sfixed_a(0.00025014003040269017)),(to_sfixed_a(-0.010990959592163563)),(to_sfixed_a(-6.433451926568523e-05)),(to_sfixed_a(-2.3392349248752e-06)),(to_sfixed_a(-0.0002858319494407624)),(to_sfixed_a(-0.0014495367649942636)),(to_sfixed_a(0.16664086282253265)),(to_sfixed_a(-5.1146253099432215e-05)),(to_sfixed_a(0.00020516121003311127)),(to_sfixed_a(-0.0001166299989563413)),(to_sfixed_a(-0.0002911769552156329)),(to_sfixed_a(-0.2177581787109375)),(to_sfixed_a(-0.005683331284672022)),(to_sfixed_a(-0.36474940180778503)),(to_sfixed_a(0.330745667219162)),(to_sfixed_a(0.1375337839126587)),(to_sfixed_a(6.765182479284704e-05)),(to_sfixed_a(0.0001542253594379872)),(to_sfixed_a(-6.944670167285949e-05)),(to_sfixed_a(-0.0049766129814088345)),(to_sfixed_a(-2.2920226911082864e-05)),(to_sfixed_a(0.0002479887625668198)),(to_sfixed_a(0.29687851667404175)),(to_sfixed_a(-0.0074127777479588985)),(to_sfixed_a(-7.523926615249366e-05)),(to_sfixed_a(4.947206616634503e-05)),(to_sfixed_a(-8.31665238365531e-05)),(to_sfixed_a(-0.004897122737020254)),(to_sfixed_a(0.0029126908630132675)),(to_sfixed_a(5.7399389334023e-05)),(to_sfixed_a(0.020524177700281143)),(to_sfixed_a(-0.2522197961807251)),(to_sfixed_a(-0.0005044634453952312)),(to_sfixed_a(-1.6839949239511043e-06)),(to_sfixed_a(-0.015693994238972664)),(to_sfixed_a(0.17031888663768768)),(to_sfixed_a(-0.004947397857904434)));

    constant weight_n2_8 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.023265564814209938)),(to_sfixed_a(0.0001370518293697387)),(to_sfixed_a(0.00015176780289039016)),(to_sfixed_a(-4.127994543523528e-06)),(to_sfixed_a(6.151638081064448e-05)),(to_sfixed_a(-0.0001669223274802789)),(to_sfixed_a(-0.00011311916750855744)),(to_sfixed_a(-0.0001168950111605227)),(to_sfixed_a(8.686819637659937e-05)),(to_sfixed_a(0.0001036181056406349)),(to_sfixed_a(-7.02120378264226e-05)),(to_sfixed_a(5.8567871747072786e-05)),(to_sfixed_a(-0.00011714365246007219)),(to_sfixed_a(-0.0003153442812617868)),(to_sfixed_a(4.86847129650414e-05)),(to_sfixed_a(2.0210398361086845e-05)),(to_sfixed_a(-0.00011251531395828351)),(to_sfixed_a(-0.00011421395174693316)),(to_sfixed_a(7.583963451907039e-06)),(to_sfixed_a(-0.00011702286428771913)),(to_sfixed_a(-3.784471482504159e-05)),(to_sfixed_a(-5.7651399401947856e-05)),(to_sfixed_a(-0.00011639873991953209)),(to_sfixed_a(4.2698167817434296e-05)),(to_sfixed_a(0.00010119019134435803)),(to_sfixed_a(-0.00011516486847540364)),(to_sfixed_a(2.7869380573974922e-05)),(to_sfixed_a(-8.782297663856298e-05)),(to_sfixed_a(0.00015173139399848878)),(to_sfixed_a(7.167721923906356e-05)),(to_sfixed_a(-0.00023136823438107967)),(to_sfixed_a(-0.00018331222236156464)),(to_sfixed_a(0.00013475862215273082)),(to_sfixed_a(-1.2846030585933477e-06)),(to_sfixed_a(-0.00010100552754011005)),(to_sfixed_a(-0.00015307989087887108)),(to_sfixed_a(5.684866482624784e-05)),(to_sfixed_a(6.560001929756254e-05)),(to_sfixed_a(0.00012882851297035813)),(to_sfixed_a(-2.9648908821400255e-06)),(to_sfixed_a(0.00010904068039963022)),(to_sfixed_a(-0.0002897362282965332)),(to_sfixed_a(0.00023728390806354582)),(to_sfixed_a(-6.172176654217765e-05)),(to_sfixed_a(-4.4122134568169713e-07)),(to_sfixed_a(-1.0202329576713964e-06)),(to_sfixed_a(-5.898913514101878e-05)),(to_sfixed_a(-0.00019161871750839055)),(to_sfixed_a(0.00011300943151582032)),(to_sfixed_a(6.078337173676118e-05)),(to_sfixed_a(-0.00016045592201408)),(to_sfixed_a(-7.464286318281665e-05)),(to_sfixed_a(-8.91669187694788e-05)),(to_sfixed_a(-8.921934204408899e-05)),(to_sfixed_a(0.00019758609414566308)),(to_sfixed_a(-0.0002384334511589259)),(to_sfixed_a(-0.00011819173232652247)),(to_sfixed_a(5.784594395663589e-05)),(to_sfixed_a(-0.00014891276077833027)),(to_sfixed_a(-8.638237341074273e-05)),(to_sfixed_a(7.016136078163981e-05)),(to_sfixed_a(-0.00017298782768193632)),(to_sfixed_a(4.02222212869674e-05)),(to_sfixed_a(-2.7885937015525997e-05)),(to_sfixed_a(-0.0004556484054774046)),(to_sfixed_a(9.177446190733463e-05)),(to_sfixed_a(-0.00010351647506467998)),(to_sfixed_a(6.847965414635837e-05)),(to_sfixed_a(1.0525500329094939e-05)),(to_sfixed_a(1.2083648471161723e-05)),(to_sfixed_a(-0.0002963297883979976)),(to_sfixed_a(-0.00013655985821969807)),(to_sfixed_a(0.00011827794514829293)),(to_sfixed_a(-6.908446812303737e-05)),(to_sfixed_a(-1.891801366582513e-05)),(to_sfixed_a(0.0001829478715080768)),(to_sfixed_a(6.251218292163685e-05)),(to_sfixed_a(1.291270018555224e-05)),(to_sfixed_a(-0.0002382933598710224)),(to_sfixed_a(-9.017906268127263e-05)),(to_sfixed_a(0.00026998695102520287)),(to_sfixed_a(-8.26683608465828e-05)),(to_sfixed_a(-4.9740665417630225e-06)),(to_sfixed_a(0.00010412832489237189)),(to_sfixed_a(0.0002478639071341604)),(to_sfixed_a(-0.0003099558234680444)),(to_sfixed_a(-7.052897854009643e-05)),(to_sfixed_a(2.934060466941446e-05)),(to_sfixed_a(6.771666812710464e-05)),(to_sfixed_a(-0.00015171279665082693)),(to_sfixed_a(7.005780207691714e-05)),(to_sfixed_a(-7.617875235155225e-05)),(to_sfixed_a(-6.693194154649973e-05)),(to_sfixed_a(-8.894572965800762e-05)),(to_sfixed_a(3.201030631316826e-05)),(to_sfixed_a(-9.544252679916099e-05)),(to_sfixed_a(-6.844475865364075e-05)),(to_sfixed_a(0.00014567014295607805)),(to_sfixed_a(-6.03724765824154e-06)),(to_sfixed_a(0.00024969837977550924)),(to_sfixed_a(-0.00011664068006211892)),(to_sfixed_a(6.14194359513931e-05)),(to_sfixed_a(0.00015717768110334873)),(to_sfixed_a(-1.6117497580125928e-05)),(to_sfixed_a(-0.00013018969912081957)),(to_sfixed_a(0.00017567379109095782)),(to_sfixed_a(3.233029565308243e-05)),(to_sfixed_a(7.59615795686841e-06)),(to_sfixed_a(-0.00021672870207112283)),(to_sfixed_a(7.738322165096179e-05)),(to_sfixed_a(-0.00018972597899846733)),(to_sfixed_a(0.00025093700969591737)),(to_sfixed_a(4.338464350439608e-06)),(to_sfixed_a(-3.0289724236354232e-05)),(to_sfixed_a(0.00018215295858681202)),(to_sfixed_a(-0.00014843295502942055)),(to_sfixed_a(-0.0001813342678360641)),(to_sfixed_a(-0.0002144057652913034)),(to_sfixed_a(0.000300272717140615)),(to_sfixed_a(4.467509643291123e-05)),(to_sfixed_a(-0.00014030415331944823)),(to_sfixed_a(0.00014681200264021754)),(to_sfixed_a(-1.8847276805900037e-05)),(to_sfixed_a(0.00010154139454243705)),(to_sfixed_a(-0.00018166657537221909)),(to_sfixed_a(2.108923945343122e-05)),(to_sfixed_a(0.0002793139428831637)),(to_sfixed_a(7.0989626692608e-05)),(to_sfixed_a(-2.0296807633712888e-05)),(to_sfixed_a(0.00011640800221357495)),(to_sfixed_a(0.00028652677428908646)),(to_sfixed_a(0.00011137343244627118)),(to_sfixed_a(2.106515967170708e-05)),(to_sfixed_a(-0.00020755015430040658)),(to_sfixed_a(0.00024295109324157238)),(to_sfixed_a(3.801527782343328e-06)),(to_sfixed_a(-0.0002061011764453724)),(to_sfixed_a(0.00014666220522485673)),(to_sfixed_a(3.776025550905615e-06)),(to_sfixed_a(6.833629595348611e-05)),(to_sfixed_a(0.00012665832764469087)),(to_sfixed_a(-6.073360418668017e-05)),(to_sfixed_a(-0.00024188903626054525)),(to_sfixed_a(7.471885328413919e-05)),(to_sfixed_a(-0.00019149991567246616)),(to_sfixed_a(-6.7790417233482e-05)),(to_sfixed_a(-0.00025322724832221866)),(to_sfixed_a(-6.500448216684163e-05)),(to_sfixed_a(-0.0001667989999987185)),(to_sfixed_a(-0.00012090589007129893)),(to_sfixed_a(0.00019310039351694286)),(to_sfixed_a(-0.0002954759111162275)),(to_sfixed_a(-0.00010149428999284282)),(to_sfixed_a(0.00021272698359098285)),(to_sfixed_a(-1.1399919458199292e-05)),(to_sfixed_a(0.0002843186666723341)),(to_sfixed_a(7.591319445054978e-05)),(to_sfixed_a(-7.339932199101895e-05)),(to_sfixed_a(-0.0002470154140610248)),(to_sfixed_a(-2.4628243409097195e-06)),(to_sfixed_a(-2.6949463062919676e-05)),(to_sfixed_a(0.00021709452266804874)),(to_sfixed_a(0.00015082306344993412)),(to_sfixed_a(5.1559651183197275e-05)),(to_sfixed_a(0.0001514749019406736)),(to_sfixed_a(-1.7694910638965666e-06)),(to_sfixed_a(1.6125319234561175e-05)),(to_sfixed_a(-0.0001703404850559309)),(to_sfixed_a(-2.1870495402254164e-05)),(to_sfixed_a(0.00010743489838205278)),(to_sfixed_a(-1.0748699423857033e-05)),(to_sfixed_a(-0.0001524780527688563)),(to_sfixed_a(-0.00015873470692895353)),(to_sfixed_a(-0.0002944343432318419)),(to_sfixed_a(0.0001174186181742698)),(to_sfixed_a(-0.000378615251975134)),(to_sfixed_a(-3.1855524866841733e-05)),(to_sfixed_a(-3.392051439732313e-07)),(to_sfixed_a(-1.494470052421093e-05)),(to_sfixed_a(-0.0001424972724635154)),(to_sfixed_a(0.00018534853006713092)),(to_sfixed_a(3.65083797078114e-05)),(to_sfixed_a(0.0001077037159120664)),(to_sfixed_a(0.00015602483472321182)),(to_sfixed_a(0.00011722554336301982)),(to_sfixed_a(-3.1286464945878834e-05)),(to_sfixed_a(0.00023696768039371818)),(to_sfixed_a(6.980355829000473e-05)),(to_sfixed_a(0.0002507712924852967)),(to_sfixed_a(-0.00016873417189344764)),(to_sfixed_a(0.00014329131226986647)),(to_sfixed_a(-4.375979187898338e-06)),(to_sfixed_a(-0.00019984600658062845)),(to_sfixed_a(1.0549792932579294e-06)),(to_sfixed_a(-3.2542691769776866e-05)),(to_sfixed_a(0.00025128558627329767)),(to_sfixed_a(-1.0534295142861083e-05)),(to_sfixed_a(-2.2050095140002668e-05)),(to_sfixed_a(7.12604378350079e-05)),(to_sfixed_a(0.00011608262138906866)),(to_sfixed_a(5.867551590199582e-05)),(to_sfixed_a(-0.00021965392807032913)),(to_sfixed_a(-0.00027259625494480133)),(to_sfixed_a(2.0942541596014053e-05)),(to_sfixed_a(-0.00011823548993561417)),(to_sfixed_a(-2.29589240916539e-05)),(to_sfixed_a(-0.00013762121670879424)),(to_sfixed_a(-0.00021819525863975286)),(to_sfixed_a(-2.724773366935551e-07)),(to_sfixed_a(-3.912312968168408e-05)),(to_sfixed_a(-5.951053026365116e-06)),(to_sfixed_a(-0.0002893878554459661)),(to_sfixed_a(-3.3405161957489327e-05)),(to_sfixed_a(6.420441786758602e-05)),(to_sfixed_a(0.0003054043627344072)),(to_sfixed_a(-0.0001688081247266382)),(to_sfixed_a(8.738797623664141e-05)),(to_sfixed_a(7.283559534698725e-05)),(to_sfixed_a(-8.273455023299903e-06)),(to_sfixed_a(0.00013417121954262257)),(to_sfixed_a(-0.00018647915567271411)),(to_sfixed_a(-2.984218008350581e-05)),(to_sfixed_a(-7.4107301770709455e-06)),(to_sfixed_a(0.00020780900376848876)),(to_sfixed_a(-0.0001081637165043503)),(to_sfixed_a(-2.0305116777308285e-05)),(to_sfixed_a(7.878267206251621e-05)),(to_sfixed_a(-0.00019090832211077213)),(to_sfixed_a(-3.584675141610205e-06)),(to_sfixed_a(-2.6160385459661484e-05)),(to_sfixed_a(6.040359221515246e-05)),(to_sfixed_a(4.524015821516514e-05)),(to_sfixed_a(2.7171212423127145e-05)),(to_sfixed_a(0.000151271146023646)),(to_sfixed_a(0.000251361692789942)),(to_sfixed_a(-0.0001369713427266106)),(to_sfixed_a(-0.00018248535343445837)),(to_sfixed_a(1.9579572835937142e-05)),(to_sfixed_a(-0.0004256590036675334)),(to_sfixed_a(0.00012776427320204675)),(to_sfixed_a(-8.550556958653033e-05)),(to_sfixed_a(-1.0239979019388556e-05)),(to_sfixed_a(-2.9124552384018898e-05)),(to_sfixed_a(-6.923059117980301e-05)),(to_sfixed_a(-0.0001386083458783105)),(to_sfixed_a(-8.879076631274074e-05)),(to_sfixed_a(-0.00011505266593303531)),(to_sfixed_a(0.00011278709280304611)),(to_sfixed_a(-5.701574991689995e-06)),(to_sfixed_a(-0.00010085157555295154)),(to_sfixed_a(0.00015726752462796867)),(to_sfixed_a(6.559814210049808e-05)),(to_sfixed_a(4.4411979615688324e-05)),(to_sfixed_a(-0.0002503157884348184)),(to_sfixed_a(-6.452416710089892e-05)),(to_sfixed_a(5.500380211742595e-05)),(to_sfixed_a(4.3990974518237635e-05)),(to_sfixed_a(-7.328970241360366e-06)),(to_sfixed_a(-0.00010116604244103655)),(to_sfixed_a(4.410039400681853e-05)),(to_sfixed_a(-0.00012998028250876814)),(to_sfixed_a(0.0001921244984259829)),(to_sfixed_a(-0.00015535447164438665)),(to_sfixed_a(0.00015445200551766902)),(to_sfixed_a(-5.604713805951178e-05)),(to_sfixed_a(-8.743397484067827e-05)),(to_sfixed_a(0.00015574926510453224)),(to_sfixed_a(-8.130627975333482e-07)),(to_sfixed_a(0.00013383483747020364)),(to_sfixed_a(-6.570066034328192e-05)),(to_sfixed_a(-0.00016811754903756082)),(to_sfixed_a(-1.759696169756353e-05)),(to_sfixed_a(4.805429125553928e-05)),(to_sfixed_a(-0.00012995673750992864)),(to_sfixed_a(-3.980768087785691e-05)),(to_sfixed_a(-1.6443082131445408e-06)),(to_sfixed_a(7.019525219220668e-05)),(to_sfixed_a(7.991075835889205e-05)),(to_sfixed_a(-0.00017250538803637028)),(to_sfixed_a(-0.00011510376498335972)),(to_sfixed_a(4.9256854254053906e-05)),(to_sfixed_a(7.339876901824027e-05)),(to_sfixed_a(-5.575013346970081e-06)),(to_sfixed_a(-0.00015921032172627747)),(to_sfixed_a(-0.00019209727179259062)),(to_sfixed_a(8.155403338605538e-05)),(to_sfixed_a(-9.806748857954517e-05)),(to_sfixed_a(-3.4372511436231434e-05)),(to_sfixed_a(3.248767461627722e-05)),(to_sfixed_a(-8.0366269685328e-05)),(to_sfixed_a(0.0001541393285151571)),(to_sfixed_a(-2.5164525141008198e-05)),(to_sfixed_a(-0.00011575799726415426)),(to_sfixed_a(-4.092129529453814e-06)),(to_sfixed_a(-7.080232171574607e-05)),(to_sfixed_a(-6.144527287688106e-05)),(to_sfixed_a(-2.794239844661206e-05)),(to_sfixed_a(0.00010842242045328021)),(to_sfixed_a(4.1464918467681855e-06)),(to_sfixed_a(5.642268661176786e-05)),(to_sfixed_a(-2.068518369924277e-06)));

    constant weight_n2_9 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.295376718044281)),(to_sfixed_a(0.6319247484207153)),(to_sfixed_a(-0.14743825793266296)),(to_sfixed_a(-3.2948511943686754e-05)),(to_sfixed_a(0.011252576485276222)),(to_sfixed_a(0.00014411813754122704)),(to_sfixed_a(0.4154655635356903)),(to_sfixed_a(-0.00015784744755364954)),(to_sfixed_a(0.00015580291801597923)),(to_sfixed_a(0.00023787903774064034)),(to_sfixed_a(6.802812276873738e-05)),(to_sfixed_a(0.26218748092651367)),(to_sfixed_a(-0.0023491759784519672)),(to_sfixed_a(-0.29180553555488586)),(to_sfixed_a(4.611618351191282e-06)),(to_sfixed_a(-0.00015349917521234602)),(to_sfixed_a(-0.009570935741066933)),(to_sfixed_a(-0.00010144786210730672)),(to_sfixed_a(0.01421418972313404)),(to_sfixed_a(-0.0014926902949810028)),(to_sfixed_a(-6.20604696450755e-05)),(to_sfixed_a(-0.00015322111721616238)),(to_sfixed_a(0.001120787812396884)),(to_sfixed_a(-0.0015405084704980254)),(to_sfixed_a(-0.0017412807792425156)),(to_sfixed_a(-0.22526857256889343)),(to_sfixed_a(2.5719200493767858e-06)),(to_sfixed_a(0.000836423016153276)),(to_sfixed_a(-0.0004261438734829426)),(to_sfixed_a(0.00016773918468970805)),(to_sfixed_a(0.24881789088249207)),(to_sfixed_a(-0.00045137040433473885)),(to_sfixed_a(-0.11244305968284607)),(to_sfixed_a(-3.066790304728784e-05)),(to_sfixed_a(0.00024703898816369474)),(to_sfixed_a(0.0002181203744839877)),(to_sfixed_a(0.013789298012852669)),(to_sfixed_a(-0.2866208255290985)),(to_sfixed_a(0.3465654253959656)),(to_sfixed_a(0.00021586967341136187)),(to_sfixed_a(-0.5310841202735901)),(to_sfixed_a(-0.0018527391366660595)),(to_sfixed_a(-0.00014791410649195313)),(to_sfixed_a(-0.00016929040430113673)),(to_sfixed_a(0.006959747988730669)),(to_sfixed_a(0.5149295926094055)),(to_sfixed_a(0.5813756585121155)),(to_sfixed_a(-0.0011859831865876913)),(to_sfixed_a(2.215297718066722e-05)),(to_sfixed_a(0.2089489847421646)),(to_sfixed_a(-0.2675689458847046)),(to_sfixed_a(-0.000759680406190455)),(to_sfixed_a(-0.0002434611669741571)),(to_sfixed_a(-0.0009637931943871081)),(to_sfixed_a(0.0018169311806559563)),(to_sfixed_a(-0.0064163291826844215)),(to_sfixed_a(0.00025620186352171004)),(to_sfixed_a(-0.010533087886869907)),(to_sfixed_a(0.00018627394456416368)),(to_sfixed_a(0.00027937343111261725)),(to_sfixed_a(0.002363660605624318)),(to_sfixed_a(0.0005074668442830443)),(to_sfixed_a(0.0004589401069097221)),(to_sfixed_a(0.3297596871852875)),(to_sfixed_a(0.00011456572246970609)),(to_sfixed_a(-0.10208987444639206)),(to_sfixed_a(0.0002503512951079756)),(to_sfixed_a(-0.006675777491182089)),(to_sfixed_a(-0.012720203027129173)),(to_sfixed_a(-4.342013198765926e-05)),(to_sfixed_a(0.02911028265953064)),(to_sfixed_a(-0.005783496890217066)),(to_sfixed_a(-0.013500421307981014)),(to_sfixed_a(-0.00012921880988869816)),(to_sfixed_a(8.931526099331677e-05)),(to_sfixed_a(5.342887743609026e-05)),(to_sfixed_a(-0.00021111223031766713)),(to_sfixed_a(-0.007968406192958355)),(to_sfixed_a(0.00012905984476674348)),(to_sfixed_a(0.35052675008773804)),(to_sfixed_a(0.07589341700077057)),(to_sfixed_a(0.0002463931741658598)),(to_sfixed_a(0.4796319007873535)),(to_sfixed_a(0.022037111222743988)),(to_sfixed_a(0.0003217074554413557)),(to_sfixed_a(0.00034806315670721233)),(to_sfixed_a(-0.09056118130683899)),(to_sfixed_a(-1.048816557158716e-05)),(to_sfixed_a(-0.0001818114542402327)),(to_sfixed_a(0.00011328820983180776)),(to_sfixed_a(0.13909423351287842)),(to_sfixed_a(0.00021200274932198226)),(to_sfixed_a(0.0014426754787564278)),(to_sfixed_a(-6.992588168941438e-06)),(to_sfixed_a(-0.00441324757412076)),(to_sfixed_a(-1.1496333172544837e-05)),(to_sfixed_a(-3.57838325726334e-05)),(to_sfixed_a(-2.9640941647812724e-05)),(to_sfixed_a(-3.17450103466399e-05)),(to_sfixed_a(4.802881448995322e-06)),(to_sfixed_a(-0.001841154065914452)),(to_sfixed_a(0.00015918634016998112)),(to_sfixed_a(0.00011332850408507511)),(to_sfixed_a(0.3661409914493561)),(to_sfixed_a(0.29584404826164246)),(to_sfixed_a(6.25679676886648e-05)),(to_sfixed_a(-0.00016827238141559064)),(to_sfixed_a(3.570392800611444e-05)),(to_sfixed_a(1.9599145161919296e-05)),(to_sfixed_a(0.23780079185962677)),(to_sfixed_a(0.009860758669674397)),(to_sfixed_a(4.002329660579562e-06)),(to_sfixed_a(0.005826189182698727)),(to_sfixed_a(-5.827505447086878e-05)),(to_sfixed_a(0.00015405636804644018)),(to_sfixed_a(-0.002656914759427309)),(to_sfixed_a(0.00165564042981714)),(to_sfixed_a(-0.006043381989002228)),(to_sfixed_a(0.0001712836092337966)),(to_sfixed_a(-0.00011298558820271865)),(to_sfixed_a(-0.00015450746286660433)),(to_sfixed_a(-2.316975951544009e-05)),(to_sfixed_a(-0.010199102573096752)),(to_sfixed_a(-7.225036097224802e-05)),(to_sfixed_a(-0.00020546924497466534)),(to_sfixed_a(5.203588807489723e-05)),(to_sfixed_a(0.000532209814991802)),(to_sfixed_a(4.070690192747861e-05)),(to_sfixed_a(-3.901678428519517e-05)),(to_sfixed_a(-1.502578379586339e-05)),(to_sfixed_a(-2.9378352337516844e-05)),(to_sfixed_a(6.192510045366362e-05)),(to_sfixed_a(0.0012394522782415152)),(to_sfixed_a(0.004809812176972628)),(to_sfixed_a(9.738343942444772e-05)),(to_sfixed_a(-6.05579734838102e-05)),(to_sfixed_a(-0.09234855324029922)),(to_sfixed_a(-0.22632984817028046)),(to_sfixed_a(0.00014971342170611024)),(to_sfixed_a(-0.00023833825252950191)),(to_sfixed_a(0.00019036441517528147)),(to_sfixed_a(-4.610772157320753e-05)),(to_sfixed_a(-0.00010827337973751128)),(to_sfixed_a(0.36798790097236633)),(to_sfixed_a(0.4185580313205719)),(to_sfixed_a(8.036859071580693e-05)),(to_sfixed_a(-0.0008567081531509757)),(to_sfixed_a(0.0002545209717936814)),(to_sfixed_a(-0.000174358268850483)),(to_sfixed_a(-0.010876634158194065)),(to_sfixed_a(-6.763108831364661e-05)),(to_sfixed_a(4.390208050608635e-05)),(to_sfixed_a(-0.01535434927791357)),(to_sfixed_a(0.00027395127108320594)),(to_sfixed_a(-3.0733528546988964e-05)),(to_sfixed_a(-0.0405123345553875)),(to_sfixed_a(8.814866305328906e-06)),(to_sfixed_a(0.0019802413880825043)),(to_sfixed_a(4.310488293413073e-05)),(to_sfixed_a(2.1405459847301245e-05)),(to_sfixed_a(5.7933117204811424e-05)),(to_sfixed_a(0.0002996508846990764)),(to_sfixed_a(0.00432888139039278)),(to_sfixed_a(5.56204431632068e-05)),(to_sfixed_a(-0.002594465622678399)),(to_sfixed_a(0.4233928322792053)),(to_sfixed_a(0.00018550257664173841)),(to_sfixed_a(-0.29632753133773804)),(to_sfixed_a(1.6087942640297115e-05)),(to_sfixed_a(5.069166581961326e-05)),(to_sfixed_a(-0.006988024339079857)),(to_sfixed_a(-0.0071854195557534695)),(to_sfixed_a(-0.0014136781683191657)),(to_sfixed_a(-1.961134694283828e-05)),(to_sfixed_a(0.004094169475138187)),(to_sfixed_a(0.00010244836448691785)),(to_sfixed_a(-0.4883648157119751)),(to_sfixed_a(-0.14723433554172516)),(to_sfixed_a(-0.001147587550804019)),(to_sfixed_a(0.15453776717185974)),(to_sfixed_a(-0.0016523487865924835)),(to_sfixed_a(-0.009542591869831085)),(to_sfixed_a(-0.00013634416973218322)),(to_sfixed_a(1.2182405043859035e-05)),(to_sfixed_a(-1.2599539331858978e-06)),(to_sfixed_a(0.005536745768040419)),(to_sfixed_a(0.0008171009831130505)),(to_sfixed_a(-0.0016450013499706984)),(to_sfixed_a(-0.0695885419845581)),(to_sfixed_a(0.09221925586462021)),(to_sfixed_a(-0.0005335601745173335)),(to_sfixed_a(0.00012965714267920703)),(to_sfixed_a(-0.22559335827827454)),(to_sfixed_a(-0.00795290619134903)),(to_sfixed_a(-1.753525430103764e-05)),(to_sfixed_a(0.006252209190279245)),(to_sfixed_a(1.7393846064805984e-05)),(to_sfixed_a(0.0621231347322464)),(to_sfixed_a(0.4413323402404785)),(to_sfixed_a(-0.00014769501285627484)),(to_sfixed_a(1.2564225471578538e-05)),(to_sfixed_a(-3.0373983463505283e-05)),(to_sfixed_a(-1.2589651305461302e-05)),(to_sfixed_a(-1.1765732779167593e-06)),(to_sfixed_a(-0.00016774266259744763)),(to_sfixed_a(0.5139986276626587)),(to_sfixed_a(0.4764069616794586)),(to_sfixed_a(0.001996018458157778)),(to_sfixed_a(-0.004992817062884569)),(to_sfixed_a(0.0008637510472908616)),(to_sfixed_a(-0.010737273842096329)),(to_sfixed_a(2.2329848434310406e-05)),(to_sfixed_a(0.00011287588131381199)),(to_sfixed_a(7.630690379301086e-05)),(to_sfixed_a(-1.722958404570818e-05)),(to_sfixed_a(-0.00011998163972748443)),(to_sfixed_a(3.232780727557838e-07)),(to_sfixed_a(-0.2378089278936386)),(to_sfixed_a(-0.015650790184736252)),(to_sfixed_a(0.00015497305139433593)),(to_sfixed_a(0.000166024750797078)),(to_sfixed_a(5.393725587055087e-06)),(to_sfixed_a(0.00029087718576192856)),(to_sfixed_a(0.0005799629143439233)),(to_sfixed_a(0.32140517234802246)),(to_sfixed_a(-6.975380529183894e-05)),(to_sfixed_a(-8.794899622444063e-05)),(to_sfixed_a(3.8296988350339234e-05)),(to_sfixed_a(0.4894195795059204)),(to_sfixed_a(0.5439329743385315)),(to_sfixed_a(-0.0028566301334649324)),(to_sfixed_a(-0.00016655099170748144)),(to_sfixed_a(3.104418283328414e-06)),(to_sfixed_a(5.9217953094048426e-05)),(to_sfixed_a(0.0038449415005743504)),(to_sfixed_a(-0.00037484674248844385)),(to_sfixed_a(0.015710581094026566)),(to_sfixed_a(1.658450491959229e-05)),(to_sfixed_a(-0.0011924176942557096)),(to_sfixed_a(-7.917564653325826e-05)),(to_sfixed_a(0.07601039856672287)),(to_sfixed_a(0.00038142129778862)),(to_sfixed_a(-0.001818404532968998)),(to_sfixed_a(2.00783324544318e-06)),(to_sfixed_a(-0.8731244206428528)),(to_sfixed_a(-0.001867590588517487)),(to_sfixed_a(0.017984844744205475)),(to_sfixed_a(0.010275484062731266)),(to_sfixed_a(-0.00011297891614958644)),(to_sfixed_a(-0.0026360435876995325)),(to_sfixed_a(0.0007868322427384555)),(to_sfixed_a(-0.00023962008708622307)),(to_sfixed_a(8.704101492185146e-05)),(to_sfixed_a(-3.0144092306727543e-05)),(to_sfixed_a(0.0004635055083781481)),(to_sfixed_a(0.0009550431277602911)),(to_sfixed_a(-0.1757456660270691)),(to_sfixed_a(-0.00020547202439047396)),(to_sfixed_a(-0.0002046778390649706)),(to_sfixed_a(0.00035079196095466614)),(to_sfixed_a(0.00010724650201154873)),(to_sfixed_a(-0.0016516833566129208)),(to_sfixed_a(9.59975368459709e-05)),(to_sfixed_a(-0.001666569383814931)),(to_sfixed_a(6.816131644882262e-05)),(to_sfixed_a(-0.5396603345870972)),(to_sfixed_a(-0.0004218144458718598)),(to_sfixed_a(0.0001564578851684928)),(to_sfixed_a(0.00014929016469977796)),(to_sfixed_a(0.004845826420933008)),(to_sfixed_a(0.2737736701965332)),(to_sfixed_a(-1.1492666089907289e-06)),(to_sfixed_a(0.0002958611003123224)),(to_sfixed_a(-1.9983399397460744e-05)),(to_sfixed_a(1.2986609362997115e-05)),(to_sfixed_a(-0.0030553035903722048)),(to_sfixed_a(-0.0028551907744258642)),(to_sfixed_a(-0.0012104986235499382)),(to_sfixed_a(0.020870277658104897)),(to_sfixed_a(0.3066520392894745)),(to_sfixed_a(0.0001465087989345193)),(to_sfixed_a(3.0354927730513737e-05)),(to_sfixed_a(1.0189150998485275e-05)),(to_sfixed_a(-0.00086678855586797)),(to_sfixed_a(0.00025054544676095247)),(to_sfixed_a(0.0003839516721200198)),(to_sfixed_a(-3.042820571863558e-05)),(to_sfixed_a(0.013050318695604801)),(to_sfixed_a(1.1071992048528045e-05)),(to_sfixed_a(0.8360999226570129)),(to_sfixed_a(-0.0017115422524511814)),(to_sfixed_a(0.30078259110450745)),(to_sfixed_a(-0.0008390639559365809)),(to_sfixed_a(-4.694944800576195e-05)),(to_sfixed_a(-0.0019021754851564765)),(to_sfixed_a(0.00016795947158243507)),(to_sfixed_a(0.008695455268025398)),(to_sfixed_a(0.00015092449029907584)),(to_sfixed_a(-0.15214575827121735)),(to_sfixed_a(-0.008376868441700935)),(to_sfixed_a(-0.30536332726478577)));

    constant weight_n2_10 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.20960234105587006)),(to_sfixed_a(-0.23156404495239258)),(to_sfixed_a(-0.7164607048034668)),(to_sfixed_a(6.306017166934907e-05)),(to_sfixed_a(0.002464896533638239)),(to_sfixed_a(0.00022154119506012648)),(to_sfixed_a(-0.0011718260357156396)),(to_sfixed_a(0.0001899505587061867)),(to_sfixed_a(-5.5487616918981075e-06)),(to_sfixed_a(-0.00041777355363592505)),(to_sfixed_a(0.0001686745381448418)),(to_sfixed_a(-0.002873701509088278)),(to_sfixed_a(0.0005468036979436874)),(to_sfixed_a(-5.372889063437469e-05)),(to_sfixed_a(0.00024086413031909615)),(to_sfixed_a(3.661678056232631e-05)),(to_sfixed_a(0.0010866258526220918)),(to_sfixed_a(7.002049096627161e-05)),(to_sfixed_a(-0.006347022019326687)),(to_sfixed_a(-0.005370498634874821)),(to_sfixed_a(-2.47634707193356e-05)),(to_sfixed_a(-0.000163591728778556)),(to_sfixed_a(-2.9118733436916955e-05)),(to_sfixed_a(0.0012558848829939961)),(to_sfixed_a(-0.0007695772219449282)),(to_sfixed_a(0.02828577719628811)),(to_sfixed_a(-0.00030806672293692827)),(to_sfixed_a(-0.0011767984833568335)),(to_sfixed_a(0.00021289440337568521)),(to_sfixed_a(0.0001518126082373783)),(to_sfixed_a(0.1149013414978981)),(to_sfixed_a(-0.00018941276357509196)),(to_sfixed_a(0.2361564040184021)),(to_sfixed_a(7.098860805854201e-05)),(to_sfixed_a(2.4989654775708914e-05)),(to_sfixed_a(9.872695954982191e-05)),(to_sfixed_a(-0.0011921296827495098)),(to_sfixed_a(-0.0002839973021764308)),(to_sfixed_a(-0.4677499830722809)),(to_sfixed_a(-1.5798432286828756e-06)),(to_sfixed_a(0.0005005376879125834)),(to_sfixed_a(0.27478063106536865)),(to_sfixed_a(-0.00010536057379795238)),(to_sfixed_a(-9.487279021413997e-05)),(to_sfixed_a(-0.009659785777330399)),(to_sfixed_a(-0.008143818937242031)),(to_sfixed_a(-0.6062712669372559)),(to_sfixed_a(-0.001010335050523281)),(to_sfixed_a(-4.519151116255671e-05)),(to_sfixed_a(0.0012679444625973701)),(to_sfixed_a(-0.00270282500423491)),(to_sfixed_a(4.8896719818003476e-05)),(to_sfixed_a(-0.00014183000894263387)),(to_sfixed_a(-0.0002473045024089515)),(to_sfixed_a(-0.002441172720864415)),(to_sfixed_a(-0.00015251703734975308)),(to_sfixed_a(-0.0002913276548497379)),(to_sfixed_a(-0.011469329707324505)),(to_sfixed_a(-7.180100510595366e-05)),(to_sfixed_a(0.0002229609526693821)),(to_sfixed_a(-0.004924374166876078)),(to_sfixed_a(-1.99371570488438e-05)),(to_sfixed_a(-0.000916309014428407)),(to_sfixed_a(0.0028719494584947824)),(to_sfixed_a(3.369331534486264e-05)),(to_sfixed_a(0.0006712275207974017)),(to_sfixed_a(-7.128887227736413e-05)),(to_sfixed_a(0.006006999406963587)),(to_sfixed_a(-0.00015882053412497044)),(to_sfixed_a(-5.4524134611710906e-05)),(to_sfixed_a(-0.1784057915210724)),(to_sfixed_a(-0.005705111660063267)),(to_sfixed_a(-2.2380243535735644e-05)),(to_sfixed_a(-1.2156728189438581e-05)),(to_sfixed_a(0.00012072641402482986)),(to_sfixed_a(0.00010479785851202905)),(to_sfixed_a(-0.007533482275903225)),(to_sfixed_a(-4.600624379236251e-05)),(to_sfixed_a(0.00013995837070979178)),(to_sfixed_a(2.265696821268648e-06)),(to_sfixed_a(-0.012048606760799885)),(to_sfixed_a(0.00014998079859651625)),(to_sfixed_a(0.00017733342247083783)),(to_sfixed_a(-0.002250327728688717)),(to_sfixed_a(-1.0188459782511927e-05)),(to_sfixed_a(-0.002044076332822442)),(to_sfixed_a(0.003539629280567169)),(to_sfixed_a(-0.0001149949966929853)),(to_sfixed_a(2.9421182262012735e-05)),(to_sfixed_a(-0.0001009928819257766)),(to_sfixed_a(-0.5643952488899231)),(to_sfixed_a(-0.00011387010454200208)),(to_sfixed_a(0.2816363275051117)),(to_sfixed_a(0.00023714501003269106)),(to_sfixed_a(-0.000848044699523598)),(to_sfixed_a(0.00024019903503358364)),(to_sfixed_a(7.173695485107601e-05)),(to_sfixed_a(0.00010318458953406662)),(to_sfixed_a(0.0002474283683113754)),(to_sfixed_a(6.694428157061338e-05)),(to_sfixed_a(0.4912737011909485)),(to_sfixed_a(-0.0009203857625834644)),(to_sfixed_a(-0.00020533186034299433)),(to_sfixed_a(-0.006200030446052551)),(to_sfixed_a(-0.009269117377698421)),(to_sfixed_a(-0.000456764071714133)),(to_sfixed_a(0.00021975001436658204)),(to_sfixed_a(-7.454689330188558e-05)),(to_sfixed_a(-0.00018604395154397935)),(to_sfixed_a(-0.003735026577487588)),(to_sfixed_a(-0.0008589091012254357)),(to_sfixed_a(0.00015462924784515053)),(to_sfixed_a(-0.0004286316398065537)),(to_sfixed_a(-6.76274357829243e-05)),(to_sfixed_a(-5.707763193640858e-05)),(to_sfixed_a(0.03136240318417549)),(to_sfixed_a(-0.00019286471069790423)),(to_sfixed_a(1.8676117178983986e-05)),(to_sfixed_a(9.535792196402326e-05)),(to_sfixed_a(0.0003723307163454592)),(to_sfixed_a(0.00015409514890052378)),(to_sfixed_a(-0.00018058647401630878)),(to_sfixed_a(-0.009884849190711975)),(to_sfixed_a(-0.00013007133384235203)),(to_sfixed_a(8.618535503046587e-07)),(to_sfixed_a(0.14498591423034668)),(to_sfixed_a(0.2544005215167999)),(to_sfixed_a(-0.00010809399100253358)),(to_sfixed_a(-0.00015794960199855268)),(to_sfixed_a(4.730900400318205e-06)),(to_sfixed_a(1.748432987369597e-05)),(to_sfixed_a(5.969575795461424e-05)),(to_sfixed_a(0.00030565191991627216)),(to_sfixed_a(-0.004087027627974749)),(to_sfixed_a(-0.0001658877299632877)),(to_sfixed_a(3.971466503571719e-05)),(to_sfixed_a(-0.010405891574919224)),(to_sfixed_a(-0.0006884575705043972)),(to_sfixed_a(-3.0166269425535575e-05)),(to_sfixed_a(-8.794477616902441e-05)),(to_sfixed_a(-0.0006567303789779544)),(to_sfixed_a(9.432152000954375e-05)),(to_sfixed_a(4.676739627029747e-05)),(to_sfixed_a(1.2659102139878087e-05)),(to_sfixed_a(8.226613863371313e-05)),(to_sfixed_a(0.00018525138148106635)),(to_sfixed_a(-5.794427124783397e-06)),(to_sfixed_a(0.00015019682177808136)),(to_sfixed_a(-3.5139964893460274e-07)),(to_sfixed_a(-0.0473775789141655)),(to_sfixed_a(-0.00014862029638607055)),(to_sfixed_a(0.00015829078620299697)),(to_sfixed_a(0.00023607659386470914)),(to_sfixed_a(-0.0001340594608336687)),(to_sfixed_a(0.0003791323397308588)),(to_sfixed_a(0.08285356312990189)),(to_sfixed_a(-0.0001793579285731539)),(to_sfixed_a(-0.002012063516303897)),(to_sfixed_a(-0.00030206225346773863)),(to_sfixed_a(-6.226076220627874e-05)),(to_sfixed_a(0.0002951185160782188)),(to_sfixed_a(0.00014917498629074544)),(to_sfixed_a(-0.0041112108156085014)),(to_sfixed_a(0.00477329408749938)),(to_sfixed_a(-6.460365693783388e-05)),(to_sfixed_a(-0.0006411880603991449)),(to_sfixed_a(7.781601743772626e-05)),(to_sfixed_a(7.644764264114201e-05)),(to_sfixed_a(-3.7744139262940735e-05)),(to_sfixed_a(-8.368001726921648e-05)),(to_sfixed_a(0.004559551365673542)),(to_sfixed_a(-0.00011093995999544859)),(to_sfixed_a(-8.917318336898461e-05)),(to_sfixed_a(6.925583875272423e-05)),(to_sfixed_a(0.0002135463582817465)),(to_sfixed_a(0.0007418913883157074)),(to_sfixed_a(-0.001573347020894289)),(to_sfixed_a(-0.001265249797143042)),(to_sfixed_a(-0.43603605031967163)),(to_sfixed_a(-0.011517203412950039)),(to_sfixed_a(-5.4460979299619794e-05)),(to_sfixed_a(-0.00019102453370578587)),(to_sfixed_a(-4.310960866860114e-05)),(to_sfixed_a(-0.00017651350935921073)),(to_sfixed_a(-2.4383043637499213e-05)),(to_sfixed_a(-3.177870166837238e-05)),(to_sfixed_a(-0.001700812834315002)),(to_sfixed_a(0.00022229418391361833)),(to_sfixed_a(-0.0014226260827854276)),(to_sfixed_a(-0.0006462481687776744)),(to_sfixed_a(-0.01321294903755188)),(to_sfixed_a(5.8775411162059754e-05)),(to_sfixed_a(-0.0009232907323166728)),(to_sfixed_a(0.0011893871705979109)),(to_sfixed_a(8.542847353965044e-05)),(to_sfixed_a(-0.001215930562466383)),(to_sfixed_a(-2.461907934048213e-05)),(to_sfixed_a(0.0015966627979651093)),(to_sfixed_a(-0.0031452502589672804)),(to_sfixed_a(-0.00018268964777234942)),(to_sfixed_a(2.751059946604073e-05)),(to_sfixed_a(6.353096250677481e-05)),(to_sfixed_a(0.00023194734239950776)),(to_sfixed_a(0.00014718377497047186)),(to_sfixed_a(-2.9079827072564512e-05)),(to_sfixed_a(-9.313742339145392e-05)),(to_sfixed_a(-0.0013079890049993992)),(to_sfixed_a(0.0011531971395015717)),(to_sfixed_a(0.0029499526135623455)),(to_sfixed_a(-0.0009917384013533592)),(to_sfixed_a(-0.001784570631571114)),(to_sfixed_a(-3.840013960143551e-07)),(to_sfixed_a(0.0001150180323747918)),(to_sfixed_a(5.5897551646921784e-05)),(to_sfixed_a(6.571195262949914e-05)),(to_sfixed_a(-8.619514846941456e-05)),(to_sfixed_a(-0.0010488313855603337)),(to_sfixed_a(-0.003754212288185954)),(to_sfixed_a(-0.014611435122787952)),(to_sfixed_a(6.637386832153425e-05)),(to_sfixed_a(-0.00011213916150154546)),(to_sfixed_a(0.00025157982599921525)),(to_sfixed_a(-1.2618227628991008e-05)),(to_sfixed_a(-0.005782066844403744)),(to_sfixed_a(-0.01728671044111252)),(to_sfixed_a(0.0003759757673833519)),(to_sfixed_a(0.00014840766380075365)),(to_sfixed_a(6.888678035466e-05)),(to_sfixed_a(-0.002503489376977086)),(to_sfixed_a(0.005089742597192526)),(to_sfixed_a(-0.5702447295188904)),(to_sfixed_a(-8.550028724130243e-05)),(to_sfixed_a(-8.48367199068889e-05)),(to_sfixed_a(-1.0470830602571368e-07)),(to_sfixed_a(0.0001265845203306526)),(to_sfixed_a(0.00023157638497650623)),(to_sfixed_a(-0.012584223411977291)),(to_sfixed_a(-5.851874448126182e-05)),(to_sfixed_a(0.0007838158635422587)),(to_sfixed_a(1.0808143997564912e-05)),(to_sfixed_a(-0.0002987014304380864)),(to_sfixed_a(-0.00019957170297857374)),(to_sfixed_a(5.136995605425909e-05)),(to_sfixed_a(0.0001023158329189755)),(to_sfixed_a(0.0020097449887543917)),(to_sfixed_a(-0.0007186115835793316)),(to_sfixed_a(0.420283704996109)),(to_sfixed_a(-0.0025966311804950237)),(to_sfixed_a(-7.04996709828265e-05)),(to_sfixed_a(-0.007257732562720776)),(to_sfixed_a(-0.007752560544759035)),(to_sfixed_a(0.00015603212523274124)),(to_sfixed_a(-0.0016657526139169931)),(to_sfixed_a(-0.00017668638611212373)),(to_sfixed_a(-2.1066274712211452e-05)),(to_sfixed_a(0.0027654743753373623)),(to_sfixed_a(-0.008962144143879414)),(to_sfixed_a(-2.8217276849318296e-05)),(to_sfixed_a(4.4574506318895146e-05)),(to_sfixed_a(0.332967072725296)),(to_sfixed_a(0.0002096310636261478)),(to_sfixed_a(-0.00024398750974796712)),(to_sfixed_a(0.00030177869484759867)),(to_sfixed_a(-2.3739437892800197e-05)),(to_sfixed_a(-0.00010487948748050258)),(to_sfixed_a(0.006333417259156704)),(to_sfixed_a(-0.00013326579937711358)),(to_sfixed_a(0.00045090983621776104)),(to_sfixed_a(-7.01967510394752e-05)),(to_sfixed_a(-0.02139207161962986)),(to_sfixed_a(-0.0018615233711898327)),(to_sfixed_a(0.00015536471619270742)),(to_sfixed_a(5.677234003087506e-05)),(to_sfixed_a(2.224092895630747e-06)),(to_sfixed_a(0.00018485287728253752)),(to_sfixed_a(0.011224490590393543)),(to_sfixed_a(-0.0015159685863181949)),(to_sfixed_a(0.0018039240967482328)),(to_sfixed_a(-0.007215374149382114)),(to_sfixed_a(-0.006956021301448345)),(to_sfixed_a(0.0002017051592702046)),(to_sfixed_a(-0.00011699362949002534)),(to_sfixed_a(0.00018152096890844405)),(to_sfixed_a(-7.850547262933105e-05)),(to_sfixed_a(-0.00021492369705811143)),(to_sfixed_a(-1.5155737855820917e-05)),(to_sfixed_a(-0.00227857637219131)),(to_sfixed_a(0.005634180270135403)),(to_sfixed_a(0.00012571687693707645)),(to_sfixed_a(9.201964712701738e-05)),(to_sfixed_a(0.18494060635566711)),(to_sfixed_a(-0.0034468574449419975)),(to_sfixed_a(0.0029838967602699995)),(to_sfixed_a(-6.953000411158428e-05)),(to_sfixed_a(0.00723045039921999)),(to_sfixed_a(-2.8263466447242536e-06)),(to_sfixed_a(-0.011445291340351105)),(to_sfixed_a(4.917019396089017e-07)),(to_sfixed_a(-0.0048229084350168705)),(to_sfixed_a(0.005849997978657484)),(to_sfixed_a(-0.003998329862952232)));

    constant weight_n2_11 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.05202234908938408)),(to_sfixed_a(-0.0021910914219915867)),(to_sfixed_a(-0.8352421522140503)),(to_sfixed_a(-6.795593071728945e-05)),(to_sfixed_a(-0.00914974045008421)),(to_sfixed_a(-0.0003797072567977011)),(to_sfixed_a(-0.013349127024412155)),(to_sfixed_a(4.667454049922526e-06)),(to_sfixed_a(-7.706748874625191e-05)),(to_sfixed_a(4.842676571570337e-05)),(to_sfixed_a(-5.734367005061358e-05)),(to_sfixed_a(0.0030661551281809807)),(to_sfixed_a(-0.0002213288244092837)),(to_sfixed_a(-0.00020198857237119228)),(to_sfixed_a(3.974066930823028e-05)),(to_sfixed_a(-3.2055031624622643e-06)),(to_sfixed_a(-0.006295270752161741)),(to_sfixed_a(-7.147734868340194e-05)),(to_sfixed_a(0.000644079758785665)),(to_sfixed_a(0.136184424161911)),(to_sfixed_a(-0.00013717316323891282)),(to_sfixed_a(-0.00019761350995395333)),(to_sfixed_a(-0.00033263248042203486)),(to_sfixed_a(0.0054120877757668495)),(to_sfixed_a(-0.005466381087899208)),(to_sfixed_a(-0.002170137595385313)),(to_sfixed_a(-2.3250737285707146e-05)),(to_sfixed_a(-0.00021861682762391865)),(to_sfixed_a(0.047812677919864655)),(to_sfixed_a(-3.922839823644608e-06)),(to_sfixed_a(0.3630439341068268)),(to_sfixed_a(0.0001814012648537755)),(to_sfixed_a(0.014824590645730495)),(to_sfixed_a(5.753092409577221e-05)),(to_sfixed_a(-7.621665281476453e-05)),(to_sfixed_a(-0.00045843308907933533)),(to_sfixed_a(-0.003156819846481085)),(to_sfixed_a(0.006943386979401112)),(to_sfixed_a(-0.003148982534185052)),(to_sfixed_a(6.750304601155221e-05)),(to_sfixed_a(-0.011909282766282558)),(to_sfixed_a(-0.39038175344467163)),(to_sfixed_a(8.510069892508909e-05)),(to_sfixed_a(5.944908480159938e-05)),(to_sfixed_a(0.004061858635395765)),(to_sfixed_a(0.3530571460723877)),(to_sfixed_a(-0.004288829863071442)),(to_sfixed_a(-0.009819055907428265)),(to_sfixed_a(-5.0920840294566005e-05)),(to_sfixed_a(-0.0064469752833247185)),(to_sfixed_a(0.009188386611640453)),(to_sfixed_a(-0.0005954933585599065)),(to_sfixed_a(-9.439785208087415e-05)),(to_sfixed_a(-0.002126189647242427)),(to_sfixed_a(-0.0025934940204024315)),(to_sfixed_a(0.307087242603302)),(to_sfixed_a(0.0003014283429365605)),(to_sfixed_a(-0.002296482678502798)),(to_sfixed_a(2.8737777029164135e-06)),(to_sfixed_a(7.750284567009658e-05)),(to_sfixed_a(7.032569556031376e-05)),(to_sfixed_a(-0.00040188070852309465)),(to_sfixed_a(0.40347087383270264)),(to_sfixed_a(-0.005268456880003214)),(to_sfixed_a(0.00015091305249370635)),(to_sfixed_a(-0.0011634397087618709)),(to_sfixed_a(5.749814590672031e-05)),(to_sfixed_a(-0.0005663862102665007)),(to_sfixed_a(-0.0003836259711533785)),(to_sfixed_a(6.400776328518987e-05)),(to_sfixed_a(0.008526856079697609)),(to_sfixed_a(-0.013915130868554115)),(to_sfixed_a(0.28369492292404175)),(to_sfixed_a(-0.00016334198880940676)),(to_sfixed_a(0.00011200781591469422)),(to_sfixed_a(-0.00017576548270881176)),(to_sfixed_a(-0.003724360838532448)),(to_sfixed_a(-0.2991935908794403)),(to_sfixed_a(0.00010460232442710549)),(to_sfixed_a(-0.38148918747901917)),(to_sfixed_a(-0.01137594599276781)),(to_sfixed_a(6.074440898373723e-05)),(to_sfixed_a(-0.0006140244076959789)),(to_sfixed_a(-0.004151216708123684)),(to_sfixed_a(-0.00018178447498939931)),(to_sfixed_a(-0.010141043923795223)),(to_sfixed_a(0.28025245666503906)),(to_sfixed_a(-0.0006116266013123095)),(to_sfixed_a(0.00013787818897981197)),(to_sfixed_a(0.00010166307765757665)),(to_sfixed_a(6.7902758019045e-05)),(to_sfixed_a(0.00028560232021845877)),(to_sfixed_a(0.37624916434288025)),(to_sfixed_a(-0.00013588499859906733)),(to_sfixed_a(0.0009829183109104633)),(to_sfixed_a(-0.00020843822858296335)),(to_sfixed_a(-5.3858919272897765e-05)),(to_sfixed_a(0.00017042031686287373)),(to_sfixed_a(-4.812044062418863e-05)),(to_sfixed_a(-0.00011305048246867955)),(to_sfixed_a(-0.002439271891489625)),(to_sfixed_a(-0.0007760850130580366)),(to_sfixed_a(-9.111743565881625e-05)),(to_sfixed_a(0.42655766010284424)),(to_sfixed_a(-0.0007243569125421345)),(to_sfixed_a(-0.003979505505412817)),(to_sfixed_a(-0.00010128474968951195)),(to_sfixed_a(-0.00014377049228642136)),(to_sfixed_a(1.87441983143799e-05)),(to_sfixed_a(-0.012632153928279877)),(to_sfixed_a(-0.004562476649880409)),(to_sfixed_a(-0.0001504069077782333)),(to_sfixed_a(0.06019919738173485)),(to_sfixed_a(4.6321001718752086e-05)),(to_sfixed_a(6.940487946849316e-05)),(to_sfixed_a(-0.011006451211869717)),(to_sfixed_a(0.0041626389138400555)),(to_sfixed_a(-0.0015236185863614082)),(to_sfixed_a(0.0004202031996101141)),(to_sfixed_a(0.0017642802558839321)),(to_sfixed_a(-0.00015695109323132783)),(to_sfixed_a(-0.00020615194807760417)),(to_sfixed_a(-0.01621847413480282)),(to_sfixed_a(7.691954670008272e-05)),(to_sfixed_a(-7.708396879024804e-06)),(to_sfixed_a(0.0088281761854887)),(to_sfixed_a(-0.09138685464859009)),(to_sfixed_a(-7.280506542883813e-05)),(to_sfixed_a(-0.00018618801550474018)),(to_sfixed_a(0.0004223703290335834)),(to_sfixed_a(0.00024642731295898557)),(to_sfixed_a(0.00011293014540569857)),(to_sfixed_a(-0.007889688946306705)),(to_sfixed_a(-0.00025317614199593663)),(to_sfixed_a(-0.00016798697470221668)),(to_sfixed_a(-0.0002931139897555113)),(to_sfixed_a(-0.541267991065979)),(to_sfixed_a(-0.00266807503066957)),(to_sfixed_a(3.36937555402983e-05)),(to_sfixed_a(4.451445784070529e-05)),(to_sfixed_a(-0.00013870885595679283)),(to_sfixed_a(0.00012043150491081178)),(to_sfixed_a(0.00011359740165062249)),(to_sfixed_a(-1.5814735888852738e-05)),(to_sfixed_a(-0.0012544282944872975)),(to_sfixed_a(-0.00037077473825775087)),(to_sfixed_a(-0.00864199735224247)),(to_sfixed_a(0.0001548910076962784)),(to_sfixed_a(4.2938256228808314e-05)),(to_sfixed_a(-0.0006786516169086099)),(to_sfixed_a(-2.385120023973286e-05)),(to_sfixed_a(-7.96201202319935e-05)),(to_sfixed_a(-0.0008464292623102665)),(to_sfixed_a(-2.5119123165495694e-05)),(to_sfixed_a(0.00023595377570018172)),(to_sfixed_a(0.02569917030632496)),(to_sfixed_a(9.580930782249197e-05)),(to_sfixed_a(-0.6522176265716553)),(to_sfixed_a(-0.00012030127254547551)),(to_sfixed_a(-0.00016917215543799102)),(to_sfixed_a(6.889023643452674e-05)),(to_sfixed_a(0.00010622521222103387)),(to_sfixed_a(-0.0004890427808277309)),(to_sfixed_a(-5.430986129795201e-05)),(to_sfixed_a(-0.008055135607719421)),(to_sfixed_a(-0.00545137096196413)),(to_sfixed_a(0.00010618737724144012)),(to_sfixed_a(-7.262607687152922e-05)),(to_sfixed_a(-0.0001046837423928082)),(to_sfixed_a(-6.993361603235826e-05)),(to_sfixed_a(-0.0016175979981198907)),(to_sfixed_a(-0.001673170831054449)),(to_sfixed_a(0.005002439487725496)),(to_sfixed_a(1.3168028090149164e-06)),(to_sfixed_a(0.01892751455307007)),(to_sfixed_a(0.00673281354829669)),(to_sfixed_a(-0.0022131099831312895)),(to_sfixed_a(-0.40466612577438354)),(to_sfixed_a(0.011793641373515129)),(to_sfixed_a(0.00928221084177494)),(to_sfixed_a(-0.0014669334050267935)),(to_sfixed_a(0.010191353969275951)),(to_sfixed_a(6.988922541495413e-05)),(to_sfixed_a(-0.00010382058098912239)),(to_sfixed_a(-2.8119618946220726e-05)),(to_sfixed_a(-0.011180880479514599)),(to_sfixed_a(0.0017132567008957267)),(to_sfixed_a(-0.0008560518035665154)),(to_sfixed_a(6.038697756594047e-05)),(to_sfixed_a(-0.012043874710798264)),(to_sfixed_a(-7.932263542898e-06)),(to_sfixed_a(0.00044800102477893233)),(to_sfixed_a(-0.015505341812968254)),(to_sfixed_a(-0.24949093163013458)),(to_sfixed_a(-6.945442146388814e-05)),(to_sfixed_a(0.13869573175907135)),(to_sfixed_a(6.143709470052272e-07)),(to_sfixed_a(0.005985608324408531)),(to_sfixed_a(-0.005544318817555904)),(to_sfixed_a(6.445273174904287e-05)),(to_sfixed_a(0.000380947079975158)),(to_sfixed_a(5.7190605730284005e-05)),(to_sfixed_a(-7.370050298050046e-06)),(to_sfixed_a(2.9248069040477276e-05)),(to_sfixed_a(-9.906617196975276e-05)),(to_sfixed_a(-0.0006869289791211486)),(to_sfixed_a(1.0681786079658195e-05)),(to_sfixed_a(-0.2757294476032257)),(to_sfixed_a(-0.013621974736452103)),(to_sfixed_a(-0.0008953934302553535)),(to_sfixed_a(-0.004083578009158373)),(to_sfixed_a(-1.4795859897276387e-06)),(to_sfixed_a(0.00010237019159831107)),(to_sfixed_a(3.461200321908109e-07)),(to_sfixed_a(-4.8146415792871267e-05)),(to_sfixed_a(-1.931914630404208e-05)),(to_sfixed_a(0.0009724164847284555)),(to_sfixed_a(-0.0023581902496516705)),(to_sfixed_a(-0.01191025786101818)),(to_sfixed_a(5.736401362810284e-07)),(to_sfixed_a(-0.0002475657674949616)),(to_sfixed_a(-6.212925654835999e-06)),(to_sfixed_a(3.555131843313575e-05)),(to_sfixed_a(-0.011907091364264488)),(to_sfixed_a(-0.0084147397428751)),(to_sfixed_a(1.2226424587424845e-05)),(to_sfixed_a(4.2710002162493765e-05)),(to_sfixed_a(0.00011465077113825828)),(to_sfixed_a(-0.014358063228428364)),(to_sfixed_a(0.00018136184371542186)),(to_sfixed_a(-0.005744322203099728)),(to_sfixed_a(4.5258726458996534e-05)),(to_sfixed_a(-0.0001621164265088737)),(to_sfixed_a(4.859694672632031e-05)),(to_sfixed_a(-0.0014314635191112757)),(to_sfixed_a(0.008166924118995667)),(to_sfixed_a(-0.413709431886673)),(to_sfixed_a(8.057919330894947e-06)),(to_sfixed_a(-6.652055162703618e-05)),(to_sfixed_a(-0.00017406800179742277)),(to_sfixed_a(0.00723636569455266)),(to_sfixed_a(3.238863428123295e-05)),(to_sfixed_a(0.45432233810424805)),(to_sfixed_a(2.928900357801467e-06)),(to_sfixed_a(0.19164034724235535)),(to_sfixed_a(0.00043805770110338926)),(to_sfixed_a(-0.01481110043823719)),(to_sfixed_a(0.020470479503273964)),(to_sfixed_a(-1.5499363144044764e-05)),(to_sfixed_a(0.006739207077771425)),(to_sfixed_a(-0.01884254440665245)),(to_sfixed_a(7.083616219460964e-05)),(to_sfixed_a(-0.0012883077142760158)),(to_sfixed_a(2.533665974624455e-05)),(to_sfixed_a(-0.0003380854323040694)),(to_sfixed_a(0.00047088245628401637)),(to_sfixed_a(-0.0033297971822321415)),(to_sfixed_a(-0.00012877979315817356)),(to_sfixed_a(-0.0001933412568178028)),(to_sfixed_a(0.5526950359344482)),(to_sfixed_a(2.941484854090959e-05)),(to_sfixed_a(-0.00783043447881937)),(to_sfixed_a(-0.00017348815163131803)),(to_sfixed_a(-0.00016694342775736004)),(to_sfixed_a(0.00026279804296791553)),(to_sfixed_a(-0.007627794053405523)),(to_sfixed_a(7.721766451140866e-05)),(to_sfixed_a(8.100494596874341e-05)),(to_sfixed_a(-3.307405495434068e-05)),(to_sfixed_a(-0.007530289702117443)),(to_sfixed_a(-0.007068052422255278)),(to_sfixed_a(-2.4341614334844053e-05)),(to_sfixed_a(-8.511693158652633e-05)),(to_sfixed_a(0.0002484761644154787)),(to_sfixed_a(-0.00028180895606055856)),(to_sfixed_a(-0.0007472626166418195)),(to_sfixed_a(-0.02170461229979992)),(to_sfixed_a(-0.26908621191978455)),(to_sfixed_a(-0.01757754012942314)),(to_sfixed_a(0.005180563312023878)),(to_sfixed_a(-8.862659160513431e-05)),(to_sfixed_a(6.283437687670812e-05)),(to_sfixed_a(-2.1284080503392033e-05)),(to_sfixed_a(0.0037360854912549257)),(to_sfixed_a(0.0001020412310026586)),(to_sfixed_a(-0.0001532787282485515)),(to_sfixed_a(0.00011362503573764116)),(to_sfixed_a(-0.0008405059343203902)),(to_sfixed_a(7.93051440268755e-05)),(to_sfixed_a(-3.2910444133449346e-05)),(to_sfixed_a(-0.010471905581653118)),(to_sfixed_a(0.35473039746284485)),(to_sfixed_a(-0.0033310898579657078)),(to_sfixed_a(-4.415983858052641e-05)),(to_sfixed_a(-0.00048095485544763505)),(to_sfixed_a(-0.30551713705062866)),(to_sfixed_a(-0.02391606569290161)),(to_sfixed_a(0.0002902456617448479)),(to_sfixed_a(-0.013418451882898808)),(to_sfixed_a(0.0012001466238871217)),(to_sfixed_a(-0.0036883819848299026)));

    constant weight_n2_12 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.40585261583328247)),(to_sfixed_a(0.600795567035675)),(to_sfixed_a(-0.48606690764427185)),(to_sfixed_a(-6.953245610930026e-05)),(to_sfixed_a(-0.0003021713928319514)),(to_sfixed_a(8.638326107757166e-05)),(to_sfixed_a(0.004615386947989464)),(to_sfixed_a(-0.0003053868131246418)),(to_sfixed_a(7.132633618311957e-05)),(to_sfixed_a(0.00016864814097061753)),(to_sfixed_a(-3.5105185816064477e-06)),(to_sfixed_a(-0.006582219153642654)),(to_sfixed_a(-0.07754028588533401)),(to_sfixed_a(-0.42706140875816345)),(to_sfixed_a(0.00014898748486302793)),(to_sfixed_a(3.703968832269311e-05)),(to_sfixed_a(0.46682968735694885)),(to_sfixed_a(-0.00015260730287991464)),(to_sfixed_a(0.15649963915348053)),(to_sfixed_a(-0.0017279975581914186)),(to_sfixed_a(2.2240194084588438e-05)),(to_sfixed_a(0.00015676161274313927)),(to_sfixed_a(3.372537685208954e-05)),(to_sfixed_a(-0.004254210740327835)),(to_sfixed_a(0.3684205114841461)),(to_sfixed_a(0.21797776222229004)),(to_sfixed_a(-6.347343150991946e-05)),(to_sfixed_a(0.0009260649676434696)),(to_sfixed_a(-0.0007475949823856354)),(to_sfixed_a(0.00010559678776189685)),(to_sfixed_a(0.004045078065246344)),(to_sfixed_a(-0.0002426103310426697)),(to_sfixed_a(-0.6845139265060425)),(to_sfixed_a(-6.787203892599791e-05)),(to_sfixed_a(0.00018136932339984924)),(to_sfixed_a(-0.0001760096929501742)),(to_sfixed_a(-0.023780403658747673)),(to_sfixed_a(0.00883009284734726)),(to_sfixed_a(-0.38881149888038635)),(to_sfixed_a(-0.00010681113053578883)),(to_sfixed_a(-0.5210239887237549)),(to_sfixed_a(-0.31851741671562195)),(to_sfixed_a(-0.0004179569659754634)),(to_sfixed_a(-0.00010855669825104997)),(to_sfixed_a(0.002848181640729308)),(to_sfixed_a(0.02369631454348564)),(to_sfixed_a(0.44619089365005493)),(to_sfixed_a(0.015627309679985046)),(to_sfixed_a(-7.737287523923442e-05)),(to_sfixed_a(0.003320542396977544)),(to_sfixed_a(-0.013255195692181587)),(to_sfixed_a(-0.0006742958794347942)),(to_sfixed_a(0.00015321349201258272)),(to_sfixed_a(0.0029202650766819715)),(to_sfixed_a(-0.018490198999643326)),(to_sfixed_a(0.007480276748538017)),(to_sfixed_a(0.00011590298527153209)),(to_sfixed_a(0.01044733077287674)),(to_sfixed_a(-0.0001817680458771065)),(to_sfixed_a(1.9371334929019213e-05)),(to_sfixed_a(0.007662413641810417)),(to_sfixed_a(-0.0005214574048295617)),(to_sfixed_a(-0.004575781989842653)),(to_sfixed_a(-0.0013151605380699039)),(to_sfixed_a(8.885755960363895e-06)),(to_sfixed_a(-0.3755348324775696)),(to_sfixed_a(-0.00045088317710906267)),(to_sfixed_a(-0.0018535088747739792)),(to_sfixed_a(0.0038808444514870644)),(to_sfixed_a(-6.945841596461833e-05)),(to_sfixed_a(0.17331528663635254)),(to_sfixed_a(-0.008146069012582302)),(to_sfixed_a(0.007134099490940571)),(to_sfixed_a(6.295504863373935e-05)),(to_sfixed_a(1.5553632692899555e-06)),(to_sfixed_a(4.69888182124123e-05)),(to_sfixed_a(0.2003687024116516)),(to_sfixed_a(0.0016200818354263902)),(to_sfixed_a(0.00016580696683377028)),(to_sfixed_a(-0.008214340545237064)),(to_sfixed_a(0.009128699079155922)),(to_sfixed_a(0.0001507025008322671)),(to_sfixed_a(0.08003903180360794)),(to_sfixed_a(0.0024623158387839794)),(to_sfixed_a(5.919524119235575e-05)),(to_sfixed_a(0.010210679844021797)),(to_sfixed_a(0.25962257385253906)),(to_sfixed_a(-3.5805605875793844e-05)),(to_sfixed_a(0.00011381376680219546)),(to_sfixed_a(-0.0001493364106863737)),(to_sfixed_a(-0.0026372517459094524)),(to_sfixed_a(-0.00012968419468961656)),(to_sfixed_a(0.01890014484524727)),(to_sfixed_a(-6.344428402371705e-05)),(to_sfixed_a(0.0002468561287969351)),(to_sfixed_a(0.00019971052824985236)),(to_sfixed_a(0.00012616634194273502)),(to_sfixed_a(0.0001302410673815757)),(to_sfixed_a(-3.7087855162099004e-05)),(to_sfixed_a(0.00014954085054341704)),(to_sfixed_a(-0.0010572189930826426)),(to_sfixed_a(0.0043642898090183735)),(to_sfixed_a(-4.834109859075397e-05)),(to_sfixed_a(0.004197047557681799)),(to_sfixed_a(0.12932147085666656)),(to_sfixed_a(0.0006025195471011102)),(to_sfixed_a(-0.00011386041296645999)),(to_sfixed_a(-3.911305248038843e-05)),(to_sfixed_a(-0.00011304221698082983)),(to_sfixed_a(0.010015299543738365)),(to_sfixed_a(0.002706627594307065)),(to_sfixed_a(-1.0479277989361435e-05)),(to_sfixed_a(0.09112495183944702)),(to_sfixed_a(-2.5578527129255235e-05)),(to_sfixed_a(2.0784927983186208e-05)),(to_sfixed_a(-0.34461894631385803)),(to_sfixed_a(0.0009193719015456736)),(to_sfixed_a(-0.07852928340435028)),(to_sfixed_a(0.0001836760202422738)),(to_sfixed_a(-0.00010164048580918461)),(to_sfixed_a(-0.00011335039744153619)),(to_sfixed_a(-4.389679088490084e-05)),(to_sfixed_a(-0.0012147420784458518)),(to_sfixed_a(-0.00010666513117030263)),(to_sfixed_a(-4.0402504964731634e-05)),(to_sfixed_a(-0.15669961273670197)),(to_sfixed_a(-0.014512860216200352)),(to_sfixed_a(-1.0613453923724592e-05)),(to_sfixed_a(-0.00012280227383598685)),(to_sfixed_a(3.239096258766949e-06)),(to_sfixed_a(-9.8830321803689e-05)),(to_sfixed_a(-6.330880569294095e-05)),(to_sfixed_a(0.001953922212123871)),(to_sfixed_a(0.18132638931274414)),(to_sfixed_a(0.00023707406944595277)),(to_sfixed_a(-0.00011517070379341021)),(to_sfixed_a(-0.0003442729648668319)),(to_sfixed_a(0.000932325201574713)),(to_sfixed_a(6.777551607228816e-05)),(to_sfixed_a(6.920152372913435e-05)),(to_sfixed_a(0.008030898869037628)),(to_sfixed_a(-0.00011339453340042382)),(to_sfixed_a(-0.00018332593026570976)),(to_sfixed_a(0.0001086320262402296)),(to_sfixed_a(0.543647825717926)),(to_sfixed_a(3.0511808290611953e-05)),(to_sfixed_a(-0.3002704381942749)),(to_sfixed_a(0.00013725752069149166)),(to_sfixed_a(3.531749825924635e-08)),(to_sfixed_a(0.0010124273831024766)),(to_sfixed_a(2.8840913728345186e-05)),(to_sfixed_a(-3.824878513114527e-05)),(to_sfixed_a(0.0010099239880219102)),(to_sfixed_a(0.0001273973612114787)),(to_sfixed_a(5.71652090002317e-05)),(to_sfixed_a(-0.0010933935409411788)),(to_sfixed_a(-6.709150329697877e-05)),(to_sfixed_a(-0.3733599781990051)),(to_sfixed_a(-9.379560651723295e-05)),(to_sfixed_a(-0.00022720370907336473)),(to_sfixed_a(0.00022854826238472015)),(to_sfixed_a(-0.0001688599877525121)),(to_sfixed_a(-0.006124892737716436)),(to_sfixed_a(-0.01964048482477665)),(to_sfixed_a(-0.0014487130101770163)),(to_sfixed_a(0.0008183233439922333)),(to_sfixed_a(8.575202082283795e-05)),(to_sfixed_a(0.005528447218239307)),(to_sfixed_a(2.0811723516089842e-05)),(to_sfixed_a(2.8441805625334382e-05)),(to_sfixed_a(-0.16742616891860962)),(to_sfixed_a(0.02288517914712429)),(to_sfixed_a(-0.006300035398453474)),(to_sfixed_a(-0.00014045272837392986)),(to_sfixed_a(0.08722030371427536)),(to_sfixed_a(-0.18940049409866333)),(to_sfixed_a(0.0012620416237041354)),(to_sfixed_a(0.1933874487876892)),(to_sfixed_a(0.011742636561393738)),(to_sfixed_a(0.25948309898376465)),(to_sfixed_a(-0.25339049100875854)),(to_sfixed_a(-0.14812703430652618)),(to_sfixed_a(1.1485477443784475e-05)),(to_sfixed_a(0.00031066752853803337)),(to_sfixed_a(4.4957134377909824e-05)),(to_sfixed_a(-0.07427316159009933)),(to_sfixed_a(-0.0046043675392866135)),(to_sfixed_a(-0.004172202665358782)),(to_sfixed_a(-0.006981961894780397)),(to_sfixed_a(-0.007878350093960762)),(to_sfixed_a(-0.2730509042739868)),(to_sfixed_a(-0.00012789903848897666)),(to_sfixed_a(-0.14295214414596558)),(to_sfixed_a(0.0098910853266716)),(to_sfixed_a(8.84009205037728e-05)),(to_sfixed_a(0.2993720471858978)),(to_sfixed_a(0.00011244531197007746)),(to_sfixed_a(0.0009442534064874053)),(to_sfixed_a(0.11616871505975723)),(to_sfixed_a(1.1725045624189079e-05)),(to_sfixed_a(-1.0263771400786936e-05)),(to_sfixed_a(-0.00017510098405182362)),(to_sfixed_a(0.00024295708863064647)),(to_sfixed_a(3.663240931928158e-05)),(to_sfixed_a(0.00013031705748289824)),(to_sfixed_a(0.29717880487442017)),(to_sfixed_a(0.3251807987689972)),(to_sfixed_a(-0.580836832523346)),(to_sfixed_a(-0.0009308477165177464)),(to_sfixed_a(-0.0016686295857653022)),(to_sfixed_a(-0.09662081301212311)),(to_sfixed_a(8.48563649924472e-06)),(to_sfixed_a(-0.00020488524751272053)),(to_sfixed_a(5.2891009545419365e-05)),(to_sfixed_a(0.00021754649060312659)),(to_sfixed_a(-3.3665637602098286e-05)),(to_sfixed_a(-0.43708157539367676)),(to_sfixed_a(-0.002078382298350334)),(to_sfixed_a(0.004692496731877327)),(to_sfixed_a(-3.0083643650868908e-05)),(to_sfixed_a(-0.0001202266284963116)),(to_sfixed_a(-0.00013669926556758583)),(to_sfixed_a(-0.00025483634090051055)),(to_sfixed_a(0.007975934073328972)),(to_sfixed_a(0.5229803323745728)),(to_sfixed_a(7.127896242309362e-05)),(to_sfixed_a(-2.1605439542327076e-05)),(to_sfixed_a(-9.743117698235437e-05)),(to_sfixed_a(0.30600422620773315)),(to_sfixed_a(-0.21941572427749634)),(to_sfixed_a(0.271657258272171)),(to_sfixed_a(-4.858018655795604e-06)),(to_sfixed_a(-0.00018522579921409488)),(to_sfixed_a(8.535238157492131e-05)),(to_sfixed_a(-0.0008415286429226398)),(to_sfixed_a(0.014405162073671818)),(to_sfixed_a(0.0017480857204645872)),(to_sfixed_a(1.3646407751366496e-05)),(to_sfixed_a(-0.002603710163384676)),(to_sfixed_a(0.00018046112381853163)),(to_sfixed_a(-0.0024902422446757555)),(to_sfixed_a(-0.00019933281873818487)),(to_sfixed_a(-0.0005220880266278982)),(to_sfixed_a(7.285900937858969e-05)),(to_sfixed_a(-0.3785243332386017)),(to_sfixed_a(-0.0056589446030557156)),(to_sfixed_a(0.5960302948951721)),(to_sfixed_a(0.009223350323736668)),(to_sfixed_a(-7.219485996756703e-05)),(to_sfixed_a(0.005861023440957069)),(to_sfixed_a(0.010549547150731087)),(to_sfixed_a(3.0863782740198076e-05)),(to_sfixed_a(-7.060520874802023e-05)),(to_sfixed_a(0.00013983127428218722)),(to_sfixed_a(0.0001845531805884093)),(to_sfixed_a(0.28243589401245117)),(to_sfixed_a(-0.5840291976928711)),(to_sfixed_a(0.00010994624608429149)),(to_sfixed_a(0.0001697651023278013)),(to_sfixed_a(0.256790429353714)),(to_sfixed_a(-0.00015704860561527312)),(to_sfixed_a(-0.0034476725850254297)),(to_sfixed_a(4.802032344741747e-05)),(to_sfixed_a(-0.0011037465883418918)),(to_sfixed_a(0.00014693092089146376)),(to_sfixed_a(-0.595452070236206)),(to_sfixed_a(-3.0031587812118232e-06)),(to_sfixed_a(0.0003138228494208306)),(to_sfixed_a(-3.058053334825672e-05)),(to_sfixed_a(0.28123530745506287)),(to_sfixed_a(0.006000157445669174)),(to_sfixed_a(-0.00019921304192394018)),(to_sfixed_a(3.531230322550982e-05)),(to_sfixed_a(0.00024250928254332393)),(to_sfixed_a(-2.207777288276702e-05)),(to_sfixed_a(0.00046514460700564086)),(to_sfixed_a(9.158419561572373e-05)),(to_sfixed_a(0.0015266406117007136)),(to_sfixed_a(0.23665864765644073)),(to_sfixed_a(0.02000284381210804)),(to_sfixed_a(0.00012058186257490888)),(to_sfixed_a(-6.421994476113468e-05)),(to_sfixed_a(1.0260220733471215e-05)),(to_sfixed_a(-0.3878748118877411)),(to_sfixed_a(6.947708607185632e-05)),(to_sfixed_a(2.4905446480261162e-05)),(to_sfixed_a(0.0009216985199600458)),(to_sfixed_a(-0.0014584949240088463)),(to_sfixed_a(-0.0003124900977127254)),(to_sfixed_a(0.5632117390632629)),(to_sfixed_a(-0.00033019750844687223)),(to_sfixed_a(0.008293000981211662)),(to_sfixed_a(-0.002905695466324687)),(to_sfixed_a(-6.316658982541412e-07)),(to_sfixed_a(-0.03564926236867905)),(to_sfixed_a(0.3766935169696808)),(to_sfixed_a(0.010967717505991459)),(to_sfixed_a(0.0001160369865829125)),(to_sfixed_a(3.379493864485994e-05)),(to_sfixed_a(0.004900223575532436)),(to_sfixed_a(0.006636017467826605)));

    constant weight_n2_13 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.5238252282142639)),(to_sfixed_a(0.010357297025620937)),(to_sfixed_a(-0.0003310128813609481)),(to_sfixed_a(-6.503918120870367e-05)),(to_sfixed_a(-0.002654639072716236)),(to_sfixed_a(-0.00013034531730227172)),(to_sfixed_a(0.16846303641796112)),(to_sfixed_a(-0.00013488769764080644)),(to_sfixed_a(0.00015443415031768382)),(to_sfixed_a(-6.900400330778211e-05)),(to_sfixed_a(3.775634468183853e-05)),(to_sfixed_a(-0.006926975212991238)),(to_sfixed_a(-0.000830307079013437)),(to_sfixed_a(0.0037071185652166605)),(to_sfixed_a(8.353278826689348e-05)),(to_sfixed_a(-2.6883601094596088e-05)),(to_sfixed_a(0.003990273457020521)),(to_sfixed_a(6.452937668655068e-06)),(to_sfixed_a(0.008178907446563244)),(to_sfixed_a(7.227614696603268e-05)),(to_sfixed_a(0.0001058827547240071)),(to_sfixed_a(-5.51971243112348e-06)),(to_sfixed_a(-0.002029085299000144)),(to_sfixed_a(5.474123827298172e-05)),(to_sfixed_a(0.004531010054051876)),(to_sfixed_a(0.0070033264346420765)),(to_sfixed_a(-0.00018153806740883738)),(to_sfixed_a(-0.0001996292849071324)),(to_sfixed_a(0.00011432907194830477)),(to_sfixed_a(0.00012931630772072822)),(to_sfixed_a(-0.0032295798882842064)),(to_sfixed_a(-0.00013970246072858572)),(to_sfixed_a(-0.0018357469234615564)),(to_sfixed_a(0.00011375157191650942)),(to_sfixed_a(1.514170435257256e-05)),(to_sfixed_a(0.00028959399787709117)),(to_sfixed_a(0.025167370215058327)),(to_sfixed_a(-0.27635619044303894)),(to_sfixed_a(-0.00753041822463274)),(to_sfixed_a(-0.00016218838572967798)),(to_sfixed_a(1.8252147128805518e-05)),(to_sfixed_a(0.001832912559621036)),(to_sfixed_a(-0.0001592871849425137)),(to_sfixed_a(2.0234656403772533e-06)),(to_sfixed_a(-0.0008067355956882238)),(to_sfixed_a(-0.00889548659324646)),(to_sfixed_a(0.003512484487146139)),(to_sfixed_a(-0.0007672765059396625)),(to_sfixed_a(-0.0002165738114854321)),(to_sfixed_a(-0.0010382587788626552)),(to_sfixed_a(0.0074837650172412395)),(to_sfixed_a(0.0019790134392678738)),(to_sfixed_a(9.84547077678144e-05)),(to_sfixed_a(0.006150225643068552)),(to_sfixed_a(-0.3442831039428711)),(to_sfixed_a(-0.007324254605919123)),(to_sfixed_a(0.00015248646377585828)),(to_sfixed_a(-0.01616857573390007)),(to_sfixed_a(6.709409353788942e-05)),(to_sfixed_a(-6.800427217967808e-05)),(to_sfixed_a(-0.004304929170757532)),(to_sfixed_a(-0.00523677933961153)),(to_sfixed_a(-0.0008198339492082596)),(to_sfixed_a(0.005005707032978535)),(to_sfixed_a(-0.00020446820417419076)),(to_sfixed_a(0.0026550767943263054)),(to_sfixed_a(0.00011302067287033424)),(to_sfixed_a(0.00018571733380667865)),(to_sfixed_a(-0.012922825291752815)),(to_sfixed_a(-0.00015729745791759342)),(to_sfixed_a(-0.0045265029184520245)),(to_sfixed_a(-0.007532894145697355)),(to_sfixed_a(0.009387992322444916)),(to_sfixed_a(-7.56367517169565e-05)),(to_sfixed_a(5.7516153901815414e-06)),(to_sfixed_a(-0.00011254558921791613)),(to_sfixed_a(-0.011834230273962021)),(to_sfixed_a(-0.01301883440464735)),(to_sfixed_a(-0.00010090431169373915)),(to_sfixed_a(0.020108668133616447)),(to_sfixed_a(0.44375476241111755)),(to_sfixed_a(0.00012069346848875284)),(to_sfixed_a(-0.0004978433717042208)),(to_sfixed_a(0.011859351769089699)),(to_sfixed_a(7.248221663758159e-05)),(to_sfixed_a(-0.0012073577381670475)),(to_sfixed_a(0.0009034264367073774)),(to_sfixed_a(0.0002736399765126407)),(to_sfixed_a(0.00018522009486332536)),(to_sfixed_a(-0.0001814570277929306)),(to_sfixed_a(-0.011334181763231754)),(to_sfixed_a(-0.00041361074545420706)),(to_sfixed_a(-0.010736110620200634)),(to_sfixed_a(0.00018521473975852132)),(to_sfixed_a(-0.005533652845770121)),(to_sfixed_a(-3.5299541195854545e-05)),(to_sfixed_a(8.565696043660864e-05)),(to_sfixed_a(-0.00013778785069007427)),(to_sfixed_a(0.00030398089438676834)),(to_sfixed_a(-7.948598795337602e-05)),(to_sfixed_a(0.000670638051815331)),(to_sfixed_a(-0.4461626708507538)),(to_sfixed_a(2.358078199904412e-05)),(to_sfixed_a(-0.012911435216665268)),(to_sfixed_a(-0.007655662950128317)),(to_sfixed_a(-0.00019145131227560341)),(to_sfixed_a(0.00015125516802072525)),(to_sfixed_a(6.395841046469286e-05)),(to_sfixed_a(2.7957081329077482e-05)),(to_sfixed_a(0.23262979090213776)),(to_sfixed_a(-0.0007540748338215053)),(to_sfixed_a(-8.43236266518943e-05)),(to_sfixed_a(-0.0016314227832481265)),(to_sfixed_a(0.00020666354976128787)),(to_sfixed_a(0.00017783672956284136)),(to_sfixed_a(-0.018160466104745865)),(to_sfixed_a(0.0001324202457908541)),(to_sfixed_a(-0.0061248550191521645)),(to_sfixed_a(0.00031139751081354916)),(to_sfixed_a(-0.28227293491363525)),(to_sfixed_a(0.00015031720977276564)),(to_sfixed_a(0.0001337225694442168)),(to_sfixed_a(-0.005061212461441755)),(to_sfixed_a(-5.114157102070749e-05)),(to_sfixed_a(-8.089029870461673e-05)),(to_sfixed_a(-0.28487828373908997)),(to_sfixed_a(0.007306961342692375)),(to_sfixed_a(-3.470828232821077e-06)),(to_sfixed_a(-7.033161091385409e-05)),(to_sfixed_a(0.0001789951929822564)),(to_sfixed_a(-2.1196159650571644e-05)),(to_sfixed_a(-0.0002899133542086929)),(to_sfixed_a(0.005787003319710493)),(to_sfixed_a(-0.016311777755618095)),(to_sfixed_a(-3.214333264622837e-05)),(to_sfixed_a(0.0002887581940740347)),(to_sfixed_a(-0.018224872648715973)),(to_sfixed_a(0.00016326358309015632)),(to_sfixed_a(6.753380876034498e-05)),(to_sfixed_a(0.0001345719792880118)),(to_sfixed_a(-0.007552043534815311)),(to_sfixed_a(-9.55604191403836e-05)),(to_sfixed_a(0.0001415625592926517)),(to_sfixed_a(1.7014550394378603e-05)),(to_sfixed_a(0.004849139600992203)),(to_sfixed_a(0.00026681445888243616)),(to_sfixed_a(-0.0003008561616297811)),(to_sfixed_a(5.647896614391357e-05)),(to_sfixed_a(0.0002548657066654414)),(to_sfixed_a(-0.0004119104123674333)),(to_sfixed_a(-0.0001025134333758615)),(to_sfixed_a(-0.00017809182463679463)),(to_sfixed_a(-0.0034015255514532328)),(to_sfixed_a(0.00010493420995771885)),(to_sfixed_a(-6.892788223922253e-05)),(to_sfixed_a(0.006130078341811895)),(to_sfixed_a(-9.543449414195493e-05)),(to_sfixed_a(-0.0007443799986504018)),(to_sfixed_a(-9.001742000691593e-06)),(to_sfixed_a(0.00030474961386062205)),(to_sfixed_a(2.420904638711363e-05)),(to_sfixed_a(-9.465882612857968e-06)),(to_sfixed_a(0.007888446561992168)),(to_sfixed_a(0.005028934683650732)),(to_sfixed_a(-0.0009270609589293599)),(to_sfixed_a(0.0008994921809062362)),(to_sfixed_a(4.315773185226135e-05)),(to_sfixed_a(-0.0054097771644592285)),(to_sfixed_a(-0.00015055641415528953)),(to_sfixed_a(-2.061135819531046e-05)),(to_sfixed_a(0.012112430296838284)),(to_sfixed_a(0.0033973813988268375)),(to_sfixed_a(0.002942791674286127)),(to_sfixed_a(3.125561124761589e-05)),(to_sfixed_a(0.0007742050802335143)),(to_sfixed_a(-7.236737292259932e-05)),(to_sfixed_a(-0.003080653492361307)),(to_sfixed_a(-0.716934084892273)),(to_sfixed_a(-0.012548149563372135)),(to_sfixed_a(-0.36767929792404175)),(to_sfixed_a(-8.874121704138815e-07)),(to_sfixed_a(0.0016231425106525421)),(to_sfixed_a(-9.861049329629168e-05)),(to_sfixed_a(0.00011568234185688198)),(to_sfixed_a(-0.00011330650886520743)),(to_sfixed_a(0.00043057918082922697)),(to_sfixed_a(0.005421456415206194)),(to_sfixed_a(-5.497210077010095e-05)),(to_sfixed_a(0.0030572013929486275)),(to_sfixed_a(0.006178179290145636)),(to_sfixed_a(0.0049566058441996574)),(to_sfixed_a(0.0001765280612744391)),(to_sfixed_a(-0.26543429493904114)),(to_sfixed_a(-0.004742820747196674)),(to_sfixed_a(0.00015325326239690185)),(to_sfixed_a(-0.493932843208313)),(to_sfixed_a(-0.00015166675439104438)),(to_sfixed_a(0.0034772700164467096)),(to_sfixed_a(0.001298836199566722)),(to_sfixed_a(3.809058398474008e-05)),(to_sfixed_a(-0.00014610824291594326)),(to_sfixed_a(5.7605328038334846e-05)),(to_sfixed_a(-0.00016618492372799665)),(to_sfixed_a(3.1740015401737764e-05)),(to_sfixed_a(-3.897592250723392e-05)),(to_sfixed_a(0.003549461718648672)),(to_sfixed_a(0.0019198363879695535)),(to_sfixed_a(-0.002252083970233798)),(to_sfixed_a(6.053813558537513e-05)),(to_sfixed_a(0.21327205002307892)),(to_sfixed_a(-0.014472379349172115)),(to_sfixed_a(-7.36637448426336e-05)),(to_sfixed_a(5.025372956879437e-06)),(to_sfixed_a(-0.00012972524564247578)),(to_sfixed_a(4.02827572543174e-06)),(to_sfixed_a(-5.618199793389067e-05)),(to_sfixed_a(0.0016714967787265778)),(to_sfixed_a(6.316610961221159e-05)),(to_sfixed_a(0.0003609294362831861)),(to_sfixed_a(4.336690835771151e-05)),(to_sfixed_a(-0.00018485421605873853)),(to_sfixed_a(-8.264565258286893e-05)),(to_sfixed_a(-0.00011346388055244461)),(to_sfixed_a(-0.0030959094874560833)),(to_sfixed_a(-0.0071101621724665165)),(to_sfixed_a(-6.89957378199324e-05)),(to_sfixed_a(-5.811134906252846e-05)),(to_sfixed_a(-6.739106174791232e-05)),(to_sfixed_a(-0.012692630290985107)),(to_sfixed_a(-0.01097177155315876)),(to_sfixed_a(0.0015716170892119408)),(to_sfixed_a(2.4820521502988413e-05)),(to_sfixed_a(3.0461895221378654e-05)),(to_sfixed_a(-3.702522371895611e-05)),(to_sfixed_a(-0.0038973428308963776)),(to_sfixed_a(-0.004180393181741238)),(to_sfixed_a(0.4823456406593323)),(to_sfixed_a(-9.745999705046415e-07)),(to_sfixed_a(0.002224898198619485)),(to_sfixed_a(-0.00018572993576526642)),(to_sfixed_a(0.005246516317129135)),(to_sfixed_a(0.0001166627262136899)),(to_sfixed_a(-0.1596403568983078)),(to_sfixed_a(-4.265975803718902e-05)),(to_sfixed_a(0.006120894104242325)),(to_sfixed_a(0.25620582699775696)),(to_sfixed_a(-0.005021102260798216)),(to_sfixed_a(0.508185625076294)),(to_sfixed_a(0.00018007932521868497)),(to_sfixed_a(-0.009750527329742908)),(to_sfixed_a(-0.002299812389537692)),(to_sfixed_a(-1.0017429303843528e-05)),(to_sfixed_a(0.0022403248585760593)),(to_sfixed_a(4.096011252840981e-05)),(to_sfixed_a(0.00011400782386772335)),(to_sfixed_a(-0.0010166154243052006)),(to_sfixed_a(0.003487295238301158)),(to_sfixed_a(-3.817454125965014e-05)),(to_sfixed_a(-6.748914893250912e-05)),(to_sfixed_a(-0.41885796189308167)),(to_sfixed_a(-6.504606426460668e-05)),(to_sfixed_a(0.0009369384497404099)),(to_sfixed_a(0.0001043175725499168)),(to_sfixed_a(3.594240843085572e-05)),(to_sfixed_a(-9.013756061904132e-05)),(to_sfixed_a(0.0037229880690574646)),(to_sfixed_a(-0.00010969342110911384)),(to_sfixed_a(-2.7539863367564976e-06)),(to_sfixed_a(8.873119077179581e-05)),(to_sfixed_a(0.003759081242606044)),(to_sfixed_a(-0.0007412026170641184)),(to_sfixed_a(-0.00024668662808835506)),(to_sfixed_a(-0.00020140144624747336)),(to_sfixed_a(0.0001642286079004407)),(to_sfixed_a(5.684298230335116e-06)),(to_sfixed_a(-0.11520011723041534)),(to_sfixed_a(-0.0005669803358614445)),(to_sfixed_a(-0.14644402265548706)),(to_sfixed_a(0.2777000069618225)),(to_sfixed_a(0.007551173679530621)),(to_sfixed_a(-0.00016982411034405231)),(to_sfixed_a(3.884374018525705e-05)),(to_sfixed_a(-0.0001788845402188599)),(to_sfixed_a(0.0002946997410617769)),(to_sfixed_a(-3.733820267370902e-05)),(to_sfixed_a(3.4177421184722334e-05)),(to_sfixed_a(-0.008767357096076012)),(to_sfixed_a(0.03549491986632347)),(to_sfixed_a(-0.000196041029994376)),(to_sfixed_a(0.00019631037139333785)),(to_sfixed_a(8.587019692640752e-06)),(to_sfixed_a(1.4969438780099154e-05)),(to_sfixed_a(0.08988982439041138)),(to_sfixed_a(6.224487151484936e-05)),(to_sfixed_a(0.5029172897338867)),(to_sfixed_a(-1.9122910089208744e-05)),(to_sfixed_a(-0.005622821394354105)),(to_sfixed_a(6.879685679450631e-05)),(to_sfixed_a(-0.012384389527142048)),(to_sfixed_a(-0.0030262176878750324)),(to_sfixed_a(-0.0066448114812374115)));

    constant weight_n2_14 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.06272605061531067)),(to_sfixed_a(-0.007951456122100353)),(to_sfixed_a(0.0003618642804212868)),(to_sfixed_a(-5.4501870181411505e-06)),(to_sfixed_a(4.601806358550675e-05)),(to_sfixed_a(0.00015635957242920995)),(to_sfixed_a(0.0023001760710030794)),(to_sfixed_a(2.7939186111325398e-05)),(to_sfixed_a(-2.3572603822685778e-05)),(to_sfixed_a(-4.122659447602928e-06)),(to_sfixed_a(0.0001755812845658511)),(to_sfixed_a(0.002627369947731495)),(to_sfixed_a(-0.0007232199423015118)),(to_sfixed_a(-0.0066957902163267136)),(to_sfixed_a(0.00015611553681083024)),(to_sfixed_a(2.4701635993551463e-05)),(to_sfixed_a(-0.004423891194164753)),(to_sfixed_a(-5.8893019740935415e-05)),(to_sfixed_a(-0.007733006030321121)),(to_sfixed_a(0.0009189262636937201)),(to_sfixed_a(3.3679389161989093e-06)),(to_sfixed_a(0.00011205598275410011)),(to_sfixed_a(0.002277674851939082)),(to_sfixed_a(0.2357354611158371)),(to_sfixed_a(0.003381588961929083)),(to_sfixed_a(-0.008698035962879658)),(to_sfixed_a(7.158234075177461e-05)),(to_sfixed_a(4.167430961388163e-05)),(to_sfixed_a(6.286051939241588e-05)),(to_sfixed_a(-6.767808372387663e-05)),(to_sfixed_a(0.005140426103025675)),(to_sfixed_a(-3.4450713428668678e-06)),(to_sfixed_a(0.0010151696624234319)),(to_sfixed_a(2.406747080385685e-05)),(to_sfixed_a(-7.008848479017615e-05)),(to_sfixed_a(1.0947842383757234e-05)),(to_sfixed_a(-0.12243378162384033)),(to_sfixed_a(0.35514554381370544)),(to_sfixed_a(-0.01097537949681282)),(to_sfixed_a(-0.00012031092046527192)),(to_sfixed_a(0.005474044010043144)),(to_sfixed_a(-0.0015441421419382095)),(to_sfixed_a(0.00011926997103728354)),(to_sfixed_a(4.165558493696153e-06)),(to_sfixed_a(0.007968412712216377)),(to_sfixed_a(0.011608107946813107)),(to_sfixed_a(-0.5405461192131042)),(to_sfixed_a(0.0011266039218753576)),(to_sfixed_a(-0.0002866168797481805)),(to_sfixed_a(0.002474614419043064)),(to_sfixed_a(0.4891692101955414)),(to_sfixed_a(-0.0074685681611299515)),(to_sfixed_a(-0.00021861903951503336)),(to_sfixed_a(-0.0002530104829929769)),(to_sfixed_a(0.0112720662727952)),(to_sfixed_a(-0.03983454406261444)),(to_sfixed_a(2.4412558559561148e-05)),(to_sfixed_a(0.007212101481854916)),(to_sfixed_a(5.966332901152782e-05)),(to_sfixed_a(-0.00022228692250791937)),(to_sfixed_a(0.004113370086997747)),(to_sfixed_a(0.004594370722770691)),(to_sfixed_a(-0.004352455027401447)),(to_sfixed_a(0.00018008827464655042)),(to_sfixed_a(-7.047048711683601e-05)),(to_sfixed_a(-0.21845762431621552)),(to_sfixed_a(-3.206266774213873e-05)),(to_sfixed_a(-0.004303992725908756)),(to_sfixed_a(3.952115366701037e-05)),(to_sfixed_a(0.0001680465938989073)),(to_sfixed_a(-0.002850044285878539)),(to_sfixed_a(-0.017251942306756973)),(to_sfixed_a(0.01128364633768797)),(to_sfixed_a(-2.9562870622612536e-05)),(to_sfixed_a(4.486877878662199e-05)),(to_sfixed_a(-6.47413544356823e-05)),(to_sfixed_a(0.18175949156284332)),(to_sfixed_a(0.002217178698629141)),(to_sfixed_a(-2.5361310690641403e-05)),(to_sfixed_a(-0.02062908560037613)),(to_sfixed_a(0.005070211365818977)),(to_sfixed_a(0.0001564965641591698)),(to_sfixed_a(-0.2258087396621704)),(to_sfixed_a(-0.0039145126938819885)),(to_sfixed_a(-9.484865586273372e-07)),(to_sfixed_a(0.0007597270305268466)),(to_sfixed_a(-0.005254553165286779)),(to_sfixed_a(0.5423086285591125)),(to_sfixed_a(-3.344528886373155e-05)),(to_sfixed_a(-0.00018540235760156065)),(to_sfixed_a(-0.0034834847319871187)),(to_sfixed_a(1.888825499918312e-05)),(to_sfixed_a(0.006146858911961317)),(to_sfixed_a(-3.749656752916053e-05)),(to_sfixed_a(-0.21791081130504608)),(to_sfixed_a(2.708401734707877e-05)),(to_sfixed_a(-1.0253628715872765e-05)),(to_sfixed_a(-0.00013586845307145268)),(to_sfixed_a(9.841436985880136e-05)),(to_sfixed_a(-9.365916412207298e-06)),(to_sfixed_a(0.0024143042974174023)),(to_sfixed_a(0.37779903411865234)),(to_sfixed_a(-2.467540616635233e-05)),(to_sfixed_a(0.011443994008004665)),(to_sfixed_a(-0.004134316463023424)),(to_sfixed_a(0.3401033580303192)),(to_sfixed_a(0.0002757097245194018)),(to_sfixed_a(2.6226109184790403e-05)),(to_sfixed_a(-4.3271757022012025e-05)),(to_sfixed_a(0.002276081359013915)),(to_sfixed_a(0.0028213253244757652)),(to_sfixed_a(-0.00029079726664349437)),(to_sfixed_a(0.0013335959520190954)),(to_sfixed_a(-0.0002509331679902971)),(to_sfixed_a(-8.544888987671584e-05)),(to_sfixed_a(0.003855412593111396)),(to_sfixed_a(0.2288137823343277)),(to_sfixed_a(0.0006118654273450375)),(to_sfixed_a(-7.261321297846735e-05)),(to_sfixed_a(0.3696531653404236)),(to_sfixed_a(7.689397898502648e-05)),(to_sfixed_a(0.00026319059543311596)),(to_sfixed_a(0.0035170570481568575)),(to_sfixed_a(0.0001686663890723139)),(to_sfixed_a(0.0003815142554230988)),(to_sfixed_a(0.0026166357565671206)),(to_sfixed_a(-0.003226728178560734)),(to_sfixed_a(-1.9661994883790612e-05)),(to_sfixed_a(2.1643354557454586e-06)),(to_sfixed_a(6.755096546839923e-05)),(to_sfixed_a(4.736168193630874e-06)),(to_sfixed_a(0.00028719374677166343)),(to_sfixed_a(-0.006428443361073732)),(to_sfixed_a(0.003216577460989356)),(to_sfixed_a(0.0003101015172433108)),(to_sfixed_a(-6.724553531967103e-05)),(to_sfixed_a(0.32954663038253784)),(to_sfixed_a(0.0004507392586674541)),(to_sfixed_a(-0.00012413891090545803)),(to_sfixed_a(-0.00023847899865359068)),(to_sfixed_a(0.0006517450674436986)),(to_sfixed_a(-3.472770913504064e-06)),(to_sfixed_a(-7.919488416519016e-05)),(to_sfixed_a(1.7384874809067696e-05)),(to_sfixed_a(-0.008265173062682152)),(to_sfixed_a(-6.72757305437699e-05)),(to_sfixed_a(0.00027442246209830046)),(to_sfixed_a(0.00013034594303462654)),(to_sfixed_a(0.0002490238402970135)),(to_sfixed_a(-0.008735350333154202)),(to_sfixed_a(-2.541405410738662e-05)),(to_sfixed_a(0.00013621276593767107)),(to_sfixed_a(0.0006804278818890452)),(to_sfixed_a(1.7633326933719218e-05)),(to_sfixed_a(-7.861004996811971e-05)),(to_sfixed_a(0.11578168720006943)),(to_sfixed_a(-0.00022202072432264686)),(to_sfixed_a(0.39508044719696045)),(to_sfixed_a(0.00022775978140998632)),(to_sfixed_a(-9.783829591469839e-05)),(to_sfixed_a(-0.00023751652042847127)),(to_sfixed_a(-3.028564970009029e-05)),(to_sfixed_a(0.4209862947463989)),(to_sfixed_a(-0.002633706433698535)),(to_sfixed_a(-0.0016876541776582599)),(to_sfixed_a(-0.00375234242528677)),(to_sfixed_a(2.954155206680298e-06)),(to_sfixed_a(-0.00837712548673153)),(to_sfixed_a(6.285191921051592e-05)),(to_sfixed_a(1.7267666407860816e-07)),(to_sfixed_a(0.005550707690417767)),(to_sfixed_a(-0.009429886005818844)),(to_sfixed_a(-0.0010933929588645697)),(to_sfixed_a(5.5824348237365484e-06)),(to_sfixed_a(0.41804206371307373)),(to_sfixed_a(0.00022524395899381489)),(to_sfixed_a(0.003931897226721048)),(to_sfixed_a(0.4698803424835205)),(to_sfixed_a(-0.022196097299456596)),(to_sfixed_a(-0.3603837192058563)),(to_sfixed_a(0.0011415291810408235)),(to_sfixed_a(-0.12400910258293152)),(to_sfixed_a(-2.3678694560658187e-05)),(to_sfixed_a(0.00021153791749384254)),(to_sfixed_a(1.7954800568986684e-05)),(to_sfixed_a(0.0023158201947808266)),(to_sfixed_a(0.2300841510295868)),(to_sfixed_a(-0.00016602504183538258)),(to_sfixed_a(-0.0005199870793148875)),(to_sfixed_a(-0.0036938178818672895)),(to_sfixed_a(-0.00012757958029396832)),(to_sfixed_a(-2.1966861822875217e-05)),(to_sfixed_a(0.0028503926005214453)),(to_sfixed_a(0.1606033742427826)),(to_sfixed_a(-6.791116902604699e-05)),(to_sfixed_a(-0.009361578151583672)),(to_sfixed_a(-0.00018168851966038346)),(to_sfixed_a(0.011374793015420437)),(to_sfixed_a(-0.002374690491706133)),(to_sfixed_a(7.114635081961751e-05)),(to_sfixed_a(-6.959297752473503e-05)),(to_sfixed_a(6.358536484185606e-05)),(to_sfixed_a(-0.00018289239960722625)),(to_sfixed_a(-6.501070311060175e-05)),(to_sfixed_a(7.019617623882368e-05)),(to_sfixed_a(-0.00232065306045115)),(to_sfixed_a(0.0016392961842939258)),(to_sfixed_a(-0.009386742487549782)),(to_sfixed_a(0.00680816825479269)),(to_sfixed_a(0.004046018701046705)),(to_sfixed_a(0.00499550998210907)),(to_sfixed_a(0.0002980594290420413)),(to_sfixed_a(0.00015659857308492064)),(to_sfixed_a(-0.00028024264611303806)),(to_sfixed_a(3.3209209505002946e-05)),(to_sfixed_a(0.00013553540338762105)),(to_sfixed_a(0.000767130870372057)),(to_sfixed_a(0.0019006783841177821)),(to_sfixed_a(0.011994262225925922)),(to_sfixed_a(-0.00014782138168811798)),(to_sfixed_a(3.775550430873409e-05)),(to_sfixed_a(0.00012829834304284304)),(to_sfixed_a(-7.036404713289812e-05)),(to_sfixed_a(-0.00015964885824359953)),(to_sfixed_a(0.008342912420630455)),(to_sfixed_a(7.082626689225435e-05)),(to_sfixed_a(-4.6162313083186746e-06)),(to_sfixed_a(0.0002123812009813264)),(to_sfixed_a(0.015013353899121284)),(to_sfixed_a(-0.19650033116340637)),(to_sfixed_a(0.0002029908064287156)),(to_sfixed_a(-0.00022357759007718414)),(to_sfixed_a(-8.5494524682872e-05)),(to_sfixed_a(0.00015191621787380427)),(to_sfixed_a(0.002752563450485468)),(to_sfixed_a(0.004160786513239145)),(to_sfixed_a(-0.013201615773141384)),(to_sfixed_a(-0.0003043117467314005)),(to_sfixed_a(-0.0009045812766999006)),(to_sfixed_a(0.00018100535089615732)),(to_sfixed_a(-0.0034409884829074144)),(to_sfixed_a(-7.247366011142731e-05)),(to_sfixed_a(0.001121583511121571)),(to_sfixed_a(6.825714081060141e-05)),(to_sfixed_a(0.20730440318584442)),(to_sfixed_a(0.0049738031812012196)),(to_sfixed_a(0.0010681048734113574)),(to_sfixed_a(-0.5818359851837158)),(to_sfixed_a(-0.00015159363101702183)),(to_sfixed_a(0.12163206189870834)),(to_sfixed_a(0.008472362533211708)),(to_sfixed_a(8.348141273017973e-05)),(to_sfixed_a(0.5065602660179138)),(to_sfixed_a(6.579258479177952e-05)),(to_sfixed_a(7.3079900175798684e-06)),(to_sfixed_a(0.0002338762569706887)),(to_sfixed_a(0.005773727782070637)),(to_sfixed_a(-0.00013673139619641006)),(to_sfixed_a(-0.00013601752289105207)),(to_sfixed_a(-0.15513430535793304)),(to_sfixed_a(-6.21684012003243e-06)),(to_sfixed_a(-0.00203521060757339)),(to_sfixed_a(0.00030565293855033815)),(to_sfixed_a(4.330131923779845e-05)),(to_sfixed_a(-0.00023631709336768836)),(to_sfixed_a(0.003449512179940939)),(to_sfixed_a(0.00013731312355957925)),(to_sfixed_a(-2.1742391254520044e-05)),(to_sfixed_a(0.0001280369033338502)),(to_sfixed_a(-0.0018317201174795628)),(to_sfixed_a(0.0005433906335383654)),(to_sfixed_a(0.0002849235024768859)),(to_sfixed_a(0.00028072044369764626)),(to_sfixed_a(-0.00019342161249369383)),(to_sfixed_a(7.358851871686056e-05)),(to_sfixed_a(-0.36903175711631775)),(to_sfixed_a(0.002185311634093523)),(to_sfixed_a(0.4930793344974518)),(to_sfixed_a(-0.03238372504711151)),(to_sfixed_a(-0.0017729722894728184)),(to_sfixed_a(3.6162473406875506e-05)),(to_sfixed_a(0.0001597956579644233)),(to_sfixed_a(5.8079822338186204e-05)),(to_sfixed_a(0.0032460824586451054)),(to_sfixed_a(-3.504855339997448e-05)),(to_sfixed_a(0.00016829048399813473)),(to_sfixed_a(0.000710479449480772)),(to_sfixed_a(0.0032247749622911215)),(to_sfixed_a(0.00015097657160367817)),(to_sfixed_a(-0.4257880747318268)),(to_sfixed_a(0.0005130816134624183)),(to_sfixed_a(-0.0004748156643472612)),(to_sfixed_a(0.02971680462360382)),(to_sfixed_a(-0.00030440191039815545)),(to_sfixed_a(-0.020967693999409676)),(to_sfixed_a(0.33834370970726013)),(to_sfixed_a(0.008119340054690838)),(to_sfixed_a(-0.00025068753166124225)),(to_sfixed_a(-0.004504924640059471)),(to_sfixed_a(-0.34664782881736755)),(to_sfixed_a(0.008323121815919876)));

    constant weight_n2_15 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.21617773175239563)),(to_sfixed_a(-0.18329694867134094)),(to_sfixed_a(-0.007796654477715492)),(to_sfixed_a(-5.714629514841363e-05)),(to_sfixed_a(0.2622179090976715)),(to_sfixed_a(0.00011247643851675093)),(to_sfixed_a(0.0008073691860772669)),(to_sfixed_a(1.0575698979664594e-05)),(to_sfixed_a(-0.0001595806097611785)),(to_sfixed_a(-0.00010231781925540417)),(to_sfixed_a(-7.935766188893467e-05)),(to_sfixed_a(-0.4143151342868805)),(to_sfixed_a(-0.011511781252920628)),(to_sfixed_a(0.38901495933532715)),(to_sfixed_a(-2.15661057154648e-05)),(to_sfixed_a(0.00016675690130796283)),(to_sfixed_a(0.1959778368473053)),(to_sfixed_a(0.00010610064782667905)),(to_sfixed_a(0.0027951658703386784)),(to_sfixed_a(-0.0030577650759369135)),(to_sfixed_a(4.7126708523137495e-05)),(to_sfixed_a(7.238134276121855e-05)),(to_sfixed_a(0.26611900329589844)),(to_sfixed_a(-0.005029743537306786)),(to_sfixed_a(-0.003748824819922447)),(to_sfixed_a(0.0006714488845318556)),(to_sfixed_a(0.00014045134594198316)),(to_sfixed_a(0.15848354995250702)),(to_sfixed_a(0.009463002905249596)),(to_sfixed_a(-4.633464777725749e-05)),(to_sfixed_a(-0.011270559392869473)),(to_sfixed_a(6.851958460174501e-06)),(to_sfixed_a(0.03336305171251297)),(to_sfixed_a(0.00011632363748503849)),(to_sfixed_a(-6.937946454854682e-05)),(to_sfixed_a(0.00016188282461371273)),(to_sfixed_a(0.07239965349435806)),(to_sfixed_a(-0.0009521108004264534)),(to_sfixed_a(0.005237935576587915)),(to_sfixed_a(-7.05861602909863e-05)),(to_sfixed_a(0.07668719440698624)),(to_sfixed_a(-0.0007326305494643748)),(to_sfixed_a(-1.2943492038175464e-06)),(to_sfixed_a(-9.599461918696761e-06)),(to_sfixed_a(0.3023549020290375)),(to_sfixed_a(0.00894679594784975)),(to_sfixed_a(-0.2547825872898102)),(to_sfixed_a(0.3368062376976013)),(to_sfixed_a(0.00022400188026949763)),(to_sfixed_a(0.005562763195484877)),(to_sfixed_a(0.28159189224243164)),(to_sfixed_a(0.0003296390932518989)),(to_sfixed_a(0.00018057650595437735)),(to_sfixed_a(0.00015015406825114042)),(to_sfixed_a(-0.009712054394185543)),(to_sfixed_a(-0.012339742854237556)),(to_sfixed_a(-0.00013607789878733456)),(to_sfixed_a(-0.004721490666270256)),(to_sfixed_a(0.0001497546472819522)),(to_sfixed_a(0.00016808223153930157)),(to_sfixed_a(0.0008658189326524734)),(to_sfixed_a(-0.00011289956455584615)),(to_sfixed_a(-0.00021109799854457378)),(to_sfixed_a(-0.00010719207784859464)),(to_sfixed_a(9.235978359356523e-05)),(to_sfixed_a(0.011057578027248383)),(to_sfixed_a(7.203778659459203e-05)),(to_sfixed_a(0.006134495604783297)),(to_sfixed_a(0.002240187954157591)),(to_sfixed_a(0.0001369712845189497)),(to_sfixed_a(0.016327014192938805)),(to_sfixed_a(0.0006265425472520292)),(to_sfixed_a(-0.007879800163209438)),(to_sfixed_a(-9.347168088424951e-07)),(to_sfixed_a(0.0002060295664705336)),(to_sfixed_a(7.617097435286269e-05)),(to_sfixed_a(-0.6301912069320679)),(to_sfixed_a(-0.002361405175179243)),(to_sfixed_a(-0.00011382811499061063)),(to_sfixed_a(-0.3634254038333893)),(to_sfixed_a(0.0002310533745912835)),(to_sfixed_a(-0.00010581589594949037)),(to_sfixed_a(-0.33758610486984253)),(to_sfixed_a(-0.009284181520342827)),(to_sfixed_a(-0.00011434676707722247)),(to_sfixed_a(-0.004777754656970501)),(to_sfixed_a(0.004292291589081287)),(to_sfixed_a(0.0020591518841683865)),(to_sfixed_a(-0.00014897945220582187)),(to_sfixed_a(-2.856719947885722e-05)),(to_sfixed_a(0.2898898124694824)),(to_sfixed_a(2.3497537767980248e-05)),(to_sfixed_a(-0.002473041880875826)),(to_sfixed_a(6.624090019613504e-06)),(to_sfixed_a(-0.2022956907749176)),(to_sfixed_a(-4.868174437433481e-05)),(to_sfixed_a(-1.134566991822794e-05)),(to_sfixed_a(3.177058897563256e-05)),(to_sfixed_a(6.151928391773254e-05)),(to_sfixed_a(1.8006612663157284e-05)),(to_sfixed_a(-0.0064446753822267056)),(to_sfixed_a(-0.008339136838912964)),(to_sfixed_a(0.00014699444000143558)),(to_sfixed_a(-0.0013054523151367903)),(to_sfixed_a(-0.22274795174598694)),(to_sfixed_a(-0.0005408723372966051)),(to_sfixed_a(0.0001872805441962555)),(to_sfixed_a(-3.379905319889076e-05)),(to_sfixed_a(-0.0001847728854045272)),(to_sfixed_a(0.015304693952202797)),(to_sfixed_a(0.1138613224029541)),(to_sfixed_a(-0.00014912635379005224)),(to_sfixed_a(0.23957152664661407)),(to_sfixed_a(-0.00045273834257386625)),(to_sfixed_a(0.00013655841758009046)),(to_sfixed_a(-0.21380649507045746)),(to_sfixed_a(-0.002681704005226493)),(to_sfixed_a(8.357145998161286e-05)),(to_sfixed_a(-6.45416002953425e-05)),(to_sfixed_a(0.007592435926198959)),(to_sfixed_a(5.6510165450163186e-05)),(to_sfixed_a(-0.00023777273599989712)),(to_sfixed_a(0.007180350366979837)),(to_sfixed_a(0.0003012878296431154)),(to_sfixed_a(-6.931393727427348e-05)),(to_sfixed_a(0.0028352453373372555)),(to_sfixed_a(-0.0004419631150085479)),(to_sfixed_a(0.00023956030781846493)),(to_sfixed_a(-3.6507433833321556e-05)),(to_sfixed_a(5.9951657021883875e-05)),(to_sfixed_a(-0.00017856081831268966)),(to_sfixed_a(-0.0001745967601891607)),(to_sfixed_a(7.388580706901848e-05)),(to_sfixed_a(-0.0004896438331343234)),(to_sfixed_a(0.0002872711920645088)),(to_sfixed_a(-0.0002273978607263416)),(to_sfixed_a(0.007060131523758173)),(to_sfixed_a(0.0002809966681525111)),(to_sfixed_a(-6.607048271689564e-05)),(to_sfixed_a(0.00016090739518404007)),(to_sfixed_a(0.3885212242603302)),(to_sfixed_a(9.875085379462689e-05)),(to_sfixed_a(-8.354133751709014e-05)),(to_sfixed_a(-4.569254815578461e-05)),(to_sfixed_a(-0.39753803610801697)),(to_sfixed_a(0.0036147336941212416)),(to_sfixed_a(0.0025439588353037834)),(to_sfixed_a(-8.382994565181434e-06)),(to_sfixed_a(2.5124551029875875e-05)),(to_sfixed_a(-0.009149712510406971)),(to_sfixed_a(0.00014864170225337148)),(to_sfixed_a(0.00017961897538043559)),(to_sfixed_a(0.00042747377301566303)),(to_sfixed_a(-4.4225205783732235e-05)),(to_sfixed_a(0.00017784093506634235)),(to_sfixed_a(-0.2206079661846161)),(to_sfixed_a(6.776977534173056e-05)),(to_sfixed_a(0.0019827450159937143)),(to_sfixed_a(-2.3322278138948604e-05)),(to_sfixed_a(6.745212886016816e-05)),(to_sfixed_a(-8.305905794259161e-07)),(to_sfixed_a(0.00021924005704931915)),(to_sfixed_a(0.003133418271318078)),(to_sfixed_a(0.13342587649822235)),(to_sfixed_a(-0.0031386285554617643)),(to_sfixed_a(-0.0043052746914327145)),(to_sfixed_a(0.00011581535363802686)),(to_sfixed_a(0.6813656687736511)),(to_sfixed_a(0.00031133179436437786)),(to_sfixed_a(3.201768049621023e-05)),(to_sfixed_a(-0.3249366879463196)),(to_sfixed_a(-0.0012556720757856965)),(to_sfixed_a(0.0001812686095945537)),(to_sfixed_a(-1.8757993530016392e-05)),(to_sfixed_a(-0.0067731281742453575)),(to_sfixed_a(0.0008749378030188382)),(to_sfixed_a(-0.002709174994379282)),(to_sfixed_a(0.0013860298786312342)),(to_sfixed_a(-0.028784777969121933)),(to_sfixed_a(-0.00037984177470207214)),(to_sfixed_a(0.00027848960598930717)),(to_sfixed_a(0.39296048879623413)),(to_sfixed_a(0.0001668366603553295)),(to_sfixed_a(5.270315159577876e-05)),(to_sfixed_a(-0.00010637041850714013)),(to_sfixed_a(-0.0423622727394104)),(to_sfixed_a(0.0058166212402284145)),(to_sfixed_a(-0.003435650607571006)),(to_sfixed_a(0.00022199952218215913)),(to_sfixed_a(0.0004981544916518033)),(to_sfixed_a(-0.010324257425963879)),(to_sfixed_a(2.8569091227836907e-05)),(to_sfixed_a(0.005286108702421188)),(to_sfixed_a(0.0002904689754359424)),(to_sfixed_a(-0.00011502618144731969)),(to_sfixed_a(0.2509915828704834)),(to_sfixed_a(-3.517384175211191e-05)),(to_sfixed_a(-0.0018635645974427462)),(to_sfixed_a(-0.23503383994102478)),(to_sfixed_a(1.1707379599101841e-07)),(to_sfixed_a(0.00015051689115352929)),(to_sfixed_a(-0.00026874305331148207)),(to_sfixed_a(0.00018435339734423906)),(to_sfixed_a(8.326134411618114e-05)),(to_sfixed_a(-2.5478158931946382e-05)),(to_sfixed_a(0.007495907600969076)),(to_sfixed_a(-0.021360529586672783)),(to_sfixed_a(0.3048698306083679)),(to_sfixed_a(0.004405953921377659)),(to_sfixed_a(0.21448449790477753)),(to_sfixed_a(0.09136087447404861)),(to_sfixed_a(-0.00011616491246968508)),(to_sfixed_a(0.0001926052791532129)),(to_sfixed_a(6.109708920121193e-06)),(to_sfixed_a(-0.00012539204908534884)),(to_sfixed_a(-0.0002725614467635751)),(to_sfixed_a(0.0029549223836511374)),(to_sfixed_a(0.10280673950910568)),(to_sfixed_a(0.020282505080103874)),(to_sfixed_a(6.679864600300789e-05)),(to_sfixed_a(-0.00030510424403473735)),(to_sfixed_a(-8.574099047109485e-05)),(to_sfixed_a(-0.00011366778198862448)),(to_sfixed_a(0.0011660507880151272)),(to_sfixed_a(0.4916321337223053)),(to_sfixed_a(0.0002384420222369954)),(to_sfixed_a(4.393245035316795e-06)),(to_sfixed_a(-0.000171195380971767)),(to_sfixed_a(0.020174620673060417)),(to_sfixed_a(-0.27929404377937317)),(to_sfixed_a(-0.30246883630752563)),(to_sfixed_a(-8.119078120216727e-05)),(to_sfixed_a(-0.00018554338021203876)),(to_sfixed_a(-6.465379556175321e-05)),(to_sfixed_a(9.621826757211238e-05)),(to_sfixed_a(-0.0026948682498186827)),(to_sfixed_a(0.014367087744176388)),(to_sfixed_a(-0.00015345080464612693)),(to_sfixed_a(-2.5037817977136e-05)),(to_sfixed_a(-0.00029674224788323045)),(to_sfixed_a(-0.2260608822107315)),(to_sfixed_a(0.00020460184896364808)),(to_sfixed_a(-0.2697025239467621)),(to_sfixed_a(0.00031629117438569665)),(to_sfixed_a(0.01104773674160242)),(to_sfixed_a(0.33307355642318726)),(to_sfixed_a(0.00018273404566571116)),(to_sfixed_a(-0.21652443706989288)),(to_sfixed_a(0.0001553082838654518)),(to_sfixed_a(6.455864786403254e-05)),(to_sfixed_a(-0.010597732849419117)),(to_sfixed_a(0.0001138033258030191)),(to_sfixed_a(-0.0003255583578720689)),(to_sfixed_a(-0.00015322284889407456)),(to_sfixed_a(0.0001439689367543906)),(to_sfixed_a(-0.12482624500989914)),(to_sfixed_a(0.0047225067391991615)),(to_sfixed_a(-3.0833074561087415e-05)),(to_sfixed_a(1.2438340490916744e-06)),(to_sfixed_a(0.006987759843468666)),(to_sfixed_a(-6.130043766461313e-05)),(to_sfixed_a(-0.2075057476758957)),(to_sfixed_a(-0.00017951075278688222)),(to_sfixed_a(-0.00010357208520872518)),(to_sfixed_a(-0.0001166721194749698)),(to_sfixed_a(0.17057082056999207)),(to_sfixed_a(0.00014972077042330056)),(to_sfixed_a(0.00015876349061727524)),(to_sfixed_a(-0.00015049769717734307)),(to_sfixed_a(-0.0029717159923166037)),(to_sfixed_a(0.18747732043266296)),(to_sfixed_a(5.0631871999939904e-05)),(to_sfixed_a(6.6975990193896e-05)),(to_sfixed_a(0.00016775575932115316)),(to_sfixed_a(6.847805343568325e-05)),(to_sfixed_a(-0.3582412600517273)),(to_sfixed_a(0.003914929460734129)),(to_sfixed_a(0.00013398299051914364)),(to_sfixed_a(-0.008788788691163063)),(to_sfixed_a(0.0029996572993695736)),(to_sfixed_a(-0.00010791290696943179)),(to_sfixed_a(2.4337019567610696e-05)),(to_sfixed_a(0.00027377187507227063)),(to_sfixed_a(-0.007589160464704037)),(to_sfixed_a(-0.00023794188746251166)),(to_sfixed_a(1.5842531865928322e-05)),(to_sfixed_a(-0.003985084593296051)),(to_sfixed_a(0.02375981956720352)),(to_sfixed_a(-0.00017456940258853137)),(to_sfixed_a(-0.0017355744494125247)),(to_sfixed_a(0.0010434665018692613)),(to_sfixed_a(-0.004551921039819717)),(to_sfixed_a(-0.0016386042116209865)),(to_sfixed_a(1.9433886336628348e-05)),(to_sfixed_a(0.006507956888526678)),(to_sfixed_a(0.0022624742705374956)),(to_sfixed_a(-0.0051207635551691055)),(to_sfixed_a(-3.0575261916965246e-05)),(to_sfixed_a(-0.002842127112671733)),(to_sfixed_a(0.2211207151412964)),(to_sfixed_a(-0.009293405339121819)));

    constant weight_n2_16 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.03856227919459343)),(to_sfixed_a(0.007489468436688185)),(to_sfixed_a(0.0028883726336061954)),(to_sfixed_a(-3.913621912943199e-05)),(to_sfixed_a(0.28517216444015503)),(to_sfixed_a(0.00013386075443122536)),(to_sfixed_a(0.0027391156181693077)),(to_sfixed_a(-7.317124982364476e-05)),(to_sfixed_a(-0.0002195091510657221)),(to_sfixed_a(-0.0001055691100191325)),(to_sfixed_a(0.00015619504847563803)),(to_sfixed_a(0.00021625161753036082)),(to_sfixed_a(-0.0013149131555110216)),(to_sfixed_a(0.004556544125080109)),(to_sfixed_a(-2.5166318664560094e-05)),(to_sfixed_a(-0.0001910541468532756)),(to_sfixed_a(0.0022206378635019064)),(to_sfixed_a(0.00015776304644532502)),(to_sfixed_a(0.006048231385648251)),(to_sfixed_a(-0.016386590898036957)),(to_sfixed_a(-0.00023788146791048348)),(to_sfixed_a(0.00018211998394690454)),(to_sfixed_a(-0.00016229241737164557)),(to_sfixed_a(-0.014103911817073822)),(to_sfixed_a(9.579697507433593e-05)),(to_sfixed_a(0.17932304739952087)),(to_sfixed_a(-7.274039671756327e-05)),(to_sfixed_a(0.000625895569100976)),(to_sfixed_a(-0.0011377552291378379)),(to_sfixed_a(-0.0001070958242053166)),(to_sfixed_a(0.3549391031265259)),(to_sfixed_a(9.651890286477283e-05)),(to_sfixed_a(-0.1177818775177002)),(to_sfixed_a(3.6547440686263144e-05)),(to_sfixed_a(-1.5739642549306154e-06)),(to_sfixed_a(0.0003072481194976717)),(to_sfixed_a(0.21129557490348816)),(to_sfixed_a(-7.821075269021094e-05)),(to_sfixed_a(0.01196333859115839)),(to_sfixed_a(-5.9560625231824815e-05)),(to_sfixed_a(-0.2966969311237335)),(to_sfixed_a(0.0003846271429210901)),(to_sfixed_a(-0.0002466453588567674)),(to_sfixed_a(-0.00013403623597696424)),(to_sfixed_a(-0.00013673990906681865)),(to_sfixed_a(0.20219686627388)),(to_sfixed_a(0.0014883847907185555)),(to_sfixed_a(-0.006371624302119017)),(to_sfixed_a(0.000232772043091245)),(to_sfixed_a(-0.004821549169719219)),(to_sfixed_a(-0.015811292454600334)),(to_sfixed_a(4.9887632485479116e-05)),(to_sfixed_a(-3.7152713048271835e-06)),(to_sfixed_a(-0.0010551335290074348)),(to_sfixed_a(-0.049962833523750305)),(to_sfixed_a(0.009781130589544773)),(to_sfixed_a(-2.0113264326937497e-05)),(to_sfixed_a(0.3346881866455078)),(to_sfixed_a(-0.0002640864986460656)),(to_sfixed_a(-0.00010133324394701049)),(to_sfixed_a(-0.00019989338761661202)),(to_sfixed_a(0.0003762476844713092)),(to_sfixed_a(-0.00016430026153102517)),(to_sfixed_a(0.003209024900570512)),(to_sfixed_a(-0.0003152851713821292)),(to_sfixed_a(0.5006456971168518)),(to_sfixed_a(-0.00015368693857453763)),(to_sfixed_a(0.011340162716805935)),(to_sfixed_a(0.0027504777535796165)),(to_sfixed_a(4.3227701098658144e-06)),(to_sfixed_a(0.3043205738067627)),(to_sfixed_a(0.6545448303222656)),(to_sfixed_a(-0.0047156186774373055)),(to_sfixed_a(3.7140191125217825e-05)),(to_sfixed_a(1.7236154235433787e-05)),(to_sfixed_a(-0.00015233982412610203)),(to_sfixed_a(-0.017726602032780647)),(to_sfixed_a(-0.003739195642992854)),(to_sfixed_a(-0.00020458368817344308)),(to_sfixed_a(-0.251812219619751)),(to_sfixed_a(-0.004201299976557493)),(to_sfixed_a(-0.0001577552466187626)),(to_sfixed_a(0.4436044692993164)),(to_sfixed_a(-0.010627789422869682)),(to_sfixed_a(0.0001531406887806952)),(to_sfixed_a(-0.0020422611851245165)),(to_sfixed_a(-0.1968413144350052)),(to_sfixed_a(0.00030944732134230435)),(to_sfixed_a(-6.263570685405284e-05)),(to_sfixed_a(-9.168379619950429e-07)),(to_sfixed_a(0.018496191129088402)),(to_sfixed_a(0.00037951100966893137)),(to_sfixed_a(0.004459022544324398)),(to_sfixed_a(5.009114829590544e-06)),(to_sfixed_a(0.004839019384235144)),(to_sfixed_a(-4.487660771701485e-05)),(to_sfixed_a(-0.00019528332632035017)),(to_sfixed_a(0.00010351072705816478)),(to_sfixed_a(7.714620005572215e-05)),(to_sfixed_a(-0.00041740055894479156)),(to_sfixed_a(-0.024366557598114014)),(to_sfixed_a(8.980461279861629e-05)),(to_sfixed_a(3.099583409493789e-05)),(to_sfixed_a(0.0017700828611850739)),(to_sfixed_a(0.3625852167606354)),(to_sfixed_a(-0.003102090209722519)),(to_sfixed_a(-8.696551230968907e-05)),(to_sfixed_a(0.00011021007958333939)),(to_sfixed_a(-0.00021905521862208843)),(to_sfixed_a(-0.0003195694007445127)),(to_sfixed_a(0.1375715136528015)),(to_sfixed_a(-8.266351505881175e-05)),(to_sfixed_a(-0.0018943754257634282)),(to_sfixed_a(-0.000212672573979944)),(to_sfixed_a(-5.7872959587257355e-05)),(to_sfixed_a(-0.005181113723665476)),(to_sfixed_a(0.0039076791144907475)),(to_sfixed_a(0.0002646562934387475)),(to_sfixed_a(0.0001376264845021069)),(to_sfixed_a(-6.863056478323415e-05)),(to_sfixed_a(-2.8660375392064452e-05)),(to_sfixed_a(-0.0003059200826101005)),(to_sfixed_a(0.00020703100017271936)),(to_sfixed_a(2.9636808903887868e-05)),(to_sfixed_a(-8.470973989460617e-05)),(to_sfixed_a(-0.2991509437561035)),(to_sfixed_a(-0.008853605017066002)),(to_sfixed_a(-8.41305372887291e-05)),(to_sfixed_a(-9.824004519032314e-05)),(to_sfixed_a(0.00015718111535534263)),(to_sfixed_a(-7.755830301903188e-05)),(to_sfixed_a(6.409803609130904e-05)),(to_sfixed_a(0.264963299036026)),(to_sfixed_a(0.24419091641902924)),(to_sfixed_a(-4.727638588519767e-05)),(to_sfixed_a(6.92551548127085e-05)),(to_sfixed_a(-0.21752797067165375)),(to_sfixed_a(0.0010646377922967076)),(to_sfixed_a(-0.00012000579590676352)),(to_sfixed_a(6.78322758176364e-05)),(to_sfixed_a(0.00685980124399066)),(to_sfixed_a(-0.00015501785674132407)),(to_sfixed_a(-2.0799285266548395e-05)),(to_sfixed_a(-6.64670515106991e-05)),(to_sfixed_a(0.0036752286832779646)),(to_sfixed_a(0.0010859499452635646)),(to_sfixed_a(-0.0011995964450761676)),(to_sfixed_a(-0.0001178680031443946)),(to_sfixed_a(0.00010613564518280327)),(to_sfixed_a(0.012899977155029774)),(to_sfixed_a(8.889779564924538e-06)),(to_sfixed_a(0.00022235164942685515)),(to_sfixed_a(0.011536423116922379)),(to_sfixed_a(-6.367731839418411e-05)),(to_sfixed_a(-0.00020075369684491307)),(to_sfixed_a(0.0026704217307269573)),(to_sfixed_a(8.560877904528752e-05)),(to_sfixed_a(-0.03219429403543472)),(to_sfixed_a(-9.71029803622514e-05)),(to_sfixed_a(5.6532007874920964e-06)),(to_sfixed_a(0.0001341134193353355)),(to_sfixed_a(-7.365211786236614e-06)),(to_sfixed_a(0.000912183488253504)),(to_sfixed_a(0.0010231522610411048)),(to_sfixed_a(0.006079909857362509)),(to_sfixed_a(0.0017228976357728243)),(to_sfixed_a(-0.0004102984967175871)),(to_sfixed_a(0.0016531080473214388)),(to_sfixed_a(-0.0001841112389229238)),(to_sfixed_a(-0.00015351886395365)),(to_sfixed_a(-0.02544516697525978)),(to_sfixed_a(0.009638968855142593)),(to_sfixed_a(0.0019145195838063955)),(to_sfixed_a(0.00015502840687986463)),(to_sfixed_a(-0.5323270559310913)),(to_sfixed_a(0.004294636193662882)),(to_sfixed_a(-0.3980433940887451)),(to_sfixed_a(-4.838863605982624e-05)),(to_sfixed_a(-0.009561918675899506)),(to_sfixed_a(0.3794918358325958)),(to_sfixed_a(0.0006444230093620718)),(to_sfixed_a(0.26741883158683777)),(to_sfixed_a(-3.28449641529005e-05)),(to_sfixed_a(-0.00011522438580868766)),(to_sfixed_a(6.740183744113892e-05)),(to_sfixed_a(0.40678855776786804)),(to_sfixed_a(0.008737108670175076)),(to_sfixed_a(0.00034085914376191795)),(to_sfixed_a(7.012066816969309e-06)),(to_sfixed_a(0.0007368158549070358)),(to_sfixed_a(0.00031307560857385397)),(to_sfixed_a(-4.647143214242533e-05)),(to_sfixed_a(-0.0032373329158872366)),(to_sfixed_a(0.0035202328581362963)),(to_sfixed_a(0.00014672655379399657)),(to_sfixed_a(0.48696181178092957)),(to_sfixed_a(0.0001004127407213673)),(to_sfixed_a(0.003316644812002778)),(to_sfixed_a(-0.009154146537184715)),(to_sfixed_a(6.791832129238173e-05)),(to_sfixed_a(-7.168691081460565e-05)),(to_sfixed_a(-1.301792508456856e-05)),(to_sfixed_a(0.00010438275785418227)),(to_sfixed_a(0.0002266496594529599)),(to_sfixed_a(-9.666291589383036e-05)),(to_sfixed_a(0.004296894650906324)),(to_sfixed_a(0.0002616747806314379)),(to_sfixed_a(0.003807453438639641)),(to_sfixed_a(0.000925689993891865)),(to_sfixed_a(-0.0049936664290726185)),(to_sfixed_a(0.00976281613111496)),(to_sfixed_a(-0.0002734690497163683)),(to_sfixed_a(0.00015682249795645475)),(to_sfixed_a(-4.167846782365814e-05)),(to_sfixed_a(-0.00011253951379330829)),(to_sfixed_a(0.00010566063428996131)),(to_sfixed_a(3.2948722946457565e-05)),(to_sfixed_a(0.0014922566479071975)),(to_sfixed_a(0.004817601293325424)),(to_sfixed_a(3.7858320865780115e-05)),(to_sfixed_a(-0.00013613482587970793)),(to_sfixed_a(0.00010909747652476653)),(to_sfixed_a(-0.00016720716666895896)),(to_sfixed_a(-0.0006110897520557046)),(to_sfixed_a(-0.00703857559710741)),(to_sfixed_a(-0.000445985933765769)),(to_sfixed_a(0.00012944646005053073)),(to_sfixed_a(4.0401340811513364e-05)),(to_sfixed_a(-2.1632095013046637e-05)),(to_sfixed_a(-0.004159578122198582)),(to_sfixed_a(0.388467013835907)),(to_sfixed_a(1.0735020623542368e-06)),(to_sfixed_a(0.0002966067404486239)),(to_sfixed_a(-0.0002013982302742079)),(to_sfixed_a(0.003793630050495267)),(to_sfixed_a(0.0027289611753076315)),(to_sfixed_a(0.3682911992073059)),(to_sfixed_a(-6.622760702157393e-05)),(to_sfixed_a(-2.552017758716829e-05)),(to_sfixed_a(0.00038391887210309505)),(to_sfixed_a(0.0016844627680256963)),(to_sfixed_a(-0.00029000442009419203)),(to_sfixed_a(-0.0012825120938941836)),(to_sfixed_a(-0.0002634371048770845)),(to_sfixed_a(-0.1799192726612091)),(to_sfixed_a(-0.36781230568885803)),(to_sfixed_a(0.1763138473033905)),(to_sfixed_a(0.00012177292228443548)),(to_sfixed_a(-8.976123353932053e-05)),(to_sfixed_a(0.00683846278116107)),(to_sfixed_a(-0.01491785142570734)),(to_sfixed_a(-0.00011352567526046187)),(to_sfixed_a(0.00046421511797234416)),(to_sfixed_a(-0.00015022153093013912)),(to_sfixed_a(0.002066107001155615)),(to_sfixed_a(0.007073548156768084)),(to_sfixed_a(-0.002029696013778448)),(to_sfixed_a(9.881724690785632e-05)),(to_sfixed_a(0.00010677886893972754)),(to_sfixed_a(0.3768545091152191)),(to_sfixed_a(-0.00018589087994769216)),(to_sfixed_a(0.0015671809669584036)),(to_sfixed_a(0.00018948694923892617)),(to_sfixed_a(-0.0005008136504329741)),(to_sfixed_a(1.3356147974263877e-06)),(to_sfixed_a(-0.17849701642990112)),(to_sfixed_a(0.00013779420987702906)),(to_sfixed_a(-0.00011370090214768425)),(to_sfixed_a(0.0001678466796875)),(to_sfixed_a(0.3402903378009796)),(to_sfixed_a(0.07215842604637146)),(to_sfixed_a(0.00019459010218270123)),(to_sfixed_a(0.00011323876969981939)),(to_sfixed_a(0.00012907428026665002)),(to_sfixed_a(-3.484587068669498e-06)),(to_sfixed_a(0.005140902008861303)),(to_sfixed_a(-0.0005501837586052716)),(to_sfixed_a(4.1532228351570666e-05)),(to_sfixed_a(0.20900002121925354)),(to_sfixed_a(0.0006467816419899464)),(to_sfixed_a(3.7415738916024566e-06)),(to_sfixed_a(-0.0001819846365833655)),(to_sfixed_a(-0.00010263738658977672)),(to_sfixed_a(-0.0005249129608273506)),(to_sfixed_a(1.9640199752757326e-05)),(to_sfixed_a(-1.845127553679049e-05)),(to_sfixed_a(-0.0002241725305793807)),(to_sfixed_a(-0.03379373252391815)),(to_sfixed_a(0.00019964843522757292)),(to_sfixed_a(0.2821856439113617)),(to_sfixed_a(-3.099679452134296e-05)),(to_sfixed_a(0.00014643864415120333)),(to_sfixed_a(0.29139289259910583)),(to_sfixed_a(-4.06342587666586e-06)),(to_sfixed_a(0.0013143903343006968)),(to_sfixed_a(-0.5211092233657837)),(to_sfixed_a(-0.013890978880226612)),(to_sfixed_a(-0.00012030614743707702)),(to_sfixed_a(0.23998449742794037)),(to_sfixed_a(-0.6737775802612305)),(to_sfixed_a(-0.0009705541306175292)));

    constant weight_n2_17 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.3116753399372101)),(to_sfixed_a(-1.9304279703646898e-05)),(to_sfixed_a(-0.174137145280838)),(to_sfixed_a(-1.948764838743955e-05)),(to_sfixed_a(-0.0013356972485780716)),(to_sfixed_a(-7.08712832420133e-05)),(to_sfixed_a(-0.0008937224629335105)),(to_sfixed_a(-0.00018014184024650604)),(to_sfixed_a(-2.5599671062082052e-05)),(to_sfixed_a(-0.00010755356925074011)),(to_sfixed_a(-9.811027121031657e-05)),(to_sfixed_a(0.020352225750684738)),(to_sfixed_a(0.004304080735892057)),(to_sfixed_a(-0.0005967895849607885)),(to_sfixed_a(4.237932444084436e-05)),(to_sfixed_a(-5.658622831106186e-05)),(to_sfixed_a(0.3122752904891968)),(to_sfixed_a(-0.00013752646918874234)),(to_sfixed_a(0.0033503458835184574)),(to_sfixed_a(-0.25483158230781555)),(to_sfixed_a(-0.000153764383867383)),(to_sfixed_a(-0.00016936907195486128)),(to_sfixed_a(5.030788452131674e-05)),(to_sfixed_a(-0.017642296850681305)),(to_sfixed_a(-0.002627883106470108)),(to_sfixed_a(0.003080653492361307)),(to_sfixed_a(-0.00011511485354276374)),(to_sfixed_a(0.00010352776735089719)),(to_sfixed_a(-0.18620960414409637)),(to_sfixed_a(1.9353989046067e-05)),(to_sfixed_a(-0.00486213993281126)),(to_sfixed_a(-0.00011950139742111787)),(to_sfixed_a(0.002783417934551835)),(to_sfixed_a(-0.0002099062839988619)),(to_sfixed_a(-0.0002866225258912891)),(to_sfixed_a(0.0001578645606059581)),(to_sfixed_a(0.00014488361193798482)),(to_sfixed_a(-0.0009891304653137922)),(to_sfixed_a(0.0005397886270657182)),(to_sfixed_a(1.9119815988233313e-05)),(to_sfixed_a(-0.3639097511768341)),(to_sfixed_a(-0.5766999125480652)),(to_sfixed_a(1.677021646173671e-05)),(to_sfixed_a(4.76127679576166e-05)),(to_sfixed_a(-0.0017647022614255548)),(to_sfixed_a(-0.006820198148488998)),(to_sfixed_a(-0.002483253600075841)),(to_sfixed_a(-0.009481063112616539)),(to_sfixed_a(0.00013541422958951443)),(to_sfixed_a(-0.0029792857822030783)),(to_sfixed_a(0.0005909015308134258)),(to_sfixed_a(-0.0007720524445176125)),(to_sfixed_a(6.0162146837683395e-05)),(to_sfixed_a(0.0005551662761718035)),(to_sfixed_a(-0.0021660933271050453)),(to_sfixed_a(0.004830631427466869)),(to_sfixed_a(0.00018234402523376048)),(to_sfixed_a(0.17293669283390045)),(to_sfixed_a(0.00014688490773551166)),(to_sfixed_a(-0.0001263693266082555)),(to_sfixed_a(-0.0007832229021005332)),(to_sfixed_a(0.25938835740089417)),(to_sfixed_a(-0.0009849440539255738)),(to_sfixed_a(5.598074494628236e-05)),(to_sfixed_a(3.9465005102101713e-05)),(to_sfixed_a(-0.0008289232500828803)),(to_sfixed_a(4.337365317041986e-05)),(to_sfixed_a(-0.0006739493692293763)),(to_sfixed_a(1.2352888006716967e-05)),(to_sfixed_a(6.698718061670661e-05)),(to_sfixed_a(0.003581611905246973)),(to_sfixed_a(-0.001061446382664144)),(to_sfixed_a(-0.005897319409996271)),(to_sfixed_a(-7.429992547258735e-05)),(to_sfixed_a(0.00022774067474529147)),(to_sfixed_a(9.919670264935121e-05)),(to_sfixed_a(0.2360561043024063)),(to_sfixed_a(-0.002670327201485634)),(to_sfixed_a(-2.3726330255158246e-05)),(to_sfixed_a(-0.3171795606613159)),(to_sfixed_a(-0.002876490820199251)),(to_sfixed_a(-4.7052253648871556e-05)),(to_sfixed_a(-0.40348654985427856)),(to_sfixed_a(-0.00196881964802742)),(to_sfixed_a(-0.0001527427084511146)),(to_sfixed_a(-0.008419033139944077)),(to_sfixed_a(0.0007064040983095765)),(to_sfixed_a(-0.00014602995361201465)),(to_sfixed_a(0.00010652732453309)),(to_sfixed_a(-7.454809383489192e-05)),(to_sfixed_a(-0.0008201863965950906)),(to_sfixed_a(7.299552817130461e-05)),(to_sfixed_a(-0.0002456216316204518)),(to_sfixed_a(-0.00011370570427970961)),(to_sfixed_a(0.01593424752354622)),(to_sfixed_a(8.831106242723763e-05)),(to_sfixed_a(-2.303815563209355e-06)),(to_sfixed_a(0.00016056702588684857)),(to_sfixed_a(1.3037933968007565e-06)),(to_sfixed_a(5.627410428132862e-05)),(to_sfixed_a(-0.001358544104732573)),(to_sfixed_a(-0.0007815485587343574)),(to_sfixed_a(-1.1065458238590509e-06)),(to_sfixed_a(-0.18977606296539307)),(to_sfixed_a(-0.00010076328180730343)),(to_sfixed_a(-0.0023006589617580175)),(to_sfixed_a(6.638078775722533e-05)),(to_sfixed_a(1.2381409760564566e-05)),(to_sfixed_a(2.7948481147177517e-06)),(to_sfixed_a(-0.004223272670060396)),(to_sfixed_a(-0.00040086027001962066)),(to_sfixed_a(0.0002395105257164687)),(to_sfixed_a(0.0007375249988399446)),(to_sfixed_a(-0.0001566167047712952)),(to_sfixed_a(-2.2018466552253813e-06)),(to_sfixed_a(-0.003474154509603977)),(to_sfixed_a(0.005351128522306681)),(to_sfixed_a(0.00021044723689556122)),(to_sfixed_a(1.1140655260533094e-06)),(to_sfixed_a(0.00015380365948658437)),(to_sfixed_a(-0.00010066651157103479)),(to_sfixed_a(6.585758819710463e-05)),(to_sfixed_a(-0.0015832718927413225)),(to_sfixed_a(-2.3744505597278476e-05)),(to_sfixed_a(-2.7513160603120923e-06)),(to_sfixed_a(0.015989985316991806)),(to_sfixed_a(-0.007353695575147867)),(to_sfixed_a(-9.404431330040097e-05)),(to_sfixed_a(-0.00010391759860794991)),(to_sfixed_a(0.00012796593364328146)),(to_sfixed_a(-1.2884644092991948e-05)),(to_sfixed_a(-2.8810158255510032e-05)),(to_sfixed_a(0.0005726541276089847)),(to_sfixed_a(0.0012795035727322102)),(to_sfixed_a(-9.988090823753737e-06)),(to_sfixed_a(2.7571513783186674e-06)),(to_sfixed_a(-0.20347784459590912)),(to_sfixed_a(0.00018729298608377576)),(to_sfixed_a(-0.00029380081105045974)),(to_sfixed_a(0.00020967237651348114)),(to_sfixed_a(0.005221793428063393)),(to_sfixed_a(0.00022380278096534312)),(to_sfixed_a(0.00020167999900877476)),(to_sfixed_a(-1.6471449271193705e-05)),(to_sfixed_a(0.0007401076145470142)),(to_sfixed_a(-0.00020821610814891756)),(to_sfixed_a(0.0004783750046044588)),(to_sfixed_a(-0.0001188889509649016)),(to_sfixed_a(0.00016741348372306675)),(to_sfixed_a(0.24769921600818634)),(to_sfixed_a(-0.00020056140783708543)),(to_sfixed_a(-4.569486918626353e-05)),(to_sfixed_a(0.011622491292655468)),(to_sfixed_a(3.68434120900929e-05)),(to_sfixed_a(-0.00015032984083518386)),(to_sfixed_a(0.0031283965799957514)),(to_sfixed_a(0.00021160041796974838)),(to_sfixed_a(0.007095877546817064)),(to_sfixed_a(-6.704162660753354e-05)),(to_sfixed_a(-0.00016770872753113508)),(to_sfixed_a(-9.254926408175379e-05)),(to_sfixed_a(0.00012924362090416253)),(to_sfixed_a(0.000688342668581754)),(to_sfixed_a(-0.0022500380873680115)),(to_sfixed_a(0.39251360297203064)),(to_sfixed_a(0.0008570348145440221)),(to_sfixed_a(0.00021927997295279056)),(to_sfixed_a(-0.30142873525619507)),(to_sfixed_a(5.074882210465148e-05)),(to_sfixed_a(-0.0002018179657170549)),(to_sfixed_a(0.008006504736840725)),(to_sfixed_a(0.2955136001110077)),(to_sfixed_a(0.001466983463615179)),(to_sfixed_a(0.00011450082092778757)),(to_sfixed_a(0.012674751691520214)),(to_sfixed_a(0.0018749024020507932)),(to_sfixed_a(-0.00022603223624173552)),(to_sfixed_a(0.37761446833610535)),(to_sfixed_a(0.004038115497678518)),(to_sfixed_a(0.2593019902706146)),(to_sfixed_a(-0.0008037491934373975)),(to_sfixed_a(0.10166795551776886)),(to_sfixed_a(9.738458174979314e-05)),(to_sfixed_a(-3.039487637579441e-06)),(to_sfixed_a(2.7050162316299975e-05)),(to_sfixed_a(0.29833969473838806)),(to_sfixed_a(0.35072973370552063)),(to_sfixed_a(-0.0005212343530729413)),(to_sfixed_a(-6.59419092698954e-05)),(to_sfixed_a(0.5145688056945801)),(to_sfixed_a(-0.6220229864120483)),(to_sfixed_a(-2.94751826004358e-05)),(to_sfixed_a(-0.005043927114456892)),(to_sfixed_a(0.000152866035932675)),(to_sfixed_a(-0.00023842082009650767)),(to_sfixed_a(0.19374682009220123)),(to_sfixed_a(7.816081051714718e-06)),(to_sfixed_a(0.2764316499233246)),(to_sfixed_a(-0.0006456926930695772)),(to_sfixed_a(-4.366436769487336e-06)),(to_sfixed_a(0.0001527372223790735)),(to_sfixed_a(6.468766514444724e-05)),(to_sfixed_a(0.0001819487806642428)),(to_sfixed_a(0.00023283250629901886)),(to_sfixed_a(-0.0002864037815015763)),(to_sfixed_a(0.004145363811403513)),(to_sfixed_a(-0.00018981385801453143)),(to_sfixed_a(-0.22808530926704407)),(to_sfixed_a(-8.514308137819171e-05)),(to_sfixed_a(0.018660705536603928)),(to_sfixed_a(0.0004142542602494359)),(to_sfixed_a(0.00014664544141851366)),(to_sfixed_a(-4.1393504943698645e-05)),(to_sfixed_a(0.0001280889700865373)),(to_sfixed_a(0.00031070312252268195)),(to_sfixed_a(0.00024644736549817026)),(to_sfixed_a(0.006668452639132738)),(to_sfixed_a(0.0036759264767169952)),(to_sfixed_a(0.003493586089462042)),(to_sfixed_a(-2.2399341105483472e-05)),(to_sfixed_a(0.00016908530960790813)),(to_sfixed_a(-7.935120811453089e-05)),(to_sfixed_a(8.67556591401808e-05)),(to_sfixed_a(-0.000212421320611611)),(to_sfixed_a(0.0019098026677966118)),(to_sfixed_a(-8.334986341651529e-05)),(to_sfixed_a(1.009448169497773e-05)),(to_sfixed_a(-1.6101490473374724e-05)),(to_sfixed_a(0.3193855285644531)),(to_sfixed_a(0.0044704582542181015)),(to_sfixed_a(0.0005411727470345795)),(to_sfixed_a(5.819733996759169e-05)),(to_sfixed_a(0.00018105782510247082)),(to_sfixed_a(-0.0004129930166527629)),(to_sfixed_a(0.002914590761065483)),(to_sfixed_a(0.014830264262855053)),(to_sfixed_a(-2.446407961542718e-06)),(to_sfixed_a(-0.0001276019320357591)),(to_sfixed_a(-0.00020797828619834036)),(to_sfixed_a(-0.0002212137042079121)),(to_sfixed_a(0.001644806587137282)),(to_sfixed_a(0.00022479379549622536)),(to_sfixed_a(0.0017466654535382986)),(to_sfixed_a(0.00012613643775694072)),(to_sfixed_a(-0.00491469306871295)),(to_sfixed_a(0.00020369910635054111)),(to_sfixed_a(-0.002484146971255541)),(to_sfixed_a(-0.5703098177909851)),(to_sfixed_a(-3.908961662091315e-05)),(to_sfixed_a(0.3631496727466583)),(to_sfixed_a(-0.008940326049923897)),(to_sfixed_a(-8.491617336403579e-05)),(to_sfixed_a(0.0005678202142007649)),(to_sfixed_a(-7.032682333374396e-05)),(to_sfixed_a(0.003448331030085683)),(to_sfixed_a(-0.0021838268730789423)),(to_sfixed_a(-0.3931964039802551)),(to_sfixed_a(4.501237708609551e-05)),(to_sfixed_a(-3.824393934337422e-05)),(to_sfixed_a(0.2898997664451599)),(to_sfixed_a(0.0001043949305312708)),(to_sfixed_a(-0.0010977275669574738)),(to_sfixed_a(-3.886516788043082e-05)),(to_sfixed_a(-0.0011413050815463066)),(to_sfixed_a(2.4532222596462816e-05)),(to_sfixed_a(-0.008909521624445915)),(to_sfixed_a(5.8363424614071846e-05)),(to_sfixed_a(0.00022359246213454753)),(to_sfixed_a(-0.0001193557764054276)),(to_sfixed_a(0.49616414308547974)),(to_sfixed_a(-0.0029653471428900957)),(to_sfixed_a(-0.0002473705681040883)),(to_sfixed_a(0.00015650723071303219)),(to_sfixed_a(-0.00023678597062826157)),(to_sfixed_a(2.9670387448277324e-05)),(to_sfixed_a(0.00642926013097167)),(to_sfixed_a(0.0005735565209761262)),(to_sfixed_a(0.021307773888111115)),(to_sfixed_a(0.35164669156074524)),(to_sfixed_a(0.014582464471459389)),(to_sfixed_a(6.581882189493626e-05)),(to_sfixed_a(-1.659239933360368e-05)),(to_sfixed_a(-3.687790012918413e-05)),(to_sfixed_a(-0.0010405025677755475)),(to_sfixed_a(4.512803570833057e-06)),(to_sfixed_a(-0.00024037410912569612)),(to_sfixed_a(-6.343857967294753e-05)),(to_sfixed_a(0.2938118875026703)),(to_sfixed_a(0.0001988779113162309)),(to_sfixed_a(-0.0006650330615229905)),(to_sfixed_a(0.0016053641447797418)),(to_sfixed_a(-0.00014820322394371033)),(to_sfixed_a(0.011854685842990875)),(to_sfixed_a(0.00023643046733923256)),(to_sfixed_a(0.0013424132484942675)),(to_sfixed_a(-0.0006723811384290457)),(to_sfixed_a(0.10522580146789551)),(to_sfixed_a(6.612854485865682e-05)),(to_sfixed_a(0.31635352969169617)),(to_sfixed_a(-0.248929962515831)),(to_sfixed_a(-0.0018602991476655006)));

    constant weight_n2_18 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.3165515065193176)),(to_sfixed_a(-0.006984710693359375)),(to_sfixed_a(-0.000371187343262136)),(to_sfixed_a(1.2762175174430013e-06)),(to_sfixed_a(-0.3968222141265869)),(to_sfixed_a(-0.00022172405442688614)),(to_sfixed_a(0.018966402858495712)),(to_sfixed_a(3.095511783612892e-05)),(to_sfixed_a(7.093425665516406e-05)),(to_sfixed_a(-0.0002555914979893714)),(to_sfixed_a(-0.0001296435366384685)),(to_sfixed_a(5.565467290580273e-06)),(to_sfixed_a(0.0017290620598942041)),(to_sfixed_a(-0.0012439708225429058)),(to_sfixed_a(-8.569463534513488e-05)),(to_sfixed_a(6.35814867564477e-05)),(to_sfixed_a(0.0003366671153344214)),(to_sfixed_a(-0.00016960158245638013)),(to_sfixed_a(-0.022235283628106117)),(to_sfixed_a(0.0005199418519623578)),(to_sfixed_a(8.016233186936006e-05)),(to_sfixed_a(-0.00022252323105931282)),(to_sfixed_a(-8.01076166681014e-05)),(to_sfixed_a(0.001072983257472515)),(to_sfixed_a(0.004922407679259777)),(to_sfixed_a(-0.0013298648409545422)),(to_sfixed_a(-1.4914636267349124e-05)),(to_sfixed_a(-4.467843973543495e-05)),(to_sfixed_a(0.0008675518911331892)),(to_sfixed_a(-1.7081321857403964e-05)),(to_sfixed_a(0.011889971792697906)),(to_sfixed_a(0.00012830208288505673)),(to_sfixed_a(0.019251776859164238)),(to_sfixed_a(0.0001014970985124819)),(to_sfixed_a(1.2080090527888387e-06)),(to_sfixed_a(0.00016542081721127033)),(to_sfixed_a(-0.001482244930230081)),(to_sfixed_a(-0.005316745489835739)),(to_sfixed_a(-0.0003072292311117053)),(to_sfixed_a(-2.3077678633853793e-05)),(to_sfixed_a(0.3693672716617584)),(to_sfixed_a(0.008933734148740768)),(to_sfixed_a(2.56938801612705e-05)),(to_sfixed_a(8.488947787554935e-05)),(to_sfixed_a(-0.004375002346932888)),(to_sfixed_a(-0.1005341038107872)),(to_sfixed_a(-0.2961474061012268)),(to_sfixed_a(-1.8495211406843737e-05)),(to_sfixed_a(0.00021632021525874734)),(to_sfixed_a(0.0006969928508624434)),(to_sfixed_a(0.2319118082523346)),(to_sfixed_a(0.0004435935115907341)),(to_sfixed_a(0.00011480834655230865)),(to_sfixed_a(0.004352307878434658)),(to_sfixed_a(0.00036771546001546085)),(to_sfixed_a(-0.009870823472738266)),(to_sfixed_a(-4.5118424168322235e-05)),(to_sfixed_a(0.0018166637746617198)),(to_sfixed_a(3.683967224787921e-05)),(to_sfixed_a(1.4930992620065808e-05)),(to_sfixed_a(-0.32127201557159424)),(to_sfixed_a(0.000881565036252141)),(to_sfixed_a(-0.7215651869773865)),(to_sfixed_a(0.09417615085840225)),(to_sfixed_a(0.00017429747094865888)),(to_sfixed_a(-0.5851141810417175)),(to_sfixed_a(0.00017012396710924804)),(to_sfixed_a(0.0019267275929450989)),(to_sfixed_a(0.0003892676322720945)),(to_sfixed_a(-7.06592109054327e-05)),(to_sfixed_a(0.00173415697645396)),(to_sfixed_a(-0.007754209451377392)),(to_sfixed_a(-0.0027675130404531956)),(to_sfixed_a(-4.4153781345812604e-05)),(to_sfixed_a(-6.455451512010768e-05)),(to_sfixed_a(0.00013064091035630554)),(to_sfixed_a(0.0007800651947036386)),(to_sfixed_a(0.005975246895104647)),(to_sfixed_a(6.072826363379136e-05)),(to_sfixed_a(-0.00866515189409256)),(to_sfixed_a(0.10116598755121231)),(to_sfixed_a(-0.00010885584924835712)),(to_sfixed_a(-0.0007976364577189088)),(to_sfixed_a(-0.0007976285414770246)),(to_sfixed_a(0.0002922946878243238)),(to_sfixed_a(0.002322861459106207)),(to_sfixed_a(0.07787099480628967)),(to_sfixed_a(0.513041615486145)),(to_sfixed_a(-3.686875061248429e-05)),(to_sfixed_a(-6.96462084306404e-05)),(to_sfixed_a(-0.32769569754600525)),(to_sfixed_a(-0.00012010219506919384)),(to_sfixed_a(-0.0002869321615435183)),(to_sfixed_a(6.985645450185984e-05)),(to_sfixed_a(-0.3097834289073944)),(to_sfixed_a(-3.2014799216995016e-05)),(to_sfixed_a(-6.36408367427066e-05)),(to_sfixed_a(-9.00163286132738e-08)),(to_sfixed_a(6.345885049086064e-05)),(to_sfixed_a(-0.00013701994612347335)),(to_sfixed_a(-0.0007913687732070684)),(to_sfixed_a(0.4452202022075653)),(to_sfixed_a(0.00015375974180642515)),(to_sfixed_a(0.0005640584859065711)),(to_sfixed_a(-0.007382253184914589)),(to_sfixed_a(-0.0003609940467868)),(to_sfixed_a(-0.00013745044998358935)),(to_sfixed_a(-8.795839676167816e-06)),(to_sfixed_a(5.877076182514429e-05)),(to_sfixed_a(0.24298934638500214)),(to_sfixed_a(0.019577965140342712)),(to_sfixed_a(4.457286195247434e-05)),(to_sfixed_a(-0.0018354319036006927)),(to_sfixed_a(0.00020144088193774223)),(to_sfixed_a(0.0001168752642115578)),(to_sfixed_a(-0.07510402053594589)),(to_sfixed_a(0.001427126582711935)),(to_sfixed_a(-0.00014374818420037627)),(to_sfixed_a(8.761639764998108e-05)),(to_sfixed_a(-0.0017184690805152059)),(to_sfixed_a(-0.0001302206510445103)),(to_sfixed_a(-0.00016421612235717475)),(to_sfixed_a(-0.0031797627452760935)),(to_sfixed_a(-7.148247095756233e-05)),(to_sfixed_a(-0.00027869766927324235)),(to_sfixed_a(-0.00713656609877944)),(to_sfixed_a(0.23616206645965576)),(to_sfixed_a(0.0001746913039823994)),(to_sfixed_a(-0.00017501924594398588)),(to_sfixed_a(2.355970354983583e-05)),(to_sfixed_a(1.3472446880768985e-05)),(to_sfixed_a(-0.00012370396871119738)),(to_sfixed_a(-0.4468441307544708)),(to_sfixed_a(0.0006821146234869957)),(to_sfixed_a(0.00022765679750591516)),(to_sfixed_a(-5.720983608625829e-06)),(to_sfixed_a(-0.15429501235485077)),(to_sfixed_a(-0.00016735524695832282)),(to_sfixed_a(3.803146682912484e-05)),(to_sfixed_a(-0.00015744075062684715)),(to_sfixed_a(-0.0001081063601304777)),(to_sfixed_a(1.0937361366814002e-05)),(to_sfixed_a(1.1909309250768274e-05)),(to_sfixed_a(2.8212274628458545e-05)),(to_sfixed_a(-0.0031753929797559977)),(to_sfixed_a(3.790441405726597e-05)),(to_sfixed_a(-0.0001354869600618258)),(to_sfixed_a(5.1687093218788505e-05)),(to_sfixed_a(-0.00014911503240000457)),(to_sfixed_a(-0.0043286047875881195)),(to_sfixed_a(3.34227952407673e-05)),(to_sfixed_a(-0.0002038691018242389)),(to_sfixed_a(0.0029109977185726166)),(to_sfixed_a(5.670394602930173e-05)),(to_sfixed_a(6.900128937559202e-05)),(to_sfixed_a(0.00881364569067955)),(to_sfixed_a(5.953483560006134e-05)),(to_sfixed_a(0.26254352927207947)),(to_sfixed_a(0.0002289988042321056)),(to_sfixed_a(6.005138857290149e-06)),(to_sfixed_a(8.813823660602793e-05)),(to_sfixed_a(0.00014794376329518855)),(to_sfixed_a(-0.0011927601881325245)),(to_sfixed_a(0.002653442556038499)),(to_sfixed_a(0.018884075805544853)),(to_sfixed_a(-0.003203592961654067)),(to_sfixed_a(0.00010188547457801178)),(to_sfixed_a(-0.001055101864039898)),(to_sfixed_a(-0.00021267072588671)),(to_sfixed_a(0.00015194551087915897)),(to_sfixed_a(0.06203185394406319)),(to_sfixed_a(-0.008408249355852604)),(to_sfixed_a(0.34289321303367615)),(to_sfixed_a(-0.00014297959569375962)),(to_sfixed_a(0.003145707305520773)),(to_sfixed_a(0.2770184874534607)),(to_sfixed_a(0.004060744307935238)),(to_sfixed_a(1.751114905346185e-05)),(to_sfixed_a(0.003036698093637824)),(to_sfixed_a(-0.046866923570632935)),(to_sfixed_a(-1.6893325664568692e-05)),(to_sfixed_a(0.007678704336285591)),(to_sfixed_a(-0.00011734679719666019)),(to_sfixed_a(-7.445453957188874e-05)),(to_sfixed_a(-0.00023712449183221906)),(to_sfixed_a(0.025222577154636383)),(to_sfixed_a(0.08624422550201416)),(to_sfixed_a(-0.469608336687088)),(to_sfixed_a(0.0034772937651723623)),(to_sfixed_a(-0.00010836955334525555)),(to_sfixed_a(0.014828936196863651)),(to_sfixed_a(0.0002462013508193195)),(to_sfixed_a(0.0259889904409647)),(to_sfixed_a(0.2966102957725525)),(to_sfixed_a(3.022122837137431e-05)),(to_sfixed_a(-0.0041954792104661465)),(to_sfixed_a(2.9612183425342664e-05)),(to_sfixed_a(0.004187165759503841)),(to_sfixed_a(-0.43000179529190063)),(to_sfixed_a(0.0001041357172653079)),(to_sfixed_a(0.00014114679652266204)),(to_sfixed_a(0.00020917298388667405)),(to_sfixed_a(-0.00024310324806720018)),(to_sfixed_a(-0.00013543825480155647)),(to_sfixed_a(-1.3888886314816773e-05)),(to_sfixed_a(0.00012178636825410649)),(to_sfixed_a(-0.07359017431735992)),(to_sfixed_a(0.0028045601211488247)),(to_sfixed_a(0.006304866634309292)),(to_sfixed_a(0.19820399582386017)),(to_sfixed_a(0.0061503248289227486)),(to_sfixed_a(-2.9517905204556882e-06)),(to_sfixed_a(0.00018111195822712034)),(to_sfixed_a(0.0001313537359237671)),(to_sfixed_a(0.00011613059905357659)),(to_sfixed_a(-3.7165882531553507e-06)),(to_sfixed_a(0.0018013805383816361)),(to_sfixed_a(0.0012740353122353554)),(to_sfixed_a(0.009079089388251305)),(to_sfixed_a(0.00013693308574147522)),(to_sfixed_a(-0.00010632853081915528)),(to_sfixed_a(0.00011694643762893975)),(to_sfixed_a(-0.00011708207603078336)),(to_sfixed_a(-0.21656183898448944)),(to_sfixed_a(0.4180038273334503)),(to_sfixed_a(6.82683166814968e-05)),(to_sfixed_a(7.043189543765038e-05)),(to_sfixed_a(-0.00017579461564309895)),(to_sfixed_a(-0.008641502819955349)),(to_sfixed_a(-0.5241380929946899)),(to_sfixed_a(-0.02294306270778179)),(to_sfixed_a(-0.00024702047812752426)),(to_sfixed_a(6.328814197331667e-05)),(to_sfixed_a(0.00024754676269367337)),(to_sfixed_a(0.40734177827835083)),(to_sfixed_a(0.00017671337991487235)),(to_sfixed_a(0.29244551062583923)),(to_sfixed_a(0.0003113001585006714)),(to_sfixed_a(0.0005520649719983339)),(to_sfixed_a(0.00022894922585692257)),(to_sfixed_a(-0.0017913791816681623)),(to_sfixed_a(-0.00020629260689020157)),(to_sfixed_a(0.0028178938664495945)),(to_sfixed_a(-6.918936560396105e-05)),(to_sfixed_a(0.03890189155936241)),(to_sfixed_a(0.00030437635723501444)),(to_sfixed_a(0.43339523673057556)),(to_sfixed_a(-0.3745378255844116)),(to_sfixed_a(0.00015457702102139592)),(to_sfixed_a(0.5567164421081543)),(to_sfixed_a(-0.00014385581016540527)),(to_sfixed_a(0.00011209452350158244)),(to_sfixed_a(0.001987193478271365)),(to_sfixed_a(2.3742733901599422e-05)),(to_sfixed_a(0.00012145684740971774)),(to_sfixed_a(0.0015074880793690681)),(to_sfixed_a(0.012864715419709682)),(to_sfixed_a(-0.00013342400779947639)),(to_sfixed_a(-3.8787227822467685e-05)),(to_sfixed_a(-3.645571996457875e-05)),(to_sfixed_a(3.700701199704781e-05)),(to_sfixed_a(-0.0021217174362391233)),(to_sfixed_a(0.0001307059428654611)),(to_sfixed_a(2.1322664906620048e-05)),(to_sfixed_a(0.00010091083095176145)),(to_sfixed_a(0.003245830535888672)),(to_sfixed_a(0.00011309992987662554)),(to_sfixed_a(3.942806870327331e-05)),(to_sfixed_a(3.0407783924601972e-05)),(to_sfixed_a(-0.0033470885828137398)),(to_sfixed_a(0.001068080309778452)),(to_sfixed_a(6.857725384179503e-05)),(to_sfixed_a(1.8433966033626348e-05)),(to_sfixed_a(7.201131666079164e-05)),(to_sfixed_a(-2.7588685043156147e-06)),(to_sfixed_a(-0.26120421290397644)),(to_sfixed_a(0.0002150143845938146)),(to_sfixed_a(0.001639647758565843)),(to_sfixed_a(-0.0033018249087035656)),(to_sfixed_a(0.0005976497777737677)),(to_sfixed_a(-5.338137270882726e-06)),(to_sfixed_a(0.00030751776648685336)),(to_sfixed_a(0.0002425355778541416)),(to_sfixed_a(0.002980974968522787)),(to_sfixed_a(0.00016807977226562798)),(to_sfixed_a(1.2641045032069087e-05)),(to_sfixed_a(0.0025607000570744276)),(to_sfixed_a(0.00043749914038926363)),(to_sfixed_a(2.4211993149947375e-05)),(to_sfixed_a(-0.0037261738907545805)),(to_sfixed_a(0.0012862918665632606)),(to_sfixed_a(-0.0011052817571908236)),(to_sfixed_a(-0.3081550896167755)),(to_sfixed_a(-5.587278792518191e-05)),(to_sfixed_a(0.0021579815074801445)),(to_sfixed_a(3.2319770980393514e-05)),(to_sfixed_a(-0.0011727079981938004)),(to_sfixed_a(6.424381717806682e-05)),(to_sfixed_a(-0.0038848326075822115)),(to_sfixed_a(0.2457418143749237)),(to_sfixed_a(-1.72312356880866e-05)));

    constant weight_n2_19 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.030354389920830727)),(to_sfixed_a(1.1503332643769681e-05)),(to_sfixed_a(2.4618408133392222e-05)),(to_sfixed_a(-0.00015173041902016848)),(to_sfixed_a(1.238757249666378e-06)),(to_sfixed_a(-3.117202140856534e-05)),(to_sfixed_a(-9.911289089359343e-05)),(to_sfixed_a(-6.94193149683997e-05)),(to_sfixed_a(-0.00013378328003454953)),(to_sfixed_a(-0.00020342535572126508)),(to_sfixed_a(-1.2022617738693953e-05)),(to_sfixed_a(0.0002938294783234596)),(to_sfixed_a(0.0002984096063300967)),(to_sfixed_a(6.567055243067443e-05)),(to_sfixed_a(-0.0001995065395021811)),(to_sfixed_a(0.00014621323498431593)),(to_sfixed_a(-7.761360029689968e-05)),(to_sfixed_a(-6.753373600076884e-05)),(to_sfixed_a(3.738015948329121e-06)),(to_sfixed_a(0.0001060142312780954)),(to_sfixed_a(-0.0001066826080204919)),(to_sfixed_a(-0.0002077385870506987)),(to_sfixed_a(-0.0001498024066677317)),(to_sfixed_a(1.1761108908103779e-05)),(to_sfixed_a(0.00018881616415455937)),(to_sfixed_a(-0.00013494878658093512)),(to_sfixed_a(-1.3121658412273973e-05)),(to_sfixed_a(-3.203153028152883e-05)),(to_sfixed_a(-0.00041445111855864525)),(to_sfixed_a(-0.0002961145364679396)),(to_sfixed_a(0.0003176068712491542)),(to_sfixed_a(0.00024000491248443723)),(to_sfixed_a(0.0002393985487287864)),(to_sfixed_a(-0.00015001845895312726)),(to_sfixed_a(8.439296652795747e-05)),(to_sfixed_a(-1.149830495705828e-06)),(to_sfixed_a(-0.00015331579197663814)),(to_sfixed_a(0.00015758773952256888)),(to_sfixed_a(-4.3016349081881344e-05)),(to_sfixed_a(-4.8122063162736595e-05)),(to_sfixed_a(0.00010866271622944623)),(to_sfixed_a(-1.3290366041474044e-05)),(to_sfixed_a(-2.9826187528669834e-05)),(to_sfixed_a(-0.00025449326494708657)),(to_sfixed_a(0.00011413544416427612)),(to_sfixed_a(-6.210010906215757e-05)),(to_sfixed_a(-0.0001681262074271217)),(to_sfixed_a(-0.0001386279909638688)),(to_sfixed_a(6.716213829349726e-05)),(to_sfixed_a(-5.022536788601428e-05)),(to_sfixed_a(-4.8718880861997604e-05)),(to_sfixed_a(6.520995520986617e-05)),(to_sfixed_a(-0.00016490957932546735)),(to_sfixed_a(-0.00015428612823598087)),(to_sfixed_a(-4.862415516981855e-05)),(to_sfixed_a(-0.0002558989799581468)),(to_sfixed_a(0.0001050726423272863)),(to_sfixed_a(5.978708577458747e-05)),(to_sfixed_a(2.270994991704356e-05)),(to_sfixed_a(-7.900466152932495e-05)),(to_sfixed_a(-7.130931771825999e-05)),(to_sfixed_a(-9.785335714695975e-05)),(to_sfixed_a(0.00015593560237903148)),(to_sfixed_a(-2.7555215638130903e-06)),(to_sfixed_a(-6.870503420941532e-05)),(to_sfixed_a(-9.048875654116273e-06)),(to_sfixed_a(-9.316577052231878e-05)),(to_sfixed_a(-0.00015567464288324118)),(to_sfixed_a(0.00017452739120926708)),(to_sfixed_a(-2.3480017262045294e-05)),(to_sfixed_a(-7.93610088294372e-05)),(to_sfixed_a(0.00011231630196562037)),(to_sfixed_a(-8.493576751789078e-05)),(to_sfixed_a(6.588128599105403e-05)),(to_sfixed_a(0.00014912454935256392)),(to_sfixed_a(6.328276504063979e-05)),(to_sfixed_a(7.030779670458287e-05)),(to_sfixed_a(-1.7574813682585955e-05)),(to_sfixed_a(0.0002843069960363209)),(to_sfixed_a(4.1942912503145635e-06)),(to_sfixed_a(7.06103746779263e-05)),(to_sfixed_a(-3.755269790417515e-05)),(to_sfixed_a(-0.00011320567864459008)),(to_sfixed_a(-1.8549355445429683e-05)),(to_sfixed_a(-3.224237298127264e-05)),(to_sfixed_a(0.00011694336717482656)),(to_sfixed_a(4.2322735680500045e-05)),(to_sfixed_a(-0.0002607146161608398)),(to_sfixed_a(0.0001835150906117633)),(to_sfixed_a(4.2782641685334966e-05)),(to_sfixed_a(7.18440132914111e-05)),(to_sfixed_a(-4.7128283767960966e-05)),(to_sfixed_a(-0.0001684640592429787)),(to_sfixed_a(-6.852390652056783e-05)),(to_sfixed_a(0.00018722336972132325)),(to_sfixed_a(-0.00011490716133266687)),(to_sfixed_a(0.00015446079487446696)),(to_sfixed_a(-0.00013909909466747195)),(to_sfixed_a(-0.00014599772111978382)),(to_sfixed_a(-4.264294693712145e-05)),(to_sfixed_a(-0.00011351686407579109)),(to_sfixed_a(-0.0001433981815353036)),(to_sfixed_a(0.0001416931045241654)),(to_sfixed_a(-7.145506970118731e-05)),(to_sfixed_a(-0.0001307434868067503)),(to_sfixed_a(0.0001966639538295567)),(to_sfixed_a(-5.72458520764485e-06)),(to_sfixed_a(-7.132376049412414e-05)),(to_sfixed_a(3.1625659175915644e-05)),(to_sfixed_a(9.553147538099438e-05)),(to_sfixed_a(8.473169873468578e-05)),(to_sfixed_a(-0.00012734670599456877)),(to_sfixed_a(0.000155641304445453)),(to_sfixed_a(8.663117478135973e-05)),(to_sfixed_a(-2.29033685172908e-05)),(to_sfixed_a(2.074041185551323e-05)),(to_sfixed_a(-0.00019547116244211793)),(to_sfixed_a(1.7227648640982807e-05)),(to_sfixed_a(-0.0001849496184149757)),(to_sfixed_a(-6.378706893883646e-05)),(to_sfixed_a(0.00013454037252813578)),(to_sfixed_a(7.410162652377039e-07)),(to_sfixed_a(-7.083226955728605e-05)),(to_sfixed_a(-0.0001473149168305099)),(to_sfixed_a(6.2398481532e-05)),(to_sfixed_a(0.00010393172124167904)),(to_sfixed_a(-0.00029499002266675234)),(to_sfixed_a(-0.00019659263489302248)),(to_sfixed_a(1.2705917470157146e-05)),(to_sfixed_a(0.00015587816596962512)),(to_sfixed_a(-0.00025638192892074585)),(to_sfixed_a(-0.00018216919852420688)),(to_sfixed_a(0.00010195496724918485)),(to_sfixed_a(-0.00031225892598740757)),(to_sfixed_a(0.00027749978471547365)),(to_sfixed_a(-0.00013617149670608342)),(to_sfixed_a(-4.700099816545844e-05)),(to_sfixed_a(6.687457789666951e-05)),(to_sfixed_a(5.9025478549301624e-06)),(to_sfixed_a(6.177095201564953e-05)),(to_sfixed_a(-7.077332702465355e-05)),(to_sfixed_a(0.00015629289555363357)),(to_sfixed_a(-4.241868737153709e-06)),(to_sfixed_a(-0.00015662792429793626)),(to_sfixed_a(0.00029693773831240833)),(to_sfixed_a(-0.00014068983728066087)),(to_sfixed_a(-2.3786689780536108e-05)),(to_sfixed_a(-1.0679927072487772e-05)),(to_sfixed_a(0.00021300320804584771)),(to_sfixed_a(9.247937850886956e-05)),(to_sfixed_a(6.058865619706921e-05)),(to_sfixed_a(1.2458694982342422e-05)),(to_sfixed_a(0.00012199316552141681)),(to_sfixed_a(0.00010057346662506461)),(to_sfixed_a(0.00013606056745629758)),(to_sfixed_a(-2.439538366161287e-05)),(to_sfixed_a(-0.00024326209677383304)),(to_sfixed_a(7.420592737616971e-06)),(to_sfixed_a(1.5609308320563287e-05)),(to_sfixed_a(-0.00011348195403115824)),(to_sfixed_a(-0.00010686731548048556)),(to_sfixed_a(-0.0002001140092033893)),(to_sfixed_a(-0.0001044836244545877)),(to_sfixed_a(5.916136797168292e-05)),(to_sfixed_a(9.233829041477293e-05)),(to_sfixed_a(-3.162426583003253e-05)),(to_sfixed_a(0.00016032400890253484)),(to_sfixed_a(-6.64121616864577e-05)),(to_sfixed_a(0.0002491131308488548)),(to_sfixed_a(0.00010616573854349554)),(to_sfixed_a(5.827502172905952e-05)),(to_sfixed_a(4.770320083480328e-05)),(to_sfixed_a(-1.7846810806076974e-05)),(to_sfixed_a(0.0001543753023725003)),(to_sfixed_a(6.895892147440463e-05)),(to_sfixed_a(3.842976730084047e-05)),(to_sfixed_a(0.00030943070305511355)),(to_sfixed_a(-0.00024351946194656193)),(to_sfixed_a(0.0001824472565203905)),(to_sfixed_a(0.00012772614718414843)),(to_sfixed_a(-0.00011346889368724078)),(to_sfixed_a(6.920999294379726e-05)),(to_sfixed_a(1.0564399417489767e-05)),(to_sfixed_a(-1.2512857210822403e-05)),(to_sfixed_a(-0.0001520538644399494)),(to_sfixed_a(-6.788087193854153e-05)),(to_sfixed_a(-2.5826477212831378e-05)),(to_sfixed_a(-1.6793062968645245e-05)),(to_sfixed_a(-2.425908314762637e-05)),(to_sfixed_a(0.0002355395699851215)),(to_sfixed_a(-0.00020034192129969597)),(to_sfixed_a(0.0002843195106834173)),(to_sfixed_a(1.3770441000815481e-05)),(to_sfixed_a(0.0001166837610071525)),(to_sfixed_a(-4.420089680934325e-06)),(to_sfixed_a(-3.144755100947805e-05)),(to_sfixed_a(0.00029510827152989805)),(to_sfixed_a(0.00022691194317303598)),(to_sfixed_a(0.00016677613893989474)),(to_sfixed_a(-2.3517233785241842e-05)),(to_sfixed_a(-1.62241849466227e-05)),(to_sfixed_a(-0.00010199873213423416)),(to_sfixed_a(7.322536839637905e-05)),(to_sfixed_a(-0.00025040912441909313)),(to_sfixed_a(1.9198632799088955e-05)),(to_sfixed_a(-2.7472902729641646e-05)),(to_sfixed_a(6.654502067249268e-05)),(to_sfixed_a(-0.00020334876899141818)),(to_sfixed_a(-5.762580985901877e-05)),(to_sfixed_a(4.32590240961872e-06)),(to_sfixed_a(6.993820716161281e-05)),(to_sfixed_a(0.0001505925611127168)),(to_sfixed_a(2.3996097297640517e-05)),(to_sfixed_a(6.817071698606014e-05)),(to_sfixed_a(0.00028365309117361903)),(to_sfixed_a(0.00016191510076168925)),(to_sfixed_a(2.43351241806522e-05)),(to_sfixed_a(0.00020498831872828305)),(to_sfixed_a(4.384433850646019e-05)),(to_sfixed_a(-0.00014022899267729372)),(to_sfixed_a(-2.2999593056738377e-06)),(to_sfixed_a(-0.000169175022165291)),(to_sfixed_a(-0.00020156842947471887)),(to_sfixed_a(-8.332085417350754e-05)),(to_sfixed_a(2.95500285574235e-07)),(to_sfixed_a(1.8632083083502948e-05)),(to_sfixed_a(-0.00030393904307857156)),(to_sfixed_a(-6.0004109400324523e-05)),(to_sfixed_a(-0.00016824026533868164)),(to_sfixed_a(-0.00024284841492772102)),(to_sfixed_a(6.316036160569638e-05)),(to_sfixed_a(-5.480393519974314e-05)),(to_sfixed_a(0.00011629384243860841)),(to_sfixed_a(-0.0002897893136832863)),(to_sfixed_a(0.00013607944129034877)),(to_sfixed_a(-0.00018180120969191194)),(to_sfixed_a(0.00011557860852917656)),(to_sfixed_a(-0.00015586716472171247)),(to_sfixed_a(6.920317537151277e-05)),(to_sfixed_a(0.00015628139954060316)),(to_sfixed_a(-0.00014820882643107325)),(to_sfixed_a(4.585417627822608e-07)),(to_sfixed_a(0.0001131839380832389)),(to_sfixed_a(-0.0002760272764135152)),(to_sfixed_a(7.403705239994451e-07)),(to_sfixed_a(-6.100473183323629e-05)),(to_sfixed_a(-6.796409434173256e-05)),(to_sfixed_a(2.1159619791433215e-05)),(to_sfixed_a(-0.00011925465514650568)),(to_sfixed_a(4.410148176248185e-05)),(to_sfixed_a(-7.883551734266803e-05)),(to_sfixed_a(3.4051205147989094e-05)),(to_sfixed_a(-4.933491436531767e-05)),(to_sfixed_a(-0.00015555947902612388)),(to_sfixed_a(-0.00010571871825959533)),(to_sfixed_a(-0.00024171939003281295)),(to_sfixed_a(0.0001486503315391019)),(to_sfixed_a(0.00011175795225426555)),(to_sfixed_a(0.0001023227086989209)),(to_sfixed_a(0.00011172040103701875)),(to_sfixed_a(3.244165418436751e-05)),(to_sfixed_a(-4.508794518187642e-06)),(to_sfixed_a(8.145150059135631e-05)),(to_sfixed_a(9.790048352442682e-05)),(to_sfixed_a(0.00015105049533303827)),(to_sfixed_a(6.94192131049931e-05)),(to_sfixed_a(2.3836983018554747e-06)),(to_sfixed_a(-0.00028669394669122994)),(to_sfixed_a(4.2802970710908994e-05)),(to_sfixed_a(0.00026598008116707206)),(to_sfixed_a(0.00018023625307250768)),(to_sfixed_a(0.0002203962067142129)),(to_sfixed_a(6.993986607994884e-05)),(to_sfixed_a(0.0001362282200716436)),(to_sfixed_a(-0.00023683623294346035)),(to_sfixed_a(4.428097599884495e-05)),(to_sfixed_a(-0.0001784935884643346)),(to_sfixed_a(4.614714998751879e-05)),(to_sfixed_a(-6.844595191068947e-05)),(to_sfixed_a(-7.656846719328314e-06)),(to_sfixed_a(8.480052929371595e-05)),(to_sfixed_a(4.007056122645736e-05)),(to_sfixed_a(-0.00011681900650728494)),(to_sfixed_a(-0.00018639134941622615)),(to_sfixed_a(0.0003224255924578756)),(to_sfixed_a(0.00011785042443079874)),(to_sfixed_a(5.935298395343125e-05)),(to_sfixed_a(4.45819714514073e-05)),(to_sfixed_a(0.00010680139530450106)),(to_sfixed_a(-1.1230982636334375e-05)),(to_sfixed_a(-1.3432276318781078e-05)),(to_sfixed_a(7.739081047475338e-05)),(to_sfixed_a(-0.00010551894956734031)),(to_sfixed_a(0.00027120683807879686)),(to_sfixed_a(-7.155630737543106e-05)),(to_sfixed_a(-0.00011362443183315918)),(to_sfixed_a(0.00018951940000988543)),(to_sfixed_a(-0.00010825772915268317)),(to_sfixed_a(6.197166658239439e-05)),(to_sfixed_a(-0.00018150036339648068)),(to_sfixed_a(0.0002315168094355613)));

    constant weight_n2_20 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.05833280459046364)),(to_sfixed_a(-0.0015068576904013753)),(to_sfixed_a(-0.00038345844950526953)),(to_sfixed_a(-5.7383193052373827e-05)),(to_sfixed_a(0.018746929243206978)),(to_sfixed_a(-2.2767137124901637e-05)),(to_sfixed_a(-0.003732645185664296)),(to_sfixed_a(-4.72497777082026e-06)),(to_sfixed_a(0.0002872672048397362)),(to_sfixed_a(6.083962944103405e-06)),(to_sfixed_a(1.1446907592471689e-05)),(to_sfixed_a(0.29532840847969055)),(to_sfixed_a(-0.6044324636459351)),(to_sfixed_a(-3.439421925577335e-05)),(to_sfixed_a(7.20290991012007e-05)),(to_sfixed_a(-6.557017331942916e-05)),(to_sfixed_a(0.005732452031224966)),(to_sfixed_a(-0.00029788960819132626)),(to_sfixed_a(-0.002391657093539834)),(to_sfixed_a(0.2502075731754303)),(to_sfixed_a(1.2027107004541904e-05)),(to_sfixed_a(-2.120773569913581e-05)),(to_sfixed_a(-0.00014841571100987494)),(to_sfixed_a(0.0018343423726037145)),(to_sfixed_a(0.002552544930949807)),(to_sfixed_a(-0.018488658592104912)),(to_sfixed_a(-0.00017844296235125512)),(to_sfixed_a(-6.491360545624048e-05)),(to_sfixed_a(-6.818564725108445e-05)),(to_sfixed_a(4.749758227262646e-05)),(to_sfixed_a(-0.003683921415358782)),(to_sfixed_a(6.5320637077093124e-06)),(to_sfixed_a(-0.007657101843506098)),(to_sfixed_a(0.00018345692660659552)),(to_sfixed_a(-0.0001277739938814193)),(to_sfixed_a(-7.895999442553148e-05)),(to_sfixed_a(-0.016133485361933708)),(to_sfixed_a(-0.2137739360332489)),(to_sfixed_a(-0.4382803738117218)),(to_sfixed_a(-0.00016826263163238764)),(to_sfixed_a(-0.47434213757514954)),(to_sfixed_a(-3.853629095829092e-05)),(to_sfixed_a(0.00017556996317580342)),(to_sfixed_a(1.4665216440334916e-05)),(to_sfixed_a(-0.015045469626784325)),(to_sfixed_a(-0.01788225583732128)),(to_sfixed_a(-0.23914285004138947)),(to_sfixed_a(-0.0013194887433201075)),(to_sfixed_a(0.00018716728664003313)),(to_sfixed_a(3.468750583124347e-05)),(to_sfixed_a(0.010240988805890083)),(to_sfixed_a(-0.00045883451821282506)),(to_sfixed_a(0.0001034827801049687)),(to_sfixed_a(-0.0007762814639136195)),(to_sfixed_a(-0.007429901044815779)),(to_sfixed_a(0.011017544195055962)),(to_sfixed_a(7.119608926586807e-05)),(to_sfixed_a(-0.007903982885181904)),(to_sfixed_a(0.0002320054773008451)),(to_sfixed_a(-7.11499887984246e-05)),(to_sfixed_a(-0.008815284818410873)),(to_sfixed_a(-0.0004357877769507468)),(to_sfixed_a(-4.126311978325248e-05)),(to_sfixed_a(-0.0043145278468728065)),(to_sfixed_a(-0.000297871622024104)),(to_sfixed_a(0.2052830308675766)),(to_sfixed_a(1.6126759874168783e-05)),(to_sfixed_a(-5.257257726043463e-06)),(to_sfixed_a(0.00021221398492343724)),(to_sfixed_a(2.255873187095858e-05)),(to_sfixed_a(0.005213416181504726)),(to_sfixed_a(0.033537011593580246)),(to_sfixed_a(-0.31361672282218933)),(to_sfixed_a(-0.0002543198934290558)),(to_sfixed_a(-4.5425233111018315e-05)),(to_sfixed_a(9.768715244717896e-06)),(to_sfixed_a(0.0006083441548980772)),(to_sfixed_a(-0.0009822164429351687)),(to_sfixed_a(-1.265540049644187e-06)),(to_sfixed_a(-0.008379537612199783)),(to_sfixed_a(-0.008605836890637875)),(to_sfixed_a(0.00014913898485247046)),(to_sfixed_a(-0.0004770748200826347)),(to_sfixed_a(-0.0011255685240030289)),(to_sfixed_a(-0.00019890557450708002)),(to_sfixed_a(0.0027159324381500483)),(to_sfixed_a(-0.010577956214547157)),(to_sfixed_a(3.867860414175084e-06)),(to_sfixed_a(-9.574090654496104e-06)),(to_sfixed_a(4.4046413677278906e-05)),(to_sfixed_a(-0.008256006985902786)),(to_sfixed_a(0.0001297735725529492)),(to_sfixed_a(-0.00875068362802267)),(to_sfixed_a(0.0002435243222862482)),(to_sfixed_a(-0.002829036908224225)),(to_sfixed_a(5.853189941262826e-05)),(to_sfixed_a(7.153532351367176e-06)),(to_sfixed_a(-0.00015558252925984561)),(to_sfixed_a(0.00011692081898218021)),(to_sfixed_a(-9.949792001862079e-06)),(to_sfixed_a(0.5258280038833618)),(to_sfixed_a(-0.003952413331717253)),(to_sfixed_a(-3.405650204513222e-06)),(to_sfixed_a(0.412801593542099)),(to_sfixed_a(0.011302361264824867)),(to_sfixed_a(-3.0488341508316807e-05)),(to_sfixed_a(-0.00029791926499456167)),(to_sfixed_a(-0.00013007139205001295)),(to_sfixed_a(0.000156334979692474)),(to_sfixed_a(-0.009081324562430382)),(to_sfixed_a(-0.002240424044430256)),(to_sfixed_a(0.00013645562285091728)),(to_sfixed_a(-0.010070535354316235)),(to_sfixed_a(7.37010850571096e-05)),(to_sfixed_a(-0.00017945480067282915)),(to_sfixed_a(0.18302571773529053)),(to_sfixed_a(-0.00026735267601907253)),(to_sfixed_a(0.25523263216018677)),(to_sfixed_a(0.00013373249385040253)),(to_sfixed_a(0.00013277391553856432)),(to_sfixed_a(0.00018045102478936315)),(to_sfixed_a(0.000238678403547965)),(to_sfixed_a(-0.030031718313694)),(to_sfixed_a(6.970307003939524e-05)),(to_sfixed_a(0.00024877398391254246)),(to_sfixed_a(0.21239984035491943)),(to_sfixed_a(0.04256918653845787)),(to_sfixed_a(6.68353313812986e-05)),(to_sfixed_a(-8.333328878507018e-06)),(to_sfixed_a(2.0632367522921413e-05)),(to_sfixed_a(3.133009158773348e-07)),(to_sfixed_a(-5.808683636132628e-05)),(to_sfixed_a(1.2153512216173112e-05)),(to_sfixed_a(-0.01101878471672535)),(to_sfixed_a(0.00018364925927016884)),(to_sfixed_a(6.948801456019282e-05)),(to_sfixed_a(-0.026591850444674492)),(to_sfixed_a(-1.3085725640848977e-06)),(to_sfixed_a(0.00015424239973071963)),(to_sfixed_a(0.00010676569945644587)),(to_sfixed_a(-0.005483683664351702)),(to_sfixed_a(0.0001994068588828668)),(to_sfixed_a(0.00010575616033747792)),(to_sfixed_a(0.5075724720954895)),(to_sfixed_a(-3.7191704905126244e-05)),(to_sfixed_a(-6.44562387606129e-05)),(to_sfixed_a(-6.830775237176567e-05)),(to_sfixed_a(1.9012244592886418e-05)),(to_sfixed_a(0.00015344312123488635)),(to_sfixed_a(-0.00013453378051053733)),(to_sfixed_a(-4.168541636317968e-06)),(to_sfixed_a(1.7149672203231603e-05)),(to_sfixed_a(0.003239395096898079)),(to_sfixed_a(2.2675827494822443e-05)),(to_sfixed_a(0.00011663679470075294)),(to_sfixed_a(-0.034393299371004105)),(to_sfixed_a(1.6929458070080727e-05)),(to_sfixed_a(9.001805301522836e-05)),(to_sfixed_a(0.00012177578901173547)),(to_sfixed_a(-9.885759936878458e-05)),(to_sfixed_a(-4.231923958286643e-05)),(to_sfixed_a(7.142439426388592e-05)),(to_sfixed_a(-0.001016368973068893)),(to_sfixed_a(-0.00021969930094201118)),(to_sfixed_a(0.002990104490891099)),(to_sfixed_a(5.104897718410939e-05)),(to_sfixed_a(5.5047436035238206e-05)),(to_sfixed_a(-0.38574397563934326)),(to_sfixed_a(-0.00011634801921900362)),(to_sfixed_a(-0.00010804138582898304)),(to_sfixed_a(0.0009522369364276528)),(to_sfixed_a(-3.0893274924892467e-06)),(to_sfixed_a(-0.33521750569343567)),(to_sfixed_a(3.0686744139529765e-05)),(to_sfixed_a(-0.002632041461765766)),(to_sfixed_a(0.002298298990353942)),(to_sfixed_a(0.0009485968039371073)),(to_sfixed_a(0.0003232004528399557)),(to_sfixed_a(0.24041426181793213)),(to_sfixed_a(-0.015240120701491833)),(to_sfixed_a(-0.001011288957670331)),(to_sfixed_a(0.0034641099628061056)),(to_sfixed_a(-0.00012883005547337234)),(to_sfixed_a(1.246358806383796e-06)),(to_sfixed_a(0.00025098654441535473)),(to_sfixed_a(-0.0003699742374010384)),(to_sfixed_a(-0.044295139610767365)),(to_sfixed_a(-0.00012457506090868264)),(to_sfixed_a(3.0317241908051074e-06)),(to_sfixed_a(-0.00014990291674621403)),(to_sfixed_a(-4.578940206556581e-06)),(to_sfixed_a(0.0001020268100546673)),(to_sfixed_a(-0.29888367652893066)),(to_sfixed_a(-0.007353680208325386)),(to_sfixed_a(0.00011467618605820462)),(to_sfixed_a(0.013667520135641098)),(to_sfixed_a(-9.754876373335719e-08)),(to_sfixed_a(-0.0027464195154607296)),(to_sfixed_a(0.6093331575393677)),(to_sfixed_a(7.1741160354577e-05)),(to_sfixed_a(-0.00016746277105994523)),(to_sfixed_a(7.087266567396e-05)),(to_sfixed_a(-3.7539692129939795e-05)),(to_sfixed_a(-0.00015261377848219126)),(to_sfixed_a(-0.00025544792879372835)),(to_sfixed_a(-0.00017296665464527905)),(to_sfixed_a(0.0002445357677061111)),(to_sfixed_a(0.015238718129694462)),(to_sfixed_a(-0.001087714685127139)),(to_sfixed_a(-0.0009410511120222509)),(to_sfixed_a(-0.00013312922965269536)),(to_sfixed_a(7.035923772491515e-05)),(to_sfixed_a(-0.00029682391323149204)),(to_sfixed_a(3.645320248324424e-05)),(to_sfixed_a(-0.00026368716498836875)),(to_sfixed_a(-0.0004560399684123695)),(to_sfixed_a(-4.503972377278842e-07)),(to_sfixed_a(-0.0029281843453645706)),(to_sfixed_a(-0.6774504780769348)),(to_sfixed_a(0.00014675241254735738)),(to_sfixed_a(-1.53512810356915e-05)),(to_sfixed_a(-0.0002366574335610494)),(to_sfixed_a(-7.984059629961848e-05)),(to_sfixed_a(8.270279067801312e-05)),(to_sfixed_a(0.12654277682304382)),(to_sfixed_a(6.874487007735297e-05)),(to_sfixed_a(-1.8708888092078269e-06)),(to_sfixed_a(6.80333178024739e-05)),(to_sfixed_a(0.3510279357433319)),(to_sfixed_a(-0.0009206623653881252)),(to_sfixed_a(-0.41489923000335693)),(to_sfixed_a(-0.00013977849448565394)),(to_sfixed_a(-0.00022266706218943)),(to_sfixed_a(0.00029112922493368387)),(to_sfixed_a(-0.01029240619391203)),(to_sfixed_a(-0.004411395639181137)),(to_sfixed_a(0.005565195344388485)),(to_sfixed_a(-7.096541958162561e-05)),(to_sfixed_a(-0.004522284027189016)),(to_sfixed_a(0.00015882967272773385)),(to_sfixed_a(-0.00459122471511364)),(to_sfixed_a(-8.74967809068039e-05)),(to_sfixed_a(0.003902989672496915)),(to_sfixed_a(-8.927301678340882e-06)),(to_sfixed_a(0.00011860043741762638)),(to_sfixed_a(-0.006347841117531061)),(to_sfixed_a(0.31301721930503845)),(to_sfixed_a(-0.0028752791695296764)),(to_sfixed_a(6.929671508260071e-05)),(to_sfixed_a(-0.017677655443549156)),(to_sfixed_a(0.0023595334496349096)),(to_sfixed_a(-8.778877963777632e-05)),(to_sfixed_a(4.137886571697891e-05)),(to_sfixed_a(-4.037559847347438e-06)),(to_sfixed_a(-0.0006360769621096551)),(to_sfixed_a(-0.0006170155829750001)),(to_sfixed_a(-0.3145052194595337)),(to_sfixed_a(-0.00022601752425543964)),(to_sfixed_a(-0.00024403762654401362)),(to_sfixed_a(-0.0088521558791399)),(to_sfixed_a(0.00028917487361468375)),(to_sfixed_a(-0.6459257006645203)),(to_sfixed_a(-0.00010913654114119709)),(to_sfixed_a(-0.001371067832224071)),(to_sfixed_a(2.1409250621218234e-06)),(to_sfixed_a(-0.26197102665901184)),(to_sfixed_a(-1.1452357284724712e-08)),(to_sfixed_a(-0.0002513169893063605)),(to_sfixed_a(8.29362979857251e-05)),(to_sfixed_a(-0.002610960975289345)),(to_sfixed_a(-0.006535954307764769)),(to_sfixed_a(0.00011422758689150214)),(to_sfixed_a(6.018214480718598e-05)),(to_sfixed_a(-0.0001562247343827039)),(to_sfixed_a(0.0001506324188085273)),(to_sfixed_a(0.0013637846568599343)),(to_sfixed_a(0.05286416783928871)),(to_sfixed_a(-0.25193002820014954)),(to_sfixed_a(-0.4215124845504761)),(to_sfixed_a(-0.00152147701010108)),(to_sfixed_a(0.0001975304912775755)),(to_sfixed_a(-0.00045566027984023094)),(to_sfixed_a(-0.00013588901492767036)),(to_sfixed_a(-0.0010904842056334019)),(to_sfixed_a(-5.725491791963577e-05)),(to_sfixed_a(-2.305045200046152e-05)),(to_sfixed_a(9.60202596616e-05)),(to_sfixed_a(0.00047670258209109306)),(to_sfixed_a(-0.0001343608892057091)),(to_sfixed_a(0.35366564989089966)),(to_sfixed_a(-0.00040356075624004006)),(to_sfixed_a(0.0006395956734195352)),(to_sfixed_a(-0.003784327767789364)),(to_sfixed_a(0.00012829310435336083)),(to_sfixed_a(-0.0015212839934974909)),(to_sfixed_a(-0.0020954543724656105)),(to_sfixed_a(-0.1366277039051056)),(to_sfixed_a(-0.00019980872457381338)),(to_sfixed_a(-0.6125065684318542)),(to_sfixed_a(0.05897027254104614)),(to_sfixed_a(-0.011088673956692219)));

    constant weight_n2_21 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.35052937269210815)),(to_sfixed_a(0.011200456880033016)),(to_sfixed_a(0.0009181358618661761)),(to_sfixed_a(-6.793495413148776e-05)),(to_sfixed_a(0.0011149777565151453)),(to_sfixed_a(-9.715491614770144e-06)),(to_sfixed_a(0.054456960409879684)),(to_sfixed_a(1.3571640010923147e-05)),(to_sfixed_a(1.5720725059509277e-05)),(to_sfixed_a(6.33781892247498e-05)),(to_sfixed_a(0.00014735983859281987)),(to_sfixed_a(-0.0011124046286568046)),(to_sfixed_a(-0.23306559026241302)),(to_sfixed_a(0.0015415949746966362)),(to_sfixed_a(6.838783156126738e-05)),(to_sfixed_a(-0.0001168213493656367)),(to_sfixed_a(0.1940128356218338)),(to_sfixed_a(-3.709793963935226e-05)),(to_sfixed_a(0.47905412316322327)),(to_sfixed_a(-0.022535083815455437)),(to_sfixed_a(0.00013646367006003857)),(to_sfixed_a(0.00015383557183668017)),(to_sfixed_a(-0.0005246838554739952)),(to_sfixed_a(-0.0002544985618442297)),(to_sfixed_a(0.04088997468352318)),(to_sfixed_a(0.010348515585064888)),(to_sfixed_a(-5.136233812663704e-05)),(to_sfixed_a(-3.271513196523301e-05)),(to_sfixed_a(0.014445382170379162)),(to_sfixed_a(-3.0029397748876363e-05)),(to_sfixed_a(-0.23518577218055725)),(to_sfixed_a(-2.533318183850497e-05)),(to_sfixed_a(0.36615607142448425)),(to_sfixed_a(0.0004459570918697864)),(to_sfixed_a(1.5953904949128628e-05)),(to_sfixed_a(-0.00018753745825961232)),(to_sfixed_a(-0.10876451432704926)),(to_sfixed_a(-0.45946362614631653)),(to_sfixed_a(0.0041037206538021564)),(to_sfixed_a(-0.0002105365856550634)),(to_sfixed_a(-0.30140358209609985)),(to_sfixed_a(0.036736343055963516)),(to_sfixed_a(6.736465002177283e-05)),(to_sfixed_a(0.0001428655523341149)),(to_sfixed_a(-0.0014612453524023294)),(to_sfixed_a(0.007118646986782551)),(to_sfixed_a(0.23293925821781158)),(to_sfixed_a(0.23662303388118744)),(to_sfixed_a(0.00019457285816315562)),(to_sfixed_a(0.04107104241847992)),(to_sfixed_a(0.002718838397413492)),(to_sfixed_a(0.004590997006744146)),(to_sfixed_a(-0.00011277874000370502)),(to_sfixed_a(0.004797728266566992)),(to_sfixed_a(-0.04811994358897209)),(to_sfixed_a(-0.0009957941947504878)),(to_sfixed_a(-0.0001530037698103115)),(to_sfixed_a(0.0004647287423722446)),(to_sfixed_a(-0.0001697663974482566)),(to_sfixed_a(-0.00010361937893321738)),(to_sfixed_a(0.00017604786262381822)),(to_sfixed_a(0.0007155153434723616)),(to_sfixed_a(-0.0058293151669204235)),(to_sfixed_a(-0.3089049458503723)),(to_sfixed_a(0.0001558964140713215)),(to_sfixed_a(0.45258113741874695)),(to_sfixed_a(3.423976886551827e-05)),(to_sfixed_a(0.3313749134540558)),(to_sfixed_a(0.0014843761455267668)),(to_sfixed_a(-0.0002614112163428217)),(to_sfixed_a(0.005523469299077988)),(to_sfixed_a(-0.005307160317897797)),(to_sfixed_a(0.003850989742204547)),(to_sfixed_a(-0.0001520620717201382)),(to_sfixed_a(0.00020116707310080528)),(to_sfixed_a(-6.38831261312589e-05)),(to_sfixed_a(-0.016466302797198296)),(to_sfixed_a(0.0017631073715165257)),(to_sfixed_a(-0.000130283588077873)),(to_sfixed_a(-0.006443470250815153)),(to_sfixed_a(-3.3617907320149243e-06)),(to_sfixed_a(0.00023881267406977713)),(to_sfixed_a(-0.31713780760765076)),(to_sfixed_a(0.003603752702474594)),(to_sfixed_a(-4.5565284381154925e-06)),(to_sfixed_a(0.006871339865028858)),(to_sfixed_a(0.008869366720318794)),(to_sfixed_a(0.0009232587763108313)),(to_sfixed_a(-0.000239825458265841)),(to_sfixed_a(-0.0001487033296143636)),(to_sfixed_a(-0.006717072334140539)),(to_sfixed_a(1.5853212971705943e-05)),(to_sfixed_a(-0.0006301947869360447)),(to_sfixed_a(-1.3925673556514084e-06)),(to_sfixed_a(0.002416996518149972)),(to_sfixed_a(-5.249139940133318e-05)),(to_sfixed_a(-0.00015416875248774886)),(to_sfixed_a(-1.3195458450354636e-06)),(to_sfixed_a(-8.582612645113841e-05)),(to_sfixed_a(0.0002900508407037705)),(to_sfixed_a(0.0005676456494256854)),(to_sfixed_a(-0.17590078711509705)),(to_sfixed_a(-3.484979970380664e-06)),(to_sfixed_a(-0.2546730637550354)),(to_sfixed_a(-0.16798372566699982)),(to_sfixed_a(-0.00017311220290139318)),(to_sfixed_a(0.0004232183564454317)),(to_sfixed_a(-0.00010017376916948706)),(to_sfixed_a(-0.00024355578352697194)),(to_sfixed_a(0.01559379044920206)),(to_sfixed_a(0.017605235800147057)),(to_sfixed_a(-6.82387180859223e-05)),(to_sfixed_a(0.003282463876530528)),(to_sfixed_a(5.877571675227955e-05)),(to_sfixed_a(-6.298987864283845e-05)),(to_sfixed_a(0.5478111505508423)),(to_sfixed_a(-0.00012361460539977998)),(to_sfixed_a(0.11689326912164688)),(to_sfixed_a(0.00022392078244592994)),(to_sfixed_a(-0.00034247327130287886)),(to_sfixed_a(-0.00023031383170746267)),(to_sfixed_a(-5.157420309842564e-05)),(to_sfixed_a(0.001058653462678194)),(to_sfixed_a(-2.372130984440446e-05)),(to_sfixed_a(-0.00030091116786934435)),(to_sfixed_a(0.3119749128818512)),(to_sfixed_a(0.006617049220949411)),(to_sfixed_a(-0.0002440180687699467)),(to_sfixed_a(0.00011596815602388233)),(to_sfixed_a(0.00012968055671080947)),(to_sfixed_a(0.00011379749048501253)),(to_sfixed_a(-0.00015701926895417273)),(to_sfixed_a(0.004231369588524103)),(to_sfixed_a(0.2594880759716034)),(to_sfixed_a(0.00015664890815969557)),(to_sfixed_a(-1.3219003449194133e-05)),(to_sfixed_a(0.2572920322418213)),(to_sfixed_a(0.28569644689559937)),(to_sfixed_a(4.779314622282982e-05)),(to_sfixed_a(0.00010025327355833724)),(to_sfixed_a(0.2592928111553192)),(to_sfixed_a(-3.0607152439188212e-06)),(to_sfixed_a(-0.000197019093320705)),(to_sfixed_a(0.00019864441128447652)),(to_sfixed_a(-0.000762835203204304)),(to_sfixed_a(-0.0006112921400927007)),(to_sfixed_a(0.00034672010224312544)),(to_sfixed_a(-0.0002522706345189363)),(to_sfixed_a(4.953682218911126e-05)),(to_sfixed_a(0.009052827022969723)),(to_sfixed_a(7.339379953918979e-05)),(to_sfixed_a(-0.0001365701900795102)),(to_sfixed_a(-0.20078130066394806)),(to_sfixed_a(3.0127339414320886e-06)),(to_sfixed_a(-2.3949891328811646e-05)),(to_sfixed_a(-0.06561176478862762)),(to_sfixed_a(0.00024329370353370905)),(to_sfixed_a(0.0032298362348228693)),(to_sfixed_a(0.00010816967551363632)),(to_sfixed_a(0.00015420389536302537)),(to_sfixed_a(-0.00010616821236908436)),(to_sfixed_a(0.0001135470301960595)),(to_sfixed_a(-0.269980251789093)),(to_sfixed_a(0.0021571435499936342)),(to_sfixed_a(0.0029593599028885365)),(to_sfixed_a(0.001384455244988203)),(to_sfixed_a(0.00031778885750100017)),(to_sfixed_a(0.30915799736976624)),(to_sfixed_a(6.959169695619494e-05)),(to_sfixed_a(2.3093427444109693e-05)),(to_sfixed_a(-0.3987101912498474)),(to_sfixed_a(0.03363632410764694)),(to_sfixed_a(-0.4538896679878235)),(to_sfixed_a(0.00017303091590292752)),(to_sfixed_a(0.5113407373428345)),(to_sfixed_a(-0.16830839216709137)),(to_sfixed_a(0.00065259711118415)),(to_sfixed_a(0.0006582866190001369)),(to_sfixed_a(-0.16767802834510803)),(to_sfixed_a(0.25882747769355774)),(to_sfixed_a(0.2776103615760803)),(to_sfixed_a(0.01044770423322916)),(to_sfixed_a(-1.1611507943598554e-05)),(to_sfixed_a(7.173239282565191e-05)),(to_sfixed_a(2.414140908513218e-06)),(to_sfixed_a(0.00025044300127774477)),(to_sfixed_a(0.005486876238137484)),(to_sfixed_a(0.0022648731246590614)),(to_sfixed_a(-0.0008259511087089777)),(to_sfixed_a(-0.36706140637397766)),(to_sfixed_a(-0.2265695482492447)),(to_sfixed_a(-0.00032258438295684755)),(to_sfixed_a(0.0024159238673746586)),(to_sfixed_a(-0.00825316458940506)),(to_sfixed_a(-0.0001580290263518691)),(to_sfixed_a(0.4182174503803253)),(to_sfixed_a(-0.00014836073387414217)),(to_sfixed_a(0.0005000420496799052)),(to_sfixed_a(-0.004328325390815735)),(to_sfixed_a(0.00015595820150338113)),(to_sfixed_a(0.00026074331253767014)),(to_sfixed_a(4.457951945369132e-05)),(to_sfixed_a(0.00014120635751169175)),(to_sfixed_a(0.00011591881047934294)),(to_sfixed_a(-7.040670607239008e-05)),(to_sfixed_a(0.003030665684491396)),(to_sfixed_a(-0.0074334172531962395)),(to_sfixed_a(-0.009776435792446136)),(to_sfixed_a(0.00027496233815327287)),(to_sfixed_a(0.0013733492232859135)),(to_sfixed_a(-0.26348572969436646)),(to_sfixed_a(0.00016657206288073212)),(to_sfixed_a(1.9395964045543224e-05)),(to_sfixed_a(2.0334340661065653e-05)),(to_sfixed_a(0.0003753296041395515)),(to_sfixed_a(6.429539644159377e-05)),(to_sfixed_a(0.020014174282550812)),(to_sfixed_a(0.2685616910457611)),(to_sfixed_a(0.009645230136811733)),(to_sfixed_a(-0.00026287988293915987)),(to_sfixed_a(-6.462173769250512e-05)),(to_sfixed_a(-0.00011988387268502265)),(to_sfixed_a(0.0001374979328829795)),(to_sfixed_a(-0.00015048476052470505)),(to_sfixed_a(-0.0006566968513652682)),(to_sfixed_a(0.00018044994794763625)),(to_sfixed_a(-9.843497537076473e-07)),(to_sfixed_a(0.00030355394119396806)),(to_sfixed_a(0.019215965643525124)),(to_sfixed_a(0.0006653736345469952)),(to_sfixed_a(0.028814589604735374)),(to_sfixed_a(0.00020461430540308356)),(to_sfixed_a(-0.00014690024545416236)),(to_sfixed_a(0.00013342767488211393)),(to_sfixed_a(-0.00047851906856521964)),(to_sfixed_a(0.00387888727709651)),(to_sfixed_a(-0.0032267607748508453)),(to_sfixed_a(6.294594641076401e-05)),(to_sfixed_a(6.948793452465907e-05)),(to_sfixed_a(1.5716224879724905e-05)),(to_sfixed_a(-0.19938619434833527)),(to_sfixed_a(-0.00022243634157348424)),(to_sfixed_a(-0.16857454180717468)),(to_sfixed_a(-2.8989079510211013e-05)),(to_sfixed_a(0.013782058842480183)),(to_sfixed_a(0.0004471816646400839)),(to_sfixed_a(0.1550057828426361)),(to_sfixed_a(0.07168850302696228)),(to_sfixed_a(6.650754949077964e-05)),(to_sfixed_a(-0.0029204359743744135)),(to_sfixed_a(0.0008595630642957985)),(to_sfixed_a(7.908592669991776e-05)),(to_sfixed_a(-0.11268499493598938)),(to_sfixed_a(7.006918895058334e-05)),(to_sfixed_a(-0.00020580073760356754)),(to_sfixed_a(0.00457785977050662)),(to_sfixed_a(-0.01884685643017292)),(to_sfixed_a(0.00010410866525489837)),(to_sfixed_a(-0.00014567113248631358)),(to_sfixed_a(0.3496951460838318)),(to_sfixed_a(-0.00013018798199482262)),(to_sfixed_a(0.0018516955897212029)),(to_sfixed_a(0.00015196064487099648)),(to_sfixed_a(0.0009906822815537453)),(to_sfixed_a(-0.00013655671500600874)),(to_sfixed_a(-0.14150460064411163)),(to_sfixed_a(0.00018689384160097688)),(to_sfixed_a(-4.126655403524637e-05)),(to_sfixed_a(4.797893780050799e-07)),(to_sfixed_a(0.007790348492562771)),(to_sfixed_a(0.025907769799232483)),(to_sfixed_a(-0.0002459873503539711)),(to_sfixed_a(-6.0386497352737933e-05)),(to_sfixed_a(4.7223555156961083e-05)),(to_sfixed_a(0.0002934869844466448)),(to_sfixed_a(0.0009069882798939943)),(to_sfixed_a(0.003329609986394644)),(to_sfixed_a(0.00029078105580992997)),(to_sfixed_a(0.028383009135723114)),(to_sfixed_a(0.5674475431442261)),(to_sfixed_a(-0.00018527224892750382)),(to_sfixed_a(2.4991799364215694e-05)),(to_sfixed_a(0.00015194391016848385)),(to_sfixed_a(-0.00028115889290347695)),(to_sfixed_a(-0.0002039668324869126)),(to_sfixed_a(-0.00017717821174301207)),(to_sfixed_a(-0.002527522621676326)),(to_sfixed_a(-0.41565245389938354)),(to_sfixed_a(-0.00011064660066040233)),(to_sfixed_a(-0.006349131930619478)),(to_sfixed_a(0.001064665149897337)),(to_sfixed_a(0.037439774721860886)),(to_sfixed_a(0.006299599073827267)),(to_sfixed_a(0.00011634860857157037)),(to_sfixed_a(0.25817039608955383)),(to_sfixed_a(-0.019908377900719643)),(to_sfixed_a(0.0008213610271923244)),(to_sfixed_a(2.932742063421756e-05)),(to_sfixed_a(-0.18363840878009796)),(to_sfixed_a(0.00106462009716779)),(to_sfixed_a(-0.18240049481391907)));

    constant weight_n2_22 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.20101702213287354)),(to_sfixed_a(0.0028365019243210554)),(to_sfixed_a(0.0008861490641720593)),(to_sfixed_a(-0.00011838739737868309)),(to_sfixed_a(-0.015426571480929852)),(to_sfixed_a(0.00029789539985358715)),(to_sfixed_a(0.014730244874954224)),(to_sfixed_a(-9.916498675011098e-05)),(to_sfixed_a(0.00015132190310396254)),(to_sfixed_a(0.00023753309505991638)),(to_sfixed_a(-0.00021047690825071186)),(to_sfixed_a(0.002758123679086566)),(to_sfixed_a(-0.28638097643852234)),(to_sfixed_a(0.0030494669917970896)),(to_sfixed_a(6.6075284848921e-05)),(to_sfixed_a(5.603647150564939e-05)),(to_sfixed_a(0.00041885103564709425)),(to_sfixed_a(8.150329813361168e-05)),(to_sfixed_a(0.04406441003084183)),(to_sfixed_a(0.060529205948114395)),(to_sfixed_a(1.736480407998897e-05)),(to_sfixed_a(-0.00017453738837502897)),(to_sfixed_a(0.19872280955314636)),(to_sfixed_a(0.3818485736846924)),(to_sfixed_a(0.2365771383047104)),(to_sfixed_a(0.0006404604064300656)),(to_sfixed_a(0.00030528282513841987)),(to_sfixed_a(3.458379796938971e-05)),(to_sfixed_a(0.0176687128841877)),(to_sfixed_a(-0.00022774614626541734)),(to_sfixed_a(0.33550864458084106)),(to_sfixed_a(-6.926980131538585e-05)),(to_sfixed_a(0.0025395164266228676)),(to_sfixed_a(1.8857659597415477e-05)),(to_sfixed_a(-0.00023894431069493294)),(to_sfixed_a(-6.003612361382693e-05)),(to_sfixed_a(-0.010037037543952465)),(to_sfixed_a(0.0011735165026038885)),(to_sfixed_a(0.013258754275739193)),(to_sfixed_a(-1.1765609087888151e-05)),(to_sfixed_a(0.004604286514222622)),(to_sfixed_a(0.0020633952226489782)),(to_sfixed_a(-0.00010161783575313166)),(to_sfixed_a(2.1283183741616085e-05)),(to_sfixed_a(0.006470490712672472)),(to_sfixed_a(0.02129466086626053)),(to_sfixed_a(0.2858729362487793)),(to_sfixed_a(0.01911098323762417)),(to_sfixed_a(-0.00018274963076692075)),(to_sfixed_a(0.0075303358025848866)),(to_sfixed_a(0.26829665899276733)),(to_sfixed_a(0.0009315633215010166)),(to_sfixed_a(-2.487487654434517e-05)),(to_sfixed_a(-0.0016554539324715734)),(to_sfixed_a(0.000467355246655643)),(to_sfixed_a(0.009974136017262936)),(to_sfixed_a(-7.189391180872917e-05)),(to_sfixed_a(0.013402671553194523)),(to_sfixed_a(-0.00014692239346913993)),(to_sfixed_a(-0.0004240071284584701)),(to_sfixed_a(0.006774956826120615)),(to_sfixed_a(0.0063052186742424965)),(to_sfixed_a(0.0001726738119032234)),(to_sfixed_a(0.008410248905420303)),(to_sfixed_a(-0.00010747602209448814)),(to_sfixed_a(0.012434788048267365)),(to_sfixed_a(-2.514842344680801e-05)),(to_sfixed_a(-0.0035163445863872766)),(to_sfixed_a(0.01235042605549097)),(to_sfixed_a(-0.0001683357113506645)),(to_sfixed_a(-0.016967330127954483)),(to_sfixed_a(0.438973993062973)),(to_sfixed_a(-0.18237069249153137)),(to_sfixed_a(-0.00012105161295039579)),(to_sfixed_a(-6.447511987062171e-05)),(to_sfixed_a(2.3007518393569626e-05)),(to_sfixed_a(0.015867307782173157)),(to_sfixed_a(0.007368152029812336)),(to_sfixed_a(-1.0631629265844822e-06)),(to_sfixed_a(0.000541534973308444)),(to_sfixed_a(0.006339037325233221)),(to_sfixed_a(-6.591177952941507e-05)),(to_sfixed_a(0.5918905735015869)),(to_sfixed_a(-0.009252545423805714)),(to_sfixed_a(-0.00013080872304271907)),(to_sfixed_a(0.0038541126996278763)),(to_sfixed_a(0.21167871356010437)),(to_sfixed_a(-0.0032638104166835546)),(to_sfixed_a(0.00025132769951596856)),(to_sfixed_a(-0.0004114631738048047)),(to_sfixed_a(0.01666264794766903)),(to_sfixed_a(7.115262269508094e-05)),(to_sfixed_a(0.013130486942827702)),(to_sfixed_a(0.00027740123914554715)),(to_sfixed_a(0.002184527926146984)),(to_sfixed_a(0.00015369727043434978)),(to_sfixed_a(1.4326375094242394e-05)),(to_sfixed_a(1.6781013982836157e-06)),(to_sfixed_a(0.0001483093510614708)),(to_sfixed_a(3.0243099899962544e-05)),(to_sfixed_a(0.0007118675857782364)),(to_sfixed_a(0.0018647026736289263)),(to_sfixed_a(-0.0002044309367192909)),(to_sfixed_a(0.004520357120782137)),(to_sfixed_a(-0.4380595088005066)),(to_sfixed_a(0.0005164170288480818)),(to_sfixed_a(5.0074304454028606e-05)),(to_sfixed_a(8.719562902115285e-05)),(to_sfixed_a(0.00015505192277487367)),(to_sfixed_a(0.19411920011043549)),(to_sfixed_a(0.0031711384654045105)),(to_sfixed_a(6.4380161347799e-05)),(to_sfixed_a(0.7686141729354858)),(to_sfixed_a(-2.9085465939715505e-05)),(to_sfixed_a(3.253668546676636e-05)),(to_sfixed_a(-0.18787071108818054)),(to_sfixed_a(-0.00011374394671292976)),(to_sfixed_a(0.006421164143830538)),(to_sfixed_a(-0.00022263819118961692)),(to_sfixed_a(0.13971446454524994)),(to_sfixed_a(-3.825976455118507e-05)),(to_sfixed_a(0.00018176813318859786)),(to_sfixed_a(0.009801249951124191)),(to_sfixed_a(-6.916309212101623e-05)),(to_sfixed_a(-1.0753252354334109e-05)),(to_sfixed_a(0.0011506122536957264)),(to_sfixed_a(-0.19612500071525574)),(to_sfixed_a(-0.00021890476637054235)),(to_sfixed_a(0.0002309172268724069)),(to_sfixed_a(-6.858802225906402e-05)),(to_sfixed_a(0.0002467409649398178)),(to_sfixed_a(6.207900878507644e-05)),(to_sfixed_a(0.000331818126142025)),(to_sfixed_a(0.0015105248894542456)),(to_sfixed_a(-5.816691555082798e-07)),(to_sfixed_a(-2.423875776003115e-05)),(to_sfixed_a(0.0240124873816967)),(to_sfixed_a(0.41245853900909424)),(to_sfixed_a(-0.0002359952195547521)),(to_sfixed_a(0.00019691379566211253)),(to_sfixed_a(0.0012395854573696852)),(to_sfixed_a(-2.5045295842573978e-05)),(to_sfixed_a(0.00013509842392522842)),(to_sfixed_a(-2.6782427084981464e-05)),(to_sfixed_a(9.118888556258753e-05)),(to_sfixed_a(0.004690897651016712)),(to_sfixed_a(0.0032038779463618994)),(to_sfixed_a(-0.0001005858212010935)),(to_sfixed_a(-0.00016895594308152795)),(to_sfixed_a(0.010052036494016647)),(to_sfixed_a(-0.00011842083767987788)),(to_sfixed_a(0.00010490859858691692)),(to_sfixed_a(0.0007870416739024222)),(to_sfixed_a(-0.00012924624024890363)),(to_sfixed_a(0.00023873356985859573)),(to_sfixed_a(0.0010297626722604036)),(to_sfixed_a(-9.111817053053528e-05)),(to_sfixed_a(0.0017993387300521135)),(to_sfixed_a(-0.0004704854218289256)),(to_sfixed_a(-1.618974783923477e-05)),(to_sfixed_a(-0.0001693356316536665)),(to_sfixed_a(2.9444065148709342e-05)),(to_sfixed_a(0.1245415061712265)),(to_sfixed_a(-0.00292026624083519)),(to_sfixed_a(0.004282280802726746)),(to_sfixed_a(0.0005943329306319356)),(to_sfixed_a(-8.781391807133332e-05)),(to_sfixed_a(0.3631129562854767)),(to_sfixed_a(0.00016840566240716726)),(to_sfixed_a(0.00012858858099207282)),(to_sfixed_a(0.03586508333683014)),(to_sfixed_a(0.005485622677952051)),(to_sfixed_a(-0.00039270147681236267)),(to_sfixed_a(7.124762487364933e-05)),(to_sfixed_a(0.014572517946362495)),(to_sfixed_a(2.744546509347856e-05)),(to_sfixed_a(0.3369388282299042)),(to_sfixed_a(3.47936074831523e-05)),(to_sfixed_a(0.002863714238628745)),(to_sfixed_a(0.1651366651058197)),(to_sfixed_a(0.0010409718379378319)),(to_sfixed_a(0.18524503707885742)),(to_sfixed_a(-2.0000923541374505e-05)),(to_sfixed_a(-3.0246737878769636e-06)),(to_sfixed_a(0.0002782806695904583)),(to_sfixed_a(0.0006231174920685589)),(to_sfixed_a(-0.49024346470832825)),(to_sfixed_a(0.0020836666226387024)),(to_sfixed_a(0.002960714977234602)),(to_sfixed_a(9.249174763681367e-05)),(to_sfixed_a(-0.019071249291300774)),(to_sfixed_a(0.00011944174184463918)),(to_sfixed_a(0.012580635026097298)),(to_sfixed_a(0.24623972177505493)),(to_sfixed_a(-6.792344356654212e-05)),(to_sfixed_a(0.0003396657120902091)),(to_sfixed_a(-0.00025202930555678904)),(to_sfixed_a(-0.0005119203706271946)),(to_sfixed_a(-0.23409192264080048)),(to_sfixed_a(0.0002377677010372281)),(to_sfixed_a(-0.00020889134611934423)),(to_sfixed_a(0.0002054994838545099)),(to_sfixed_a(9.451039659325033e-05)),(to_sfixed_a(-3.2435877074021846e-05)),(to_sfixed_a(-9.038299322128296e-05)),(to_sfixed_a(0.0009107080986723304)),(to_sfixed_a(0.0008312214631587267)),(to_sfixed_a(-0.3257569372653961)),(to_sfixed_a(0.004527722951024771)),(to_sfixed_a(0.008528308011591434)),(to_sfixed_a(0.00695052882656455)),(to_sfixed_a(-0.00019557597988750786)),(to_sfixed_a(0.00025650381576269865)),(to_sfixed_a(-5.275898729451001e-06)),(to_sfixed_a(0.0002990041975863278)),(to_sfixed_a(-0.00041815382428467274)),(to_sfixed_a(0.001335430657491088)),(to_sfixed_a(-9.264916297979653e-05)),(to_sfixed_a(0.24066758155822754)),(to_sfixed_a(-1.925208925968036e-05)),(to_sfixed_a(-6.325013237074018e-05)),(to_sfixed_a(0.00011375168833183125)),(to_sfixed_a(-7.233706128317863e-05)),(to_sfixed_a(-8.379949576919898e-05)),(to_sfixed_a(0.011514756828546524)),(to_sfixed_a(-0.00010848901001736522)),(to_sfixed_a(3.230729271308519e-05)),(to_sfixed_a(-7.436989835696295e-05)),(to_sfixed_a(-0.010251108556985855)),(to_sfixed_a(0.04229378700256348)),(to_sfixed_a(0.004795231390744448)),(to_sfixed_a(-0.0002985927276313305)),(to_sfixed_a(-0.00042350913281552494)),(to_sfixed_a(-0.00020583963487297297)),(to_sfixed_a(0.0033558134455233812)),(to_sfixed_a(0.0016990762669593096)),(to_sfixed_a(-0.0004053401935379952)),(to_sfixed_a(8.46067487145774e-05)),(to_sfixed_a(0.000809891615062952)),(to_sfixed_a(0.00020968701574020088)),(to_sfixed_a(-0.00029070256277918816)),(to_sfixed_a(-4.385699867270887e-06)),(to_sfixed_a(0.24171662330627441)),(to_sfixed_a(0.0001660720445215702)),(to_sfixed_a(-0.25494384765625)),(to_sfixed_a(0.00462593138217926)),(to_sfixed_a(0.18951807916164398)),(to_sfixed_a(0.012312016449868679)),(to_sfixed_a(-0.00015588408859912306)),(to_sfixed_a(0.01181337982416153)),(to_sfixed_a(0.003686053678393364)),(to_sfixed_a(-1.8930686564999633e-05)),(to_sfixed_a(0.007550792768597603)),(to_sfixed_a(7.07143044564873e-05)),(to_sfixed_a(-0.00022506546520162374)),(to_sfixed_a(0.023600473999977112)),(to_sfixed_a(0.02282271906733513)),(to_sfixed_a(5.880822573089972e-05)),(to_sfixed_a(1.406863157171756e-05)),(to_sfixed_a(0.006809015292674303)),(to_sfixed_a(-7.333621033467352e-05)),(to_sfixed_a(-0.03652460128068924)),(to_sfixed_a(-0.00015336857177317142)),(to_sfixed_a(0.0010592928156256676)),(to_sfixed_a(-3.953051054850221e-05)),(to_sfixed_a(-0.4075872004032135)),(to_sfixed_a(0.00015646254178136587)),(to_sfixed_a(-0.00018851208733394742)),(to_sfixed_a(-8.508354221703485e-05)),(to_sfixed_a(0.0033640973269939423)),(to_sfixed_a(-0.005744559690356255)),(to_sfixed_a(0.000224695832002908)),(to_sfixed_a(-2.4408931494690478e-05)),(to_sfixed_a(0.00010245812882203609)),(to_sfixed_a(1.3357501302380115e-05)),(to_sfixed_a(-0.004828369710594416)),(to_sfixed_a(0.01674274541437626)),(to_sfixed_a(0.20559754967689514)),(to_sfixed_a(0.009556571952998638)),(to_sfixed_a(-0.0004200286930426955)),(to_sfixed_a(-5.217334546614438e-06)),(to_sfixed_a(0.00023990521731320769)),(to_sfixed_a(0.00016861526819411665)),(to_sfixed_a(0.16688449680805206)),(to_sfixed_a(-0.00018277518393006176)),(to_sfixed_a(0.00011662359611364082)),(to_sfixed_a(0.17239730060100555)),(to_sfixed_a(0.00038205718738026917)),(to_sfixed_a(6.227575067896396e-05)),(to_sfixed_a(-0.20823752880096436)),(to_sfixed_a(-0.000748691032640636)),(to_sfixed_a(-0.3279157280921936)),(to_sfixed_a(0.006449245847761631)),(to_sfixed_a(-9.282326573156752e-06)),(to_sfixed_a(0.0044906605035066605)),(to_sfixed_a(0.004440579097718)),(to_sfixed_a(0.007946956902742386)),(to_sfixed_a(-0.0001484660169808194)),(to_sfixed_a(0.253019779920578)),(to_sfixed_a(-0.004704222548753023)),(to_sfixed_a(0.013370883651077747)));

    constant weight_n2_23 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.027909686788916588)),(to_sfixed_a(0.00015137612354010344)),(to_sfixed_a(2.497301102266647e-05)),(to_sfixed_a(-7.330744119826704e-05)),(to_sfixed_a(3.2736930734245107e-05)),(to_sfixed_a(0.00012600906484294683)),(to_sfixed_a(0.00013543502427637577)),(to_sfixed_a(-0.0001270062493858859)),(to_sfixed_a(-2.0753679564222693e-05)),(to_sfixed_a(6.711750756949186e-05)),(to_sfixed_a(2.88514893327374e-05)),(to_sfixed_a(0.0004236869572196156)),(to_sfixed_a(-7.083135278662667e-05)),(to_sfixed_a(9.829147165874019e-05)),(to_sfixed_a(-0.00017230582307092845)),(to_sfixed_a(0.00010905280942097306)),(to_sfixed_a(-0.00011834659380838275)),(to_sfixed_a(-0.00018401682609692216)),(to_sfixed_a(-0.00029995146906003356)),(to_sfixed_a(0.00017847266281023622)),(to_sfixed_a(-6.190673593664542e-05)),(to_sfixed_a(-1.70085986610502e-05)),(to_sfixed_a(-9.489068906987086e-05)),(to_sfixed_a(2.0052530089742504e-05)),(to_sfixed_a(-8.968886686488986e-05)),(to_sfixed_a(-4.445901868166402e-05)),(to_sfixed_a(0.00010878073226194829)),(to_sfixed_a(0.00011017722135875374)),(to_sfixed_a(-7.073321467032656e-05)),(to_sfixed_a(4.432069545146078e-05)),(to_sfixed_a(1.038682967191562e-05)),(to_sfixed_a(-9.170662087853998e-05)),(to_sfixed_a(-0.00018004314915742725)),(to_sfixed_a(-1.1845197150250897e-05)),(to_sfixed_a(-0.0004137326031923294)),(to_sfixed_a(-0.00015643975348211825)),(to_sfixed_a(-0.00020400798530317843)),(to_sfixed_a(-3.680132431327365e-05)),(to_sfixed_a(-1.833326678024605e-06)),(to_sfixed_a(-0.00022936987807042897)),(to_sfixed_a(2.4797900550765917e-05)),(to_sfixed_a(1.2123186024837196e-05)),(to_sfixed_a(-2.0925825083395466e-05)),(to_sfixed_a(1.8883538359659724e-05)),(to_sfixed_a(2.0790030248463154e-06)),(to_sfixed_a(-7.123398245312274e-05)),(to_sfixed_a(-0.00029545952565968037)),(to_sfixed_a(-2.376825432293117e-05)),(to_sfixed_a(5.8258625358575955e-05)),(to_sfixed_a(-6.03889930061996e-07)),(to_sfixed_a(2.9359729524003342e-05)),(to_sfixed_a(8.93384130904451e-05)),(to_sfixed_a(7.083882519509643e-05)),(to_sfixed_a(-7.84762087278068e-05)),(to_sfixed_a(1.1760661436710507e-05)),(to_sfixed_a(-1.2448035704437643e-06)),(to_sfixed_a(-2.571981167420745e-05)),(to_sfixed_a(-2.353965101065114e-05)),(to_sfixed_a(2.0926090655848384e-06)),(to_sfixed_a(-0.00011226551578147337)),(to_sfixed_a(0.00011586353502934799)),(to_sfixed_a(-0.00010045826638815925)),(to_sfixed_a(-5.457790393847972e-06)),(to_sfixed_a(-0.00011211063247174025)),(to_sfixed_a(2.7036163373850286e-05)),(to_sfixed_a(-6.949628004804254e-05)),(to_sfixed_a(-0.00045211860560812056)),(to_sfixed_a(0.0001041116047417745)),(to_sfixed_a(5.859904922544956e-05)),(to_sfixed_a(1.577362127136439e-06)),(to_sfixed_a(-0.00015116319991648197)),(to_sfixed_a(0.00044928808347322047)),(to_sfixed_a(0.00011397586786188185)),(to_sfixed_a(0.0002381765516474843)),(to_sfixed_a(-5.108865298097953e-05)),(to_sfixed_a(-7.264017767738551e-05)),(to_sfixed_a(-3.886858394253068e-05)),(to_sfixed_a(-0.0001827071828301996)),(to_sfixed_a(3.7874982808716595e-05)),(to_sfixed_a(0.00041176044032908976)),(to_sfixed_a(-0.0001667326141614467)),(to_sfixed_a(5.405292904470116e-05)),(to_sfixed_a(-1.5681136574130505e-05)),(to_sfixed_a(-0.00011394407920306548)),(to_sfixed_a(0.00011617610289249569)),(to_sfixed_a(0.00011641768651315942)),(to_sfixed_a(3.52314964402467e-06)),(to_sfixed_a(-0.00011254155833739787)),(to_sfixed_a(1.3215452781878412e-05)),(to_sfixed_a(-0.0001300904550589621)),(to_sfixed_a(-7.177088264143094e-05)),(to_sfixed_a(0.0002628086367622018)),(to_sfixed_a(3.179382474627346e-06)),(to_sfixed_a(-0.00010228062456008047)),(to_sfixed_a(7.315463153645396e-05)),(to_sfixed_a(6.37606717646122e-05)),(to_sfixed_a(2.6646150217857212e-05)),(to_sfixed_a(0.0002473464410286397)),(to_sfixed_a(4.769096267409623e-05)),(to_sfixed_a(-0.0002369297726545483)),(to_sfixed_a(-5.719110049540177e-06)),(to_sfixed_a(0.00025097219622693956)),(to_sfixed_a(-7.18350347597152e-05)),(to_sfixed_a(-0.0001638189860386774)),(to_sfixed_a(-6.851699436083436e-05)),(to_sfixed_a(-0.0001525694679003209)),(to_sfixed_a(0.00011390555300749838)),(to_sfixed_a(4.7976984205888584e-05)),(to_sfixed_a(6.020273576723412e-05)),(to_sfixed_a(-3.0120336305117235e-05)),(to_sfixed_a(-9.691204468254e-05)),(to_sfixed_a(-4.64574623038061e-06)),(to_sfixed_a(6.56614065519534e-05)),(to_sfixed_a(-0.00015715076006017625)),(to_sfixed_a(-0.00013801106251776218)),(to_sfixed_a(-9.184443115373142e-06)),(to_sfixed_a(0.00010494436719454825)),(to_sfixed_a(5.344993405742571e-05)),(to_sfixed_a(4.6718378143850714e-05)),(to_sfixed_a(-8.554405940230936e-05)),(to_sfixed_a(-7.050145359244198e-05)),(to_sfixed_a(-0.0001139590167440474)),(to_sfixed_a(-6.65212282910943e-05)),(to_sfixed_a(-0.00010515988833503798)),(to_sfixed_a(0.0002878757659345865)),(to_sfixed_a(1.4864010154269636e-05)),(to_sfixed_a(0.00011734232248272747)),(to_sfixed_a(0.0001838989119278267)),(to_sfixed_a(-6.504688644781709e-05)),(to_sfixed_a(-0.00013619184028357267)),(to_sfixed_a(2.3356300516752526e-05)),(to_sfixed_a(-0.00021219084737822413)),(to_sfixed_a(-6.938666047062725e-05)),(to_sfixed_a(-0.00014673522673547268)),(to_sfixed_a(-0.00013515836326405406)),(to_sfixed_a(-1.66265235748142e-05)),(to_sfixed_a(0.0004150182649027556)),(to_sfixed_a(0.00029593458748422563)),(to_sfixed_a(7.23088305676356e-07)),(to_sfixed_a(-2.855540515156463e-06)),(to_sfixed_a(0.00015161755436565727)),(to_sfixed_a(0.0001165315552498214)),(to_sfixed_a(4.931673174723983e-06)),(to_sfixed_a(7.153697515605018e-05)),(to_sfixed_a(1.9720398995559663e-05)),(to_sfixed_a(-1.1235770216444507e-05)),(to_sfixed_a(0.0003023374592885375)),(to_sfixed_a(7.129392179194838e-05)),(to_sfixed_a(-0.0001359357702312991)),(to_sfixed_a(9.066719212569296e-05)),(to_sfixed_a(0.00012838827387895435)),(to_sfixed_a(0.00014941570407245308)),(to_sfixed_a(5.917670932831243e-05)),(to_sfixed_a(-1.913493179017678e-05)),(to_sfixed_a(-6.727204890921712e-05)),(to_sfixed_a(-0.00015639342018403113)),(to_sfixed_a(-2.2284970327746123e-05)),(to_sfixed_a(4.039502528030425e-05)),(to_sfixed_a(-4.35273141192738e-05)),(to_sfixed_a(0.00010922525689238682)),(to_sfixed_a(-0.00014453806215897202)),(to_sfixed_a(0.00019535867613740265)),(to_sfixed_a(0.000300844490993768)),(to_sfixed_a(-2.4797525838948786e-05)),(to_sfixed_a(-0.00015300976519938558)),(to_sfixed_a(4.86716307932511e-05)),(to_sfixed_a(-2.3348809918388724e-05)),(to_sfixed_a(-0.0001130825185100548)),(to_sfixed_a(0.00015965619240887463)),(to_sfixed_a(3.951245889766142e-05)),(to_sfixed_a(8.617120329290628e-06)),(to_sfixed_a(-0.00011621628073044121)),(to_sfixed_a(-6.38464480289258e-05)),(to_sfixed_a(-7.943141099531204e-05)),(to_sfixed_a(5.6707271141931415e-05)),(to_sfixed_a(-0.0001203979627462104)),(to_sfixed_a(-7.234801887534559e-05)),(to_sfixed_a(-5.944350778008811e-05)),(to_sfixed_a(6.116828444646671e-05)),(to_sfixed_a(0.00023567810421809554)),(to_sfixed_a(-3.559862307156436e-06)),(to_sfixed_a(-4.009265103377402e-05)),(to_sfixed_a(8.400975639233366e-05)),(to_sfixed_a(-0.00010141155507881194)),(to_sfixed_a(6.043834946467541e-05)),(to_sfixed_a(-0.000446068326709792)),(to_sfixed_a(-0.00010408920934423804)),(to_sfixed_a(0.00016153970500454307)),(to_sfixed_a(-0.000291670294245705)),(to_sfixed_a(0.00018817429372575134)),(to_sfixed_a(-7.135189662221819e-05)),(to_sfixed_a(0.00010088293493026868)),(to_sfixed_a(4.125807390664704e-05)),(to_sfixed_a(-0.00019858003361150622)),(to_sfixed_a(-0.00018828583415597677)),(to_sfixed_a(-2.2136810002848506e-06)),(to_sfixed_a(0.000173383901710622)),(to_sfixed_a(-2.5649627787061036e-05)),(to_sfixed_a(4.8768877604743466e-05)),(to_sfixed_a(1.788920781109482e-05)),(to_sfixed_a(-0.00024227604444604367)),(to_sfixed_a(9.586803935235366e-05)),(to_sfixed_a(-1.0291179933119565e-05)),(to_sfixed_a(0.00014857797941658646)),(to_sfixed_a(0.00029231823282316327)),(to_sfixed_a(6.706315616611391e-06)),(to_sfixed_a(0.00010516286420170218)),(to_sfixed_a(9.720341040519997e-05)),(to_sfixed_a(0.00010098623897647485)),(to_sfixed_a(-6.0549999034265056e-05)),(to_sfixed_a(-1.911350409500301e-06)),(to_sfixed_a(2.0433835743460804e-05)),(to_sfixed_a(-9.606989624444395e-05)),(to_sfixed_a(-7.105409167706966e-05)),(to_sfixed_a(-1.2079217412974685e-06)),(to_sfixed_a(-4.411070767673664e-05)),(to_sfixed_a(6.529044185299426e-05)),(to_sfixed_a(-6.626917456742376e-05)),(to_sfixed_a(4.5698179746977985e-06)),(to_sfixed_a(-0.00016600702656432986)),(to_sfixed_a(2.9551236366387457e-05)),(to_sfixed_a(6.963835039641708e-05)),(to_sfixed_a(-0.00011688281665556133)),(to_sfixed_a(-6.944406050024554e-05)),(to_sfixed_a(-0.00011277305020485073)),(to_sfixed_a(-6.265832053031772e-05)),(to_sfixed_a(-0.00012821656127925962)),(to_sfixed_a(3.182256477884948e-05)),(to_sfixed_a(0.00016645762661937624)),(to_sfixed_a(-6.276328349485993e-06)),(to_sfixed_a(-8.902260742615908e-05)),(to_sfixed_a(-0.00015399375115521252)),(to_sfixed_a(-8.283014904009178e-05)),(to_sfixed_a(0.00019059467012993991)),(to_sfixed_a(0.00015310199523810297)),(to_sfixed_a(0.00020403569214977324)),(to_sfixed_a(6.233529711607844e-05)),(to_sfixed_a(-0.00012903951574116945)),(to_sfixed_a(-0.00017433791072107852)),(to_sfixed_a(5.8274876209907234e-05)),(to_sfixed_a(-5.3907278925180435e-06)),(to_sfixed_a(0.00010866535740206018)),(to_sfixed_a(-0.00023217870329972357)),(to_sfixed_a(-0.00010628635936882347)),(to_sfixed_a(-3.0049621273064986e-05)),(to_sfixed_a(0.00012804620200768113)),(to_sfixed_a(4.73861291538924e-06)),(to_sfixed_a(-0.00010085532267112285)),(to_sfixed_a(1.2484924809541553e-06)),(to_sfixed_a(0.00016645049618091434)),(to_sfixed_a(3.867522900691256e-05)),(to_sfixed_a(8.61442822497338e-06)),(to_sfixed_a(0.0002102718863170594)),(to_sfixed_a(4.612202610587701e-05)),(to_sfixed_a(-0.0001535981282358989)),(to_sfixed_a(0.00010456895688548684)),(to_sfixed_a(5.547440377995372e-05)),(to_sfixed_a(8.972470823209733e-06)),(to_sfixed_a(7.34684435883537e-05)),(to_sfixed_a(-5.680662434315309e-05)),(to_sfixed_a(0.00017860892694443464)),(to_sfixed_a(-0.00023968018649611622)),(to_sfixed_a(-0.0002884076093323529)),(to_sfixed_a(2.658292942214757e-06)),(to_sfixed_a(4.6073910198174417e-07)),(to_sfixed_a(9.100473835133016e-05)),(to_sfixed_a(6.912702519912273e-05)),(to_sfixed_a(-7.833114068489522e-06)),(to_sfixed_a(-4.05147293349728e-05)),(to_sfixed_a(0.00015499943401664495)),(to_sfixed_a(-0.0001390292018186301)),(to_sfixed_a(0.00021558970911428332)),(to_sfixed_a(-3.7703346606576815e-05)),(to_sfixed_a(7.470000127796084e-05)),(to_sfixed_a(-3.899409784935415e-05)),(to_sfixed_a(-0.00010575648047961295)),(to_sfixed_a(-0.00011564228043425828)),(to_sfixed_a(8.969887130660936e-05)),(to_sfixed_a(-0.0002346701658098027)),(to_sfixed_a(-5.45491639059037e-06)),(to_sfixed_a(-0.00022040403564460576)),(to_sfixed_a(-6.225518154678866e-05)),(to_sfixed_a(-3.360771370353177e-05)),(to_sfixed_a(6.431695510400459e-06)),(to_sfixed_a(-2.2214302589418367e-05)),(to_sfixed_a(-0.00015132765111047775)),(to_sfixed_a(0.00014831224689260125)),(to_sfixed_a(-5.571361543843523e-05)),(to_sfixed_a(0.0004593153716996312)),(to_sfixed_a(0.00015694832836743444)),(to_sfixed_a(6.702209793729708e-05)),(to_sfixed_a(7.666178862564266e-05)),(to_sfixed_a(0.00020440848311409354)),(to_sfixed_a(1.861571945482865e-07)),(to_sfixed_a(2.7233967557549477e-05)),(to_sfixed_a(-0.00018361269030719995)),(to_sfixed_a(0.0001502792874816805)),(to_sfixed_a(-3.622944132075645e-05)),(to_sfixed_a(2.8820533771067858e-05)),(to_sfixed_a(0.00018511794041842222)),(to_sfixed_a(7.44401550036855e-05)));

    constant weight_n2_24 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.0590708926320076)),(to_sfixed_a(-0.007424648385494947)),(to_sfixed_a(-0.00235198182053864)),(to_sfixed_a(6.433880480471998e-05)),(to_sfixed_a(-0.00043634380563162267)),(to_sfixed_a(-6.639446655754e-05)),(to_sfixed_a(-0.0015988253289833665)),(to_sfixed_a(3.5408018447924405e-05)),(to_sfixed_a(-4.824685674975626e-05)),(to_sfixed_a(-0.00038196294917725027)),(to_sfixed_a(-0.00022006324434187263)),(to_sfixed_a(-0.0023993700742721558)),(to_sfixed_a(0.0008346748072654009)),(to_sfixed_a(-0.15597045421600342)),(to_sfixed_a(4.424538929015398e-05)),(to_sfixed_a(6.261540693230927e-05)),(to_sfixed_a(0.41187742352485657)),(to_sfixed_a(-0.00022101525973994285)),(to_sfixed_a(-0.052325233817100525)),(to_sfixed_a(0.004091391805559397)),(to_sfixed_a(2.4278262571897358e-05)),(to_sfixed_a(0.0001528184802737087)),(to_sfixed_a(-4.145708226133138e-05)),(to_sfixed_a(-0.0006547524244524539)),(to_sfixed_a(0.47644439339637756)),(to_sfixed_a(0.40123721957206726)),(to_sfixed_a(5.83188229938969e-05)),(to_sfixed_a(-6.10543429502286e-05)),(to_sfixed_a(-4.9705689889378846e-05)),(to_sfixed_a(0.00010546707198955119)),(to_sfixed_a(-0.002485192148014903)),(to_sfixed_a(-2.918546670116484e-06)),(to_sfixed_a(0.009764987975358963)),(to_sfixed_a(3.3530668588355184e-06)),(to_sfixed_a(-0.00014689433737657964)),(to_sfixed_a(3.721733810380101e-05)),(to_sfixed_a(-0.0054280441254377365)),(to_sfixed_a(0.45581120252609253)),(to_sfixed_a(-0.0029877249617129564)),(to_sfixed_a(5.0229165935888886e-05)),(to_sfixed_a(0.00014944697613827884)),(to_sfixed_a(-0.000951093970797956)),(to_sfixed_a(5.861739919055253e-05)),(to_sfixed_a(5.7111159549094737e-05)),(to_sfixed_a(-0.005522590130567551)),(to_sfixed_a(0.5561497807502747)),(to_sfixed_a(-0.00289949681609869)),(to_sfixed_a(0.01197306253015995)),(to_sfixed_a(-0.0003075014683417976)),(to_sfixed_a(-0.22265079617500305)),(to_sfixed_a(0.16762107610702515)),(to_sfixed_a(0.0007483570370823145)),(to_sfixed_a(3.91344801755622e-05)),(to_sfixed_a(-0.0012054177932441235)),(to_sfixed_a(0.009956935420632362)),(to_sfixed_a(-0.3582395017147064)),(to_sfixed_a(-6.625770765822381e-05)),(to_sfixed_a(-0.008628809824585915)),(to_sfixed_a(4.168396117165685e-06)),(to_sfixed_a(-0.0002987876068800688)),(to_sfixed_a(-0.008672011084854603)),(to_sfixed_a(-0.0020710641983896494)),(to_sfixed_a(5.3828858654014766e-05)),(to_sfixed_a(-0.009891651570796967)),(to_sfixed_a(-0.00018164725042879581)),(to_sfixed_a(-0.0014300545444712043)),(to_sfixed_a(0.00022926002566237003)),(to_sfixed_a(0.005457645282149315)),(to_sfixed_a(0.00011600468860706314)),(to_sfixed_a(-0.00019995582988485694)),(to_sfixed_a(0.5986126661300659)),(to_sfixed_a(0.20387957990169525)),(to_sfixed_a(0.023038554936647415)),(to_sfixed_a(0.00011262798943789676)),(to_sfixed_a(8.498769602738321e-05)),(to_sfixed_a(2.2000240278430283e-05)),(to_sfixed_a(-0.6207098364830017)),(to_sfixed_a(0.0014990366762503982)),(to_sfixed_a(2.4364413548028097e-05)),(to_sfixed_a(-0.008735956624150276)),(to_sfixed_a(-0.008825716562569141)),(to_sfixed_a(0.000133632798679173)),(to_sfixed_a(-0.002525895368307829)),(to_sfixed_a(-0.004249706398695707)),(to_sfixed_a(-0.0002371462614974007)),(to_sfixed_a(0.3685876429080963)),(to_sfixed_a(-0.009383628144860268)),(to_sfixed_a(-0.0007709068013355136)),(to_sfixed_a(7.338091381825507e-05)),(to_sfixed_a(-0.0001542674144729972)),(to_sfixed_a(-0.23833118379116058)),(to_sfixed_a(0.00015572833945043385)),(to_sfixed_a(-0.001439245999790728)),(to_sfixed_a(-6.862953887321055e-05)),(to_sfixed_a(0.00092216458870098)),(to_sfixed_a(0.0001771360111888498)),(to_sfixed_a(7.670201739529148e-05)),(to_sfixed_a(-0.00024905853206291795)),(to_sfixed_a(-4.016206366941333e-05)),(to_sfixed_a(-0.00010556009510764852)),(to_sfixed_a(-0.004089174326509237)),(to_sfixed_a(0.1168941855430603)),(to_sfixed_a(-0.00017857100465334952)),(to_sfixed_a(-0.0034771498758345842)),(to_sfixed_a(-0.00772574357688427)),(to_sfixed_a(-0.0018678288906812668)),(to_sfixed_a(4.812987754121423e-05)),(to_sfixed_a(-7.163180271163583e-05)),(to_sfixed_a(-6.697513163089752e-05)),(to_sfixed_a(-0.006738561205565929)),(to_sfixed_a(0.002435801550745964)),(to_sfixed_a(-0.00011258300219196826)),(to_sfixed_a(0.34728533029556274)),(to_sfixed_a(-1.0783867764985189e-05)),(to_sfixed_a(-0.00016681471606716514)),(to_sfixed_a(0.0002713938301894814)),(to_sfixed_a(-4.0621835069032386e-05)),(to_sfixed_a(0.10653361678123474)),(to_sfixed_a(0.00017982663121074438)),(to_sfixed_a(0.016139835119247437)),(to_sfixed_a(-6.602045323234051e-05)),(to_sfixed_a(-4.686835745815188e-05)),(to_sfixed_a(-0.0015544717898592353)),(to_sfixed_a(0.0002141063887393102)),(to_sfixed_a(-0.0002033460041275248)),(to_sfixed_a(0.19485773146152496)),(to_sfixed_a(0.4109900891780853)),(to_sfixed_a(-3.59692785423249e-06)),(to_sfixed_a(0.00045595946721732616)),(to_sfixed_a(-1.0647459930623882e-05)),(to_sfixed_a(-0.00015926289779599756)),(to_sfixed_a(-2.388664142927155e-05)),(to_sfixed_a(-0.007383468095213175)),(to_sfixed_a(-0.00313379243016243)),(to_sfixed_a(0.00014824709796812385)),(to_sfixed_a(8.159878780134022e-05)),(to_sfixed_a(-0.29484814405441284)),(to_sfixed_a(-0.0009610339184291661)),(to_sfixed_a(-0.0002041292900685221)),(to_sfixed_a(-0.00018026292673312128)),(to_sfixed_a(-0.0018627388635650277)),(to_sfixed_a(-5.9200880059506744e-05)),(to_sfixed_a(0.00021951261442154646)),(to_sfixed_a(-3.6155746784061193e-05)),(to_sfixed_a(-0.003084699623286724)),(to_sfixed_a(0.0004354623379185796)),(to_sfixed_a(-0.0002437312068650499)),(to_sfixed_a(-0.00016641156980767846)),(to_sfixed_a(0.0002678119344636798)),(to_sfixed_a(-0.00946077425032854)),(to_sfixed_a(6.850197678431869e-05)),(to_sfixed_a(2.9136666853446513e-05)),(to_sfixed_a(0.01105524506419897)),(to_sfixed_a(0.00024690382997505367)),(to_sfixed_a(-2.5728288164827973e-05)),(to_sfixed_a(-0.01544303260743618)),(to_sfixed_a(0.00010773746180348098)),(to_sfixed_a(0.2725464105606079)),(to_sfixed_a(-9.217687875207048e-06)),(to_sfixed_a(0.0001527147978777066)),(to_sfixed_a(1.5031393559183925e-05)),(to_sfixed_a(5.735524609917775e-05)),(to_sfixed_a(-0.01306064147502184)),(to_sfixed_a(-0.14463426172733307)),(to_sfixed_a(0.0006487774662673473)),(to_sfixed_a(-0.0023428495042026043)),(to_sfixed_a(6.930597010068595e-05)),(to_sfixed_a(-0.0028383927419781685)),(to_sfixed_a(-2.660058089531958e-05)),(to_sfixed_a(0.00025038758758455515)),(to_sfixed_a(0.022440966218709946)),(to_sfixed_a(-0.005014393012970686)),(to_sfixed_a(0.2144973874092102)),(to_sfixed_a(-0.0001496670302003622)),(to_sfixed_a(-0.3263079822063446)),(to_sfixed_a(0.002610051305964589)),(to_sfixed_a(-0.014528017491102219)),(to_sfixed_a(0.5686203241348267)),(to_sfixed_a(0.005336398724466562)),(to_sfixed_a(0.5708157420158386)),(to_sfixed_a(-0.0013053251896053553)),(to_sfixed_a(0.3106392025947571)),(to_sfixed_a(-0.00010981281957356259)),(to_sfixed_a(-0.00013513531303033233)),(to_sfixed_a(0.00010127086716238409)),(to_sfixed_a(-0.007114870939403772)),(to_sfixed_a(0.164879709482193)),(to_sfixed_a(-0.0016627503791823983)),(to_sfixed_a(-0.000504982890561223)),(to_sfixed_a(0.0023900577798485756)),(to_sfixed_a(0.05127459391951561)),(to_sfixed_a(-0.0001022517099045217)),(to_sfixed_a(0.04300256446003914)),(to_sfixed_a(0.8589792847633362)),(to_sfixed_a(-0.00024605204816907644)),(to_sfixed_a(0.22087708115577698)),(to_sfixed_a(1.934784813784063e-05)),(to_sfixed_a(-0.0024650900159031153)),(to_sfixed_a(-0.35493072867393494)),(to_sfixed_a(-0.00012907445488963276)),(to_sfixed_a(-2.9497525247279555e-05)),(to_sfixed_a(7.159746019169688e-05)),(to_sfixed_a(0.00022855821589473635)),(to_sfixed_a(0.00011205676855752245)),(to_sfixed_a(0.00011382062803022563)),(to_sfixed_a(0.001040955656208098)),(to_sfixed_a(-0.005220034159719944)),(to_sfixed_a(0.0006657622870989144)),(to_sfixed_a(-0.00047540635569021106)),(to_sfixed_a(0.0008414684562012553)),(to_sfixed_a(0.001752527547068894)),(to_sfixed_a(-0.00010206384467892349)),(to_sfixed_a(4.7012981667649e-06)),(to_sfixed_a(-4.729527063318528e-07)),(to_sfixed_a(0.00013334950199350715)),(to_sfixed_a(0.0001523162063676864)),(to_sfixed_a(-0.0004134805058129132)),(to_sfixed_a(-0.0009143078350462019)),(to_sfixed_a(0.04143020883202553)),(to_sfixed_a(1.797145523596555e-05)),(to_sfixed_a(0.000114310416392982)),(to_sfixed_a(5.087217141408473e-05)),(to_sfixed_a(-0.00010213847417617217)),(to_sfixed_a(-8.466149301966652e-05)),(to_sfixed_a(-0.006268705241382122)),(to_sfixed_a(0.00015697386697866023)),(to_sfixed_a(-0.0001562699762871489)),(to_sfixed_a(-2.808934368658811e-06)),(to_sfixed_a(0.12520337104797363)),(to_sfixed_a(0.00010550805018283427)),(to_sfixed_a(0.35643449425697327)),(to_sfixed_a(3.1298783142119646e-05)),(to_sfixed_a(-0.00010329947690479457)),(to_sfixed_a(0.00012710466398857534)),(to_sfixed_a(0.0018887600162997842)),(to_sfixed_a(-0.0063262986950576305)),(to_sfixed_a(-0.327739953994751)),(to_sfixed_a(-0.0002188713406212628)),(to_sfixed_a(-0.007089283317327499)),(to_sfixed_a(0.00018496123084332794)),(to_sfixed_a(-0.0038371486589312553)),(to_sfixed_a(0.0002546425967011601)),(to_sfixed_a(-0.0018011742504313588)),(to_sfixed_a(0.00010760745499283075)),(to_sfixed_a(0.27926602959632874)),(to_sfixed_a(-0.16011837124824524)),(to_sfixed_a(0.6544234752655029)),(to_sfixed_a(-0.15444201231002808)),(to_sfixed_a(-7.153092883527279e-05)),(to_sfixed_a(-0.0050894999876618385)),(to_sfixed_a(0.35051029920578003)),(to_sfixed_a(-0.0003121210902463645)),(to_sfixed_a(0.02743520587682724)),(to_sfixed_a(-0.0001898403570521623)),(to_sfixed_a(-5.124092785990797e-05)),(to_sfixed_a(0.01441105268895626)),(to_sfixed_a(-0.31547772884368896)),(to_sfixed_a(1.110518496716395e-06)),(to_sfixed_a(-2.3715107090538368e-05)),(to_sfixed_a(0.0002866737195290625)),(to_sfixed_a(-8.552592771593481e-05)),(to_sfixed_a(-0.0004375509452074766)),(to_sfixed_a(-6.644320819759741e-05)),(to_sfixed_a(0.00018927236669696867)),(to_sfixed_a(0.00010126369306817651)),(to_sfixed_a(0.032989148050546646)),(to_sfixed_a(-7.162358815548941e-05)),(to_sfixed_a(-0.00012897266424261034)),(to_sfixed_a(-0.00022420461755245924)),(to_sfixed_a(-0.009083881974220276)),(to_sfixed_a(0.2582983374595642)),(to_sfixed_a(-8.463135600322857e-05)),(to_sfixed_a(7.147174619603902e-05)),(to_sfixed_a(1.4550023479387164e-05)),(to_sfixed_a(4.6118970203679055e-05)),(to_sfixed_a(0.005072717554867268)),(to_sfixed_a(-0.0013570144074037671)),(to_sfixed_a(-0.0031695072539150715)),(to_sfixed_a(-0.27563008666038513)),(to_sfixed_a(0.29249078035354614)),(to_sfixed_a(4.8378511564806104e-05)),(to_sfixed_a(-0.0001502070517744869)),(to_sfixed_a(-1.1576004908420146e-05)),(to_sfixed_a(0.0002499710244592279)),(to_sfixed_a(-0.0002517577086109668)),(to_sfixed_a(-7.744766480755061e-05)),(to_sfixed_a(7.797535363351926e-05)),(to_sfixed_a(0.004307487513870001)),(to_sfixed_a(-0.0002954292867798358)),(to_sfixed_a(-0.032857123762369156)),(to_sfixed_a(0.0013111305888742208)),(to_sfixed_a(-0.005054905079305172)),(to_sfixed_a(-0.22358866035938263)),(to_sfixed_a(-0.00012728874571621418)),(to_sfixed_a(-0.3585370182991028)),(to_sfixed_a(0.032951951026916504)),(to_sfixed_a(-0.008690509013831615)),(to_sfixed_a(0.00018347424338571727)),(to_sfixed_a(-0.008506666868925095)),(to_sfixed_a(0.16056282818317413)),(to_sfixed_a(-0.0023817250039428473)));

    constant weight_n2_25 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.22908887267112732)),(to_sfixed_a(-0.0054564750753343105)),(to_sfixed_a(0.0021839826367795467)),(to_sfixed_a(0.00011471040488686413)),(to_sfixed_a(0.0035078527871519327)),(to_sfixed_a(-2.3576350940857083e-05)),(to_sfixed_a(-0.006442875135689974)),(to_sfixed_a(0.00031537419999949634)),(to_sfixed_a(-2.5592184101697057e-05)),(to_sfixed_a(0.0001313475368078798)),(to_sfixed_a(-0.00024035823298618197)),(to_sfixed_a(0.0007094548782333732)),(to_sfixed_a(-0.00041595182847231627)),(to_sfixed_a(-0.3662119507789612)),(to_sfixed_a(0.00020034135377500206)),(to_sfixed_a(0.00021950394148007035)),(to_sfixed_a(0.002192101441323757)),(to_sfixed_a(-0.0002039372338913381)),(to_sfixed_a(0.005742703098803759)),(to_sfixed_a(-0.0007459074258804321)),(to_sfixed_a(0.00012681499356403947)),(to_sfixed_a(-0.00014228688087314367)),(to_sfixed_a(0.0007738901767879725)),(to_sfixed_a(0.004559989552944899)),(to_sfixed_a(-0.0014315618900582194)),(to_sfixed_a(0.004794507287442684)),(to_sfixed_a(0.00012800171680282801)),(to_sfixed_a(0.000993158551864326)),(to_sfixed_a(-0.0003772139607463032)),(to_sfixed_a(-6.761113763786852e-05)),(to_sfixed_a(-0.009772188030183315)),(to_sfixed_a(-2.4950713850557804e-07)),(to_sfixed_a(-0.08730515837669373)),(to_sfixed_a(0.00010171016765525565)),(to_sfixed_a(-0.00016745677567087114)),(to_sfixed_a(-0.00015707846614532173)),(to_sfixed_a(0.44031304121017456)),(to_sfixed_a(0.0019132659072056413)),(to_sfixed_a(0.21389925479888916)),(to_sfixed_a(6.931422103662044e-05)),(to_sfixed_a(-0.008100013248622417)),(to_sfixed_a(-0.18306376039981842)),(to_sfixed_a(-0.00020238840079400688)),(to_sfixed_a(-4.5024782593827695e-05)),(to_sfixed_a(-0.012631318531930447)),(to_sfixed_a(0.15875844657421112)),(to_sfixed_a(0.008065213449299335)),(to_sfixed_a(-0.00949055515229702)),(to_sfixed_a(-3.622781514422968e-05)),(to_sfixed_a(-0.005159047432243824)),(to_sfixed_a(-0.004051427356898785)),(to_sfixed_a(-1.6432180927949958e-05)),(to_sfixed_a(-0.00015628288383595645)),(to_sfixed_a(0.2480953484773636)),(to_sfixed_a(-0.3998611271381378)),(to_sfixed_a(0.0025684675201773643)),(to_sfixed_a(0.00015281932428479195)),(to_sfixed_a(-0.01412036083638668)),(to_sfixed_a(1.2365089787635952e-06)),(to_sfixed_a(-6.952178955543786e-05)),(to_sfixed_a(-0.007438825909048319)),(to_sfixed_a(-0.0024633107241243124)),(to_sfixed_a(0.0006629124982282519)),(to_sfixed_a(-0.0015692553715780377)),(to_sfixed_a(-8.724729559617117e-05)),(to_sfixed_a(0.0023032338358461857)),(to_sfixed_a(-0.0001886385289253667)),(to_sfixed_a(-0.27936166524887085)),(to_sfixed_a(0.0011831086594611406)),(to_sfixed_a(0.00018283766985405236)),(to_sfixed_a(0.2355106621980667)),(to_sfixed_a(-0.00023826338292565197)),(to_sfixed_a(-0.011969671584665775)),(to_sfixed_a(8.725142106413841e-05)),(to_sfixed_a(8.405770495301113e-05)),(to_sfixed_a(-3.204419408575632e-05)),(to_sfixed_a(-0.010198628529906273)),(to_sfixed_a(0.1535019427537918)),(to_sfixed_a(-3.7866640923311934e-05)),(to_sfixed_a(-0.019157694652676582)),(to_sfixed_a(-0.015042931772768497)),(to_sfixed_a(6.250301521504298e-05)),(to_sfixed_a(0.0001716826664051041)),(to_sfixed_a(0.0007815977442078292)),(to_sfixed_a(-4.8610003432258964e-05)),(to_sfixed_a(0.08476261794567108)),(to_sfixed_a(-0.007411366794258356)),(to_sfixed_a(-0.3810429275035858)),(to_sfixed_a(-2.6688889192882925e-05)),(to_sfixed_a(0.0001504574902355671)),(to_sfixed_a(-0.29660311341285706)),(to_sfixed_a(-5.994362072669901e-05)),(to_sfixed_a(-0.00330339465290308)),(to_sfixed_a(0.00010403061605757102)),(to_sfixed_a(-0.0002902280248235911)),(to_sfixed_a(4.2752209992613643e-05)),(to_sfixed_a(-0.0003164074441883713)),(to_sfixed_a(0.00011502404231578112)),(to_sfixed_a(4.7772235120646656e-05)),(to_sfixed_a(-7.065344834700227e-05)),(to_sfixed_a(-0.030339384451508522)),(to_sfixed_a(-0.004237711895257235)),(to_sfixed_a(-6.257370114326477e-05)),(to_sfixed_a(-0.004226064775139093)),(to_sfixed_a(0.21249130368232727)),(to_sfixed_a(-0.005985627416521311)),(to_sfixed_a(-0.0001519415236543864)),(to_sfixed_a(7.175150676630437e-05)),(to_sfixed_a(-2.9571117920568213e-05)),(to_sfixed_a(0.4357320964336395)),(to_sfixed_a(-0.005448195151984692)),(to_sfixed_a(-0.00016596975910943002)),(to_sfixed_a(0.30367156863212585)),(to_sfixed_a(4.454445661394857e-05)),(to_sfixed_a(-7.097599882399663e-05)),(to_sfixed_a(0.35098883509635925)),(to_sfixed_a(0.007386626675724983)),(to_sfixed_a(0.17765012383460999)),(to_sfixed_a(0.00012812550994567573)),(to_sfixed_a(-0.00024219317128881812)),(to_sfixed_a(-1.973274993360974e-05)),(to_sfixed_a(-0.00012954085832461715)),(to_sfixed_a(0.0022934735752642155)),(to_sfixed_a(-1.5960009477566928e-05)),(to_sfixed_a(-2.7994014089927077e-05)),(to_sfixed_a(-0.0014986175810918212)),(to_sfixed_a(-0.010062376968562603)),(to_sfixed_a(-6.769434548914433e-05)),(to_sfixed_a(0.0002312685683136806)),(to_sfixed_a(-0.00014591269427910447)),(to_sfixed_a(7.803246262483299e-05)),(to_sfixed_a(0.00025467269006185234)),(to_sfixed_a(-0.0013205134309828281)),(to_sfixed_a(-0.0035843881778419018)),(to_sfixed_a(-0.00021465659665409476)),(to_sfixed_a(-0.00019880807667504996)),(to_sfixed_a(-0.11054351180791855)),(to_sfixed_a(0.00021638484031427652)),(to_sfixed_a(0.00028272782219573855)),(to_sfixed_a(1.6547484847251326e-05)),(to_sfixed_a(0.002360597951337695)),(to_sfixed_a(0.00015349246677942574)),(to_sfixed_a(0.00022723941947333515)),(to_sfixed_a(0.0038336748257279396)),(to_sfixed_a(-0.0013717253459617496)),(to_sfixed_a(0.0003158029867336154)),(to_sfixed_a(0.000542360998224467)),(to_sfixed_a(0.000178095608134754)),(to_sfixed_a(2.198218135163188e-05)),(to_sfixed_a(-0.001382395625114441)),(to_sfixed_a(-6.36213953839615e-05)),(to_sfixed_a(0.00025171582819893956)),(to_sfixed_a(0.013117838650941849)),(to_sfixed_a(-0.00017401372315362096)),(to_sfixed_a(0.0001672574580879882)),(to_sfixed_a(-0.014417284168303013)),(to_sfixed_a(-9.958484588423744e-05)),(to_sfixed_a(-0.3658658564090729)),(to_sfixed_a(0.00014013810141477734)),(to_sfixed_a(1.0884505172725767e-06)),(to_sfixed_a(8.5665044025518e-05)),(to_sfixed_a(0.00015647217514924705)),(to_sfixed_a(-0.03996562957763672)),(to_sfixed_a(0.0001574325142428279)),(to_sfixed_a(-0.0026101183611899614)),(to_sfixed_a(0.004186027683317661)),(to_sfixed_a(8.002617687452585e-05)),(to_sfixed_a(-0.3625428378582001)),(to_sfixed_a(-0.00016732298536226153)),(to_sfixed_a(0.0002466518199071288)),(to_sfixed_a(-0.2371986210346222)),(to_sfixed_a(0.0027192106936126947)),(to_sfixed_a(-0.002583342371508479)),(to_sfixed_a(0.00016109587159007788)),(to_sfixed_a(-0.36020320653915405)),(to_sfixed_a(0.0005205305642448366)),(to_sfixed_a(-0.00323665258474648)),(to_sfixed_a(-0.0022252569906413555)),(to_sfixed_a(0.0024212144780904055)),(to_sfixed_a(0.025282640010118484)),(to_sfixed_a(-0.0016933886799961329)),(to_sfixed_a(-0.0006532333209179342)),(to_sfixed_a(9.612303983885795e-07)),(to_sfixed_a(3.238274439354427e-05)),(to_sfixed_a(-0.0001680447458056733)),(to_sfixed_a(-0.016150547191500664)),(to_sfixed_a(-0.008637518621981144)),(to_sfixed_a(0.006045751739293337)),(to_sfixed_a(-0.00019818302826024592)),(to_sfixed_a(0.003658619709312916)),(to_sfixed_a(0.0002382617094554007)),(to_sfixed_a(0.0001974753977265209)),(to_sfixed_a(-0.007024062797427177)),(to_sfixed_a(-0.0020366059616208076)),(to_sfixed_a(2.0817813492612913e-05)),(to_sfixed_a(0.009685062803328037)),(to_sfixed_a(-7.190606265794486e-05)),(to_sfixed_a(-0.013907943852245808)),(to_sfixed_a(-0.0003218345227651298)),(to_sfixed_a(-2.7291607693769038e-05)),(to_sfixed_a(-0.00015545345377177)),(to_sfixed_a(-0.00024293683236464858)),(to_sfixed_a(-0.00022201221145223826)),(to_sfixed_a(0.00013617021613754332)),(to_sfixed_a(0.00011827429989352822)),(to_sfixed_a(0.0009028201457113028)),(to_sfixed_a(0.4336002767086029)),(to_sfixed_a(0.0006489657680504024)),(to_sfixed_a(-0.002139573683962226)),(to_sfixed_a(-0.0010722798760980368)),(to_sfixed_a(-0.0017388842534273863)),(to_sfixed_a(0.0003839307464659214)),(to_sfixed_a(-4.449206608114764e-05)),(to_sfixed_a(0.00018357791122980416)),(to_sfixed_a(0.00013592702453024685)),(to_sfixed_a(0.00011244734923820943)),(to_sfixed_a(-0.0029736533761024475)),(to_sfixed_a(0.005169199779629707)),(to_sfixed_a(-0.00022376692504622042)),(to_sfixed_a(-2.8061462217010558e-05)),(to_sfixed_a(-0.00010187839507125318)),(to_sfixed_a(-0.00011633911344688386)),(to_sfixed_a(0.00022373348474502563)),(to_sfixed_a(0.008056213147938251)),(to_sfixed_a(0.4064154028892517)),(to_sfixed_a(-0.00024240394122898579)),(to_sfixed_a(-0.00016745508764870465)),(to_sfixed_a(0.00020174961537122726)),(to_sfixed_a(0.0018479895079508424)),(to_sfixed_a(-0.0018173661082983017)),(to_sfixed_a(0.0010313724633306265)),(to_sfixed_a(-0.0002739891642704606)),(to_sfixed_a(-0.00032321488833986223)),(to_sfixed_a(-7.160750101320446e-05)),(to_sfixed_a(-0.0014370118733495474)),(to_sfixed_a(-0.0019389030057936907)),(to_sfixed_a(-0.002871623495593667)),(to_sfixed_a(0.0001281403237953782)),(to_sfixed_a(-0.0061820209957659245)),(to_sfixed_a(6.499643495772034e-05)),(to_sfixed_a(-0.011478143744170666)),(to_sfixed_a(0.00017921249673236161)),(to_sfixed_a(-0.009048733860254288)),(to_sfixed_a(-6.063302862457931e-06)),(to_sfixed_a(0.16862079501152039)),(to_sfixed_a(0.00040171589353121817)),(to_sfixed_a(-0.1706760823726654)),(to_sfixed_a(-0.004296215251088142)),(to_sfixed_a(0.0001901151263155043)),(to_sfixed_a(-0.0031535623129457235)),(to_sfixed_a(-0.02119571529328823)),(to_sfixed_a(9.784513531485572e-05)),(to_sfixed_a(-0.00015748391160741448)),(to_sfixed_a(-2.7941163352807052e-05)),(to_sfixed_a(-0.0003631055005826056)),(to_sfixed_a(0.005671270657330751)),(to_sfixed_a(-0.3686721920967102)),(to_sfixed_a(0.00024075205146800727)),(to_sfixed_a(-0.00017044477863237262)),(to_sfixed_a(-0.322306364774704)),(to_sfixed_a(-6.043697430868633e-05)),(to_sfixed_a(0.00029914037440903485)),(to_sfixed_a(-0.00015845980669837445)),(to_sfixed_a(-0.0006423743907362223)),(to_sfixed_a(2.1964562620269135e-05)),(to_sfixed_a(-0.005648287944495678)),(to_sfixed_a(1.8154518329538405e-05)),(to_sfixed_a(6.979958561714739e-05)),(to_sfixed_a(7.687544712098315e-05)),(to_sfixed_a(-0.008601787500083447)),(to_sfixed_a(-0.00820598192512989)),(to_sfixed_a(6.246486736927181e-05)),(to_sfixed_a(-0.00028478758758865297)),(to_sfixed_a(-1.538598007755354e-05)),(to_sfixed_a(7.801854371791705e-05)),(to_sfixed_a(0.0020917130168527365)),(to_sfixed_a(-0.012204010970890522)),(to_sfixed_a(-0.005805215332657099)),(to_sfixed_a(-0.012340179644525051)),(to_sfixed_a(0.0019275123486295342)),(to_sfixed_a(-8.613162935944274e-05)),(to_sfixed_a(0.00015804977738298476)),(to_sfixed_a(0.00018943767645396292)),(to_sfixed_a(-0.0006542212795466185)),(to_sfixed_a(-5.7750632549868897e-05)),(to_sfixed_a(0.00016708450857549906)),(to_sfixed_a(-6.462451710831374e-05)),(to_sfixed_a(-0.0016793133690953255)),(to_sfixed_a(-8.452514884993434e-05)),(to_sfixed_a(0.6577464938163757)),(to_sfixed_a(-0.00022107359836809337)),(to_sfixed_a(-0.0067246584221720695)),(to_sfixed_a(0.2240648865699768)),(to_sfixed_a(4.761855598189868e-05)),(to_sfixed_a(0.0007873408030718565)),(to_sfixed_a(-5.974393570795655e-05)),(to_sfixed_a(-0.01701628975570202)),(to_sfixed_a(1.2833552318625152e-05)),(to_sfixed_a(-0.1379455327987671)),(to_sfixed_a(0.007007647305727005)),(to_sfixed_a(-0.01380130648612976)));

    constant weight_n2_26 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.021776597946882248)),(to_sfixed_a(0.0017841795925050974)),(to_sfixed_a(0.0011494741775095463)),(to_sfixed_a(7.584603736177087e-07)),(to_sfixed_a(0.0010069875279441476)),(to_sfixed_a(-0.00015535650891251862)),(to_sfixed_a(0.0008552999352104962)),(to_sfixed_a(-0.00011381899821572006)),(to_sfixed_a(-0.00010337097046431154)),(to_sfixed_a(-0.0001369499950669706)),(to_sfixed_a(-0.00029706419445574284)),(to_sfixed_a(0.003992440644651651)),(to_sfixed_a(-0.0033624358475208282)),(to_sfixed_a(0.0014317861059680581)),(to_sfixed_a(-6.423273589462042e-06)),(to_sfixed_a(-1.800331665435806e-05)),(to_sfixed_a(0.0031986499670892954)),(to_sfixed_a(6.707872671540827e-05)),(to_sfixed_a(0.16780595481395721)),(to_sfixed_a(-0.008408678695559502)),(to_sfixed_a(0.0001192386043840088)),(to_sfixed_a(-6.833251245552674e-05)),(to_sfixed_a(9.32245166040957e-05)),(to_sfixed_a(0.0031321337446570396)),(to_sfixed_a(0.402463436126709)),(to_sfixed_a(0.005123774986714125)),(to_sfixed_a(1.0827738151419908e-05)),(to_sfixed_a(0.001152532291598618)),(to_sfixed_a(0.0013106337282806635)),(to_sfixed_a(0.0002474552602507174)),(to_sfixed_a(-0.002250035060569644)),(to_sfixed_a(-7.340918091358617e-05)),(to_sfixed_a(-0.006580764893442392)),(to_sfixed_a(-0.00010009811376221478)),(to_sfixed_a(2.476633744663559e-05)),(to_sfixed_a(0.0002184579207096249)),(to_sfixed_a(0.00879125390201807)),(to_sfixed_a(0.002177075482904911)),(to_sfixed_a(0.0075420052744448185)),(to_sfixed_a(0.00018386486044619232)),(to_sfixed_a(-0.004065193701535463)),(to_sfixed_a(-0.0025128074921667576)),(to_sfixed_a(-0.00021585123613476753)),(to_sfixed_a(5.7426252169534564e-05)),(to_sfixed_a(-0.008784604258835316)),(to_sfixed_a(-0.008302433416247368)),(to_sfixed_a(0.011069243773818016)),(to_sfixed_a(-0.003474793629720807)),(to_sfixed_a(-1.6013806089176796e-05)),(to_sfixed_a(-0.6579181551933289)),(to_sfixed_a(0.0002607267815619707)),(to_sfixed_a(0.0003180591156706214)),(to_sfixed_a(-0.00017475835920777172)),(to_sfixed_a(0.004714962560683489)),(to_sfixed_a(-0.013142582960426807)),(to_sfixed_a(0.005417496431618929)),(to_sfixed_a(0.00020062396652065217)),(to_sfixed_a(-0.005126284435391426)),(to_sfixed_a(5.4398969950852916e-05)),(to_sfixed_a(5.71870623389259e-05)),(to_sfixed_a(-0.0013964733807370067)),(to_sfixed_a(3.329625178594142e-05)),(to_sfixed_a(0.002147993305698037)),(to_sfixed_a(0.005829667206853628)),(to_sfixed_a(0.00030520843574777246)),(to_sfixed_a(0.0002575037651695311)),(to_sfixed_a(2.171382584492676e-05)),(to_sfixed_a(-0.004880223888903856)),(to_sfixed_a(0.004600990563631058)),(to_sfixed_a(-4.000324406661093e-05)),(to_sfixed_a(0.267440527677536)),(to_sfixed_a(0.001663879374973476)),(to_sfixed_a(-0.00021099903096910566)),(to_sfixed_a(3.972927515860647e-05)),(to_sfixed_a(0.0001895792520372197)),(to_sfixed_a(1.1126685421913862e-06)),(to_sfixed_a(0.007677823770791292)),(to_sfixed_a(0.0033899054396897554)),(to_sfixed_a(-1.1965323210461065e-05)),(to_sfixed_a(0.007140756584703922)),(to_sfixed_a(-0.002052535070106387)),(to_sfixed_a(-2.943087019957602e-05)),(to_sfixed_a(0.00383395585231483)),(to_sfixed_a(-0.0010765264742076397)),(to_sfixed_a(-0.0001674321829341352)),(to_sfixed_a(0.0012156144948676229)),(to_sfixed_a(-0.0079996008425951)),(to_sfixed_a(0.003965808544307947)),(to_sfixed_a(0.00021549421944655478)),(to_sfixed_a(-0.00022036988229956478)),(to_sfixed_a(-0.013427896425127983)),(to_sfixed_a(6.3702646002639085e-06)),(to_sfixed_a(0.0003264604602009058)),(to_sfixed_a(2.449868043186143e-05)),(to_sfixed_a(6.903967005200684e-05)),(to_sfixed_a(0.0001394017308484763)),(to_sfixed_a(-1.6285324818454683e-05)),(to_sfixed_a(-0.0001992170000448823)),(to_sfixed_a(6.096804645494558e-05)),(to_sfixed_a(-0.00016403812333010137)),(to_sfixed_a(-0.002594137331470847)),(to_sfixed_a(0.0002967806067317724)),(to_sfixed_a(-0.00020574158406816423)),(to_sfixed_a(0.0023582158610224724)),(to_sfixed_a(0.24678684771060944)),(to_sfixed_a(0.0011443805415183306)),(to_sfixed_a(-2.6326575607527047e-05)),(to_sfixed_a(-2.0826730178669095e-05)),(to_sfixed_a(0.00010761411977000535)),(to_sfixed_a(0.28047096729278564)),(to_sfixed_a(-0.002592534525319934)),(to_sfixed_a(0.00011593222006922588)),(to_sfixed_a(0.20077736675739288)),(to_sfixed_a(4.309884388931096e-06)),(to_sfixed_a(-7.042322249617428e-05)),(to_sfixed_a(0.009732292033731937)),(to_sfixed_a(-0.0003648572019301355)),(to_sfixed_a(-0.0006164031801745296)),(to_sfixed_a(0.000460665236460045)),(to_sfixed_a(-0.002126254141330719)),(to_sfixed_a(-0.00010903614747803658)),(to_sfixed_a(4.267050462658517e-05)),(to_sfixed_a(0.0033251189161092043)),(to_sfixed_a(0.0001301220036111772)),(to_sfixed_a(-2.0788296751561575e-05)),(to_sfixed_a(-0.005045880563557148)),(to_sfixed_a(0.016186799854040146)),(to_sfixed_a(-0.00010054469748865813)),(to_sfixed_a(0.0002708836691454053)),(to_sfixed_a(2.377669807174243e-05)),(to_sfixed_a(-0.0002483384741935879)),(to_sfixed_a(-3.605811798479408e-05)),(to_sfixed_a(0.0035976471845060587)),(to_sfixed_a(0.0014495623763650656)),(to_sfixed_a(-2.0471452444326133e-06)),(to_sfixed_a(0.00015417163376696408)),(to_sfixed_a(0.0023750904947519302)),(to_sfixed_a(0.0023510728497058153)),(to_sfixed_a(0.00017451427993364632)),(to_sfixed_a(0.00030132741085253656)),(to_sfixed_a(0.0035163331776857376)),(to_sfixed_a(-3.3739790524123237e-05)),(to_sfixed_a(-0.0002854603808373213)),(to_sfixed_a(-0.00028036447474732995)),(to_sfixed_a(-0.0002319652121514082)),(to_sfixed_a(-0.0005421589594334364)),(to_sfixed_a(0.008873991668224335)),(to_sfixed_a(-0.00015652697766199708)),(to_sfixed_a(-6.27471599727869e-05)),(to_sfixed_a(-0.0003024313773494214)),(to_sfixed_a(5.849735316587612e-05)),(to_sfixed_a(1.5809520846232772e-05)),(to_sfixed_a(0.007888483814895153)),(to_sfixed_a(2.232371480204165e-05)),(to_sfixed_a(-5.682138362317346e-05)),(to_sfixed_a(0.0012783356942236423)),(to_sfixed_a(0.00011542998254299164)),(to_sfixed_a(3.530579851940274e-05)),(to_sfixed_a(-3.736191865755245e-05)),(to_sfixed_a(-0.00016209244495257735)),(to_sfixed_a(0.0001119118242058903)),(to_sfixed_a(-0.0001499366044299677)),(to_sfixed_a(-0.04906325042247772)),(to_sfixed_a(-0.0005160677246749401)),(to_sfixed_a(0.0006866347976028919)),(to_sfixed_a(0.005763010121881962)),(to_sfixed_a(-2.4573069822508842e-05)),(to_sfixed_a(0.007809040602296591)),(to_sfixed_a(6.650872091995552e-05)),(to_sfixed_a(0.0002391050657024607)),(to_sfixed_a(-0.34749504923820496)),(to_sfixed_a(0.005267228931188583)),(to_sfixed_a(-0.00030761578818783164)),(to_sfixed_a(2.3971017071744427e-05)),(to_sfixed_a(-0.0353008396923542)),(to_sfixed_a(-0.00028045845101587474)),(to_sfixed_a(-0.01913396082818508)),(to_sfixed_a(0.0012562114279717207)),(to_sfixed_a(-0.004589605610817671)),(to_sfixed_a(-0.0059991939924657345)),(to_sfixed_a(0.00031654458143748343)),(to_sfixed_a(0.35200318694114685)),(to_sfixed_a(-6.713056791340932e-06)),(to_sfixed_a(-9.601717465557158e-06)),(to_sfixed_a(1.9538951164577156e-05)),(to_sfixed_a(-0.0036487041506916285)),(to_sfixed_a(0.0016682149143889546)),(to_sfixed_a(0.008027319796383381)),(to_sfixed_a(-0.00015793388593010604)),(to_sfixed_a(0.00527891144156456)),(to_sfixed_a(-0.018513960763812065)),(to_sfixed_a(-8.281676127808169e-05)),(to_sfixed_a(0.000681049597915262)),(to_sfixed_a(0.0005061063566245139)),(to_sfixed_a(-0.00029797005117870867)),(to_sfixed_a(0.0040320889092981815)),(to_sfixed_a(6.995821604505181e-05)),(to_sfixed_a(0.01651817001402378)),(to_sfixed_a(-0.2550760805606842)),(to_sfixed_a(-3.34442884195596e-05)),(to_sfixed_a(-1.101009183912538e-05)),(to_sfixed_a(0.00010888907127082348)),(to_sfixed_a(-0.00011484952847240493)),(to_sfixed_a(6.162298086564988e-05)),(to_sfixed_a(-0.0001793049304978922)),(to_sfixed_a(0.0026666277553886175)),(to_sfixed_a(-0.006662403699010611)),(to_sfixed_a(-0.003001728095114231)),(to_sfixed_a(0.001714246696792543)),(to_sfixed_a(0.001791816670447588)),(to_sfixed_a(-0.003463378408923745)),(to_sfixed_a(-6.744932034052908e-05)),(to_sfixed_a(0.00019184699340257794)),(to_sfixed_a(-1.4658100553788245e-05)),(to_sfixed_a(0.0001518595963716507)),(to_sfixed_a(-0.0003896860289387405)),(to_sfixed_a(-0.00175719172693789)),(to_sfixed_a(0.0004349874798208475)),(to_sfixed_a(0.0025870823301374912)),(to_sfixed_a(4.5289722038432956e-05)),(to_sfixed_a(1.6716148820705712e-05)),(to_sfixed_a(-6.977262091822922e-05)),(to_sfixed_a(-6.575811130460352e-05)),(to_sfixed_a(0.0030637148302048445)),(to_sfixed_a(-0.0003741166146937758)),(to_sfixed_a(1.792408511391841e-05)),(to_sfixed_a(6.729083543177694e-05)),(to_sfixed_a(-0.00030410493491217494)),(to_sfixed_a(0.002142622834071517)),(to_sfixed_a(-0.4294225871562958)),(to_sfixed_a(0.01041337102651596)),(to_sfixed_a(1.165449430118315e-05)),(to_sfixed_a(0.00018422806169837713)),(to_sfixed_a(-0.00022076811001170427)),(to_sfixed_a(-0.0010965504916384816)),(to_sfixed_a(0.0004384409112390131)),(to_sfixed_a(0.002963010687381029)),(to_sfixed_a(-0.00017989129992201924)),(to_sfixed_a(0.0011549690971150994)),(to_sfixed_a(-8.504577272105962e-05)),(to_sfixed_a(0.004481269512325525)),(to_sfixed_a(-0.00010544410906732082)),(to_sfixed_a(-0.7089309096336365)),(to_sfixed_a(4.460480704437941e-05)),(to_sfixed_a(0.3644261658191681)),(to_sfixed_a(-3.4256663639098406e-05)),(to_sfixed_a(-0.005467666313052177)),(to_sfixed_a(0.0020404579117894173)),(to_sfixed_a(0.0002259578468510881)),(to_sfixed_a(-0.0040612476877868176)),(to_sfixed_a(-0.010637267492711544)),(to_sfixed_a(2.811285958159715e-05)),(to_sfixed_a(-0.0009912926470860839)),(to_sfixed_a(-5.568601409322582e-05)),(to_sfixed_a(-0.00021085049957036972)),(to_sfixed_a(0.007314430084079504)),(to_sfixed_a(-0.2548344135284424)),(to_sfixed_a(0.00015776744112372398)),(to_sfixed_a(0.00020565729937516153)),(to_sfixed_a(1.927014091052115e-05)),(to_sfixed_a(0.00010432115232106298)),(to_sfixed_a(-0.00038563026464544237)),(to_sfixed_a(0.00018054993415717036)),(to_sfixed_a(-0.00011164296302013099)),(to_sfixed_a(0.00011426466517150402)),(to_sfixed_a(-0.003552217036485672)),(to_sfixed_a(-2.9469854780472815e-05)),(to_sfixed_a(-2.054107426374685e-05)),(to_sfixed_a(1.141789834946394e-05)),(to_sfixed_a(0.00014905496209394187)),(to_sfixed_a(0.004556911066174507)),(to_sfixed_a(-4.764823825098574e-05)),(to_sfixed_a(7.031227141851559e-05)),(to_sfixed_a(-0.00023746714578010142)),(to_sfixed_a(0.00031503470381721854)),(to_sfixed_a(0.0055690729059278965)),(to_sfixed_a(0.0003472113166935742)),(to_sfixed_a(0.0003864557947963476)),(to_sfixed_a(0.02193610928952694)),(to_sfixed_a(0.0002790904836729169)),(to_sfixed_a(2.46259369305335e-05)),(to_sfixed_a(-0.00020046619465574622)),(to_sfixed_a(-0.0001173273049062118)),(to_sfixed_a(-0.013265428133308887)),(to_sfixed_a(-0.00011620323493843898)),(to_sfixed_a(8.636301208753139e-05)),(to_sfixed_a(-0.00803012028336525)),(to_sfixed_a(9.144106297753751e-05)),(to_sfixed_a(6.526104698423296e-05)),(to_sfixed_a(2.9774848371744156e-05)),(to_sfixed_a(0.0015765102580189705)),(to_sfixed_a(-0.002411839086562395)),(to_sfixed_a(0.24469149112701416)),(to_sfixed_a(0.00023915016208775342)),(to_sfixed_a(0.0035604943986982107)),(to_sfixed_a(0.0009816100355237722)),(to_sfixed_a(-0.004052609670907259)),(to_sfixed_a(-1.0502320947125554e-05)),(to_sfixed_a(-0.0008541597053408623)),(to_sfixed_a(-0.06872319430112839)),(to_sfixed_a(-0.008504407480359077)));

    constant weight_n2_27 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.3945747911930084)),(to_sfixed_a(0.002678975462913513)),(to_sfixed_a(5.647700163535774e-06)),(to_sfixed_a(8.352406439371407e-05)),(to_sfixed_a(-0.0010481131030246615)),(to_sfixed_a(-0.00012902787420898676)),(to_sfixed_a(-0.006054192315787077)),(to_sfixed_a(4.2616899008862674e-05)),(to_sfixed_a(5.325578968040645e-06)),(to_sfixed_a(4.935952165396884e-05)),(to_sfixed_a(-0.00030941603472456336)),(to_sfixed_a(-0.00028335078968666494)),(to_sfixed_a(-0.00015048834029585123)),(to_sfixed_a(0.0033157896250486374)),(to_sfixed_a(0.00022039300529286265)),(to_sfixed_a(-0.00023067645088303834)),(to_sfixed_a(1.844398502726108e-05)),(to_sfixed_a(5.1562401495175436e-05)),(to_sfixed_a(0.006898511201143265)),(to_sfixed_a(0.0022202422842383385)),(to_sfixed_a(0.00017721632320899516)),(to_sfixed_a(4.944644388160668e-05)),(to_sfixed_a(-0.0036940108984708786)),(to_sfixed_a(-0.0002832530881278217)),(to_sfixed_a(-0.004193633329123259)),(to_sfixed_a(0.0024833427742123604)),(to_sfixed_a(0.00011430876475060359)),(to_sfixed_a(5.203930049901828e-05)),(to_sfixed_a(0.00017217136337421834)),(to_sfixed_a(-1.8529550288803875e-05)),(to_sfixed_a(-0.23520368337631226)),(to_sfixed_a(-9.519479499431327e-05)),(to_sfixed_a(-0.0012267085257917643)),(to_sfixed_a(9.529784438200295e-05)),(to_sfixed_a(-0.00013191477046348155)),(to_sfixed_a(9.536610741633922e-05)),(to_sfixed_a(0.00242648646235466)),(to_sfixed_a(0.00020612127264030278)),(to_sfixed_a(-0.014088072814047337)),(to_sfixed_a(-4.276793333701789e-06)),(to_sfixed_a(-0.0006502943579107523)),(to_sfixed_a(0.00024178664898499846)),(to_sfixed_a(7.171643665060401e-05)),(to_sfixed_a(1.8627571989782155e-05)),(to_sfixed_a(-0.011780851520597935)),(to_sfixed_a(-0.01830378547310829)),(to_sfixed_a(0.004547119606286287)),(to_sfixed_a(-7.895694579929113e-06)),(to_sfixed_a(-2.741160278674215e-05)),(to_sfixed_a(-0.0008084827568382025)),(to_sfixed_a(-0.0017027115682139993)),(to_sfixed_a(-0.0008688982925377786)),(to_sfixed_a(-0.00026800986961461604)),(to_sfixed_a(0.001901485724374652)),(to_sfixed_a(-0.31533920764923096)),(to_sfixed_a(-0.0028343666344881058)),(to_sfixed_a(-0.00015669240383431315)),(to_sfixed_a(-0.011457514017820358)),(to_sfixed_a(0.00013675828813575208)),(to_sfixed_a(-2.3628050257684663e-05)),(to_sfixed_a(-0.007643624674528837)),(to_sfixed_a(-0.005934292450547218)),(to_sfixed_a(3.580521297408268e-05)),(to_sfixed_a(-0.0035029808059334755)),(to_sfixed_a(5.921746196690947e-05)),(to_sfixed_a(-0.28057974576950073)),(to_sfixed_a(1.9382929167477414e-05)),(to_sfixed_a(-0.017417408525943756)),(to_sfixed_a(-0.005782690364867449)),(to_sfixed_a(-0.00014872806787025183)),(to_sfixed_a(0.0011577900731936097)),(to_sfixed_a(-0.0019532882142812014)),(to_sfixed_a(0.0017467649886384606)),(to_sfixed_a(1.849301224865485e-05)),(to_sfixed_a(3.407601616345346e-05)),(to_sfixed_a(6.848287011962384e-05)),(to_sfixed_a(-0.008229807019233704)),(to_sfixed_a(-0.003305082442238927)),(to_sfixed_a(7.167353760451078e-05)),(to_sfixed_a(0.011228539049625397)),(to_sfixed_a(-0.005356526002287865)),(to_sfixed_a(-0.00020498523372225463)),(to_sfixed_a(-0.0004697589611168951)),(to_sfixed_a(0.0028813902754336596)),(to_sfixed_a(-6.455342372646555e-06)),(to_sfixed_a(-0.0027784158010035753)),(to_sfixed_a(0.006038884166628122)),(to_sfixed_a(-7.873345020925626e-05)),(to_sfixed_a(0.00013630202738568187)),(to_sfixed_a(-3.8332673284457996e-05)),(to_sfixed_a(-0.0076779574155807495)),(to_sfixed_a(-1.3679098628927022e-05)),(to_sfixed_a(-0.01163195725530386)),(to_sfixed_a(7.80942355049774e-06)),(to_sfixed_a(-0.0024883602745831013)),(to_sfixed_a(6.162810313981026e-05)),(to_sfixed_a(-2.3853881430113688e-05)),(to_sfixed_a(-0.00015329004963859916)),(to_sfixed_a(2.2466909285867587e-05)),(to_sfixed_a(1.1409538274165243e-05)),(to_sfixed_a(-0.00015465937030967325)),(to_sfixed_a(-0.0015813976060599089)),(to_sfixed_a(-2.1375517462729476e-05)),(to_sfixed_a(-0.0064525422640144825)),(to_sfixed_a(-0.006561228074133396)),(to_sfixed_a(-5.849204171681777e-06)),(to_sfixed_a(0.00010311471851309761)),(to_sfixed_a(-3.299106901977211e-05)),(to_sfixed_a(4.3628690036712214e-05)),(to_sfixed_a(-0.0032752426341176033)),(to_sfixed_a(0.3203054368495941)),(to_sfixed_a(0.00011246032227063552)),(to_sfixed_a(-0.22746826708316803)),(to_sfixed_a(-3.97861294914037e-05)),(to_sfixed_a(6.939256854820997e-05)),(to_sfixed_a(-0.029720844700932503)),(to_sfixed_a(-7.417535380227491e-05)),(to_sfixed_a(-0.0014992662472650409)),(to_sfixed_a(0.00041858546319417655)),(to_sfixed_a(-0.49700039625167847)),(to_sfixed_a(-0.00015182344941422343)),(to_sfixed_a(6.76584750181064e-05)),(to_sfixed_a(-0.006694457959383726)),(to_sfixed_a(0.000166009966051206)),(to_sfixed_a(-0.00011784253001678735)),(to_sfixed_a(-0.0008847907884046435)),(to_sfixed_a(0.21878787875175476)),(to_sfixed_a(4.85443088109605e-05)),(to_sfixed_a(-0.00022545702813658863)),(to_sfixed_a(0.00023807062825653702)),(to_sfixed_a(0.00014822445518802851)),(to_sfixed_a(9.218116247211583e-06)),(to_sfixed_a(-1.6444508219137788e-05)),(to_sfixed_a(0.21310050785541534)),(to_sfixed_a(4.823332346859388e-05)),(to_sfixed_a(1.221153070218861e-06)),(to_sfixed_a(-0.013159768655896187)),(to_sfixed_a(-5.777166006737389e-05)),(to_sfixed_a(0.00011835931945824996)),(to_sfixed_a(-2.9466886189766228e-05)),(to_sfixed_a(-0.0035101445391774178)),(to_sfixed_a(-8.412000897806138e-05)),(to_sfixed_a(0.0002436190115986392)),(to_sfixed_a(3.4964035876328126e-05)),(to_sfixed_a(0.0011842899257317185)),(to_sfixed_a(-8.238392183557153e-05)),(to_sfixed_a(-0.0014110232004895806)),(to_sfixed_a(4.683396764448844e-05)),(to_sfixed_a(-0.00011235734564252198)),(to_sfixed_a(-0.30170944333076477)),(to_sfixed_a(-0.00018226589600089937)),(to_sfixed_a(-4.4141983380541205e-05)),(to_sfixed_a(-9.413794032298028e-05)),(to_sfixed_a(0.00023940458777360618)),(to_sfixed_a(-0.00042089540511369705)),(to_sfixed_a(0.0007292110240086913)),(to_sfixed_a(0.00017611427756492049)),(to_sfixed_a(-0.0028879919555038214)),(to_sfixed_a(2.5931049094651826e-05)),(to_sfixed_a(0.00014690466923639178)),(to_sfixed_a(-1.510561560280621e-06)),(to_sfixed_a(-4.028093826491386e-06)),(to_sfixed_a(0.0010390359675511718)),(to_sfixed_a(0.0005966742755845189)),(to_sfixed_a(-0.00035443244269117713)),(to_sfixed_a(-0.0005518483812920749)),(to_sfixed_a(2.618201688164845e-05)),(to_sfixed_a(-0.5067739486694336)),(to_sfixed_a(6.552630657097325e-05)),(to_sfixed_a(-2.208107616752386e-06)),(to_sfixed_a(-0.10808759182691574)),(to_sfixed_a(0.0011569017078727484)),(to_sfixed_a(-0.00022110072313807905)),(to_sfixed_a(-0.0003080377937294543)),(to_sfixed_a(-0.00033056316897273064)),(to_sfixed_a(-3.995973020209931e-05)),(to_sfixed_a(0.0005078878602944314)),(to_sfixed_a(-7.8778357419651e-06)),(to_sfixed_a(-0.48801398277282715)),(to_sfixed_a(-0.010963665321469307)),(to_sfixed_a(-7.045390520943329e-05)),(to_sfixed_a(-0.0023348797112703323)),(to_sfixed_a(-0.0001076374901458621)),(to_sfixed_a(-0.00011971628555329517)),(to_sfixed_a(-0.0001738895516609773)),(to_sfixed_a(3.3172596886288375e-05)),(to_sfixed_a(-0.0011362722143530846)),(to_sfixed_a(-0.0007072364678606391)),(to_sfixed_a(0.0017171099316328764)),(to_sfixed_a(0.0072283209301531315)),(to_sfixed_a(0.00811983272433281)),(to_sfixed_a(-2.968954504467547e-07)),(to_sfixed_a(-0.0026285359635949135)),(to_sfixed_a(-0.010268473997712135)),(to_sfixed_a(-0.00014810469292569906)),(to_sfixed_a(-0.00022312965302262455)),(to_sfixed_a(0.00015023717423900962)),(to_sfixed_a(-0.016070181503891945)),(to_sfixed_a(-0.0009386481833644211)),(to_sfixed_a(-0.00016875960864126682)),(to_sfixed_a(5.137342668604106e-06)),(to_sfixed_a(-0.00015017417899798602)),(to_sfixed_a(-2.0202605810482055e-05)),(to_sfixed_a(-0.00017761434719432145)),(to_sfixed_a(1.738710852805525e-05)),(to_sfixed_a(0.0014361431822180748)),(to_sfixed_a(-9.446934564039111e-05)),(to_sfixed_a(0.003741001943126321)),(to_sfixed_a(0.15699037909507751)),(to_sfixed_a(-0.0012102436739951372)),(to_sfixed_a(0.0007285326719284058)),(to_sfixed_a(-0.0001491512666689232)),(to_sfixed_a(-9.771336772246286e-05)),(to_sfixed_a(7.109741272870451e-05)),(to_sfixed_a(-6.76937197567895e-05)),(to_sfixed_a(7.67353194532916e-05)),(to_sfixed_a(0.0004916305770166218)),(to_sfixed_a(-0.0018443920416757464)),(to_sfixed_a(-0.00033952019293792546)),(to_sfixed_a(-0.0001354933192487806)),(to_sfixed_a(6.728289008606225e-05)),(to_sfixed_a(-8.322895155288279e-07)),(to_sfixed_a(-4.333784818300046e-05)),(to_sfixed_a(-1.2065816918038763e-05)),(to_sfixed_a(-0.008322183042764664)),(to_sfixed_a(5.765722744399682e-05)),(to_sfixed_a(-4.8100308049470186e-05)),(to_sfixed_a(-0.0004458497860468924)),(to_sfixed_a(-0.006683585699647665)),(to_sfixed_a(-0.004359838552772999)),(to_sfixed_a(0.005424456670880318)),(to_sfixed_a(-5.802288433187641e-05)),(to_sfixed_a(0.00013659156684298068)),(to_sfixed_a(-0.0001973019097931683)),(to_sfixed_a(-0.007775625679641962)),(to_sfixed_a(-0.004314923658967018)),(to_sfixed_a(-0.005146995652467012)),(to_sfixed_a(-0.00012843958393204957)),(to_sfixed_a(0.0022400766611099243)),(to_sfixed_a(-0.0002877078950405121)),(to_sfixed_a(0.004745206795632839)),(to_sfixed_a(-1.1748488759621978e-07)),(to_sfixed_a(-0.2648521065711975)),(to_sfixed_a(-0.00010627335723256692)),(to_sfixed_a(0.196771040558815)),(to_sfixed_a(0.0007090161670930684)),(to_sfixed_a(-0.010841228067874908)),(to_sfixed_a(-0.0038280778098851442)),(to_sfixed_a(0.00014861903036944568)),(to_sfixed_a(-0.017789600417017937)),(to_sfixed_a(0.0005630620289593935)),(to_sfixed_a(-6.755820504622534e-05)),(to_sfixed_a(0.0002085115120280534)),(to_sfixed_a(1.8559268937679008e-05)),(to_sfixed_a(-2.6810068447957747e-05)),(to_sfixed_a(-0.006234811153262854)),(to_sfixed_a(0.005582098849117756)),(to_sfixed_a(-4.922670268570073e-05)),(to_sfixed_a(6.1758270021528e-05)),(to_sfixed_a(8.484508725814521e-06)),(to_sfixed_a(0.0002811008598655462)),(to_sfixed_a(0.00010612922051222995)),(to_sfixed_a(1.1458920198492706e-05)),(to_sfixed_a(0.00018169338000006974)),(to_sfixed_a(2.3615539248567075e-05)),(to_sfixed_a(-3.377949178684503e-05)),(to_sfixed_a(0.0002140251745004207)),(to_sfixed_a(-3.869244392262772e-05)),(to_sfixed_a(0.00018687243573367596)),(to_sfixed_a(-0.0010395750869065523)),(to_sfixed_a(0.0025098216719925404)),(to_sfixed_a(-0.00012462338781915605)),(to_sfixed_a(0.00030116175184957683)),(to_sfixed_a(0.0001862348581198603)),(to_sfixed_a(0.00011172172526130453)),(to_sfixed_a(-0.00536264618858695)),(to_sfixed_a(-0.0020441352389752865)),(to_sfixed_a(-0.13592815399169922)),(to_sfixed_a(-0.002194294473156333)),(to_sfixed_a(0.0018864823505282402)),(to_sfixed_a(6.449406646424904e-05)),(to_sfixed_a(-2.2865497157908976e-05)),(to_sfixed_a(-0.0002516281383577734)),(to_sfixed_a(0.001850197440944612)),(to_sfixed_a(-1.4199395081959665e-06)),(to_sfixed_a(0.00018144688510801643)),(to_sfixed_a(0.0017438243376091123)),(to_sfixed_a(-0.0011082583805546165)),(to_sfixed_a(-0.00010318773274775594)),(to_sfixed_a(3.524088970152661e-05)),(to_sfixed_a(-0.0005490445182658732)),(to_sfixed_a(0.17048688232898712)),(to_sfixed_a(-0.008019988425076008)),(to_sfixed_a(2.5551016733516008e-06)),(to_sfixed_a(-0.0018655144376680255)),(to_sfixed_a(6.36367331026122e-05)),(to_sfixed_a(-0.009237980470061302)),(to_sfixed_a(-0.00013302027946338058)),(to_sfixed_a(-0.008761080913245678)),(to_sfixed_a(0.4774526357650757)),(to_sfixed_a(-0.017631765455007553)));

    constant weight_n2_28 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.1396181583404541)),(to_sfixed_a(0.0012213055742904544)),(to_sfixed_a(0.0004084015963599086)),(to_sfixed_a(-0.000171108782524243)),(to_sfixed_a(0.17084182798862457)),(to_sfixed_a(7.671496132388711e-05)),(to_sfixed_a(0.0034967774990946054)),(to_sfixed_a(1.9603212422225624e-06)),(to_sfixed_a(0.00015649254783056676)),(to_sfixed_a(-3.770920739043504e-05)),(to_sfixed_a(-0.00015466850891243666)),(to_sfixed_a(0.00019833685655612499)),(to_sfixed_a(-0.00832045916467905)),(to_sfixed_a(0.009437683038413525)),(to_sfixed_a(3.204375389032066e-06)),(to_sfixed_a(0.00015828352479729801)),(to_sfixed_a(-0.5068323612213135)),(to_sfixed_a(7.605871360283345e-05)),(to_sfixed_a(0.29754358530044556)),(to_sfixed_a(0.0011058590607717633)),(to_sfixed_a(-0.00010560686496319249)),(to_sfixed_a(7.528760761488229e-06)),(to_sfixed_a(-0.0005179743748158216)),(to_sfixed_a(0.0037300889380276203)),(to_sfixed_a(-0.006112344563007355)),(to_sfixed_a(0.0008847886929288507)),(to_sfixed_a(-0.00011407829879317433)),(to_sfixed_a(-0.00010368691437179223)),(to_sfixed_a(-0.0009379631374031305)),(to_sfixed_a(-0.00015952804824337363)),(to_sfixed_a(-0.0020800866186618805)),(to_sfixed_a(-0.00010689436749089509)),(to_sfixed_a(0.002038128674030304)),(to_sfixed_a(2.057322853943333e-05)),(to_sfixed_a(-0.00019305750902276486)),(to_sfixed_a(-9.733445767778903e-05)),(to_sfixed_a(-0.025001544505357742)),(to_sfixed_a(0.013843764550983906)),(to_sfixed_a(-0.2920585870742798)),(to_sfixed_a(0.00021771145111415535)),(to_sfixed_a(0.031484898179769516)),(to_sfixed_a(0.0014191147638484836)),(to_sfixed_a(-5.0624239520402625e-05)),(to_sfixed_a(0.00011118005204480141)),(to_sfixed_a(0.23233471810817719)),(to_sfixed_a(-0.010518782772123814)),(to_sfixed_a(0.0016041755443438888)),(to_sfixed_a(-0.010370871052145958)),(to_sfixed_a(-0.00019896247249562293)),(to_sfixed_a(-0.0040463292971253395)),(to_sfixed_a(-0.012076782993972301)),(to_sfixed_a(0.28456273674964905)),(to_sfixed_a(0.0004111723101232201)),(to_sfixed_a(0.0010168339358642697)),(to_sfixed_a(-0.008044159039855003)),(to_sfixed_a(-0.0068946173414587975)),(to_sfixed_a(0.00023796138702891767)),(to_sfixed_a(-0.005775582045316696)),(to_sfixed_a(-0.00010402061889180914)),(to_sfixed_a(6.933954864507541e-05)),(to_sfixed_a(-0.00011075561633333564)),(to_sfixed_a(0.0015707224374637008)),(to_sfixed_a(-0.0012093388941138983)),(to_sfixed_a(-0.0059240213595330715)),(to_sfixed_a(0.00024214065342675894)),(to_sfixed_a(0.00169561302755028)),(to_sfixed_a(-6.540038157254457e-05)),(to_sfixed_a(0.26093214750289917)),(to_sfixed_a(-0.00036259344778954983)),(to_sfixed_a(6.738974479958415e-05)),(to_sfixed_a(0.03654303774237633)),(to_sfixed_a(0.00034595493343658745)),(to_sfixed_a(0.0007889201515354216)),(to_sfixed_a(3.8933445466682315e-05)),(to_sfixed_a(3.8271580706350505e-05)),(to_sfixed_a(-1.4140343409962952e-05)),(to_sfixed_a(0.006906557362526655)),(to_sfixed_a(-0.0019996047485619783)),(to_sfixed_a(-0.00017946148000191897)),(to_sfixed_a(-0.0076257530599832535)),(to_sfixed_a(0.0008798405760899186)),(to_sfixed_a(4.594199708662927e-06)),(to_sfixed_a(0.03247736021876335)),(to_sfixed_a(0.0005714254803024232)),(to_sfixed_a(-3.900037336279638e-05)),(to_sfixed_a(0.0019533359445631504)),(to_sfixed_a(0.00731235183775425)),(to_sfixed_a(0.0017002519452944398)),(to_sfixed_a(7.207602175185457e-05)),(to_sfixed_a(2.392436726950109e-06)),(to_sfixed_a(0.4552931487560272)),(to_sfixed_a(-3.7291549233486876e-05)),(to_sfixed_a(-0.014969353564083576)),(to_sfixed_a(0.00016698919353075325)),(to_sfixed_a(0.016535025089979172)),(to_sfixed_a(5.3821040637558326e-05)),(to_sfixed_a(0.00023660734586883336)),(to_sfixed_a(0.00010176563955610618)),(to_sfixed_a(6.762361590517685e-05)),(to_sfixed_a(7.904483936727047e-05)),(to_sfixed_a(-0.0114089110866189)),(to_sfixed_a(-0.003054323373362422)),(to_sfixed_a(-0.00018941942835226655)),(to_sfixed_a(-0.012540651485323906)),(to_sfixed_a(0.0011514873476698995)),(to_sfixed_a(-0.0018767138244584203)),(to_sfixed_a(0.00013140957162249833)),(to_sfixed_a(0.00011231019016122445)),(to_sfixed_a(0.00017982185818254948)),(to_sfixed_a(-0.005355113185942173)),(to_sfixed_a(-0.0087936632335186)),(to_sfixed_a(8.5452564235311e-05)),(to_sfixed_a(-0.0011220461456105113)),(to_sfixed_a(0.0001145887072198093)),(to_sfixed_a(-2.440023308736272e-05)),(to_sfixed_a(0.014963651075959206)),(to_sfixed_a(0.0005884958081878722)),(to_sfixed_a(-0.00021427747560665011)),(to_sfixed_a(-8.441526733804494e-05)),(to_sfixed_a(0.00037512643029913306)),(to_sfixed_a(-5.7589706557337195e-05)),(to_sfixed_a(-5.890654938411899e-05)),(to_sfixed_a(-0.0016629266319796443)),(to_sfixed_a(-0.00016746504115872085)),(to_sfixed_a(-0.00010024869698099792)),(to_sfixed_a(-0.0017826742259785533)),(to_sfixed_a(-0.018887115642428398)),(to_sfixed_a(0.00027931557269766927)),(to_sfixed_a(-0.00031358757405541837)),(to_sfixed_a(2.5511006242595613e-05)),(to_sfixed_a(0.00010701864812290296)),(to_sfixed_a(0.00013313023373484612)),(to_sfixed_a(-0.00014960765838623047)),(to_sfixed_a(0.0053934333845973015)),(to_sfixed_a(1.665690797381103e-05)),(to_sfixed_a(2.120858698617667e-05)),(to_sfixed_a(0.0005110778147354722)),(to_sfixed_a(0.0006056437850929797)),(to_sfixed_a(-3.4868280636146665e-05)),(to_sfixed_a(0.00017013688920997083)),(to_sfixed_a(0.00020390894496813416)),(to_sfixed_a(0.00010565081902313977)),(to_sfixed_a(-0.00015356589574366808)),(to_sfixed_a(-9.663639502832666e-05)),(to_sfixed_a(0.0008425968699157238)),(to_sfixed_a(9.072971442947164e-05)),(to_sfixed_a(-0.0019327247282490134)),(to_sfixed_a(-0.00014654977712780237)),(to_sfixed_a(0.0002537665714044124)),(to_sfixed_a(0.005332122556865215)),(to_sfixed_a(-2.7968126232735813e-06)),(to_sfixed_a(5.927679012529552e-05)),(to_sfixed_a(-0.004964440129697323)),(to_sfixed_a(0.00022367150813806802)),(to_sfixed_a(9.85333463177085e-06)),(to_sfixed_a(-0.06664910167455673)),(to_sfixed_a(-8.960880222730339e-05)),(to_sfixed_a(0.002031586365774274)),(to_sfixed_a(-4.902907312498428e-05)),(to_sfixed_a(1.3574725016951561e-05)),(to_sfixed_a(0.00016741572471801192)),(to_sfixed_a(0.0001553594775032252)),(to_sfixed_a(-0.01326053962111473)),(to_sfixed_a(-0.3529176115989685)),(to_sfixed_a(-0.012103228829801083)),(to_sfixed_a(0.005972560029476881)),(to_sfixed_a(0.00011295820877421647)),(to_sfixed_a(0.5330820679664612)),(to_sfixed_a(-0.0001745241752360016)),(to_sfixed_a(7.290480425581336e-06)),(to_sfixed_a(0.2801356017589569)),(to_sfixed_a(0.0021880818530917168)),(to_sfixed_a(-0.001474652555771172)),(to_sfixed_a(-0.00011334215378155932)),(to_sfixed_a(-0.0004273719678167254)),(to_sfixed_a(0.00014011353778187186)),(to_sfixed_a(0.0018878330010920763)),(to_sfixed_a(-6.591719284188002e-05)),(to_sfixed_a(0.00090839306358248)),(to_sfixed_a(-0.0015150457620620728)),(to_sfixed_a(-3.0528779461747035e-05)),(to_sfixed_a(0.013117445632815361)),(to_sfixed_a(-4.235764208715409e-06)),(to_sfixed_a(0.00019441574113443494)),(to_sfixed_a(0.0001740763254929334)),(to_sfixed_a(-0.005563780199736357)),(to_sfixed_a(-0.0009912934619933367)),(to_sfixed_a(0.12752848863601685)),(to_sfixed_a(0.00041424736264161766)),(to_sfixed_a(0.6062530279159546)),(to_sfixed_a(0.008893477730453014)),(to_sfixed_a(3.0079318094067276e-05)),(to_sfixed_a(-0.0014858122449368238)),(to_sfixed_a(0.0005282765487208962)),(to_sfixed_a(6.820060661993921e-06)),(to_sfixed_a(-0.22905832529067993)),(to_sfixed_a(9.833202057052404e-05)),(to_sfixed_a(-0.012681239284574986)),(to_sfixed_a(-0.006659320555627346)),(to_sfixed_a(-0.0001763436885084957)),(to_sfixed_a(-3.676906635519117e-05)),(to_sfixed_a(-3.152425051666796e-05)),(to_sfixed_a(2.0053648768225685e-06)),(to_sfixed_a(-0.00017471579485572875)),(to_sfixed_a(0.0001546390849398449)),(to_sfixed_a(0.00020578652038238943)),(to_sfixed_a(0.007925011217594147)),(to_sfixed_a(0.011649630032479763)),(to_sfixed_a(-0.0005907166632823646)),(to_sfixed_a(-0.0050287083722651005)),(to_sfixed_a(0.6169032454490662)),(to_sfixed_a(-7.001751509960741e-05)),(to_sfixed_a(-0.00023714388953521848)),(to_sfixed_a(0.00016166025307029486)),(to_sfixed_a(-0.00014811269647907466)),(to_sfixed_a(0.00014047115109860897)),(to_sfixed_a(-0.38642677664756775)),(to_sfixed_a(0.0018952462123706937)),(to_sfixed_a(-0.004880488850176334)),(to_sfixed_a(-1.9736966351047158e-05)),(to_sfixed_a(8.676011202624068e-05)),(to_sfixed_a(0.00011216150596737862)),(to_sfixed_a(0.00015065929619595408)),(to_sfixed_a(-0.003543959930539131)),(to_sfixed_a(-0.0028643691912293434)),(to_sfixed_a(6.280378147494048e-05)),(to_sfixed_a(0.0001566229184390977)),(to_sfixed_a(0.00020037285867147148)),(to_sfixed_a(-0.0007200978579930961)),(to_sfixed_a(-0.0004570427699945867)),(to_sfixed_a(0.0013257942628115416)),(to_sfixed_a(0.00010947513510473073)),(to_sfixed_a(8.741066267248243e-05)),(to_sfixed_a(0.00010279544949298725)),(to_sfixed_a(-0.001246530213393271)),(to_sfixed_a(0.008119492791593075)),(to_sfixed_a(0.18520468473434448)),(to_sfixed_a(-1.87696423381567e-06)),(to_sfixed_a(0.00013838664744980633)),(to_sfixed_a(-2.4542532628402114e-05)),(to_sfixed_a(-0.0017770257545635104)),(to_sfixed_a(-0.00022240464750211686)),(to_sfixed_a(0.004675713367760181)),(to_sfixed_a(-0.00020470740855671465)),(to_sfixed_a(-0.3404686748981476)),(to_sfixed_a(0.00046721185208298266)),(to_sfixed_a(-0.4207470417022705)),(to_sfixed_a(-0.006719781551510096)),(to_sfixed_a(3.605925303418189e-05)),(to_sfixed_a(-0.003036681329831481)),(to_sfixed_a(-0.011808391660451889)),(to_sfixed_a(0.00018295453628525138)),(to_sfixed_a(0.0011716751614585519)),(to_sfixed_a(7.049560372252017e-05)),(to_sfixed_a(-0.0001413310965290293)),(to_sfixed_a(-0.199205219745636)),(to_sfixed_a(0.16712217032909393)),(to_sfixed_a(7.3569390224292874e-06)),(to_sfixed_a(-0.00015155179426074028)),(to_sfixed_a(0.0020393035374581814)),(to_sfixed_a(-2.4380351533181965e-05)),(to_sfixed_a(-0.00618555024266243)),(to_sfixed_a(0.00023685020278207958)),(to_sfixed_a(0.00038806803058832884)),(to_sfixed_a(-0.00020653118554037064)),(to_sfixed_a(-0.019919661805033684)),(to_sfixed_a(-0.00018629623809829354)),(to_sfixed_a(-0.0002477607340551913)),(to_sfixed_a(-2.6305948267690837e-05)),(to_sfixed_a(0.005648574326187372)),(to_sfixed_a(0.26814839243888855)),(to_sfixed_a(-5.615357804344967e-05)),(to_sfixed_a(-0.00017722498159855604)),(to_sfixed_a(-0.000119275129691232)),(to_sfixed_a(-0.00010090766591019928)),(to_sfixed_a(-0.44686082005500793)),(to_sfixed_a(-0.012091506272554398)),(to_sfixed_a(0.15693624317646027)),(to_sfixed_a(0.06869406253099442)),(to_sfixed_a(-0.00255345506593585)),(to_sfixed_a(0.00015298239304684103)),(to_sfixed_a(-4.6701414248673245e-05)),(to_sfixed_a(-0.00022982610971666873)),(to_sfixed_a(0.0029211982619017363)),(to_sfixed_a(9.29415546124801e-06)),(to_sfixed_a(0.00011475123028503731)),(to_sfixed_a(0.2523277997970581)),(to_sfixed_a(-0.012307550758123398)),(to_sfixed_a(-0.00015046804037410766)),(to_sfixed_a(-0.00015414318477269262)),(to_sfixed_a(0.16467052698135376)),(to_sfixed_a(-0.011813831515610218)),(to_sfixed_a(-0.23207399249076843)),(to_sfixed_a(5.0465299864299595e-05)),(to_sfixed_a(-0.0033043138682842255)),(to_sfixed_a(0.003445050911977887)),(to_sfixed_a(0.2641240656375885)),(to_sfixed_a(9.09978843992576e-05)),(to_sfixed_a(0.0680234432220459)),(to_sfixed_a(0.40796324610710144)),(to_sfixed_a(-0.015909047797322273)));

    constant weight_n2_29 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.1886346936225891)),(to_sfixed_a(-9.794760262593627e-05)),(to_sfixed_a(-0.45873597264289856)),(to_sfixed_a(-0.00021605368237942457)),(to_sfixed_a(-0.005974547937512398)),(to_sfixed_a(-2.2306732716970146e-05)),(to_sfixed_a(-0.0023085607681423426)),(to_sfixed_a(-7.005862426012754e-05)),(to_sfixed_a(-0.0001166767324320972)),(to_sfixed_a(-1.6019883332774043e-05)),(to_sfixed_a(-0.00024564852355979383)),(to_sfixed_a(0.015640797093510628)),(to_sfixed_a(0.1593257039785385)),(to_sfixed_a(0.0040280637331306934)),(to_sfixed_a(-5.916597729083151e-06)),(to_sfixed_a(0.0001300169969908893)),(to_sfixed_a(-0.035437703132629395)),(to_sfixed_a(0.00010157293581869453)),(to_sfixed_a(0.005627037957310677)),(to_sfixed_a(0.3543590307235718)),(to_sfixed_a(-5.879503441974521e-05)),(to_sfixed_a(-0.0001409813412465155)),(to_sfixed_a(0.0008943973225541413)),(to_sfixed_a(0.004295276012271643)),(to_sfixed_a(-0.005616846960037947)),(to_sfixed_a(-0.001427796552889049)),(to_sfixed_a(0.0001546338462503627)),(to_sfixed_a(-0.001090467325411737)),(to_sfixed_a(-0.0051674204878509045)),(to_sfixed_a(-0.00018380532856099308)),(to_sfixed_a(0.011735028587281704)),(to_sfixed_a(-0.0002890007453970611)),(to_sfixed_a(0.14632943272590637)),(to_sfixed_a(0.0004140334203839302)),(to_sfixed_a(-2.780579961836338e-05)),(to_sfixed_a(0.0001432380231563002)),(to_sfixed_a(-0.07788018137216568)),(to_sfixed_a(0.015242730267345905)),(to_sfixed_a(0.008442189544439316)),(to_sfixed_a(7.708849443588406e-05)),(to_sfixed_a(-0.5064061284065247)),(to_sfixed_a(0.350050151348114)),(to_sfixed_a(6.927407230250537e-05)),(to_sfixed_a(1.8643011571839452e-05)),(to_sfixed_a(-0.015507293865084648)),(to_sfixed_a(-0.004118715412914753)),(to_sfixed_a(-0.3266949951648712)),(to_sfixed_a(-0.16725118458271027)),(to_sfixed_a(2.5091852876357734e-05)),(to_sfixed_a(0.31365346908569336)),(to_sfixed_a(-0.030335096642374992)),(to_sfixed_a(-0.0011511852499097586)),(to_sfixed_a(-1.0268988262396306e-05)),(to_sfixed_a(-0.0015073930844664574)),(to_sfixed_a(0.294001966714859)),(to_sfixed_a(0.00048430211609229445)),(to_sfixed_a(-7.060762436594814e-05)),(to_sfixed_a(-0.002677589189261198)),(to_sfixed_a(-0.00010193274647463113)),(to_sfixed_a(-3.918290894944221e-05)),(to_sfixed_a(-0.001933942548930645)),(to_sfixed_a(0.0012898354325443506)),(to_sfixed_a(0.24017377197742462)),(to_sfixed_a(0.13633286952972412)),(to_sfixed_a(-4.321339656598866e-05)),(to_sfixed_a(0.0024133112747222185)),(to_sfixed_a(-5.745723319705576e-05)),(to_sfixed_a(0.19369487464427948)),(to_sfixed_a(-0.004468641243875027)),(to_sfixed_a(0.00011962158896494657)),(to_sfixed_a(-0.2421727329492569)),(to_sfixed_a(-0.6946342587471008)),(to_sfixed_a(-0.011577890254557133)),(to_sfixed_a(1.3949334970675409e-05)),(to_sfixed_a(0.00024424653383903205)),(to_sfixed_a(2.9203833037172444e-05)),(to_sfixed_a(0.0027947539929300547)),(to_sfixed_a(-0.0006794423097744584)),(to_sfixed_a(-3.813311195699498e-07)),(to_sfixed_a(-0.008202405646443367)),(to_sfixed_a(-0.0011206412455067039)),(to_sfixed_a(6.98221629136242e-05)),(to_sfixed_a(-0.001622926676645875)),(to_sfixed_a(-0.0006385893793776631)),(to_sfixed_a(4.8119374696398154e-05)),(to_sfixed_a(-0.0037638144567608833)),(to_sfixed_a(0.0007440642802976072)),(to_sfixed_a(7.930635183583945e-05)),(to_sfixed_a(-0.0001817768206819892)),(to_sfixed_a(-0.0001542168902233243)),(to_sfixed_a(-0.27523675560951233)),(to_sfixed_a(-6.481191667262465e-05)),(to_sfixed_a(-0.001423144363798201)),(to_sfixed_a(1.884698576759547e-06)),(to_sfixed_a(0.0007881501223891973)),(to_sfixed_a(0.15419884026050568)),(to_sfixed_a(0.00012758831144310534)),(to_sfixed_a(0.00011540805280674249)),(to_sfixed_a(4.464600351639092e-06)),(to_sfixed_a(0.0001529828878119588)),(to_sfixed_a(0.001647208002395928)),(to_sfixed_a(5.1970797358080745e-05)),(to_sfixed_a(-4.953762982040644e-07)),(to_sfixed_a(0.28185415267944336)),(to_sfixed_a(-0.0051505351439118385)),(to_sfixed_a(2.2219204765860923e-05)),(to_sfixed_a(-0.0001687743642833084)),(to_sfixed_a(2.9768809326924384e-05)),(to_sfixed_a(-5.42117704753764e-05)),(to_sfixed_a(0.0011599051067605615)),(to_sfixed_a(0.001996654085814953)),(to_sfixed_a(3.78555414499715e-05)),(to_sfixed_a(0.00016466749366372824)),(to_sfixed_a(-1.189437898574397e-05)),(to_sfixed_a(-0.00010400912287877873)),(to_sfixed_a(0.17325200140476227)),(to_sfixed_a(0.0034806986805051565)),(to_sfixed_a(0.026237545534968376)),(to_sfixed_a(-0.00019161103409714997)),(to_sfixed_a(0.6268605589866638)),(to_sfixed_a(6.921536987647414e-05)),(to_sfixed_a(0.00019822298781946301)),(to_sfixed_a(-0.003984049428254366)),(to_sfixed_a(7.002470374573022e-05)),(to_sfixed_a(-0.00024095980916172266)),(to_sfixed_a(-0.0066518220119178295)),(to_sfixed_a(-0.0017039960948750377)),(to_sfixed_a(0.00019995718321297318)),(to_sfixed_a(5.104106094222516e-06)),(to_sfixed_a(-0.0002613175311125815)),(to_sfixed_a(-7.30697502149269e-05)),(to_sfixed_a(-7.165219722082838e-05)),(to_sfixed_a(-0.0011827501002699137)),(to_sfixed_a(-0.04250284284353256)),(to_sfixed_a(0.0002088354085572064)),(to_sfixed_a(-4.38901552115567e-05)),(to_sfixed_a(-0.005414028186351061)),(to_sfixed_a(0.00036287124385125935)),(to_sfixed_a(-0.0001058978377841413)),(to_sfixed_a(-7.985523552633822e-06)),(to_sfixed_a(0.01580602116882801)),(to_sfixed_a(-0.0002177520509576425)),(to_sfixed_a(1.93131563719362e-06)),(to_sfixed_a(2.435628994135186e-05)),(to_sfixed_a(0.21598728001117706)),(to_sfixed_a(-5.747294926550239e-05)),(to_sfixed_a(0.18102847039699554)),(to_sfixed_a(0.0001883282675407827)),(to_sfixed_a(0.0001758198777679354)),(to_sfixed_a(0.00451328931376338)),(to_sfixed_a(-0.00016524732927791774)),(to_sfixed_a(6.150254921521991e-05)),(to_sfixed_a(-9.838808909989893e-05)),(to_sfixed_a(-6.664796819677576e-05)),(to_sfixed_a(-0.00010287044278811663)),(to_sfixed_a(0.0031021786853671074)),(to_sfixed_a(6.805811426602304e-05)),(to_sfixed_a(-0.0009808341274037957)),(to_sfixed_a(0.23368202149868011)),(to_sfixed_a(-0.000124762489576824)),(to_sfixed_a(0.0001996686332859099)),(to_sfixed_a(0.00023008060816209763)),(to_sfixed_a(-0.009439797140657902)),(to_sfixed_a(-0.0008358171908184886)),(to_sfixed_a(0.0018806305015459657)),(to_sfixed_a(0.2110069990158081)),(to_sfixed_a(0.00010991178714903072)),(to_sfixed_a(-0.2603316009044647)),(to_sfixed_a(0.00014861844829283655)),(to_sfixed_a(-6.33889067103155e-05)),(to_sfixed_a(0.41930511593818665)),(to_sfixed_a(0.00011981265561189502)),(to_sfixed_a(-0.013337102718651295)),(to_sfixed_a(6.120491889305413e-05)),(to_sfixed_a(0.022704247385263443)),(to_sfixed_a(-0.014398206025362015)),(to_sfixed_a(0.3107595443725586)),(to_sfixed_a(0.0014156292891129851)),(to_sfixed_a(-0.02081771194934845)),(to_sfixed_a(-0.6660894155502319)),(to_sfixed_a(-0.0011076590744778514)),(to_sfixed_a(-0.003907420206815004)),(to_sfixed_a(-3.604764424380846e-05)),(to_sfixed_a(-0.0001521637022960931)),(to_sfixed_a(0.0001495939795859158)),(to_sfixed_a(-8.58712701301556e-06)),(to_sfixed_a(-0.009238491766154766)),(to_sfixed_a(-0.0015796700026839972)),(to_sfixed_a(0.0013238933170214295)),(to_sfixed_a(-0.00014509219909086823)),(to_sfixed_a(0.00658858846873045)),(to_sfixed_a(9.570501424605027e-05)),(to_sfixed_a(0.3423340320587158)),(to_sfixed_a(-0.4560575783252716)),(to_sfixed_a(0.0002658785379026085)),(to_sfixed_a(-0.0038164122961461544)),(to_sfixed_a(-0.0001400239416398108)),(to_sfixed_a(-0.18483079969882965)),(to_sfixed_a(0.0005615099216811359)),(to_sfixed_a(3.621713403845206e-05)),(to_sfixed_a(5.367901030695066e-05)),(to_sfixed_a(7.118899520719424e-05)),(to_sfixed_a(-0.00014709567767567933)),(to_sfixed_a(0.00013887429668102413)),(to_sfixed_a(-7.940776413306594e-06)),(to_sfixed_a(0.18856078386306763)),(to_sfixed_a(0.0037761053536087275)),(to_sfixed_a(0.13790838420391083)),(to_sfixed_a(0.0035529157612472773)),(to_sfixed_a(-0.2296907752752304)),(to_sfixed_a(0.005408419296145439)),(to_sfixed_a(7.296837429748848e-05)),(to_sfixed_a(0.0001564731210237369)),(to_sfixed_a(6.32711744401604e-05)),(to_sfixed_a(0.00016696358215995133)),(to_sfixed_a(-9.774507634574547e-05)),(to_sfixed_a(0.0024705331306904554)),(to_sfixed_a(-0.0001730779476929456)),(to_sfixed_a(0.0012596654705703259)),(to_sfixed_a(3.510088208713569e-05)),(to_sfixed_a(3.1052040867507458e-06)),(to_sfixed_a(0.00013372446119319648)),(to_sfixed_a(3.901234595105052e-05)),(to_sfixed_a(-0.00024826612207107246)),(to_sfixed_a(-0.002623752923682332)),(to_sfixed_a(-6.52250018902123e-05)),(to_sfixed_a(4.099641955690458e-06)),(to_sfixed_a(-0.000178378468262963)),(to_sfixed_a(0.00023399016936309636)),(to_sfixed_a(0.0908854752779007)),(to_sfixed_a(-0.7702196836471558)),(to_sfixed_a(5.812477320432663e-05)),(to_sfixed_a(0.0001513844617875293)),(to_sfixed_a(2.4745273549342528e-05)),(to_sfixed_a(4.67325808131136e-05)),(to_sfixed_a(0.366769939661026)),(to_sfixed_a(-0.022766083478927612)),(to_sfixed_a(0.00010718392150010914)),(to_sfixed_a(-6.870373908895999e-05)),(to_sfixed_a(0.00013345896149985492)),(to_sfixed_a(-0.0003451109805610031)),(to_sfixed_a(0.00015081383753567934)),(to_sfixed_a(0.3267803192138672)),(to_sfixed_a(-6.279542139964178e-05)),(to_sfixed_a(0.4808956980705261)),(to_sfixed_a(0.005484503693878651)),(to_sfixed_a(-0.04060407355427742)),(to_sfixed_a(-0.005744162946939468)),(to_sfixed_a(-0.00010849709360627457)),(to_sfixed_a(0.0021690567955374718)),(to_sfixed_a(-0.0001117758802138269)),(to_sfixed_a(-1.4831923181191087e-05)),(to_sfixed_a(-0.004980935715138912)),(to_sfixed_a(9.671039879322052e-05)),(to_sfixed_a(-6.14841264905408e-05)),(to_sfixed_a(0.5557140707969666)),(to_sfixed_a(0.37377190589904785)),(to_sfixed_a(2.0231527741998434e-06)),(to_sfixed_a(-0.00010320852743461728)),(to_sfixed_a(-0.01015950832515955)),(to_sfixed_a(0.0001533480390207842)),(to_sfixed_a(0.6797201633453369)),(to_sfixed_a(-0.00018862583965528756)),(to_sfixed_a(-0.0004579908272717148)),(to_sfixed_a(6.0579623095691204e-05)),(to_sfixed_a(-0.010127020999789238)),(to_sfixed_a(-0.00017953835777007043)),(to_sfixed_a(-3.384106094017625e-06)),(to_sfixed_a(-0.0002046094450633973)),(to_sfixed_a(-0.0022861019242554903)),(to_sfixed_a(-0.003011049935594201)),(to_sfixed_a(0.00019827061623800546)),(to_sfixed_a(3.804649168159813e-05)),(to_sfixed_a(-7.423843635478988e-05)),(to_sfixed_a(1.591173349879682e-05)),(to_sfixed_a(0.002125590108335018)),(to_sfixed_a(-0.009773463010787964)),(to_sfixed_a(0.003194741904735565)),(to_sfixed_a(-0.0016426639631390572)),(to_sfixed_a(-0.38949859142303467)),(to_sfixed_a(-0.00014896919310558587)),(to_sfixed_a(-0.0002250557445222512)),(to_sfixed_a(7.737611304037273e-05)),(to_sfixed_a(0.009251507930457592)),(to_sfixed_a(-6.056488928152248e-05)),(to_sfixed_a(-9.005255560623482e-05)),(to_sfixed_a(0.0038946366403251886)),(to_sfixed_a(-0.007013358175754547)),(to_sfixed_a(5.954105290584266e-06)),(to_sfixed_a(-0.4717573821544647)),(to_sfixed_a(0.0025254094507545233)),(to_sfixed_a(-0.000665551982820034)),(to_sfixed_a(-0.1387626677751541)),(to_sfixed_a(-0.00013900891644880176)),(to_sfixed_a(-0.0021320683881640434)),(to_sfixed_a(-0.015232497826218605)),(to_sfixed_a(-0.003953700419515371)),(to_sfixed_a(-0.000135012945975177)),(to_sfixed_a(0.0038563301786780357)),(to_sfixed_a(0.004321754910051823)),(to_sfixed_a(0.1224716305732727)));

    constant weight_n2_30 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.07320483028888702)),(to_sfixed_a(0.006029918789863586)),(to_sfixed_a(-0.0009704566327854991)),(to_sfixed_a(4.421756602823734e-05)),(to_sfixed_a(-0.174605131149292)),(to_sfixed_a(-6.098760786699131e-05)),(to_sfixed_a(-0.0006044055917300284)),(to_sfixed_a(-0.00038792198756709695)),(to_sfixed_a(-0.00010295714309904724)),(to_sfixed_a(-3.836453834082931e-05)),(to_sfixed_a(-0.0001669071934884414)),(to_sfixed_a(0.2297046035528183)),(to_sfixed_a(-0.47582030296325684)),(to_sfixed_a(-0.0013120385119691491)),(to_sfixed_a(0.00030973294633440673)),(to_sfixed_a(-3.1571944418828934e-05)),(to_sfixed_a(0.19603686034679413)),(to_sfixed_a(-9.52133268583566e-05)),(to_sfixed_a(0.0636497214436531)),(to_sfixed_a(-0.0026755090802907944)),(to_sfixed_a(0.00024661130737513304)),(to_sfixed_a(-0.00011027353320969269)),(to_sfixed_a(-0.0008213223773054779)),(to_sfixed_a(-0.001953410217538476)),(to_sfixed_a(-0.00030440607224591076)),(to_sfixed_a(-0.0011198464781045914)),(to_sfixed_a(-0.00017223358736373484)),(to_sfixed_a(4.3256084609311074e-05)),(to_sfixed_a(5.338156915968284e-05)),(to_sfixed_a(-3.7520163459703326e-05)),(to_sfixed_a(-0.005011881235986948)),(to_sfixed_a(1.1478095984784886e-05)),(to_sfixed_a(0.007561102043837309)),(to_sfixed_a(1.2300930393394083e-05)),(to_sfixed_a(-4.4202741264598444e-05)),(to_sfixed_a(0.00018066956545226276)),(to_sfixed_a(0.2045067846775055)),(to_sfixed_a(-0.38453495502471924)),(to_sfixed_a(-0.6933136582374573)),(to_sfixed_a(-0.00015685221296735108)),(to_sfixed_a(-0.5118781328201294)),(to_sfixed_a(-0.003243028186261654)),(to_sfixed_a(-5.7273617130704224e-05)),(to_sfixed_a(0.00011233296390855685)),(to_sfixed_a(0.001990492455661297)),(to_sfixed_a(2.658621087903157e-05)),(to_sfixed_a(-0.0012357421219348907)),(to_sfixed_a(-0.002509782323613763)),(to_sfixed_a(4.7116787754930556e-05)),(to_sfixed_a(0.000262997840764001)),(to_sfixed_a(-0.00462116627022624)),(to_sfixed_a(-0.0004264452727511525)),(to_sfixed_a(-4.31091248174198e-05)),(to_sfixed_a(-0.010353079065680504)),(to_sfixed_a(-0.044229257851839066)),(to_sfixed_a(0.024445489048957825)),(to_sfixed_a(-1.0337938874727115e-05)),(to_sfixed_a(-0.00993480533361435)),(to_sfixed_a(3.299624950159341e-06)),(to_sfixed_a(3.799409023486078e-05)),(to_sfixed_a(-0.0013402047334238887)),(to_sfixed_a(-0.0020097449887543917)),(to_sfixed_a(0.00015943658945616335)),(to_sfixed_a(0.004228521604090929)),(to_sfixed_a(-2.8475915314629674e-07)),(to_sfixed_a(0.4445156753063202)),(to_sfixed_a(0.0001733474782668054)),(to_sfixed_a(-0.13339334726333618)),(to_sfixed_a(-2.7722877348423935e-05)),(to_sfixed_a(-8.149698260240257e-06)),(to_sfixed_a(-0.0007529286085627973)),(to_sfixed_a(-0.0006350260809995234)),(to_sfixed_a(0.045683424919843674)),(to_sfixed_a(0.00018068037752527744)),(to_sfixed_a(-0.0001803779450710863)),(to_sfixed_a(1.0193358320975676e-05)),(to_sfixed_a(0.44223839044570923)),(to_sfixed_a(-0.00041438336484134197)),(to_sfixed_a(-1.0777650459203869e-05)),(to_sfixed_a(-0.6167783737182617)),(to_sfixed_a(4.983419057680294e-05)),(to_sfixed_a(0.0004182170087005943)),(to_sfixed_a(-0.011034694500267506)),(to_sfixed_a(0.3066003620624542)),(to_sfixed_a(-0.00011281004117336124)),(to_sfixed_a(0.00024676183238625526)),(to_sfixed_a(-0.24143637716770172)),(to_sfixed_a(1.0037429092335515e-06)),(to_sfixed_a(6.573151040356606e-05)),(to_sfixed_a(-0.00016867261729203165)),(to_sfixed_a(-0.01756972447037697)),(to_sfixed_a(-1.7883634427562356e-05)),(to_sfixed_a(-0.0001277058618143201)),(to_sfixed_a(-0.00020132283680140972)),(to_sfixed_a(0.017079241573810577)),(to_sfixed_a(6.471942469943315e-05)),(to_sfixed_a(6.28259003860876e-05)),(to_sfixed_a(2.3815679014660418e-05)),(to_sfixed_a(-6.740115350112319e-05)),(to_sfixed_a(-0.0001476798643125221)),(to_sfixed_a(-0.002530294004827738)),(to_sfixed_a(-0.000139990181196481)),(to_sfixed_a(-2.9356218874454498e-05)),(to_sfixed_a(0.27095869183540344)),(to_sfixed_a(0.0033515288960188627)),(to_sfixed_a(2.7871727070305496e-05)),(to_sfixed_a(-0.0001878630428109318)),(to_sfixed_a(6.730911991326138e-06)),(to_sfixed_a(5.7313394790980965e-05)),(to_sfixed_a(-0.019741499796509743)),(to_sfixed_a(-0.02667245827615261)),(to_sfixed_a(-7.157709478633478e-05)),(to_sfixed_a(0.01734348013997078)),(to_sfixed_a(6.918743019923568e-05)),(to_sfixed_a(-0.00013693617074750364)),(to_sfixed_a(-0.0051818471401929855)),(to_sfixed_a(0.0025101418141275644)),(to_sfixed_a(0.00014810884022153914)),(to_sfixed_a(2.5546964025124907e-05)),(to_sfixed_a(-0.026832837611436844)),(to_sfixed_a(-0.00015153930871747434)),(to_sfixed_a(-7.937354530440643e-05)),(to_sfixed_a(-0.0005195480771362782)),(to_sfixed_a(-1.4013327017892152e-05)),(to_sfixed_a(3.03072010865435e-06)),(to_sfixed_a(0.2627924382686615)),(to_sfixed_a(-3.719739106600173e-05)),(to_sfixed_a(-7.122381794033572e-05)),(to_sfixed_a(-1.4145407476462424e-05)),(to_sfixed_a(0.00015136264846660197)),(to_sfixed_a(-3.083056435571052e-05)),(to_sfixed_a(-1.0702686267904937e-05)),(to_sfixed_a(-0.0003894797118846327)),(to_sfixed_a(0.10489556938409805)),(to_sfixed_a(0.00010531723091844469)),(to_sfixed_a(-4.3368127080611885e-05)),(to_sfixed_a(-0.40828263759613037)),(to_sfixed_a(6.331024633254856e-05)),(to_sfixed_a(-9.357725502923131e-06)),(to_sfixed_a(0.00010266176832374185)),(to_sfixed_a(4.619437822839245e-05)),(to_sfixed_a(-1.2326643627602607e-05)),(to_sfixed_a(6.707786815240979e-05)),(to_sfixed_a(-1.686339601292275e-07)),(to_sfixed_a(-0.000265526759903878)),(to_sfixed_a(2.1322797692846507e-05)),(to_sfixed_a(-0.000401013734517619)),(to_sfixed_a(-1.0872216080315411e-05)),(to_sfixed_a(-0.0002995422692038119)),(to_sfixed_a(-0.00048647611401975155)),(to_sfixed_a(-0.00014520081458613276)),(to_sfixed_a(-4.1284627513960004e-05)),(to_sfixed_a(0.001122002024203539)),(to_sfixed_a(4.7079061914701015e-05)),(to_sfixed_a(-0.00017623029998503625)),(to_sfixed_a(-0.0052285450510680676)),(to_sfixed_a(4.269153578206897e-06)),(to_sfixed_a(-0.29416024684906006)),(to_sfixed_a(-8.009666635189205e-05)),(to_sfixed_a(-2.881964792322833e-05)),(to_sfixed_a(-3.8381247577490285e-05)),(to_sfixed_a(1.2951801181770861e-05)),(to_sfixed_a(-0.5633900165557861)),(to_sfixed_a(-0.016334032639861107)),(to_sfixed_a(-0.323839396238327)),(to_sfixed_a(0.003948770463466644)),(to_sfixed_a(0.00015198549954220653)),(to_sfixed_a(-0.5674560070037842)),(to_sfixed_a(-0.00018340516544412822)),(to_sfixed_a(-2.68472358584404e-05)),(to_sfixed_a(-0.027771512046456337)),(to_sfixed_a(0.0035845492966473103)),(to_sfixed_a(3.345404547872022e-05)),(to_sfixed_a(0.00018216072930954397)),(to_sfixed_a(0.004203916992992163)),(to_sfixed_a(3.6348683352116495e-06)),(to_sfixed_a(-0.005443713627755642)),(to_sfixed_a(-4.8603658797219396e-05)),(to_sfixed_a(0.009135918691754341)),(to_sfixed_a(0.21143941581249237)),(to_sfixed_a(-0.0010681692510843277)),(to_sfixed_a(-0.001228333916515112)),(to_sfixed_a(2.557138941483572e-05)),(to_sfixed_a(6.794861110392958e-05)),(to_sfixed_a(0.00013495341408997774)),(to_sfixed_a(-0.000712691224180162)),(to_sfixed_a(0.00759460311383009)),(to_sfixed_a(0.024264751002192497)),(to_sfixed_a(-0.0005986898904666305)),(to_sfixed_a(-0.00032565355650149286)),(to_sfixed_a(-1.7007318092510104e-05)),(to_sfixed_a(0.0002498044050298631)),(to_sfixed_a(-0.5985386967658997)),(to_sfixed_a(0.00022048423124942929)),(to_sfixed_a(-2.347279223613441e-05)),(to_sfixed_a(0.0898100882768631)),(to_sfixed_a(-6.634873716393486e-05)),(to_sfixed_a(0.0028589542489498854)),(to_sfixed_a(-0.002984865102916956)),(to_sfixed_a(-3.3022079151123762e-06)),(to_sfixed_a(5.785336543340236e-05)),(to_sfixed_a(4.018966865260154e-05)),(to_sfixed_a(0.0003113221318926662)),(to_sfixed_a(1.0393798220320605e-05)),(to_sfixed_a(-3.1803938327357173e-06)),(to_sfixed_a(-0.000472064595669508)),(to_sfixed_a(0.32071736454963684)),(to_sfixed_a(-0.15412865579128265)),(to_sfixed_a(-0.0032095680944621563)),(to_sfixed_a(-0.0009389867773279548)),(to_sfixed_a(-0.4805132746696472)),(to_sfixed_a(-8.109920599963516e-05)),(to_sfixed_a(7.132803148124367e-06)),(to_sfixed_a(6.246802513487637e-05)),(to_sfixed_a(-0.00013095322356093675)),(to_sfixed_a(-3.6798031942453235e-05)),(to_sfixed_a(6.966438377276063e-06)),(to_sfixed_a(0.0003980615292675793)),(to_sfixed_a(-0.3676552176475525)),(to_sfixed_a(0.00015410708147101104)),(to_sfixed_a(0.00038100036908872426)),(to_sfixed_a(8.485320722684264e-05)),(to_sfixed_a(-0.00010725420725066215)),(to_sfixed_a(0.2864137887954712)),(to_sfixed_a(0.5522801280021667)),(to_sfixed_a(6.175486487336457e-05)),(to_sfixed_a(7.086216646712273e-05)),(to_sfixed_a(-5.703445276594721e-05)),(to_sfixed_a(0.5377973318099976)),(to_sfixed_a(-0.007321212440729141)),(to_sfixed_a(0.02177293598651886)),(to_sfixed_a(0.0002395782939856872)),(to_sfixed_a(-0.0003122266207356006)),(to_sfixed_a(-5.556947144214064e-06)),(to_sfixed_a(4.643336797016673e-05)),(to_sfixed_a(0.004051883239299059)),(to_sfixed_a(-0.48295173048973083)),(to_sfixed_a(0.00016922972281463444)),(to_sfixed_a(-8.246539800893515e-05)),(to_sfixed_a(-4.408171298564412e-05)),(to_sfixed_a(-0.00013623059203382581)),(to_sfixed_a(-0.0003800565027631819)),(to_sfixed_a(-0.0016950223362073302)),(to_sfixed_a(6.73429312882945e-05)),(to_sfixed_a(-0.005220444407314062)),(to_sfixed_a(-0.4956059753894806)),(to_sfixed_a(0.00835002027451992)),(to_sfixed_a(-0.30095037817955017)),(to_sfixed_a(-0.00011367993283784017)),(to_sfixed_a(0.01829151250422001)),(to_sfixed_a(0.0003234410542063415)),(to_sfixed_a(0.00017483085684943944)),(to_sfixed_a(0.00032472569728270173)),(to_sfixed_a(0.000289984600385651)),(to_sfixed_a(0.0015739744994789362)),(to_sfixed_a(-0.7267874479293823)),(to_sfixed_a(-0.0024528794456273317)),(to_sfixed_a(-4.529741272563115e-05)),(to_sfixed_a(5.733288708142936e-05)),(to_sfixed_a(-0.0033928523771464825)),(to_sfixed_a(-0.00012692628661170602)),(to_sfixed_a(-0.0021326406858861446)),(to_sfixed_a(-4.334681580075994e-05)),(to_sfixed_a(-0.0013570962473750114)),(to_sfixed_a(-0.00021197502792347223)),(to_sfixed_a(-0.008171251974999905)),(to_sfixed_a(2.3878237698227167e-06)),(to_sfixed_a(-1.7373196897096932e-05)),(to_sfixed_a(0.0001918467169161886)),(to_sfixed_a(0.007510661613196135)),(to_sfixed_a(-0.023194564506411552)),(to_sfixed_a(0.00010101807856699452)),(to_sfixed_a(-2.082498394884169e-05)),(to_sfixed_a(-6.930299423402175e-05)),(to_sfixed_a(2.372993913013488e-05)),(to_sfixed_a(0.004594911355525255)),(to_sfixed_a(-0.34350770711898804)),(to_sfixed_a(-0.3278695046901703)),(to_sfixed_a(0.0018829815089702606)),(to_sfixed_a(0.03820609673857689)),(to_sfixed_a(6.067328286007978e-05)),(to_sfixed_a(0.00025224487762898207)),(to_sfixed_a(1.6128920833580196e-05)),(to_sfixed_a(-0.001023103715851903)),(to_sfixed_a(-5.019173113396391e-05)),(to_sfixed_a(-0.00011305423686280847)),(to_sfixed_a(-0.0001556935312692076)),(to_sfixed_a(0.0005017957300879061)),(to_sfixed_a(-7.300503784790635e-05)),(to_sfixed_a(0.0036594269331544638)),(to_sfixed_a(-0.0005074344808235765)),(to_sfixed_a(0.0012104535708203912)),(to_sfixed_a(0.18222440779209137)),(to_sfixed_a(5.6956312619149685e-05)),(to_sfixed_a(0.3246150314807892)),(to_sfixed_a(-0.3417186737060547)),(to_sfixed_a(-0.0010961152147501707)),(to_sfixed_a(-0.00011403484677430242)),(to_sfixed_a(-0.15987354516983032)),(to_sfixed_a(0.07631361484527588)),(to_sfixed_a(-0.3737998902797699)));

    constant weight_n2_31 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.1681174337863922)),(to_sfixed_a(0.41477760672569275)),(to_sfixed_a(0.5252810120582581)),(to_sfixed_a(2.696242881938815e-05)),(to_sfixed_a(0.004831918515264988)),(to_sfixed_a(0.00021147506777197123)),(to_sfixed_a(-0.0008760052733123302)),(to_sfixed_a(-1.467180481995456e-05)),(to_sfixed_a(7.088048732839525e-06)),(to_sfixed_a(-0.00014963740250095725)),(to_sfixed_a(5.9311019867891446e-05)),(to_sfixed_a(-0.005852707661688328)),(to_sfixed_a(0.012339489534497261)),(to_sfixed_a(0.00591582665219903)),(to_sfixed_a(1.853401045082137e-05)),(to_sfixed_a(0.00038095322088338435)),(to_sfixed_a(0.018356282263994217)),(to_sfixed_a(-0.00020973689970560372)),(to_sfixed_a(-0.00016950786812230945)),(to_sfixed_a(-0.5341242551803589)),(to_sfixed_a(-0.00029193039517849684)),(to_sfixed_a(-0.00011211341916350648)),(to_sfixed_a(9.064878395292908e-05)),(to_sfixed_a(0.2220507264137268)),(to_sfixed_a(-0.0009334611822851002)),(to_sfixed_a(0.002231159945949912)),(to_sfixed_a(0.0001526323612779379)),(to_sfixed_a(-0.000825042836368084)),(to_sfixed_a(0.011030150577425957)),(to_sfixed_a(0.00016894290456548333)),(to_sfixed_a(0.011989319697022438)),(to_sfixed_a(2.243810740765184e-05)),(to_sfixed_a(-0.006559593603014946)),(to_sfixed_a(-7.075469329720363e-05)),(to_sfixed_a(0.00010057584586320445)),(to_sfixed_a(0.0001123273468692787)),(to_sfixed_a(0.0034596475306898355)),(to_sfixed_a(0.49102330207824707)),(to_sfixed_a(0.007775787729769945)),(to_sfixed_a(0.0001207280729431659)),(to_sfixed_a(0.010237431153655052)),(to_sfixed_a(0.46631571650505066)),(to_sfixed_a(-4.375940261525102e-05)),(to_sfixed_a(5.512172356247902e-05)),(to_sfixed_a(0.013440595008432865)),(to_sfixed_a(0.017307449132204056)),(to_sfixed_a(0.03647415712475777)),(to_sfixed_a(0.016650324687361717)),(to_sfixed_a(9.870190115179867e-05)),(to_sfixed_a(0.03459538519382477)),(to_sfixed_a(0.0011586463078856468)),(to_sfixed_a(-0.0008796277106739581)),(to_sfixed_a(0.00016808474902063608)),(to_sfixed_a(-0.000788794772233814)),(to_sfixed_a(-0.02219865284860134)),(to_sfixed_a(-0.3739585280418396)),(to_sfixed_a(-6.791104533476755e-05)),(to_sfixed_a(0.002951292088255286)),(to_sfixed_a(0.00018355276552028954)),(to_sfixed_a(-3.3789052395150065e-05)),(to_sfixed_a(0.004787816666066647)),(to_sfixed_a(-0.00016291523934341967)),(to_sfixed_a(0.001562034711241722)),(to_sfixed_a(0.016820615157485008)),(to_sfixed_a(9.912633686326444e-06)),(to_sfixed_a(-0.7160270810127258)),(to_sfixed_a(-3.764063512790017e-05)),(to_sfixed_a(0.0032290169037878513)),(to_sfixed_a(-0.0009403703734278679)),(to_sfixed_a(8.295826410176232e-05)),(to_sfixed_a(-0.17305321991443634)),(to_sfixed_a(0.0007297557312995195)),(to_sfixed_a(0.005854979157447815)),(to_sfixed_a(-1.886558675323613e-05)),(to_sfixed_a(5.054011126048863e-06)),(to_sfixed_a(-9.220873835147358e-06)),(to_sfixed_a(-0.01150980219244957)),(to_sfixed_a(-7.92648279457353e-05)),(to_sfixed_a(1.5521174645982683e-05)),(to_sfixed_a(0.5377054214477539)),(to_sfixed_a(0.003888548817485571)),(to_sfixed_a(-6.980515900067985e-05)),(to_sfixed_a(0.36590108275413513)),(to_sfixed_a(-0.22551138699054718)),(to_sfixed_a(8.55181206134148e-05)),(to_sfixed_a(0.0013342465972527862)),(to_sfixed_a(-0.3456294536590576)),(to_sfixed_a(5.630700252368115e-05)),(to_sfixed_a(-3.804429798037745e-05)),(to_sfixed_a(0.00023906436399556696)),(to_sfixed_a(-0.22646398842334747)),(to_sfixed_a(-0.00024537547142244875)),(to_sfixed_a(0.0052382745780050755)),(to_sfixed_a(-0.00029538743547163904)),(to_sfixed_a(0.009147089906036854)),(to_sfixed_a(6.378830585163087e-05)),(to_sfixed_a(-1.8536644347477704e-05)),(to_sfixed_a(-0.0003815614036284387)),(to_sfixed_a(9.209084964822978e-05)),(to_sfixed_a(-1.8691520381253213e-05)),(to_sfixed_a(0.0017635038821026683)),(to_sfixed_a(-0.00024882768047973514)),(to_sfixed_a(0.00023666514607612044)),(to_sfixed_a(0.0029620984569191933)),(to_sfixed_a(0.01655511185526848)),(to_sfixed_a(-4.894263838650659e-05)),(to_sfixed_a(-0.00015934236580505967)),(to_sfixed_a(4.977900243829936e-05)),(to_sfixed_a(-5.7767647376749665e-06)),(to_sfixed_a(-0.0022245359141379595)),(to_sfixed_a(0.023848816752433777)),(to_sfixed_a(6.630385905737057e-05)),(to_sfixed_a(0.11656289547681808)),(to_sfixed_a(3.893699613399804e-06)),(to_sfixed_a(6.615927850361913e-05)),(to_sfixed_a(-0.003794665914028883)),(to_sfixed_a(-0.00021674924937542528)),(to_sfixed_a(-0.00048009908641688526)),(to_sfixed_a(-1.638346293475479e-05)),(to_sfixed_a(0.009860806167125702)),(to_sfixed_a(-1.8925857148133218e-06)),(to_sfixed_a(1.4633216778747737e-05)),(to_sfixed_a(0.007345704361796379)),(to_sfixed_a(-4.944314787280746e-05)),(to_sfixed_a(0.00018916703993454576)),(to_sfixed_a(-0.2999378442764282)),(to_sfixed_a(0.45833441615104675)),(to_sfixed_a(7.026840467005968e-05)),(to_sfixed_a(0.0002727775718085468)),(to_sfixed_a(3.728306182892993e-05)),(to_sfixed_a(4.3100335460621864e-05)),(to_sfixed_a(-5.264382343739271e-05)),(to_sfixed_a(0.00017866308917291462)),(to_sfixed_a(0.04668104276061058)),(to_sfixed_a(7.885818922659382e-05)),(to_sfixed_a(-1.179121682071127e-05)),(to_sfixed_a(0.014140674844384193)),(to_sfixed_a(-0.00017681173630990088)),(to_sfixed_a(-6.75030896672979e-05)),(to_sfixed_a(6.543096242239699e-05)),(to_sfixed_a(0.000296791666187346)),(to_sfixed_a(0.0001053128216881305)),(to_sfixed_a(-0.0002023745037149638)),(to_sfixed_a(2.3755841539241374e-05)),(to_sfixed_a(-0.0009211503784172237)),(to_sfixed_a(-0.0004300300788599998)),(to_sfixed_a(-0.0005955861415714025)),(to_sfixed_a(0.00015244573296513408)),(to_sfixed_a(-3.843141166726127e-05)),(to_sfixed_a(-0.0010121169034391642)),(to_sfixed_a(6.201244832482189e-05)),(to_sfixed_a(-7.103654934326187e-05)),(to_sfixed_a(0.13848581910133362)),(to_sfixed_a(-0.00019820773741230369)),(to_sfixed_a(-9.264094842365012e-05)),(to_sfixed_a(0.1967398226261139)),(to_sfixed_a(-1.228085602633655e-05)),(to_sfixed_a(-0.012390420772135258)),(to_sfixed_a(8.017208529054187e-06)),(to_sfixed_a(0.00010034658771473914)),(to_sfixed_a(-6.428142660297453e-05)),(to_sfixed_a(-4.258159606251866e-06)),(to_sfixed_a(0.003728081937879324)),(to_sfixed_a(-0.00014419946819543839)),(to_sfixed_a(-0.0026673756074160337)),(to_sfixed_a(0.003514355979859829)),(to_sfixed_a(-0.000244542898144573)),(to_sfixed_a(0.0012703753309324384)),(to_sfixed_a(3.4252225304953754e-06)),(to_sfixed_a(-2.8082124117645435e-05)),(to_sfixed_a(0.0017481989925727248)),(to_sfixed_a(-0.0007057514158077538)),(to_sfixed_a(0.00024553906405344605)),(to_sfixed_a(0.00017667346401140094)),(to_sfixed_a(0.0006789917824789882)),(to_sfixed_a(-3.0200069886632264e-05)),(to_sfixed_a(0.5525357127189636)),(to_sfixed_a(-0.004287682939320803)),(to_sfixed_a(-0.0005810746224597096)),(to_sfixed_a(-0.1251550167798996)),(to_sfixed_a(-1.2260832590982318e-05)),(to_sfixed_a(0.004690712317824364)),(to_sfixed_a(0.0002430592867312953)),(to_sfixed_a(2.7474728995002806e-05)),(to_sfixed_a(-8.163329039234668e-05)),(to_sfixed_a(0.0018674199236556888)),(to_sfixed_a(-0.20422925055027008)),(to_sfixed_a(0.004217867739498615)),(to_sfixed_a(9.293686889577657e-05)),(to_sfixed_a(0.001066490076482296)),(to_sfixed_a(0.005824333522468805)),(to_sfixed_a(1.0688512702472508e-05)),(to_sfixed_a(0.007409216836094856)),(to_sfixed_a(0.0053366306237876415)),(to_sfixed_a(-0.00012064458860550076)),(to_sfixed_a(0.011064887046813965)),(to_sfixed_a(4.1048406274057925e-07)),(to_sfixed_a(0.2855238914489746)),(to_sfixed_a(0.0029405183158814907)),(to_sfixed_a(-1.8686736439121887e-05)),(to_sfixed_a(-0.00016857493028510362)),(to_sfixed_a(-0.00015571212861686945)),(to_sfixed_a(0.00020141733693890274)),(to_sfixed_a(2.442896948195994e-05)),(to_sfixed_a(0.00012163615610916167)),(to_sfixed_a(-0.0026872812304645777)),(to_sfixed_a(0.3023281395435333)),(to_sfixed_a(0.028042789548635483)),(to_sfixed_a(0.00667995773255825)),(to_sfixed_a(-0.0008277160231955349)),(to_sfixed_a(-0.0016821443568915129)),(to_sfixed_a(0.00019582232926040888)),(to_sfixed_a(-0.0002999178832396865)),(to_sfixed_a(6.1440041463356465e-06)),(to_sfixed_a(6.907580973347649e-05)),(to_sfixed_a(0.0001821581245167181)),(to_sfixed_a(-0.011318551376461983)),(to_sfixed_a(0.000477376626804471)),(to_sfixed_a(-0.03663671761751175)),(to_sfixed_a(-4.432738933246583e-05)),(to_sfixed_a(-9.442200826015323e-05)),(to_sfixed_a(-3.0652692657895386e-05)),(to_sfixed_a(0.00023084350686986)),(to_sfixed_a(-0.00010574851330602542)),(to_sfixed_a(0.009791622869670391)),(to_sfixed_a(-0.0001569720625411719)),(to_sfixed_a(-0.000118804513476789)),(to_sfixed_a(3.631839717854746e-05)),(to_sfixed_a(0.00892963632941246)),(to_sfixed_a(-1.0273832231177948e-05)),(to_sfixed_a(-0.000728740356862545)),(to_sfixed_a(-4.2596297134878114e-05)),(to_sfixed_a(0.00013324720202945173)),(to_sfixed_a(-7.380698662018403e-05)),(to_sfixed_a(0.0013479964109137654)),(to_sfixed_a(-0.02020934969186783)),(to_sfixed_a(0.4328567087650299)),(to_sfixed_a(-8.700050238985568e-05)),(to_sfixed_a(0.002295475220307708)),(to_sfixed_a(0.00028240247047506273)),(to_sfixed_a(-0.004937156569212675)),(to_sfixed_a(5.901959229959175e-05)),(to_sfixed_a(2.329337803530507e-06)),(to_sfixed_a(-0.0001367777877021581)),(to_sfixed_a(-0.0022229626774787903)),(to_sfixed_a(-0.004020872991532087)),(to_sfixed_a(0.0003880648873746395)),(to_sfixed_a(0.09442649036645889)),(to_sfixed_a(0.00044788216473534703)),(to_sfixed_a(0.3265324532985687)),(to_sfixed_a(0.011523604393005371)),(to_sfixed_a(-0.00019077086471952498)),(to_sfixed_a(0.009211338125169277)),(to_sfixed_a(-7.307711348403245e-05)),(to_sfixed_a(0.24866139888763428)),(to_sfixed_a(0.5801444053649902)),(to_sfixed_a(0.0009217750048264861)),(to_sfixed_a(-5.6510354625061154e-05)),(to_sfixed_a(7.08117731846869e-05)),(to_sfixed_a(0.01566728763282299)),(to_sfixed_a(-0.00023779505863785744)),(to_sfixed_a(0.0004571815952658653)),(to_sfixed_a(-8.536810491932556e-05)),(to_sfixed_a(-0.2402481585741043)),(to_sfixed_a(4.418312892084941e-05)),(to_sfixed_a(0.006454689893871546)),(to_sfixed_a(7.351643580477685e-05)),(to_sfixed_a(-7.180465036071837e-05)),(to_sfixed_a(6.948700320208445e-05)),(to_sfixed_a(-0.15417487919330597)),(to_sfixed_a(0.29275715351104736)),(to_sfixed_a(-0.00018324691336601973)),(to_sfixed_a(0.00020252687681932002)),(to_sfixed_a(-0.00023713904374744743)),(to_sfixed_a(-8.226757927332073e-06)),(to_sfixed_a(0.7135456204414368)),(to_sfixed_a(0.01293040532618761)),(to_sfixed_a(-0.0020544833969324827)),(to_sfixed_a(0.004772009328007698)),(to_sfixed_a(0.0005270622204989195)),(to_sfixed_a(0.00014827953418716788)),(to_sfixed_a(6.276075873756781e-05)),(to_sfixed_a(0.00015984405763447285)),(to_sfixed_a(-0.4058627784252167)),(to_sfixed_a(-0.00018885673489421606)),(to_sfixed_a(0.00022366347548086196)),(to_sfixed_a(-0.0001638357643969357)),(to_sfixed_a(-0.2720576524734497)),(to_sfixed_a(0.00013221940025687218)),(to_sfixed_a(0.3590484857559204)),(to_sfixed_a(-0.0011708837701007724)),(to_sfixed_a(0.0012386735761538148)),(to_sfixed_a(-0.1351425051689148)),(to_sfixed_a(0.00014781983918510377)),(to_sfixed_a(-0.03118249773979187)),(to_sfixed_a(0.011784634552896023)),(to_sfixed_a(0.009093984961509705)),(to_sfixed_a(0.00010262746945954859)),(to_sfixed_a(-0.00749607989564538)),(to_sfixed_a(0.00785914808511734)),(to_sfixed_a(0.07750404626131058)));

    constant weight_n2_32 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.23386311531066895)),(to_sfixed_a(0.3468918800354004)),(to_sfixed_a(-0.0003919939626939595)),(to_sfixed_a(0.0002522245922591537)),(to_sfixed_a(-0.005148277152329683)),(to_sfixed_a(-0.0003085704520344734)),(to_sfixed_a(0.0006323991692624986)),(to_sfixed_a(-0.0003065630153287202)),(to_sfixed_a(-6.598696927540004e-05)),(to_sfixed_a(-3.6919256672263145e-05)),(to_sfixed_a(4.609508323483169e-06)),(to_sfixed_a(-0.0008401916129514575)),(to_sfixed_a(0.45405343174934387)),(to_sfixed_a(0.29745423793792725)),(to_sfixed_a(0.00010659120744094253)),(to_sfixed_a(0.00023651192896068096)),(to_sfixed_a(0.4532288908958435)),(to_sfixed_a(0.0002759587951004505)),(to_sfixed_a(0.1366972029209137)),(to_sfixed_a(-0.03812994062900543)),(to_sfixed_a(8.965635061031207e-07)),(to_sfixed_a(-7.168445881688967e-05)),(to_sfixed_a(0.0014463603729382157)),(to_sfixed_a(-0.005607669707387686)),(to_sfixed_a(-0.0009873607195913792)),(to_sfixed_a(0.0026740289758890867)),(to_sfixed_a(-0.00016684058937244117)),(to_sfixed_a(3.1659030355513096e-05)),(to_sfixed_a(-0.00030440124101005495)),(to_sfixed_a(0.00015189015539363027)),(to_sfixed_a(-0.0032843395601958036)),(to_sfixed_a(5.576985131483525e-05)),(to_sfixed_a(-0.001088741235435009)),(to_sfixed_a(0.00017632555682212114)),(to_sfixed_a(4.252942744642496e-07)),(to_sfixed_a(0.00041093461913987994)),(to_sfixed_a(-0.14739243686199188)),(to_sfixed_a(-0.00015071920643094927)),(to_sfixed_a(-0.007592829875648022)),(to_sfixed_a(-0.00017749394464772195)),(to_sfixed_a(-0.6298837661743164)),(to_sfixed_a(-0.0018045527394860983)),(to_sfixed_a(0.00011560214625205845)),(to_sfixed_a(2.7311187295708805e-05)),(to_sfixed_a(0.0001546718558529392)),(to_sfixed_a(0.00247454596683383)),(to_sfixed_a(-0.003958248533308506)),(to_sfixed_a(-0.005325545556843281)),(to_sfixed_a(0.00011836957128252834)),(to_sfixed_a(-0.0007883039652369916)),(to_sfixed_a(0.0024831576738506556)),(to_sfixed_a(-0.0020750691182911396)),(to_sfixed_a(-1.8681959772948176e-05)),(to_sfixed_a(0.00127803860232234)),(to_sfixed_a(-0.0008773371228016913)),(to_sfixed_a(-0.007975969463586807)),(to_sfixed_a(0.00011193923273822293)),(to_sfixed_a(0.00023999062250368297)),(to_sfixed_a(-0.00011755893501685932)),(to_sfixed_a(1.022260585159529e-05)),(to_sfixed_a(0.00034357435652054846)),(to_sfixed_a(0.003987031988799572)),(to_sfixed_a(-0.006787085440009832)),(to_sfixed_a(-0.3022192418575287)),(to_sfixed_a(-0.00021582678891718388)),(to_sfixed_a(0.1952333152294159)),(to_sfixed_a(0.00018207053653895855)),(to_sfixed_a(-0.009694140404462814)),(to_sfixed_a(9.197137842420489e-07)),(to_sfixed_a(5.917381349718198e-05)),(to_sfixed_a(-0.14980995655059814)),(to_sfixed_a(-0.14529313147068024)),(to_sfixed_a(0.004415587522089481)),(to_sfixed_a(0.00016834454436320812)),(to_sfixed_a(0.0002574794925749302)),(to_sfixed_a(-6.947244401089847e-05)),(to_sfixed_a(0.07918054610490799)),(to_sfixed_a(-0.4708138704299927)),(to_sfixed_a(-0.0001431844721082598)),(to_sfixed_a(0.3321264386177063)),(to_sfixed_a(-0.00032383567304350436)),(to_sfixed_a(-0.00018157088197767735)),(to_sfixed_a(-0.008877214044332504)),(to_sfixed_a(0.0007645590812899172)),(to_sfixed_a(0.00010674932127585635)),(to_sfixed_a(-0.0001913156738737598)),(to_sfixed_a(0.00029363343492150307)),(to_sfixed_a(0.0011560085695236921)),(to_sfixed_a(-7.626145088579506e-05)),(to_sfixed_a(8.606628398410976e-06)),(to_sfixed_a(-0.012881500646471977)),(to_sfixed_a(-8.666668145451695e-05)),(to_sfixed_a(-0.4384428858757019)),(to_sfixed_a(6.258487701416016e-06)),(to_sfixed_a(-0.005046462174504995)),(to_sfixed_a(3.3316911867586896e-05)),(to_sfixed_a(-0.00016839738236740232)),(to_sfixed_a(9.916852286551148e-05)),(to_sfixed_a(-7.165245187934488e-05)),(to_sfixed_a(2.2142503439681605e-05)),(to_sfixed_a(-0.4377104341983795)),(to_sfixed_a(0.002509712241590023)),(to_sfixed_a(0.00014686680515296757)),(to_sfixed_a(-0.45496925711631775)),(to_sfixed_a(0.010404680855572224)),(to_sfixed_a(0.002165726153180003)),(to_sfixed_a(4.988891305401921e-06)),(to_sfixed_a(-3.8552068872377276e-05)),(to_sfixed_a(0.0001336618443019688)),(to_sfixed_a(0.0005990889621898532)),(to_sfixed_a(-0.6957160234451294)),(to_sfixed_a(-0.0002369680441915989)),(to_sfixed_a(0.0017664388287812471)),(to_sfixed_a(-4.394122152007185e-05)),(to_sfixed_a(0.00017515290528535843)),(to_sfixed_a(-0.322132408618927)),(to_sfixed_a(0.00018219894263893366)),(to_sfixed_a(-6.441672303481027e-05)),(to_sfixed_a(9.507901268079877e-06)),(to_sfixed_a(-0.0005091309431008995)),(to_sfixed_a(-3.13405689666979e-05)),(to_sfixed_a(0.00027006235904991627)),(to_sfixed_a(-0.595757782459259)),(to_sfixed_a(0.00012315096682868898)),(to_sfixed_a(-0.00014655374980065972)),(to_sfixed_a(0.3702468276023865)),(to_sfixed_a(-0.49314793944358826)),(to_sfixed_a(2.587145718280226e-05)),(to_sfixed_a(-0.00018289378203917295)),(to_sfixed_a(0.00010629891767166555)),(to_sfixed_a(6.436595867853612e-05)),(to_sfixed_a(-1.8562714103609324e-05)),(to_sfixed_a(0.5367227792739868)),(to_sfixed_a(0.014671865850687027)),(to_sfixed_a(-0.0001481048675486818)),(to_sfixed_a(-0.0001894365414045751)),(to_sfixed_a(-0.00031018085428513587)),(to_sfixed_a(0.0009647745173424482)),(to_sfixed_a(-2.9921902751084417e-05)),(to_sfixed_a(6.170821870910004e-05)),(to_sfixed_a(0.00015459612768609077)),(to_sfixed_a(0.00011772345897043124)),(to_sfixed_a(-3.2072141038952395e-05)),(to_sfixed_a(-0.0021957603748887777)),(to_sfixed_a(0.0006701115053147078)),(to_sfixed_a(1.672439248068258e-05)),(to_sfixed_a(0.0013211109908297658)),(to_sfixed_a(-0.00014829530846327543)),(to_sfixed_a(0.00027038087137043476)),(to_sfixed_a(0.0067582158371806145)),(to_sfixed_a(-0.00015558894665446132)),(to_sfixed_a(-0.0002560263383202255)),(to_sfixed_a(1.5302728570532054e-05)),(to_sfixed_a(-0.00010040542838396505)),(to_sfixed_a(-0.0001160049723694101)),(to_sfixed_a(0.0034572866279631853)),(to_sfixed_a(-2.930426853708923e-05)),(to_sfixed_a(-0.13036595284938812)),(to_sfixed_a(-0.32934480905532837)),(to_sfixed_a(-2.405943814665079e-05)),(to_sfixed_a(0.00021558729349635541)),(to_sfixed_a(3.988319804193452e-06)),(to_sfixed_a(0.0021144093479961157)),(to_sfixed_a(0.0024825637228786945)),(to_sfixed_a(0.00120492500718683)),(to_sfixed_a(0.003055686829611659)),(to_sfixed_a(6.796953675802797e-05)),(to_sfixed_a(-0.009641841985285282)),(to_sfixed_a(0.0002138806157745421)),(to_sfixed_a(0.0003004720201715827)),(to_sfixed_a(-0.0013688317267224193)),(to_sfixed_a(0.00607643835246563)),(to_sfixed_a(0.0036570727825164795)),(to_sfixed_a(0.00023668981157243252)),(to_sfixed_a(-0.00295400433242321)),(to_sfixed_a(-0.00011887364235008135)),(to_sfixed_a(0.00019461293413769454)),(to_sfixed_a(0.0006851368816569448)),(to_sfixed_a(-0.00883458275347948)),(to_sfixed_a(-0.0256631001830101)),(to_sfixed_a(0.0011762462090700865)),(to_sfixed_a(0.013444291427731514)),(to_sfixed_a(1.8266777260578237e-05)),(to_sfixed_a(5.620549200102687e-05)),(to_sfixed_a(-0.0002053465141216293)),(to_sfixed_a(9.961629984900355e-06)),(to_sfixed_a(0.40039676427841187)),(to_sfixed_a(-0.007186823524534702)),(to_sfixed_a(0.00013862739433534443)),(to_sfixed_a(-0.0031641810201108456)),(to_sfixed_a(-0.0019330515060573816)),(to_sfixed_a(0.00022420057212002575)),(to_sfixed_a(-0.0001459653867641464)),(to_sfixed_a(-7.474219455616549e-05)),(to_sfixed_a(8.530114428140223e-06)),(to_sfixed_a(-0.0023167524486780167)),(to_sfixed_a(-0.00044750774395652115)),(to_sfixed_a(0.003495521377772093)),(to_sfixed_a(-0.00577166024595499)),(to_sfixed_a(0.0001738355786073953)),(to_sfixed_a(0.00020479533122852445)),(to_sfixed_a(-2.9972579795867205e-05)),(to_sfixed_a(-0.00013416912406682968)),(to_sfixed_a(-0.00015404818987008184)),(to_sfixed_a(6.244606629479676e-05)),(to_sfixed_a(0.00025319369160570204)),(to_sfixed_a(0.4023877680301666)),(to_sfixed_a(0.025197921320796013)),(to_sfixed_a(-0.0006947548245079815)),(to_sfixed_a(-0.0029077581129968166)),(to_sfixed_a(-0.0006292054313234985)),(to_sfixed_a(5.7277204177808017e-05)),(to_sfixed_a(-0.0001061654620571062)),(to_sfixed_a(-4.071521107107401e-05)),(to_sfixed_a(0.000199696805793792)),(to_sfixed_a(-3.221909355488606e-05)),(to_sfixed_a(-7.176924555096775e-05)),(to_sfixed_a(0.364998459815979)),(to_sfixed_a(-0.018263861536979675)),(to_sfixed_a(-2.2183081455295905e-05)),(to_sfixed_a(-4.4237625843379647e-05)),(to_sfixed_a(0.0002559049753472209)),(to_sfixed_a(0.0001349483645753935)),(to_sfixed_a(9.318994852947071e-05)),(to_sfixed_a(-2.433597546769306e-05)),(to_sfixed_a(-1.691468969511334e-05)),(to_sfixed_a(0.0002272286219522357)),(to_sfixed_a(-0.00014115909289103001)),(to_sfixed_a(0.08701600879430771)),(to_sfixed_a(0.00273543200455606)),(to_sfixed_a(0.003609149716794491)),(to_sfixed_a(0.00022069155238568783)),(to_sfixed_a(-9.740727546159178e-05)),(to_sfixed_a(-6.134863360784948e-05)),(to_sfixed_a(-0.0015755228232592344)),(to_sfixed_a(0.00010848480451386422)),(to_sfixed_a(-0.003939267247915268)),(to_sfixed_a(-0.00018507358618080616)),(to_sfixed_a(-0.0013735266402363777)),(to_sfixed_a(0.0001825487706810236)),(to_sfixed_a(-0.20649632811546326)),(to_sfixed_a(-8.531208004569635e-05)),(to_sfixed_a(-0.21139556169509888)),(to_sfixed_a(0.00024365526041947305)),(to_sfixed_a(-0.0029104610439389944)),(to_sfixed_a(0.0012350749457255006)),(to_sfixed_a(0.001238555763848126)),(to_sfixed_a(-0.3374927341938019)),(to_sfixed_a(2.4384702555835247e-05)),(to_sfixed_a(0.00039774959441274405)),(to_sfixed_a(9.679874892754015e-07)),(to_sfixed_a(5.284228245727718e-05)),(to_sfixed_a(-0.00040577491745352745)),(to_sfixed_a(5.447026342153549e-05)),(to_sfixed_a(-3.0382652767002583e-05)),(to_sfixed_a(-0.007897933945059776)),(to_sfixed_a(-0.004808157682418823)),(to_sfixed_a(-4.508328856900334e-06)),(to_sfixed_a(-0.0001982375542866066)),(to_sfixed_a(-0.013909033499658108)),(to_sfixed_a(-4.5872344344388694e-05)),(to_sfixed_a(0.0019709111656993628)),(to_sfixed_a(-3.36140365106985e-05)),(to_sfixed_a(-0.00010837026638910174)),(to_sfixed_a(0.0001394679129589349)),(to_sfixed_a(-0.00011980754061369225)),(to_sfixed_a(-0.00012892557424493134)),(to_sfixed_a(-0.000315165234496817)),(to_sfixed_a(-3.1367184419650584e-05)),(to_sfixed_a(0.005271403584629297)),(to_sfixed_a(-0.009751614183187485)),(to_sfixed_a(-0.0002676948788575828)),(to_sfixed_a(0.00015740242088213563)),(to_sfixed_a(6.952369585633278e-05)),(to_sfixed_a(-5.617829447146505e-05)),(to_sfixed_a(-0.00013206237053964287)),(to_sfixed_a(-0.008341233246028423)),(to_sfixed_a(0.003836100921034813)),(to_sfixed_a(0.2659883201122284)),(to_sfixed_a(0.00537278363481164)),(to_sfixed_a(-4.37939670518972e-05)),(to_sfixed_a(-0.0001583691337145865)),(to_sfixed_a(-0.00016469690308440477)),(to_sfixed_a(-1.246407555299811e-05)),(to_sfixed_a(0.0003926199278794229)),(to_sfixed_a(-4.377138247946277e-05)),(to_sfixed_a(-0.00022509763948619366)),(to_sfixed_a(-0.0037834623362869024)),(to_sfixed_a(-0.00011256287689320743)),(to_sfixed_a(-0.0008262177580036223)),(to_sfixed_a(-0.0002846182615030557)),(to_sfixed_a(0.005092712119221687)),(to_sfixed_a(-0.00012919158325530589)),(to_sfixed_a(-6.305626448011026e-05)),(to_sfixed_a(-0.015675637871026993)),(to_sfixed_a(0.5275757908821106)),(to_sfixed_a(0.0007508140988647938)),(to_sfixed_a(-0.00026742444606497884)),(to_sfixed_a(0.15962985157966614)),(to_sfixed_a(-0.08185356110334396)),(to_sfixed_a(-0.199735626578331)));

    constant weight_n2_33 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.007427520118653774)),(to_sfixed_a(0.00461966497823596)),(to_sfixed_a(0.019370580092072487)),(to_sfixed_a(1.9850582248182036e-05)),(to_sfixed_a(0.26179322600364685)),(to_sfixed_a(-2.3044049157761037e-05)),(to_sfixed_a(-0.00825275108218193)),(to_sfixed_a(-3.691941674333066e-05)),(to_sfixed_a(-0.00013991803280077875)),(to_sfixed_a(-0.00017749723338056356)),(to_sfixed_a(-0.000216468091821298)),(to_sfixed_a(0.015200330875813961)),(to_sfixed_a(-0.014930814504623413)),(to_sfixed_a(-0.007856893353164196)),(to_sfixed_a(-0.00010381735773989931)),(to_sfixed_a(0.00010717154509620741)),(to_sfixed_a(0.4735255837440491)),(to_sfixed_a(4.5222313929116353e-05)),(to_sfixed_a(0.08867008239030838)),(to_sfixed_a(-0.002646160777658224)),(to_sfixed_a(1.3106429832987487e-05)),(to_sfixed_a(0.00016794820840004832)),(to_sfixed_a(0.0003390230122022331)),(to_sfixed_a(0.001116513041779399)),(to_sfixed_a(0.003643761621788144)),(to_sfixed_a(0.4865841865539551)),(to_sfixed_a(4.561828973237425e-05)),(to_sfixed_a(-6.475287591456436e-06)),(to_sfixed_a(0.010673721320927143)),(to_sfixed_a(3.0629664252046496e-05)),(to_sfixed_a(-0.019642900675535202)),(to_sfixed_a(0.00024351227330043912)),(to_sfixed_a(-0.0006494002300314605)),(to_sfixed_a(0.00018018033006228507)),(to_sfixed_a(-0.00021565103088505566)),(to_sfixed_a(7.629711763001978e-05)),(to_sfixed_a(0.00337015138939023)),(to_sfixed_a(-0.0013152116443961859)),(to_sfixed_a(0.002527601784095168)),(to_sfixed_a(-6.475309783127159e-05)),(to_sfixed_a(0.0006088716327212751)),(to_sfixed_a(-0.008199858479201794)),(to_sfixed_a(0.00011694525892380625)),(to_sfixed_a(-5.534123920369893e-05)),(to_sfixed_a(0.007218693383038044)),(to_sfixed_a(0.024076346307992935)),(to_sfixed_a(-0.00017171836225315928)),(to_sfixed_a(-0.003076291410252452)),(to_sfixed_a(0.00044785719364881516)),(to_sfixed_a(-0.003065395401790738)),(to_sfixed_a(-0.0017341276397928596)),(to_sfixed_a(4.993783659301698e-05)),(to_sfixed_a(0.0001376405416522175)),(to_sfixed_a(-0.0014231287641450763)),(to_sfixed_a(-0.00405400525778532)),(to_sfixed_a(0.0019509999547153711)),(to_sfixed_a(0.00015453266678377986)),(to_sfixed_a(0.005189346149563789)),(to_sfixed_a(0.0002620580489747226)),(to_sfixed_a(0.0001582805998623371)),(to_sfixed_a(0.1924615502357483)),(to_sfixed_a(-0.0012175095034763217)),(to_sfixed_a(-0.0006273866747505963)),(to_sfixed_a(-0.653071939945221)),(to_sfixed_a(-9.506364585831761e-05)),(to_sfixed_a(-0.0016975936014205217)),(to_sfixed_a(8.65008041728288e-06)),(to_sfixed_a(0.4329850971698761)),(to_sfixed_a(0.003382530529052019)),(to_sfixed_a(0.00022264815925154835)),(to_sfixed_a(0.04418649151921272)),(to_sfixed_a(0.017453841865062714)),(to_sfixed_a(-0.21757203340530396)),(to_sfixed_a(-9.399739792570472e-05)),(to_sfixed_a(1.6896439774427563e-05)),(to_sfixed_a(6.940669845789671e-05)),(to_sfixed_a(0.050378043204545975)),(to_sfixed_a(0.015018457546830177)),(to_sfixed_a(-7.07331346347928e-05)),(to_sfixed_a(-0.08558513969182968)),(to_sfixed_a(0.18984587490558624)),(to_sfixed_a(0.0001078013883670792)),(to_sfixed_a(0.00847066193819046)),(to_sfixed_a(-0.005256948061287403)),(to_sfixed_a(0.00023087047156877816)),(to_sfixed_a(0.01603606715798378)),(to_sfixed_a(0.020300811156630516)),(to_sfixed_a(-0.027933677658438683)),(to_sfixed_a(-2.07592238439247e-05)),(to_sfixed_a(-0.00010615508654154837)),(to_sfixed_a(0.2897983491420746)),(to_sfixed_a(-3.053478940273635e-05)),(to_sfixed_a(0.022160494700074196)),(to_sfixed_a(0.00014992509386502206)),(to_sfixed_a(0.012637819163501263)),(to_sfixed_a(8.945668378146365e-05)),(to_sfixed_a(-0.00011382282536942512)),(to_sfixed_a(-4.623143468052149e-06)),(to_sfixed_a(0.0002728625840973109)),(to_sfixed_a(0.00022754842939320952)),(to_sfixed_a(-0.010094397701323032)),(to_sfixed_a(0.002321638399735093)),(to_sfixed_a(8.471295586787164e-06)),(to_sfixed_a(0.00878140702843666)),(to_sfixed_a(0.3018495440483093)),(to_sfixed_a(-0.02944795973598957)),(to_sfixed_a(1.0664472938515246e-05)),(to_sfixed_a(0.00017844478134065866)),(to_sfixed_a(0.00038901285734027624)),(to_sfixed_a(0.3099714517593384)),(to_sfixed_a(0.3123913109302521)),(to_sfixed_a(-6.565482181031257e-05)),(to_sfixed_a(0.03388773649930954)),(to_sfixed_a(1.7292950360570103e-06)),(to_sfixed_a(0.00015305775741580874)),(to_sfixed_a(0.20631720125675201)),(to_sfixed_a(-0.0006113947601988912)),(to_sfixed_a(0.00012828040053136647)),(to_sfixed_a(0.00022082283976487815)),(to_sfixed_a(-0.004617034923285246)),(to_sfixed_a(5.955036613158882e-05)),(to_sfixed_a(-4.379138772492297e-05)),(to_sfixed_a(0.006235670298337936)),(to_sfixed_a(-0.0003046025522053242)),(to_sfixed_a(-0.00011183024616912007)),(to_sfixed_a(0.0007418274763040245)),(to_sfixed_a(-0.0007953408057801425)),(to_sfixed_a(-0.00013663273421116173)),(to_sfixed_a(6.171033601276577e-05)),(to_sfixed_a(3.849726635962725e-05)),(to_sfixed_a(-2.7147019864059985e-05)),(to_sfixed_a(7.61734918341972e-05)),(to_sfixed_a(-0.0005788196576759219)),(to_sfixed_a(0.06465430557727814)),(to_sfixed_a(7.416515290969983e-05)),(to_sfixed_a(1.7548809410072863e-06)),(to_sfixed_a(0.011241043917834759)),(to_sfixed_a(1.1072026609326713e-05)),(to_sfixed_a(-1.905678800540045e-06)),(to_sfixed_a(-6.415866664610803e-05)),(to_sfixed_a(0.03337894380092621)),(to_sfixed_a(-9.589343244442716e-05)),(to_sfixed_a(-8.083377178991213e-05)),(to_sfixed_a(-0.004614853300154209)),(to_sfixed_a(-0.003666040487587452)),(to_sfixed_a(-0.0003226637782063335)),(to_sfixed_a(-0.0034904819913208485)),(to_sfixed_a(7.052955334074795e-05)),(to_sfixed_a(-6.996859156060964e-05)),(to_sfixed_a(-0.0011529214680194855)),(to_sfixed_a(-3.1871197279542685e-05)),(to_sfixed_a(-7.142321555875242e-05)),(to_sfixed_a(-0.0008634068653918803)),(to_sfixed_a(-0.00015602201165165752)),(to_sfixed_a(0.00015435168461408466)),(to_sfixed_a(-0.38059064745903015)),(to_sfixed_a(0.00021973028196953237)),(to_sfixed_a(-0.2759671211242676)),(to_sfixed_a(0.00019390322268009186)),(to_sfixed_a(0.00024310995650012046)),(to_sfixed_a(-0.0001533488102722913)),(to_sfixed_a(-6.126644439063966e-05)),(to_sfixed_a(-0.5862839221954346)),(to_sfixed_a(0.4128992259502411)),(to_sfixed_a(-0.05683104693889618)),(to_sfixed_a(-0.01977076195180416)),(to_sfixed_a(6.920613668626174e-05)),(to_sfixed_a(0.6520460844039917)),(to_sfixed_a(-8.788946433924139e-05)),(to_sfixed_a(-7.099434151314199e-05)),(to_sfixed_a(-0.5699521899223328)),(to_sfixed_a(-0.2392658293247223)),(to_sfixed_a(-0.0024552112445235252)),(to_sfixed_a(0.00024596427101641893)),(to_sfixed_a(-0.02237764187157154)),(to_sfixed_a(-0.5223709940910339)),(to_sfixed_a(-0.00489156786352396)),(to_sfixed_a(0.002620725193992257)),(to_sfixed_a(0.0027032210491597652)),(to_sfixed_a(0.350947767496109)),(to_sfixed_a(0.0003662863455247134)),(to_sfixed_a(0.3537726402282715)),(to_sfixed_a(1.933637395268306e-05)),(to_sfixed_a(6.753011257387698e-05)),(to_sfixed_a(-1.1093812645412982e-05)),(to_sfixed_a(-0.0073080467991530895)),(to_sfixed_a(-0.00307467277161777)),(to_sfixed_a(-0.005680456757545471)),(to_sfixed_a(0.1349201798439026)),(to_sfixed_a(-0.0064310235902667046)),(to_sfixed_a(-0.05155001953244209)),(to_sfixed_a(9.069579391507432e-05)),(to_sfixed_a(-0.0033015653025358915)),(to_sfixed_a(-0.012866497039794922)),(to_sfixed_a(-5.740371852880344e-05)),(to_sfixed_a(0.5081615447998047)),(to_sfixed_a(1.3815406418871135e-05)),(to_sfixed_a(-0.6562125086784363)),(to_sfixed_a(-0.05388430133461952)),(to_sfixed_a(6.134891009423882e-06)),(to_sfixed_a(7.188173913164064e-05)),(to_sfixed_a(4.535322659648955e-06)),(to_sfixed_a(6.707319698762149e-05)),(to_sfixed_a(3.919802111340687e-05)),(to_sfixed_a(2.981388388434425e-05)),(to_sfixed_a(-0.02597089856863022)),(to_sfixed_a(0.04398816078901291)),(to_sfixed_a(0.0176584180444479)),(to_sfixed_a(-0.012126348912715912)),(to_sfixed_a(-0.02927487902343273)),(to_sfixed_a(-0.02086731046438217)),(to_sfixed_a(-3.2696589187253267e-05)),(to_sfixed_a(0.00022712929057888687)),(to_sfixed_a(2.182374009862542e-05)),(to_sfixed_a(-2.46828276431188e-05)),(to_sfixed_a(-0.00025568262208253145)),(to_sfixed_a(-0.001496730837970972)),(to_sfixed_a(-0.03105863556265831)),(to_sfixed_a(-0.014433132484555244)),(to_sfixed_a(-1.7999293049797416e-05)),(to_sfixed_a(-0.00018039648421108723)),(to_sfixed_a(4.358548540039919e-05)),(to_sfixed_a(-0.00012640305794775486)),(to_sfixed_a(-7.293948328879196e-06)),(to_sfixed_a(0.01883425936102867)),(to_sfixed_a(-4.596106009557843e-06)),(to_sfixed_a(-0.00010822276817634702)),(to_sfixed_a(-6.91033637849614e-05)),(to_sfixed_a(-0.003849429776892066)),(to_sfixed_a(-0.19994047284126282)),(to_sfixed_a(0.0001831354747992009)),(to_sfixed_a(-3.891432425007224e-05)),(to_sfixed_a(0.00014457803627010435)),(to_sfixed_a(3.69284680346027e-06)),(to_sfixed_a(0.0001742475142236799)),(to_sfixed_a(0.00361171318218112)),(to_sfixed_a(-0.1730749011039734)),(to_sfixed_a(-0.00023836939362809062)),(to_sfixed_a(-0.002275241771712899)),(to_sfixed_a(-1.0675939847715199e-05)),(to_sfixed_a(-0.0046708788722753525)),(to_sfixed_a(0.0002907445887103677)),(to_sfixed_a(0.19253945350646973)),(to_sfixed_a(-0.0003128510434180498)),(to_sfixed_a(0.21381399035453796)),(to_sfixed_a(-6.157161260489374e-05)),(to_sfixed_a(0.3002978563308716)),(to_sfixed_a(0.004177771974354982)),(to_sfixed_a(0.0001572242472320795)),(to_sfixed_a(0.013824752531945705)),(to_sfixed_a(-0.01323089748620987)),(to_sfixed_a(3.727634248207323e-05)),(to_sfixed_a(-0.0009378762915730476)),(to_sfixed_a(-5.974383384454995e-06)),(to_sfixed_a(-3.355017543071881e-05)),(to_sfixed_a(0.012134659104049206)),(to_sfixed_a(-0.009732773527503014)),(to_sfixed_a(6.38448545942083e-05)),(to_sfixed_a(-0.00011302130587864667)),(to_sfixed_a(0.6221993565559387)),(to_sfixed_a(-0.00011696148430928588)),(to_sfixed_a(-0.008122291415929794)),(to_sfixed_a(-0.00028408755315467715)),(to_sfixed_a(4.077117773704231e-05)),(to_sfixed_a(-0.0001948846474988386)),(to_sfixed_a(-0.2944170832633972)),(to_sfixed_a(-3.770567127503455e-05)),(to_sfixed_a(-1.7381258658133447e-05)),(to_sfixed_a(-0.00010621668479871005)),(to_sfixed_a(-0.0338602140545845)),(to_sfixed_a(0.37060368061065674)),(to_sfixed_a(-4.781992174685001e-06)),(to_sfixed_a(0.00016803760081529617)),(to_sfixed_a(-0.00011379885108908638)),(to_sfixed_a(5.932248313911259e-06)),(to_sfixed_a(0.4005368947982788)),(to_sfixed_a(0.15326625108718872)),(to_sfixed_a(-0.000525249692145735)),(to_sfixed_a(-0.007672138512134552)),(to_sfixed_a(-0.0014152019284665585)),(to_sfixed_a(-0.00011254505079705268)),(to_sfixed_a(-0.00022803823230788112)),(to_sfixed_a(-0.0003040350857190788)),(to_sfixed_a(-0.0005584100144915283)),(to_sfixed_a(4.3388714402681217e-05)),(to_sfixed_a(-0.00021388279856182635)),(to_sfixed_a(-0.029390856623649597)),(to_sfixed_a(0.005413792096078396)),(to_sfixed_a(3.1139155908022076e-05)),(to_sfixed_a(0.19037485122680664)),(to_sfixed_a(0.000491224869620055)),(to_sfixed_a(-0.26353198289871216)),(to_sfixed_a(0.26358461380004883)),(to_sfixed_a(7.41457988624461e-05)),(to_sfixed_a(-0.03415736183524132)),(to_sfixed_a(0.0012459103018045425)),(to_sfixed_a(0.3145664632320404)),(to_sfixed_a(-5.770285497419536e-05)),(to_sfixed_a(-0.7938746213912964)),(to_sfixed_a(0.3361350893974304)),(to_sfixed_a(-0.6949283480644226)));

    constant weight_n2_34 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.007765611167997122)),(to_sfixed_a(5.3264677262632176e-05)),(to_sfixed_a(0.0001023020813590847)),(to_sfixed_a(-0.00011583839659579098)),(to_sfixed_a(-2.0915118511766195e-05)),(to_sfixed_a(7.209678733488545e-05)),(to_sfixed_a(9.974202839657664e-06)),(to_sfixed_a(-3.234177711419761e-06)),(to_sfixed_a(-1.5130237443372607e-05)),(to_sfixed_a(0.00015020612045191228)),(to_sfixed_a(6.715510971844196e-05)),(to_sfixed_a(-0.0001639665279071778)),(to_sfixed_a(-0.0002715138252824545)),(to_sfixed_a(-0.00010834928980330005)),(to_sfixed_a(-0.00028797000413760543)),(to_sfixed_a(1.1307129170745611e-06)),(to_sfixed_a(-6.554863648489118e-05)),(to_sfixed_a(-0.0002553072990849614)),(to_sfixed_a(-3.358911635586992e-05)),(to_sfixed_a(0.00013571821909863502)),(to_sfixed_a(0.0002989581262227148)),(to_sfixed_a(-0.00011177315900567919)),(to_sfixed_a(2.9901537345722318e-05)),(to_sfixed_a(-7.175866630859673e-05)),(to_sfixed_a(-2.3456726921722293e-05)),(to_sfixed_a(2.8102367650717497e-06)),(to_sfixed_a(-1.4368706615641713e-06)),(to_sfixed_a(7.945744437165558e-05)),(to_sfixed_a(-2.491635677870363e-05)),(to_sfixed_a(6.139795004855841e-06)),(to_sfixed_a(7.044224184937775e-05)),(to_sfixed_a(0.00020436143677216023)),(to_sfixed_a(2.359048812650144e-05)),(to_sfixed_a(-3.874504182022065e-05)),(to_sfixed_a(3.7606427213177085e-05)),(to_sfixed_a(-2.75167403742671e-05)),(to_sfixed_a(-0.00024040217977017164)),(to_sfixed_a(6.885817856527865e-05)),(to_sfixed_a(2.8053182177245617e-05)),(to_sfixed_a(7.10224558133632e-05)),(to_sfixed_a(0.00013784525799565017)),(to_sfixed_a(3.862704033963382e-06)),(to_sfixed_a(0.00011580322461668402)),(to_sfixed_a(0.00021661647770088166)),(to_sfixed_a(7.67033634474501e-05)),(to_sfixed_a(4.994407208869234e-05)),(to_sfixed_a(-3.5007105907425284e-06)),(to_sfixed_a(1.220872945850715e-06)),(to_sfixed_a(-2.2615204215981066e-05)),(to_sfixed_a(-0.00011821352381957695)),(to_sfixed_a(5.002191028324887e-05)),(to_sfixed_a(1.033609441947192e-05)),(to_sfixed_a(9.798633982427418e-06)),(to_sfixed_a(-0.00023703383340034634)),(to_sfixed_a(-2.8367023332975805e-05)),(to_sfixed_a(5.7993071095552295e-05)),(to_sfixed_a(-0.00013485015369951725)),(to_sfixed_a(-0.00010966676927637309)),(to_sfixed_a(0.00011207378702238202)),(to_sfixed_a(2.725741796893999e-05)),(to_sfixed_a(-0.00024807031149975955)),(to_sfixed_a(7.240075501613319e-05)),(to_sfixed_a(2.45669434661977e-06)),(to_sfixed_a(-6.094723357819021e-05)),(to_sfixed_a(0.00010353197285439819)),(to_sfixed_a(-1.2256132322363555e-06)),(to_sfixed_a(-0.00016751624934840947)),(to_sfixed_a(2.4673241568962112e-05)),(to_sfixed_a(-6.606688839383423e-05)),(to_sfixed_a(-0.00010386107169324532)),(to_sfixed_a(-4.88349178340286e-05)),(to_sfixed_a(0.00021905182802584022)),(to_sfixed_a(-0.00015814228390809149)),(to_sfixed_a(-0.00021902147273067385)),(to_sfixed_a(6.345879228319973e-05)),(to_sfixed_a(-0.00026621471624821424)),(to_sfixed_a(-0.0001308958453591913)),(to_sfixed_a(-4.075831384398043e-06)),(to_sfixed_a(-0.00010619076783768833)),(to_sfixed_a(-0.0001242480066139251)),(to_sfixed_a(0.00010413672862341627)),(to_sfixed_a(-6.83675316395238e-05)),(to_sfixed_a(-0.00011481012916192412)),(to_sfixed_a(-2.1476109395734966e-05)),(to_sfixed_a(0.00018141811597160995)),(to_sfixed_a(0.0002356650511501357)),(to_sfixed_a(-2.914288779720664e-05)),(to_sfixed_a(0.00013424460485111922)),(to_sfixed_a(0.00025561207439750433)),(to_sfixed_a(0.00022420051391236484)),(to_sfixed_a(2.2990585421212018e-05)),(to_sfixed_a(-8.011759200599045e-05)),(to_sfixed_a(-3.455417390796356e-05)),(to_sfixed_a(-0.00014433282194659114)),(to_sfixed_a(8.461211109533906e-07)),(to_sfixed_a(5.938755930401385e-05)),(to_sfixed_a(6.79979202686809e-05)),(to_sfixed_a(-4.702310252469033e-05)),(to_sfixed_a(-0.00020515955111477524)),(to_sfixed_a(-8.181687007891014e-07)),(to_sfixed_a(-1.577928924234584e-05)),(to_sfixed_a(1.5006968169473112e-05)),(to_sfixed_a(6.524252239614725e-05)),(to_sfixed_a(-6.212729203980416e-05)),(to_sfixed_a(0.000229474957450293)),(to_sfixed_a(7.131898018997163e-05)),(to_sfixed_a(-0.0004504291864577681)),(to_sfixed_a(2.3366374080069363e-05)),(to_sfixed_a(-1.0712094081100076e-05)),(to_sfixed_a(8.306240488309413e-06)),(to_sfixed_a(-1.8460035789757967e-05)),(to_sfixed_a(8.53178498800844e-05)),(to_sfixed_a(-9.749750461196527e-05)),(to_sfixed_a(-3.236533302697353e-05)),(to_sfixed_a(-6.551637488882989e-05)),(to_sfixed_a(6.288137228693813e-05)),(to_sfixed_a(-0.0001467126130592078)),(to_sfixed_a(-0.0002361536317039281)),(to_sfixed_a(0.00021316533093340695)),(to_sfixed_a(0.00015521817840635777)),(to_sfixed_a(-9.231003787135705e-05)),(to_sfixed_a(-3.7163696106290445e-05)),(to_sfixed_a(-3.679093060782179e-05)),(to_sfixed_a(0.00022003565391059965)),(to_sfixed_a(-3.7760924897156656e-05)),(to_sfixed_a(7.171418110374361e-05)),(to_sfixed_a(-0.0001302993478020653)),(to_sfixed_a(-6.567907985299826e-05)),(to_sfixed_a(0.00010695883975131437)),(to_sfixed_a(1.6905090888030827e-05)),(to_sfixed_a(1.4474891941063106e-05)),(to_sfixed_a(-9.66863299254328e-05)),(to_sfixed_a(-0.0002372068411204964)),(to_sfixed_a(3.903720062226057e-05)),(to_sfixed_a(-0.00010170943278353661)),(to_sfixed_a(-9.552933988743462e-06)),(to_sfixed_a(9.807624155655503e-05)),(to_sfixed_a(-0.00014640529116149992)),(to_sfixed_a(-6.429741915781051e-05)),(to_sfixed_a(-7.403342169709504e-05)),(to_sfixed_a(-0.00017714250134304166)),(to_sfixed_a(2.9997374440426938e-05)),(to_sfixed_a(-0.00016077994951047003)),(to_sfixed_a(-0.00017816823674365878)),(to_sfixed_a(0.0001743239554343745)),(to_sfixed_a(-3.0531555239576846e-05)),(to_sfixed_a(-2.4582586775068194e-05)),(to_sfixed_a(7.13229674147442e-05)),(to_sfixed_a(6.482032767962664e-05)),(to_sfixed_a(-0.00010267547622788697)),(to_sfixed_a(1.3274911907501519e-05)),(to_sfixed_a(-0.00017487190780229867)),(to_sfixed_a(0.00021909041970502585)),(to_sfixed_a(-0.00013022810162510723)),(to_sfixed_a(4.4382446503732353e-05)),(to_sfixed_a(-0.00012090984091628343)),(to_sfixed_a(0.00021376422955654562)),(to_sfixed_a(-0.00015365694707725197)),(to_sfixed_a(-1.2658907508011907e-05)),(to_sfixed_a(-0.000168655562447384)),(to_sfixed_a(-6.855087849544361e-05)),(to_sfixed_a(-1.939760841196403e-05)),(to_sfixed_a(4.38140268670395e-05)),(to_sfixed_a(-0.000273020938038826)),(to_sfixed_a(-0.00041038059862330556)),(to_sfixed_a(-0.00019995725597254932)),(to_sfixed_a(-0.00013736374967265874)),(to_sfixed_a(0.00015092674584593624)),(to_sfixed_a(0.00022312677174340934)),(to_sfixed_a(0.00023081974359229207)),(to_sfixed_a(0.00021365370776038617)),(to_sfixed_a(-9.205887181451544e-06)),(to_sfixed_a(-0.0001478493504691869)),(to_sfixed_a(-9.933569526765496e-05)),(to_sfixed_a(0.00014702323824167252)),(to_sfixed_a(-5.855525523656979e-05)),(to_sfixed_a(6.822584691690281e-05)),(to_sfixed_a(0.00010053992446046323)),(to_sfixed_a(1.3337048585526645e-06)),(to_sfixed_a(-0.00020379586203489453)),(to_sfixed_a(6.58759381622076e-05)),(to_sfixed_a(-5.027032966609113e-05)),(to_sfixed_a(4.593968333210796e-05)),(to_sfixed_a(-0.00014794257003813982)),(to_sfixed_a(9.885936015052721e-05)),(to_sfixed_a(6.7486209445633e-05)),(to_sfixed_a(0.00018789201567415148)),(to_sfixed_a(-9.813129145186394e-05)),(to_sfixed_a(8.57507111504674e-05)),(to_sfixed_a(-1.1460651876404881e-06)),(to_sfixed_a(0.00013532009324990213)),(to_sfixed_a(0.00045910265180282295)),(to_sfixed_a(-0.000160182811669074)),(to_sfixed_a(0.00016695796512067318)),(to_sfixed_a(-7.103084499249235e-05)),(to_sfixed_a(0.00020151784701738507)),(to_sfixed_a(2.0191808289382607e-05)),(to_sfixed_a(-2.1484513126779348e-05)),(to_sfixed_a(-3.221472798031755e-05)),(to_sfixed_a(-7.177675433922559e-05)),(to_sfixed_a(0.0001161086474894546)),(to_sfixed_a(0.0001984386908588931)),(to_sfixed_a(-5.3654221119359136e-06)),(to_sfixed_a(5.6614720961079e-05)),(to_sfixed_a(1.580883690621704e-08)),(to_sfixed_a(0.00024719833163544536)),(to_sfixed_a(0.000315631739795208)),(to_sfixed_a(-0.00010687822941690683)),(to_sfixed_a(1.2318949302425608e-05)),(to_sfixed_a(-0.0001261538127437234)),(to_sfixed_a(0.00010196266521234065)),(to_sfixed_a(0.00013486196985468268)),(to_sfixed_a(5.670636164722964e-05)),(to_sfixed_a(6.919393490534276e-05)),(to_sfixed_a(0.00023951703042257577)),(to_sfixed_a(-3.3505639294162393e-06)),(to_sfixed_a(0.00019695449736900628)),(to_sfixed_a(0.00011263399210292846)),(to_sfixed_a(0.00024255836615338922)),(to_sfixed_a(-0.00019585069094318897)),(to_sfixed_a(-0.0002618785365484655)),(to_sfixed_a(0.00011593430826906115)),(to_sfixed_a(-0.00018259095668327063)),(to_sfixed_a(0.0001394545251969248)),(to_sfixed_a(0.00020992050122004002)),(to_sfixed_a(6.769933679606766e-05)),(to_sfixed_a(8.105755114229396e-05)),(to_sfixed_a(4.114345938432962e-05)),(to_sfixed_a(0.00012804035213775933)),(to_sfixed_a(5.247049557510763e-06)),(to_sfixed_a(-0.00021588838717434555)),(to_sfixed_a(-0.00024692603619769216)),(to_sfixed_a(2.549404962337576e-05)),(to_sfixed_a(8.88686699909158e-05)),(to_sfixed_a(0.00019473560678306967)),(to_sfixed_a(3.9454243960790336e-05)),(to_sfixed_a(-0.00017953114002011716)),(to_sfixed_a(0.00016796450654510409)),(to_sfixed_a(-0.00021997056319378316)),(to_sfixed_a(-0.00013560762454289943)),(to_sfixed_a(-5.704862269340083e-05)),(to_sfixed_a(-6.0898186347913e-05)),(to_sfixed_a(-0.00029679856379516423)),(to_sfixed_a(7.278996054083109e-05)),(to_sfixed_a(0.00021731603192165494)),(to_sfixed_a(0.00016814352420624346)),(to_sfixed_a(-2.1715650291298516e-05)),(to_sfixed_a(2.4237684556283057e-05)),(to_sfixed_a(-2.8566186301759444e-05)),(to_sfixed_a(-6.13446973147802e-05)),(to_sfixed_a(0.00010425738582853228)),(to_sfixed_a(-4.494448148761876e-05)),(to_sfixed_a(-4.096602788195014e-05)),(to_sfixed_a(-0.0001458938786527142)),(to_sfixed_a(-5.049518222222105e-06)),(to_sfixed_a(6.74518960295245e-05)),(to_sfixed_a(-0.0001204604996019043)),(to_sfixed_a(-0.00015925962361507118)),(to_sfixed_a(-5.9785063058370724e-05)),(to_sfixed_a(1.0097995982505381e-05)),(to_sfixed_a(0.00014124991139397025)),(to_sfixed_a(2.7236819732934237e-05)),(to_sfixed_a(-0.00014621129957959056)),(to_sfixed_a(-8.413419709540904e-05)),(to_sfixed_a(-2.4482178559992462e-05)),(to_sfixed_a(-0.00010823279444593936)),(to_sfixed_a(-0.00022059892944525927)),(to_sfixed_a(5.24066126672551e-06)),(to_sfixed_a(-3.748037852346897e-05)),(to_sfixed_a(-7.11842585587874e-05)),(to_sfixed_a(-1.5555662685073912e-05)),(to_sfixed_a(-3.0746887205168605e-05)),(to_sfixed_a(-4.491842264542356e-05)),(to_sfixed_a(-0.0001350170496152714)),(to_sfixed_a(0.00010459952318342403)),(to_sfixed_a(-2.1790390746900812e-05)),(to_sfixed_a(2.6179346605204046e-05)),(to_sfixed_a(-1.1207954230485484e-05)),(to_sfixed_a(-0.00021352140174712986)),(to_sfixed_a(-1.0696712706703693e-05)),(to_sfixed_a(-0.00010882128844968975)),(to_sfixed_a(-0.0001268786727450788)),(to_sfixed_a(-9.685174154583365e-05)),(to_sfixed_a(-6.58450007904321e-05)),(to_sfixed_a(-0.00015445597819052637)),(to_sfixed_a(0.00020933570340275764)),(to_sfixed_a(-6.231560837477446e-05)),(to_sfixed_a(-3.0832889024168253e-06)),(to_sfixed_a(-4.4494550820672885e-05)),(to_sfixed_a(-0.00012967796646989882)),(to_sfixed_a(4.0459381125401706e-05)),(to_sfixed_a(3.5382763599045575e-05)),(to_sfixed_a(-4.779821028932929e-05)),(to_sfixed_a(6.202564691193402e-06)),(to_sfixed_a(-4.4405787775758654e-05)),(to_sfixed_a(-0.00032371506677009165)),(to_sfixed_a(-1.795322896214202e-05)),(to_sfixed_a(-0.0002154648391297087)),(to_sfixed_a(-1.1546137102413923e-05)),(to_sfixed_a(-7.027147512417287e-05)),(to_sfixed_a(-1.7262864275835454e-05)));

    constant weight_n2_35 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.24961994588375092)),(to_sfixed_a(0.48884156346321106)),(to_sfixed_a(0.0012587885139510036)),(to_sfixed_a(-4.4814994907937944e-05)),(to_sfixed_a(-0.8717231750488281)),(to_sfixed_a(-0.00031237772782333195)),(to_sfixed_a(0.00042583720642142)),(to_sfixed_a(8.933345816330984e-05)),(to_sfixed_a(6.997634773142636e-05)),(to_sfixed_a(0.00017909743473865092)),(to_sfixed_a(3.1885658245300874e-05)),(to_sfixed_a(0.00030745496042072773)),(to_sfixed_a(-0.10236390680074692)),(to_sfixed_a(7.737553823972121e-05)),(to_sfixed_a(0.00015310815069824457)),(to_sfixed_a(3.888251376338303e-05)),(to_sfixed_a(-0.0015660385834053159)),(to_sfixed_a(0.0001556359202368185)),(to_sfixed_a(-0.005341212265193462)),(to_sfixed_a(2.0244558982085437e-05)),(to_sfixed_a(0.00010711689537856728)),(to_sfixed_a(0.00024724495597183704)),(to_sfixed_a(-0.00011223632463952526)),(to_sfixed_a(0.0007050548447296023)),(to_sfixed_a(0.38373926281929016)),(to_sfixed_a(3.2148936952580698e-06)),(to_sfixed_a(-0.00016675176448188722)),(to_sfixed_a(5.928127393417526e-06)),(to_sfixed_a(2.2889955289429054e-05)),(to_sfixed_a(-7.131033635232598e-05)),(to_sfixed_a(0.002083780709654093)),(to_sfixed_a(-2.3427404812537134e-05)),(to_sfixed_a(0.00014837720664218068)),(to_sfixed_a(0.00014706389629282057)),(to_sfixed_a(0.0002002684195758775)),(to_sfixed_a(-0.0002973819791804999)),(to_sfixed_a(-0.00042905096779577434)),(to_sfixed_a(0.0033987020142376423)),(to_sfixed_a(-0.0013204924762248993)),(to_sfixed_a(-8.991489448817447e-05)),(to_sfixed_a(0.00018016992544289678)),(to_sfixed_a(-0.007540538907051086)),(to_sfixed_a(-1.3980534276925027e-05)),(to_sfixed_a(-0.00011282514606136829)),(to_sfixed_a(0.00045501443673856556)),(to_sfixed_a(0.002549282042309642)),(to_sfixed_a(-0.0015751540195196867)),(to_sfixed_a(4.573138721752912e-05)),(to_sfixed_a(-0.0004538946959655732)),(to_sfixed_a(-0.12036100029945374)),(to_sfixed_a(0.5208691954612732)),(to_sfixed_a(0.0005951590719632804)),(to_sfixed_a(-0.00030178550514392555)),(to_sfixed_a(-0.24864619970321655)),(to_sfixed_a(0.0010114092146977782)),(to_sfixed_a(-0.3342495560646057)),(to_sfixed_a(2.5821718736551702e-05)),(to_sfixed_a(-0.000984259182587266)),(to_sfixed_a(0.00019151667947880924)),(to_sfixed_a(-0.0001144974012277089)),(to_sfixed_a(5.4241932957665995e-05)),(to_sfixed_a(0.13031618297100067)),(to_sfixed_a(7.872045534895733e-05)),(to_sfixed_a(0.22577403485774994)),(to_sfixed_a(-0.0003057505236938596)),(to_sfixed_a(5.8646317484090105e-05)),(to_sfixed_a(-0.00041309246444143355)),(to_sfixed_a(-0.0037073635030537844)),(to_sfixed_a(7.14797861292027e-05)),(to_sfixed_a(-6.557349115610123e-05)),(to_sfixed_a(-0.010160313919186592)),(to_sfixed_a(-0.004063200205564499)),(to_sfixed_a(-0.001205763197503984)),(to_sfixed_a(0.00018133051344193518)),(to_sfixed_a(0.0002730154665187001)),(to_sfixed_a(-2.646858774824068e-05)),(to_sfixed_a(0.06718023866415024)),(to_sfixed_a(-4.149108463025186e-06)),(to_sfixed_a(4.285346221877262e-06)),(to_sfixed_a(-0.004259779583662748)),(to_sfixed_a(0.00028142431983724236)),(to_sfixed_a(0.00017651828238740563)),(to_sfixed_a(0.00014588263002224267)),(to_sfixed_a(-0.0016127392882481217)),(to_sfixed_a(-5.738078471040353e-05)),(to_sfixed_a(0.0010794405825436115)),(to_sfixed_a(0.0023713461123406887)),(to_sfixed_a(0.00022917245223652571)),(to_sfixed_a(1.2446234904928133e-05)),(to_sfixed_a(-0.00019851085380651057)),(to_sfixed_a(-0.44614794850349426)),(to_sfixed_a(0.00017592076619621366)),(to_sfixed_a(0.0006648826529271901)),(to_sfixed_a(2.6154943043366075e-05)),(to_sfixed_a(0.00016498954209964722)),(to_sfixed_a(5.139756467542611e-05)),(to_sfixed_a(4.669932241085917e-05)),(to_sfixed_a(-0.0002008661103900522)),(to_sfixed_a(0.00011238895240239799)),(to_sfixed_a(0.0004503997042775154)),(to_sfixed_a(0.011486616916954517)),(to_sfixed_a(3.8580503314733505e-05)),(to_sfixed_a(-0.00029594270745292306)),(to_sfixed_a(0.2294463813304901)),(to_sfixed_a(-0.0002044205612037331)),(to_sfixed_a(9.935277194017544e-05)),(to_sfixed_a(2.4385706637986004e-05)),(to_sfixed_a(-7.652718340978026e-05)),(to_sfixed_a(-4.174595233052969e-06)),(to_sfixed_a(0.34215566515922546)),(to_sfixed_a(-0.3030516803264618)),(to_sfixed_a(-8.887495641829446e-05)),(to_sfixed_a(0.0034737985115498304)),(to_sfixed_a(-0.00011265256762271747)),(to_sfixed_a(-3.193671000190079e-05)),(to_sfixed_a(-0.3235040307044983)),(to_sfixed_a(2.155571746698115e-05)),(to_sfixed_a(2.251247497042641e-05)),(to_sfixed_a(0.0001996166247408837)),(to_sfixed_a(-0.00029944576090201735)),(to_sfixed_a(-4.507688572630286e-06)),(to_sfixed_a(-0.00016845317441038787)),(to_sfixed_a(-1.908410013129469e-06)),(to_sfixed_a(2.7159665478393435e-05)),(to_sfixed_a(4.6439901780104265e-05)),(to_sfixed_a(-0.0006495062843896449)),(to_sfixed_a(-0.007970509119331837)),(to_sfixed_a(3.710822420543991e-05)),(to_sfixed_a(-0.0001453560689697042)),(to_sfixed_a(0.000324983149766922)),(to_sfixed_a(-1.6672493075020611e-06)),(to_sfixed_a(1.159423845820129e-06)),(to_sfixed_a(-0.002365588443353772)),(to_sfixed_a(-0.05054296553134918)),(to_sfixed_a(-5.7127959735225886e-05)),(to_sfixed_a(0.00013049677363596857)),(to_sfixed_a(0.1098051369190216)),(to_sfixed_a(0.00013364361075218767)),(to_sfixed_a(-0.00011597572301980108)),(to_sfixed_a(0.00011771984281949699)),(to_sfixed_a(-8.410483133047819e-05)),(to_sfixed_a(0.00027168128872290254)),(to_sfixed_a(-2.4898965421016328e-05)),(to_sfixed_a(-8.25706374598667e-05)),(to_sfixed_a(-0.000620292907115072)),(to_sfixed_a(6.748661689925939e-06)),(to_sfixed_a(-2.5064040528377518e-05)),(to_sfixed_a(1.854914444265887e-05)),(to_sfixed_a(-0.0004543148388620466)),(to_sfixed_a(-0.004487532190978527)),(to_sfixed_a(1.785897620720789e-05)),(to_sfixed_a(0.00030182115733623505)),(to_sfixed_a(0.001892292988486588)),(to_sfixed_a(-1.207599780173041e-05)),(to_sfixed_a(-5.969251651549712e-05)),(to_sfixed_a(0.12395667284727097)),(to_sfixed_a(-3.19686732836999e-05)),(to_sfixed_a(-0.003594022709876299)),(to_sfixed_a(2.1490062863449566e-05)),(to_sfixed_a(-0.0002237481385236606)),(to_sfixed_a(-5.48841489944607e-06)),(to_sfixed_a(-0.00015415159577969462)),(to_sfixed_a(0.2873677909374237)),(to_sfixed_a(-0.0009229840943589807)),(to_sfixed_a(0.00020407343981787562)),(to_sfixed_a(0.2322043627500534)),(to_sfixed_a(-0.00014976623060647398)),(to_sfixed_a(2.0679297449532896e-05)),(to_sfixed_a(-7.197494414867833e-05)),(to_sfixed_a(2.58167419815436e-05)),(to_sfixed_a(0.006675341632217169)),(to_sfixed_a(-0.003611598629504442)),(to_sfixed_a(0.37280401587486267)),(to_sfixed_a(0.0002626572677399963)),(to_sfixed_a(-0.0052338652312755585)),(to_sfixed_a(-0.00021697729243896902)),(to_sfixed_a(-0.0001396554580423981)),(to_sfixed_a(0.3879815340042114)),(to_sfixed_a(-0.08737540245056152)),(to_sfixed_a(-0.04710576310753822)),(to_sfixed_a(2.8813003154937178e-05)),(to_sfixed_a(-0.004300205036997795)),(to_sfixed_a(-0.00022817360877525061)),(to_sfixed_a(-0.00022320865537039936)),(to_sfixed_a(-4.7080739022931084e-05)),(to_sfixed_a(4.7446301323361695e-05)),(to_sfixed_a(0.09996675699949265)),(to_sfixed_a(-0.00019403506303206086)),(to_sfixed_a(-4.837189771933481e-05)),(to_sfixed_a(0.0002627211797516793)),(to_sfixed_a(-0.0001947289565578103)),(to_sfixed_a(0.00015499387518502772)),(to_sfixed_a(0.0009928988292813301)),(to_sfixed_a(1.8618618923937902e-05)),(to_sfixed_a(4.7436980821657926e-05)),(to_sfixed_a(-0.004474497865885496)),(to_sfixed_a(-9.80372351477854e-05)),(to_sfixed_a(-0.001970263896510005)),(to_sfixed_a(0.0013264347799122334)),(to_sfixed_a(1.385077484883368e-05)),(to_sfixed_a(0.00012879515998065472)),(to_sfixed_a(-1.1687145160976797e-05)),(to_sfixed_a(0.00014024754636920989)),(to_sfixed_a(1.679475826676935e-05)),(to_sfixed_a(-0.00014030918828211725)),(to_sfixed_a(-0.010326571762561798)),(to_sfixed_a(0.00027530285296961665)),(to_sfixed_a(-0.4364073574542999)),(to_sfixed_a(0.0009186725947074592)),(to_sfixed_a(1.7679536540526897e-05)),(to_sfixed_a(-0.00043100822949782014)),(to_sfixed_a(0.00023237444111146033)),(to_sfixed_a(-0.0001121495442930609)),(to_sfixed_a(-0.00020671289530582726)),(to_sfixed_a(3.733459016075358e-05)),(to_sfixed_a(-7.105151598807424e-05)),(to_sfixed_a(-0.006191853433847427)),(to_sfixed_a(-0.000808968092314899)),(to_sfixed_a(-0.01367000862956047)),(to_sfixed_a(0.00023655517725273967)),(to_sfixed_a(-7.060127973090857e-05)),(to_sfixed_a(0.0001719656283967197)),(to_sfixed_a(0.00016990127915050834)),(to_sfixed_a(-8.490671461913735e-05)),(to_sfixed_a(-0.008241785690188408)),(to_sfixed_a(5.526597669813782e-05)),(to_sfixed_a(2.777461486402899e-05)),(to_sfixed_a(2.9969642127980478e-05)),(to_sfixed_a(-0.016166500747203827)),(to_sfixed_a(0.0011775735765695572)),(to_sfixed_a(-0.001093233935534954)),(to_sfixed_a(-2.5639223167672753e-05)),(to_sfixed_a(-0.00010102165106218308)),(to_sfixed_a(1.3143864634912461e-05)),(to_sfixed_a(0.0020969295874238014)),(to_sfixed_a(-0.00044550816528499126)),(to_sfixed_a(0.0005001971148885787)),(to_sfixed_a(-8.521582640241832e-05)),(to_sfixed_a(-7.92821665527299e-05)),(to_sfixed_a(-0.00015982706099748611)),(to_sfixed_a(0.00302535155788064)),(to_sfixed_a(7.943860691739246e-05)),(to_sfixed_a(0.0002636041899677366)),(to_sfixed_a(-1.0852381819859147e-06)),(to_sfixed_a(-0.006186866667121649)),(to_sfixed_a(-2.2412617909139954e-05)),(to_sfixed_a(-0.0013998141512274742)),(to_sfixed_a(-0.5336822271347046)),(to_sfixed_a(-0.00044892641017213464)),(to_sfixed_a(0.00368110672570765)),(to_sfixed_a(-2.297647370141931e-07)),(to_sfixed_a(-1.9123952370136976e-05)),(to_sfixed_a(-0.0007477287435904145)),(to_sfixed_a(-9.789733303477988e-05)),(to_sfixed_a(-0.00012937880819663405)),(to_sfixed_a(0.0005740200285799801)),(to_sfixed_a(0.0015147430822253227)),(to_sfixed_a(-2.3836124455556273e-05)),(to_sfixed_a(0.00013516204489860684)),(to_sfixed_a(-4.2145984480157495e-05)),(to_sfixed_a(-6.6862121457234025e-06)),(to_sfixed_a(-0.000515719351824373)),(to_sfixed_a(-0.00014779780758544803)),(to_sfixed_a(-7.685463788220659e-05)),(to_sfixed_a(1.8901730072684586e-05)),(to_sfixed_a(0.0024957589339464903)),(to_sfixed_a(-0.0004504687385633588)),(to_sfixed_a(0.00011548816837603226)),(to_sfixed_a(0.000196376015082933)),(to_sfixed_a(-0.002379473764449358)),(to_sfixed_a(-0.39661264419555664)),(to_sfixed_a(-0.000383209902793169)),(to_sfixed_a(2.73755140369758e-05)),(to_sfixed_a(0.00017040043894667178)),(to_sfixed_a(-2.868169394787401e-05)),(to_sfixed_a(0.0036156955175101757)),(to_sfixed_a(0.0028481108602136374)),(to_sfixed_a(0.0004902424989268184)),(to_sfixed_a(-0.020420165732502937)),(to_sfixed_a(-0.0006415003444999456)),(to_sfixed_a(1.0727522749220952e-05)),(to_sfixed_a(4.716413241112605e-05)),(to_sfixed_a(-7.144399569369853e-05)),(to_sfixed_a(8.937592792790383e-05)),(to_sfixed_a(6.794622458983213e-05)),(to_sfixed_a(-5.068931932328269e-05)),(to_sfixed_a(3.4700948162935674e-05)),(to_sfixed_a(-0.011440051719546318)),(to_sfixed_a(-6.525059143314138e-05)),(to_sfixed_a(-0.00025319517590105534)),(to_sfixed_a(0.0001665637391852215)),(to_sfixed_a(-0.0011274628341197968)),(to_sfixed_a(-0.01674564741551876)),(to_sfixed_a(-0.00016819030861370265)),(to_sfixed_a(4.628370516002178e-05)),(to_sfixed_a(-4.51075311502791e-06)),(to_sfixed_a(-0.0009438868146389723)),(to_sfixed_a(-6.255708285607398e-05)),(to_sfixed_a(0.0006949887028895319)),(to_sfixed_a(0.0022623019758611917)),(to_sfixed_a(0.2891712188720703)));

    constant weight_n2_36 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.27648162841796875)),(to_sfixed_a(-0.005116987973451614)),(to_sfixed_a(-0.3025364875793457)),(to_sfixed_a(6.128758832346648e-05)),(to_sfixed_a(-0.009116563946008682)),(to_sfixed_a(0.00022133962193038315)),(to_sfixed_a(-0.00014896527864038944)),(to_sfixed_a(-6.766132719349116e-05)),(to_sfixed_a(-4.137065843679011e-05)),(to_sfixed_a(5.798527126898989e-05)),(to_sfixed_a(-3.970650868723169e-05)),(to_sfixed_a(-0.00017922744154930115)),(to_sfixed_a(-0.0148966945707798)),(to_sfixed_a(-0.005528370849788189)),(to_sfixed_a(4.8883972340263426e-05)),(to_sfixed_a(4.733436071546748e-05)),(to_sfixed_a(-0.005282024387270212)),(to_sfixed_a(-4.736693517770618e-05)),(to_sfixed_a(-0.0036114556714892387)),(to_sfixed_a(-0.00015133011038415134)),(to_sfixed_a(1.3580847735283896e-06)),(to_sfixed_a(-0.00011621323210420087)),(to_sfixed_a(6.298310472629964e-05)),(to_sfixed_a(0.0023994676303118467)),(to_sfixed_a(-0.0017624989850446582)),(to_sfixed_a(-0.003685667645186186)),(to_sfixed_a(0.00012962684559170157)),(to_sfixed_a(1.4255008863983676e-05)),(to_sfixed_a(-0.00616412702947855)),(to_sfixed_a(0.00020013589528389275)),(to_sfixed_a(-0.0018190834671258926)),(to_sfixed_a(-2.2278363758232445e-06)),(to_sfixed_a(-0.008533522486686707)),(to_sfixed_a(0.0004506015975493938)),(to_sfixed_a(-1.9085673557128757e-05)),(to_sfixed_a(0.00011999981506960467)),(to_sfixed_a(0.3844660222530365)),(to_sfixed_a(0.16727159917354584)),(to_sfixed_a(0.005746711976826191)),(to_sfixed_a(0.00010283621668349952)),(to_sfixed_a(0.28065425157546997)),(to_sfixed_a(0.00012085348134860396)),(to_sfixed_a(-3.8889324059709907e-05)),(to_sfixed_a(0.0001346825301880017)),(to_sfixed_a(-0.00800062995404005)),(to_sfixed_a(-0.01797066442668438)),(to_sfixed_a(-0.00264258636161685)),(to_sfixed_a(-0.011226894333958626)),(to_sfixed_a(0.00017731628031469882)),(to_sfixed_a(-0.00975853018462658)),(to_sfixed_a(-0.007186423521488905)),(to_sfixed_a(0.0003252592287026346)),(to_sfixed_a(-0.0002818738576024771)),(to_sfixed_a(-0.0006139979232102633)),(to_sfixed_a(-0.005651930812746286)),(to_sfixed_a(-0.002697655465453863)),(to_sfixed_a(0.0002787247358355671)),(to_sfixed_a(-0.0007092201267369092)),(to_sfixed_a(-0.00017528038006275892)),(to_sfixed_a(-5.690066609531641e-05)),(to_sfixed_a(0.00022950241691432893)),(to_sfixed_a(8.807775157038122e-05)),(to_sfixed_a(-4.58846589026507e-05)),(to_sfixed_a(-0.002565397648140788)),(to_sfixed_a(6.13317679380998e-05)),(to_sfixed_a(-0.0019552120938897133)),(to_sfixed_a(0.00017542045679874718)),(to_sfixed_a(-0.007560305297374725)),(to_sfixed_a(-0.0017618617275729775)),(to_sfixed_a(0.00010583353287074715)),(to_sfixed_a(-0.00304311141371727)),(to_sfixed_a(-0.002150757936760783)),(to_sfixed_a(0.0014015210326761007)),(to_sfixed_a(-0.00022716830426361412)),(to_sfixed_a(-0.0001125894850702025)),(to_sfixed_a(0.00017545573064126074)),(to_sfixed_a(-0.1674080640077591)),(to_sfixed_a(1.8836153685697354e-06)),(to_sfixed_a(-0.00016820619930513203)),(to_sfixed_a(-0.009430835023522377)),(to_sfixed_a(-3.2948271837085485e-05)),(to_sfixed_a(-7.006266969256103e-05)),(to_sfixed_a(-0.0007346495985984802)),(to_sfixed_a(-0.0013903460931032896)),(to_sfixed_a(-8.082880958681926e-05)),(to_sfixed_a(-0.005507109686732292)),(to_sfixed_a(0.0148124098777771)),(to_sfixed_a(8.023780537769198e-05)),(to_sfixed_a(-0.00018823539721779525)),(to_sfixed_a(-0.00011464783165138215)),(to_sfixed_a(-0.006183736026287079)),(to_sfixed_a(7.738661952316761e-05)),(to_sfixed_a(-3.8336103898473084e-05)),(to_sfixed_a(0.00012895329564344138)),(to_sfixed_a(-0.0022912530694156885)),(to_sfixed_a(2.478049100318458e-05)),(to_sfixed_a(-0.00042071309871971607)),(to_sfixed_a(-0.00015681955846957862)),(to_sfixed_a(0.00015172670828178525)),(to_sfixed_a(-6.507483340101317e-05)),(to_sfixed_a(0.0017928654560819268)),(to_sfixed_a(-0.0010018439497798681)),(to_sfixed_a(-0.00015152301057241857)),(to_sfixed_a(-0.0006571806152351201)),(to_sfixed_a(-0.0028736658859997988)),(to_sfixed_a(-0.000258027168456465)),(to_sfixed_a(0.00024227386165875942)),(to_sfixed_a(7.420623296638951e-05)),(to_sfixed_a(-0.00015748999430797994)),(to_sfixed_a(-0.006965308915823698)),(to_sfixed_a(-0.0008024901035241783)),(to_sfixed_a(3.5530571039998904e-05)),(to_sfixed_a(-0.005746831651777029)),(to_sfixed_a(0.00011228431685594842)),(to_sfixed_a(-8.510227780789137e-05)),(to_sfixed_a(-0.0062981960363686085)),(to_sfixed_a(1.578953924763482e-05)),(to_sfixed_a(6.218114867806435e-05)),(to_sfixed_a(-0.00017252667748834938)),(to_sfixed_a(-0.008757713250815868)),(to_sfixed_a(6.271510210353881e-05)),(to_sfixed_a(-1.3752323866356164e-05)),(to_sfixed_a(-1.0509204003028572e-05)),(to_sfixed_a(-6.135590956546366e-05)),(to_sfixed_a(0.00010765697516035289)),(to_sfixed_a(0.01869690977036953)),(to_sfixed_a(0.001427017035894096)),(to_sfixed_a(-4.43702083430253e-05)),(to_sfixed_a(4.1566891013644636e-06)),(to_sfixed_a(6.402307190001011e-05)),(to_sfixed_a(-0.0002862729597836733)),(to_sfixed_a(-4.6649001887999475e-06)),(to_sfixed_a(-0.0014166292967274785)),(to_sfixed_a(-0.0023832074366509914)),(to_sfixed_a(-0.00010586230928311124)),(to_sfixed_a(0.00016621837858110666)),(to_sfixed_a(0.0037686252035200596)),(to_sfixed_a(0.00016226849402301013)),(to_sfixed_a(-0.0002426877326797694)),(to_sfixed_a(1.2540571333374828e-05)),(to_sfixed_a(0.002936962293460965)),(to_sfixed_a(-3.255573028582148e-05)),(to_sfixed_a(7.117839413695037e-05)),(to_sfixed_a(-6.921511521795765e-05)),(to_sfixed_a(-0.0016677621752023697)),(to_sfixed_a(-0.00045424283598549664)),(to_sfixed_a(-0.0008399350917898118)),(to_sfixed_a(5.9878879255848005e-05)),(to_sfixed_a(0.00012073605466866866)),(to_sfixed_a(-0.00525179598480463)),(to_sfixed_a(-5.7599761930759996e-05)),(to_sfixed_a(-0.00015320298552978784)),(to_sfixed_a(-3.607167673180811e-05)),(to_sfixed_a(3.635250322986394e-07)),(to_sfixed_a(-0.00023816575412638485)),(to_sfixed_a(-0.0016418491723015904)),(to_sfixed_a(-6.895548722241074e-06)),(to_sfixed_a(0.0036418752279132605)),(to_sfixed_a(8.650121162645519e-05)),(to_sfixed_a(6.24240783508867e-06)),(to_sfixed_a(5.222248364589177e-05)),(to_sfixed_a(0.00017662154277786613)),(to_sfixed_a(0.0049650645814836025)),(to_sfixed_a(-0.004365622531622648)),(to_sfixed_a(-0.00548909604549408)),(to_sfixed_a(-0.0059603918343782425)),(to_sfixed_a(-0.00011698879825416952)),(to_sfixed_a(0.021526450291275978)),(to_sfixed_a(-0.0001057551708072424)),(to_sfixed_a(0.0003170559066347778)),(to_sfixed_a(-0.0019947595428675413)),(to_sfixed_a(-0.002887614071369171)),(to_sfixed_a(-0.004201866220682859)),(to_sfixed_a(-6.471600499935448e-07)),(to_sfixed_a(0.008232724852859974)),(to_sfixed_a(0.00034125568345189095)),(to_sfixed_a(-0.0005277948803268373)),(to_sfixed_a(-0.00062053237343207)),(to_sfixed_a(-0.00357270915992558)),(to_sfixed_a(0.2989380359649658)),(to_sfixed_a(0.00042993901297450066)),(to_sfixed_a(-0.016756778582930565)),(to_sfixed_a(6.835159729234874e-05)),(to_sfixed_a(-3.1792278605280444e-05)),(to_sfixed_a(-4.85076816403307e-06)),(to_sfixed_a(-0.0010811041574925184)),(to_sfixed_a(0.03153520077466965)),(to_sfixed_a(-0.002111786510795355)),(to_sfixed_a(-7.45114084566012e-06)),(to_sfixed_a(1.052171501214616e-05)),(to_sfixed_a(-0.0032379585318267345)),(to_sfixed_a(0.00028718746034428477)),(to_sfixed_a(-0.0024770854506641626)),(to_sfixed_a(-4.320190055295825e-05)),(to_sfixed_a(-0.0003019258438143879)),(to_sfixed_a(0.2693368196487427)),(to_sfixed_a(-6.196739559527487e-05)),(to_sfixed_a(0.004536382853984833)),(to_sfixed_a(0.00021738599753007293)),(to_sfixed_a(3.495874989312142e-05)),(to_sfixed_a(-5.7885394198819995e-05)),(to_sfixed_a(-0.00015542576147709042)),(to_sfixed_a(-5.555964889936149e-06)),(to_sfixed_a(-0.00016187339497264475)),(to_sfixed_a(-7.152769831009209e-05)),(to_sfixed_a(1.724396861391142e-05)),(to_sfixed_a(-0.5383073091506958)),(to_sfixed_a(-0.5562257170677185)),(to_sfixed_a(-0.00018993030244018883)),(to_sfixed_a(-0.0006860829889774323)),(to_sfixed_a(-0.0005773617886006832)),(to_sfixed_a(3.941437171306461e-05)),(to_sfixed_a(-0.00017950327310245484)),(to_sfixed_a(-0.0002696684969123453)),(to_sfixed_a(-0.0001730516378302127)),(to_sfixed_a(6.37766279396601e-05)),(to_sfixed_a(0.000350208196323365)),(to_sfixed_a(-0.0002785550314001739)),(to_sfixed_a(-0.0010498762130737305)),(to_sfixed_a(0.0001493987801950425)),(to_sfixed_a(0.00015447399346157908)),(to_sfixed_a(4.4243206502869725e-06)),(to_sfixed_a(5.63951107324101e-06)),(to_sfixed_a(-4.486172110773623e-05)),(to_sfixed_a(-0.3345175087451935)),(to_sfixed_a(3.0724331736564636e-05)),(to_sfixed_a(0.00011752748105209321)),(to_sfixed_a(2.4489418137818575e-07)),(to_sfixed_a(-0.00011728572280844674)),(to_sfixed_a(0.0017371518770232797)),(to_sfixed_a(-0.004105179104954004)),(to_sfixed_a(0.00012972891272511333)),(to_sfixed_a(0.0001070195939973928)),(to_sfixed_a(-9.588220564182848e-06)),(to_sfixed_a(0.00030627386877313256)),(to_sfixed_a(-0.0011637385468930006)),(to_sfixed_a(-0.24228456616401672)),(to_sfixed_a(0.0004489345592446625)),(to_sfixed_a(-6.736510840710253e-05)),(to_sfixed_a(-0.0001868469116743654)),(to_sfixed_a(-0.003540129866451025)),(to_sfixed_a(-5.580821743933484e-05)),(to_sfixed_a(0.34473100304603577)),(to_sfixed_a(6.801368726883084e-05)),(to_sfixed_a(-0.026718901470303535)),(to_sfixed_a(0.00012306174903642386)),(to_sfixed_a(-0.0003769222821574658)),(to_sfixed_a(-0.007210109382867813)),(to_sfixed_a(6.617620965698734e-05)),(to_sfixed_a(-0.0014315956505015492)),(to_sfixed_a(-0.00407134834676981)),(to_sfixed_a(-2.545188181102276e-06)),(to_sfixed_a(-0.004557743202894926)),(to_sfixed_a(-0.0002406547573627904)),(to_sfixed_a(0.0002641181636136025)),(to_sfixed_a(-0.010509357787668705)),(to_sfixed_a(-0.005726469215005636)),(to_sfixed_a(0.0003103688941337168)),(to_sfixed_a(-0.00017189423670060933)),(to_sfixed_a(-0.0014033684274181724)),(to_sfixed_a(0.00023739035532344133)),(to_sfixed_a(-0.0002628379734233022)),(to_sfixed_a(-0.00015520758461207151)),(to_sfixed_a(0.024096740409731865)),(to_sfixed_a(7.155768980737776e-05)),(to_sfixed_a(-0.00926783587783575)),(to_sfixed_a(6.590570410480723e-05)),(to_sfixed_a(-1.5726778656244278e-05)),(to_sfixed_a(-9.529713861411437e-05)),(to_sfixed_a(-0.002002360997721553)),(to_sfixed_a(-0.0028556110337376595)),(to_sfixed_a(-0.0002642713370732963)),(to_sfixed_a(-5.8490019000601023e-05)),(to_sfixed_a(-5.471774784382433e-06)),(to_sfixed_a(3.84849299734924e-05)),(to_sfixed_a(-2.8591268346644938e-05)),(to_sfixed_a(-0.008263138122856617)),(to_sfixed_a(-0.0014866403071209788)),(to_sfixed_a(-0.002126738429069519)),(to_sfixed_a(-0.0021973310504108667)),(to_sfixed_a(0.00019588421855587512)),(to_sfixed_a(4.491943400353193e-06)),(to_sfixed_a(-0.00011289474787190557)),(to_sfixed_a(0.00035156181547790766)),(to_sfixed_a(-6.084734559408389e-05)),(to_sfixed_a(-0.00017900607781484723)),(to_sfixed_a(0.0005810749717056751)),(to_sfixed_a(-0.0005702708149328828)),(to_sfixed_a(6.288157601375133e-05)),(to_sfixed_a(0.0001285721082240343)),(to_sfixed_a(0.00010282621951773763)),(to_sfixed_a(-0.004750709980726242)),(to_sfixed_a(-0.000585462839808315)),(to_sfixed_a(2.2583299141842872e-05)),(to_sfixed_a(-0.000998787465505302)),(to_sfixed_a(-0.011806660331785679)),(to_sfixed_a(-0.00020194108947180212)),(to_sfixed_a(-1.1433439794927835e-07)),(to_sfixed_a(-0.0006407320033758879)),(to_sfixed_a(-0.06636574864387512)),(to_sfixed_a(-0.005180599633604288)));

    constant weight_n2_37 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.4300774335861206)),(to_sfixed_a(0.2714555263519287)),(to_sfixed_a(0.6456983685493469)),(to_sfixed_a(3.0120520023046993e-05)),(to_sfixed_a(0.0011979301925748587)),(to_sfixed_a(-0.0001549583103042096)),(to_sfixed_a(-0.0016639442183077335)),(to_sfixed_a(-0.00012596746091730893)),(to_sfixed_a(2.407748979749158e-05)),(to_sfixed_a(2.3399326892104e-05)),(to_sfixed_a(0.0004168543382547796)),(to_sfixed_a(0.001321951043792069)),(to_sfixed_a(0.002948251087218523)),(to_sfixed_a(0.0035614653024822474)),(to_sfixed_a(3.0621173209510744e-05)),(to_sfixed_a(5.792640149593353e-05)),(to_sfixed_a(-0.005183367989957333)),(to_sfixed_a(1.2695832992903888e-05)),(to_sfixed_a(0.31930312514305115)),(to_sfixed_a(-0.0011545747984200716)),(to_sfixed_a(5.563822924159467e-06)),(to_sfixed_a(-0.0002929636975750327)),(to_sfixed_a(0.28796035051345825)),(to_sfixed_a(0.0057478491216897964)),(to_sfixed_a(-0.0017476327484473586)),(to_sfixed_a(-0.005740202497690916)),(to_sfixed_a(-0.00018236304458696395)),(to_sfixed_a(-6.287058931775391e-05)),(to_sfixed_a(0.0034759510308504105)),(to_sfixed_a(0.0001909688435262069)),(to_sfixed_a(0.00027789187151938677)),(to_sfixed_a(0.00024276608019135892)),(to_sfixed_a(-0.0005443572881631553)),(to_sfixed_a(-4.298162821214646e-06)),(to_sfixed_a(-3.802882201853208e-05)),(to_sfixed_a(1.6002843040041625e-05)),(to_sfixed_a(-0.03564673289656639)),(to_sfixed_a(-0.01094555389136076)),(to_sfixed_a(-0.0023510304745286703)),(to_sfixed_a(-0.0002763835364021361)),(to_sfixed_a(-0.002769967308267951)),(to_sfixed_a(-0.0030715966131538153)),(to_sfixed_a(0.0003857543633785099)),(to_sfixed_a(-2.1681848011212423e-05)),(to_sfixed_a(-0.011808803305029869)),(to_sfixed_a(-0.0018924137111753225)),(to_sfixed_a(0.3533097803592682)),(to_sfixed_a(0.011840399354696274)),(to_sfixed_a(0.0002900488907471299)),(to_sfixed_a(0.024098515510559082)),(to_sfixed_a(0.25991082191467285)),(to_sfixed_a(-0.0021682926453649998)),(to_sfixed_a(-5.126887117512524e-06)),(to_sfixed_a(-0.003985448740422726)),(to_sfixed_a(-0.002954483265057206)),(to_sfixed_a(0.39127621054649353)),(to_sfixed_a(-7.745067705400288e-06)),(to_sfixed_a(-0.020330721512436867)),(to_sfixed_a(-2.0551466150209308e-05)),(to_sfixed_a(6.516333087347448e-05)),(to_sfixed_a(0.2064337432384491)),(to_sfixed_a(0.005226767156273127)),(to_sfixed_a(-0.00036967344931326807)),(to_sfixed_a(-0.004555533640086651)),(to_sfixed_a(9.919384319800884e-05)),(to_sfixed_a(-0.31231385469436646)),(to_sfixed_a(0.00015436136163771152)),(to_sfixed_a(0.000923962623346597)),(to_sfixed_a(-0.017751634120941162)),(to_sfixed_a(-5.722107016481459e-05)),(to_sfixed_a(-0.008691624738276005)),(to_sfixed_a(0.35930877923965454)),(to_sfixed_a(-0.07763175666332245)),(to_sfixed_a(0.00010048150579677895)),(to_sfixed_a(7.018737960606813e-05)),(to_sfixed_a(-0.00011069144966313615)),(to_sfixed_a(-0.001499050296843052)),(to_sfixed_a(-0.00019114218594040722)),(to_sfixed_a(-4.89373633172363e-07)),(to_sfixed_a(0.4654812514781952)),(to_sfixed_a(-1.4916415238985792e-05)),(to_sfixed_a(-2.8771602956112474e-05)),(to_sfixed_a(0.5902872085571289)),(to_sfixed_a(-0.026327870786190033)),(to_sfixed_a(-2.3711745598120615e-05)),(to_sfixed_a(0.0004709938366431743)),(to_sfixed_a(-0.02292606234550476)),(to_sfixed_a(0.212922140955925)),(to_sfixed_a(-3.0515333492076024e-05)),(to_sfixed_a(8.416057971771806e-05)),(to_sfixed_a(0.1635514348745346)),(to_sfixed_a(-6.444453174481168e-05)),(to_sfixed_a(0.0030872011557221413)),(to_sfixed_a(-0.00014625751646235585)),(to_sfixed_a(0.0025089436676353216)),(to_sfixed_a(7.36500951461494e-05)),(to_sfixed_a(-8.037820225581527e-05)),(to_sfixed_a(4.2194005800411105e-06)),(to_sfixed_a(-0.00013414121349342167)),(to_sfixed_a(0.0001305976911680773)),(to_sfixed_a(0.0008503644494339824)),(to_sfixed_a(0.000680965487845242)),(to_sfixed_a(4.761442687595263e-05)),(to_sfixed_a(-0.0004890080308541656)),(to_sfixed_a(-0.009536805562675)),(to_sfixed_a(0.2646929621696472)),(to_sfixed_a(-3.682188980747014e-05)),(to_sfixed_a(5.5352156778099015e-05)),(to_sfixed_a(7.371265382971615e-05)),(to_sfixed_a(-0.377773255109787)),(to_sfixed_a(-0.004092112183570862)),(to_sfixed_a(-0.00028864271007478237)),(to_sfixed_a(0.08049057424068451)),(to_sfixed_a(-8.920126856537536e-05)),(to_sfixed_a(-0.00012056517880409956)),(to_sfixed_a(-0.41400036215782166)),(to_sfixed_a(1.256416999240173e-05)),(to_sfixed_a(1.842066558310762e-05)),(to_sfixed_a(-2.8825204935856164e-05)),(to_sfixed_a(0.002315336372703314)),(to_sfixed_a(0.0001673004444455728)),(to_sfixed_a(2.1247324184514582e-06)),(to_sfixed_a(0.004642239771783352)),(to_sfixed_a(5.009874075767584e-05)),(to_sfixed_a(-0.00011612437083385885)),(to_sfixed_a(-0.001971043646335602)),(to_sfixed_a(-0.010990236885845661)),(to_sfixed_a(2.6861802325583994e-05)),(to_sfixed_a(1.6179466911125928e-05)),(to_sfixed_a(-0.00015701338998042047)),(to_sfixed_a(-0.00018985643691848963)),(to_sfixed_a(2.366798435105011e-05)),(to_sfixed_a(-0.08371812850236893)),(to_sfixed_a(-0.44683605432510376)),(to_sfixed_a(-0.0001861228229245171)),(to_sfixed_a(-0.00016431554104201496)),(to_sfixed_a(0.333806574344635)),(to_sfixed_a(0.000221459791646339)),(to_sfixed_a(-2.337361001991667e-05)),(to_sfixed_a(0.00011358755000401288)),(to_sfixed_a(8.62830420373939e-05)),(to_sfixed_a(8.00159978098236e-05)),(to_sfixed_a(1.7986822058446705e-06)),(to_sfixed_a(-0.00023216484987642616)),(to_sfixed_a(-0.003024583449587226)),(to_sfixed_a(-1.4980801097408403e-05)),(to_sfixed_a(-0.00026432800223119557)),(to_sfixed_a(-2.1285814000293612e-07)),(to_sfixed_a(-0.00011723465286195278)),(to_sfixed_a(-0.012168453074991703)),(to_sfixed_a(0.00022950168931856751)),(to_sfixed_a(7.084882236085832e-05)),(to_sfixed_a(0.0010263314470648766)),(to_sfixed_a(0.00017562380526214838)),(to_sfixed_a(5.099544068798423e-06)),(to_sfixed_a(-0.01012637559324503)),(to_sfixed_a(-9.066786151379347e-05)),(to_sfixed_a(0.0006083886255510151)),(to_sfixed_a(-0.00012891803635284305)),(to_sfixed_a(3.6889934563077986e-05)),(to_sfixed_a(-1.0770450899144635e-05)),(to_sfixed_a(-0.0001574328780407086)),(to_sfixed_a(0.058615267276763916)),(to_sfixed_a(-0.4822750389575958)),(to_sfixed_a(-0.13108043372631073)),(to_sfixed_a(-0.0011281260522082448)),(to_sfixed_a(-2.459943061694503e-06)),(to_sfixed_a(-0.00018625067605171353)),(to_sfixed_a(-9.868534107226878e-05)),(to_sfixed_a(-2.561474684625864e-05)),(to_sfixed_a(0.04819127544760704)),(to_sfixed_a(-0.005951764993369579)),(to_sfixed_a(-0.008147102780640125)),(to_sfixed_a(5.466485163196921e-06)),(to_sfixed_a(0.10677406936883926)),(to_sfixed_a(-0.004650570452213287)),(to_sfixed_a(-0.0027766365092247725)),(to_sfixed_a(-0.0006445186445489526)),(to_sfixed_a(0.2406671643257141)),(to_sfixed_a(0.011637572199106216)),(to_sfixed_a(0.0017953976057469845)),(to_sfixed_a(-0.3605160415172577)),(to_sfixed_a(4.73293403047137e-06)),(to_sfixed_a(-0.0001541180827189237)),(to_sfixed_a(-2.499337642802857e-05)),(to_sfixed_a(0.00048542366130277514)),(to_sfixed_a(-0.002766849473118782)),(to_sfixed_a(0.0018842784920707345)),(to_sfixed_a(0.00016648965538479388)),(to_sfixed_a(-0.006325291004031897)),(to_sfixed_a(-0.007545127999037504)),(to_sfixed_a(-5.610709195025265e-06)),(to_sfixed_a(0.009123511612415314)),(to_sfixed_a(0.0005824110121466219)),(to_sfixed_a(-0.00010298617416992784)),(to_sfixed_a(0.002170444931834936)),(to_sfixed_a(-0.00012844322191085666)),(to_sfixed_a(-0.006815331522375345)),(to_sfixed_a(0.0007428221288137138)),(to_sfixed_a(6.800542905693874e-06)),(to_sfixed_a(-3.9540896977996454e-05)),(to_sfixed_a(4.796303255716339e-05)),(to_sfixed_a(-8.241311297751963e-05)),(to_sfixed_a(-7.041175558697432e-05)),(to_sfixed_a(-0.0002479851245880127)),(to_sfixed_a(-0.0043524145148694515)),(to_sfixed_a(0.000464390468550846)),(to_sfixed_a(-0.19128753244876862)),(to_sfixed_a(0.015430830419063568)),(to_sfixed_a(0.5267689824104309)),(to_sfixed_a(0.4300582706928253)),(to_sfixed_a(5.26912699569948e-05)),(to_sfixed_a(-0.000251411838689819)),(to_sfixed_a(2.7481413781060837e-05)),(to_sfixed_a(0.0001922696828842163)),(to_sfixed_a(-0.00028713318170048296)),(to_sfixed_a(0.020393865182995796)),(to_sfixed_a(-0.00045481076813302934)),(to_sfixed_a(0.43504923582077026)),(to_sfixed_a(-6.707098509650677e-05)),(to_sfixed_a(-0.00013687281170859933)),(to_sfixed_a(-0.00014961979468353093)),(to_sfixed_a(0.00022071501007303596)),(to_sfixed_a(-0.3010515868663788)),(to_sfixed_a(0.005745226982980967)),(to_sfixed_a(-1.083856841432862e-05)),(to_sfixed_a(1.0050716809928417e-06)),(to_sfixed_a(-0.00022740807617083192)),(to_sfixed_a(0.10758522897958755)),(to_sfixed_a(0.029940078034996986)),(to_sfixed_a(0.36294665932655334)),(to_sfixed_a(1.7786202079150826e-05)),(to_sfixed_a(0.0001400660548824817)),(to_sfixed_a(4.446343518793583e-05)),(to_sfixed_a(0.0030676056630909443)),(to_sfixed_a(-0.0005219197482801974)),(to_sfixed_a(0.06265446543693542)),(to_sfixed_a(-1.301168231293559e-05)),(to_sfixed_a(-0.003306630300357938)),(to_sfixed_a(7.877872849348933e-05)),(to_sfixed_a(-0.46555018424987793)),(to_sfixed_a(0.0002469325845595449)),(to_sfixed_a(0.20703773200511932)),(to_sfixed_a(-0.0003104470088146627)),(to_sfixed_a(-0.3231271505355835)),(to_sfixed_a(-0.00016017364396248013)),(to_sfixed_a(0.00989573448896408)),(to_sfixed_a(-0.007143126334995031)),(to_sfixed_a(-0.00011336391617078334)),(to_sfixed_a(-0.0012897063279524446)),(to_sfixed_a(0.0026370128616690636)),(to_sfixed_a(-0.00014974338409956545)),(to_sfixed_a(0.0030182041227817535)),(to_sfixed_a(5.7142060541082174e-05)),(to_sfixed_a(0.00015113492554519325)),(to_sfixed_a(0.008075564168393612)),(to_sfixed_a(0.020222438499331474)),(to_sfixed_a(-0.00029760421602986753)),(to_sfixed_a(3.0374492780538276e-05)),(to_sfixed_a(0.004994897171854973)),(to_sfixed_a(-0.00010733550880104303)),(to_sfixed_a(0.4606230854988098)),(to_sfixed_a(-0.0002477039524819702)),(to_sfixed_a(0.001287365099415183)),(to_sfixed_a(-4.364044070825912e-05)),(to_sfixed_a(-0.2970168888568878)),(to_sfixed_a(-0.00023739731113892049)),(to_sfixed_a(-7.822319457773119e-05)),(to_sfixed_a(0.0001799896126613021)),(to_sfixed_a(-0.003911698702722788)),(to_sfixed_a(-0.43949902057647705)),(to_sfixed_a(-1.9086073734797537e-05)),(to_sfixed_a(0.00011908862506970763)),(to_sfixed_a(-0.00017157295951619744)),(to_sfixed_a(9.052831592271104e-05)),(to_sfixed_a(0.0019318313570693135)),(to_sfixed_a(-0.007691392675042152)),(to_sfixed_a(0.41774114966392517)),(to_sfixed_a(-0.15843303501605988)),(to_sfixed_a(0.234071746468544)),(to_sfixed_a(-0.00011646159691736102)),(to_sfixed_a(8.487331797368824e-05)),(to_sfixed_a(-0.00016881147166714072)),(to_sfixed_a(-0.0020884349942207336)),(to_sfixed_a(0.0002876659273169935)),(to_sfixed_a(8.897575753508136e-05)),(to_sfixed_a(0.5090522170066833)),(to_sfixed_a(0.020734932273626328)),(to_sfixed_a(-0.00011534743680385873)),(to_sfixed_a(-0.018004879355430603)),(to_sfixed_a(-0.4655189514160156)),(to_sfixed_a(-0.2564712166786194)),(to_sfixed_a(-0.016121545806527138)),(to_sfixed_a(2.3801338102202863e-05)),(to_sfixed_a(0.18957637250423431)),(to_sfixed_a(-0.1555054932832718)),(to_sfixed_a(0.0020483240950852633)),(to_sfixed_a(-0.00010411784023744985)),(to_sfixed_a(0.005210563074797392)),(to_sfixed_a(-0.006608407478779554)),(to_sfixed_a(-0.004320124164223671)));

    constant weight_n2_38 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.1781398355960846)),(to_sfixed_a(1.713747769827023e-05)),(to_sfixed_a(1.6863159544300288e-05)),(to_sfixed_a(0.0002367128327023238)),(to_sfixed_a(0.018234234303236008)),(to_sfixed_a(0.00011508471652632579)),(to_sfixed_a(0.003230961738154292)),(to_sfixed_a(8.463526319246739e-05)),(to_sfixed_a(-1.3364915503188968e-06)),(to_sfixed_a(-7.138607907108963e-05)),(to_sfixed_a(0.00011744527000701055)),(to_sfixed_a(-0.37713342905044556)),(to_sfixed_a(-0.3048027455806732)),(to_sfixed_a(-0.0020329931285232306)),(to_sfixed_a(1.8676902982406318e-05)),(to_sfixed_a(-0.00014824273239355534)),(to_sfixed_a(-0.001671729376539588)),(to_sfixed_a(0.00017400839715264738)),(to_sfixed_a(0.0016739551210775971)),(to_sfixed_a(-0.012776629067957401)),(to_sfixed_a(3.371023922227323e-06)),(to_sfixed_a(0.00011664346675388515)),(to_sfixed_a(-0.000149845756823197)),(to_sfixed_a(-0.0019802337046712637)),(to_sfixed_a(0.004883176647126675)),(to_sfixed_a(0.000753612257540226)),(to_sfixed_a(-7.054393063299358e-05)),(to_sfixed_a(-0.00023180486459750682)),(to_sfixed_a(-0.0004157398361712694)),(to_sfixed_a(-0.00020627265621442348)),(to_sfixed_a(0.2750088572502136)),(to_sfixed_a(-0.0003811113128904253)),(to_sfixed_a(-0.002620919141918421)),(to_sfixed_a(-2.349919668631628e-05)),(to_sfixed_a(6.252258026506752e-05)),(to_sfixed_a(-2.936893724836409e-05)),(to_sfixed_a(0.005355400964617729)),(to_sfixed_a(0.0005597359267994761)),(to_sfixed_a(0.005267810076475143)),(to_sfixed_a(-0.00015026688924990594)),(to_sfixed_a(-0.0033509009517729282)),(to_sfixed_a(0.0005071828491054475)),(to_sfixed_a(0.00011196772538824007)),(to_sfixed_a(-7.51427432987839e-06)),(to_sfixed_a(-0.0001099661021726206)),(to_sfixed_a(9.700434020487592e-06)),(to_sfixed_a(0.00769858667626977)),(to_sfixed_a(7.030311098787934e-05)),(to_sfixed_a(0.00024786824360489845)),(to_sfixed_a(0.0065429736860096455)),(to_sfixed_a(-4.4600303226616234e-05)),(to_sfixed_a(-0.00032404903322458267)),(to_sfixed_a(0.00029892774182371795)),(to_sfixed_a(0.006019468419253826)),(to_sfixed_a(0.015321783721446991)),(to_sfixed_a(0.005816182121634483)),(to_sfixed_a(-4.186402657069266e-05)),(to_sfixed_a(-0.003854342270642519)),(to_sfixed_a(6.280493835220113e-05)),(to_sfixed_a(0.00023703202896285802)),(to_sfixed_a(0.0019516292959451675)),(to_sfixed_a(-0.0030842358246445656)),(to_sfixed_a(0.0004492498410400003)),(to_sfixed_a(0.0015790063189342618)),(to_sfixed_a(-0.00038045382825657725)),(to_sfixed_a(-0.3415650725364685)),(to_sfixed_a(0.00023236875131260604)),(to_sfixed_a(0.002097601071000099)),(to_sfixed_a(0.005089850164949894)),(to_sfixed_a(-2.99902749247849e-05)),(to_sfixed_a(-0.011129157617688179)),(to_sfixed_a(0.008258731104433537)),(to_sfixed_a(-0.0015350159956142306)),(to_sfixed_a(-7.143742550397292e-05)),(to_sfixed_a(-6.519598537124693e-05)),(to_sfixed_a(7.100557559169829e-05)),(to_sfixed_a(-0.0021383839193731546)),(to_sfixed_a(0.0038655735552310944)),(to_sfixed_a(0.00012902509479317814)),(to_sfixed_a(-0.00282505271025002)),(to_sfixed_a(-0.0014450044836848974)),(to_sfixed_a(3.74760857084766e-05)),(to_sfixed_a(0.002625963417813182)),(to_sfixed_a(-0.004061995539814234)),(to_sfixed_a(0.00010603276314213872)),(to_sfixed_a(4.633411663235165e-06)),(to_sfixed_a(0.3324185013771057)),(to_sfixed_a(-0.0001691188372205943)),(to_sfixed_a(0.00014910723257344216)),(to_sfixed_a(1.3861754268873483e-06)),(to_sfixed_a(0.0008638645522296429)),(to_sfixed_a(0.0002504950971342623)),(to_sfixed_a(2.9578946850961074e-05)),(to_sfixed_a(-0.0001746740599628538)),(to_sfixed_a(-0.23724175989627838)),(to_sfixed_a(4.554905171971768e-05)),(to_sfixed_a(5.6949382269522175e-05)),(to_sfixed_a(7.442155038006604e-06)),(to_sfixed_a(2.5104642190854065e-05)),(to_sfixed_a(7.540928345406428e-05)),(to_sfixed_a(7.014930815785192e-06)),(to_sfixed_a(0.20755718648433685)),(to_sfixed_a(-0.0004562248068396002)),(to_sfixed_a(-0.0006594897713512182)),(to_sfixed_a(-0.14052517712116241)),(to_sfixed_a(0.32215607166290283)),(to_sfixed_a(0.00029650077340193093)),(to_sfixed_a(4.991452078684233e-05)),(to_sfixed_a(1.4672306861029938e-05)),(to_sfixed_a(1.3113008208165411e-05)),(to_sfixed_a(-0.014321364462375641)),(to_sfixed_a(-9.07313878997229e-05)),(to_sfixed_a(-0.0010396289872005582)),(to_sfixed_a(-0.00011477935913717374)),(to_sfixed_a(6.547091470565647e-05)),(to_sfixed_a(0.005346772260963917)),(to_sfixed_a(-0.0019127210834994912)),(to_sfixed_a(2.657311961229425e-05)),(to_sfixed_a(-0.0001815737341530621)),(to_sfixed_a(-0.03808758035302162)),(to_sfixed_a(-2.2425752831622958e-05)),(to_sfixed_a(-0.00015602284111082554)),(to_sfixed_a(-9.161502384813502e-05)),(to_sfixed_a(-6.814644439145923e-05)),(to_sfixed_a(2.4633336579427123e-06)),(to_sfixed_a(0.003958491142839193)),(to_sfixed_a(0.18906502425670624)),(to_sfixed_a(0.0002656698925420642)),(to_sfixed_a(-0.00015174326836131513)),(to_sfixed_a(0.0001713037199806422)),(to_sfixed_a(0.00013021804625168443)),(to_sfixed_a(-4.2776398913701996e-05)),(to_sfixed_a(8.176897244993597e-05)),(to_sfixed_a(-0.0035078043583780527)),(to_sfixed_a(0.00027658656472340226)),(to_sfixed_a(5.95218880334869e-05)),(to_sfixed_a(-0.00022062522475607693)),(to_sfixed_a(-0.0005804160609841347)),(to_sfixed_a(-0.00013817033322993666)),(to_sfixed_a(-0.00021000606648158282)),(to_sfixed_a(7.535869372077286e-06)),(to_sfixed_a(-6.885033508297056e-05)),(to_sfixed_a(-0.00013548573770094663)),(to_sfixed_a(-0.00010816360008902848)),(to_sfixed_a(-0.0009761433466337621)),(to_sfixed_a(3.242859020247124e-05)),(to_sfixed_a(0.003987930715084076)),(to_sfixed_a(5.984197196085006e-05)),(to_sfixed_a(-2.4456185201415792e-05)),(to_sfixed_a(0.001005574595183134)),(to_sfixed_a(7.791537791490555e-05)),(to_sfixed_a(-0.0002250336983706802)),(to_sfixed_a(-2.9810695195919834e-05)),(to_sfixed_a(4.812339102500118e-05)),(to_sfixed_a(0.00010566302808001637)),(to_sfixed_a(-0.5181431770324707)),(to_sfixed_a(-0.0001466039102524519)),(to_sfixed_a(0.07921624183654785)),(to_sfixed_a(0.0001158844243036583)),(to_sfixed_a(1.42212666105479e-05)),(to_sfixed_a(0.0002459872339386493)),(to_sfixed_a(0.00011391800944693387)),(to_sfixed_a(-0.001193301985040307)),(to_sfixed_a(-0.25302374362945557)),(to_sfixed_a(0.0001275045215152204)),(to_sfixed_a(-0.0012899964349344373)),(to_sfixed_a(-6.203946395544335e-05)),(to_sfixed_a(0.005656267981976271)),(to_sfixed_a(-6.299332017078996e-05)),(to_sfixed_a(0.00015492053353227675)),(to_sfixed_a(0.001684349263086915)),(to_sfixed_a(-0.0006298889056779444)),(to_sfixed_a(-0.00020591498469002545)),(to_sfixed_a(7.124459079932421e-05)),(to_sfixed_a(0.2694460451602936)),(to_sfixed_a(0.00010264747106702998)),(to_sfixed_a(-0.0042920405976474285)),(to_sfixed_a(0.282401442527771)),(to_sfixed_a(-0.007509391754865646)),(to_sfixed_a(0.009511704556643963)),(to_sfixed_a(-0.0007046814425848424)),(to_sfixed_a(-0.004402628634124994)),(to_sfixed_a(0.00021826440934091806)),(to_sfixed_a(-0.00038350227987393737)),(to_sfixed_a(6.499965093098581e-05)),(to_sfixed_a(-2.9634175007231534e-05)),(to_sfixed_a(-0.0017057334771379828)),(to_sfixed_a(-0.14286409318447113)),(to_sfixed_a(-0.0019410636741667986)),(to_sfixed_a(-0.0001015214147628285)),(to_sfixed_a(-0.01843622326850891)),(to_sfixed_a(-0.00013420106552075595)),(to_sfixed_a(0.009047073312103748)),(to_sfixed_a(-2.510075137251988e-05)),(to_sfixed_a(0.0001998770167119801)),(to_sfixed_a(0.00013427971862256527)),(to_sfixed_a(0.00010208429011981934)),(to_sfixed_a(0.0037588211707770824)),(to_sfixed_a(0.0011981530115008354)),(to_sfixed_a(9.709208097774535e-05)),(to_sfixed_a(8.426250133197755e-07)),(to_sfixed_a(-1.5757577784825116e-05)),(to_sfixed_a(0.00018317594367545098)),(to_sfixed_a(6.678529462078586e-05)),(to_sfixed_a(2.260148903587833e-05)),(to_sfixed_a(0.0024928986094892025)),(to_sfixed_a(-0.005489910487085581)),(to_sfixed_a(-0.010052917525172234)),(to_sfixed_a(0.5278164148330688)),(to_sfixed_a(0.007833583280444145)),(to_sfixed_a(-0.004597322084009647)),(to_sfixed_a(-6.818550173193216e-05)),(to_sfixed_a(0.00011330722190905362)),(to_sfixed_a(0.00040786451427266)),(to_sfixed_a(-0.00013318966375663877)),(to_sfixed_a(-3.613336230046116e-05)),(to_sfixed_a(0.3782392144203186)),(to_sfixed_a(0.0007217573584057391)),(to_sfixed_a(0.3634849786758423)),(to_sfixed_a(-6.394074443960562e-05)),(to_sfixed_a(-0.00018026636098511517)),(to_sfixed_a(-0.00016328232595697045)),(to_sfixed_a(0.00016723650333005935)),(to_sfixed_a(-4.241627175360918e-05)),(to_sfixed_a(0.006382550112903118)),(to_sfixed_a(-3.729266609298065e-05)),(to_sfixed_a(2.1531013771891594e-07)),(to_sfixed_a(6.434252281906083e-05)),(to_sfixed_a(-0.29757413268089294)),(to_sfixed_a(0.010416333563625813)),(to_sfixed_a(0.0070745921693742275)),(to_sfixed_a(-2.2395906853489578e-06)),(to_sfixed_a(8.210126543417573e-05)),(to_sfixed_a(2.8555135941132903e-05)),(to_sfixed_a(1.398947188135935e-05)),(to_sfixed_a(0.0003823611477855593)),(to_sfixed_a(-0.0112895667552948)),(to_sfixed_a(-5.351787694962695e-05)),(to_sfixed_a(0.00015846738824620843)),(to_sfixed_a(0.0001774767297320068)),(to_sfixed_a(0.002471545012667775)),(to_sfixed_a(8.509154577041045e-05)),(to_sfixed_a(0.01044990960508585)),(to_sfixed_a(1.7405080143362284e-05)),(to_sfixed_a(-0.1932229846715927)),(to_sfixed_a(0.00012091945973224938)),(to_sfixed_a(-0.0015795259969308972)),(to_sfixed_a(-0.007987004704773426)),(to_sfixed_a(0.0001541036181151867)),(to_sfixed_a(-0.000407595798606053)),(to_sfixed_a(0.0003476917336229235)),(to_sfixed_a(8.238033478846774e-05)),(to_sfixed_a(-0.00259456317871809)),(to_sfixed_a(2.0206760382279754e-05)),(to_sfixed_a(-0.0002788773854263127)),(to_sfixed_a(0.014509356580674648)),(to_sfixed_a(-0.009522095322608948)),(to_sfixed_a(6.284627306740731e-05)),(to_sfixed_a(6.046375347068533e-05)),(to_sfixed_a(0.0029579754918813705)),(to_sfixed_a(7.694079249631613e-05)),(to_sfixed_a(-2.2091990103945136e-05)),(to_sfixed_a(-0.0001679171109572053)),(to_sfixed_a(-2.7428981411503628e-05)),(to_sfixed_a(-6.426544860005379e-05)),(to_sfixed_a(-0.20254218578338623)),(to_sfixed_a(6.721507816109806e-05)),(to_sfixed_a(-1.4944256690796465e-05)),(to_sfixed_a(-6.912842945894226e-05)),(to_sfixed_a(-0.0012235520407557487)),(to_sfixed_a(0.0028428679797798395)),(to_sfixed_a(1.912413426907733e-05)),(to_sfixed_a(6.109301466494799e-05)),(to_sfixed_a(0.00017506364383734763)),(to_sfixed_a(2.5054821890080348e-05)),(to_sfixed_a(0.008005807176232338)),(to_sfixed_a(0.011051397770643234)),(to_sfixed_a(0.3623215854167938)),(to_sfixed_a(0.006233472377061844)),(to_sfixed_a(-0.0016910219565033913)),(to_sfixed_a(-6.225726247066632e-05)),(to_sfixed_a(-0.00011663397162919864)),(to_sfixed_a(1.087944838218391e-06)),(to_sfixed_a(-0.011195109225809574)),(to_sfixed_a(0.00028932123677805066)),(to_sfixed_a(0.00010454747098265216)),(to_sfixed_a(-0.002674769377335906)),(to_sfixed_a(0.01014622300863266)),(to_sfixed_a(0.0001561274257255718)),(to_sfixed_a(-0.0015346209984272718)),(to_sfixed_a(-0.00031975164893083274)),(to_sfixed_a(-2.985825267387554e-05)),(to_sfixed_a(-0.2541644275188446)),(to_sfixed_a(-7.3920091381296515e-06)),(to_sfixed_a(0.0037798876874148846)),(to_sfixed_a(-4.0476017602486536e-05)),(to_sfixed_a(0.004680941812694073)),(to_sfixed_a(6.843649316579103e-05)),(to_sfixed_a(-0.0018935399129986763)),(to_sfixed_a(0.37994763255119324)),(to_sfixed_a(-1.741166488500312e-05)));

    constant weight_n2_39 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.22061628103256226)),(to_sfixed_a(0.19922266900539398)),(to_sfixed_a(-0.005033341236412525)),(to_sfixed_a(0.00023861072259023786)),(to_sfixed_a(-0.0015905607724562287)),(to_sfixed_a(0.0001440891355741769)),(to_sfixed_a(0.00041274455725215375)),(to_sfixed_a(-0.00021607826056424528)),(to_sfixed_a(-0.00015903692110441625)),(to_sfixed_a(-7.073479355312884e-05)),(to_sfixed_a(5.762238288298249e-05)),(to_sfixed_a(-0.0014570173807442188)),(to_sfixed_a(-0.0020289693493396044)),(to_sfixed_a(0.001998616149649024)),(to_sfixed_a(6.808572652516887e-05)),(to_sfixed_a(-5.797675112262368e-05)),(to_sfixed_a(-0.003210916416719556)),(to_sfixed_a(0.00015538626757916063)),(to_sfixed_a(-0.003630709368735552)),(to_sfixed_a(-0.006580887828022242)),(to_sfixed_a(6.343192944768816e-05)),(to_sfixed_a(-0.00015263458772096783)),(to_sfixed_a(3.874862159136683e-06)),(to_sfixed_a(0.21491557359695435)),(to_sfixed_a(-0.012486716732382774)),(to_sfixed_a(-0.0022430524695664644)),(to_sfixed_a(-8.2326507254038e-05)),(to_sfixed_a(0.0008840416558086872)),(to_sfixed_a(0.00011462887050583959)),(to_sfixed_a(6.549173849634826e-05)),(to_sfixed_a(0.02575128898024559)),(to_sfixed_a(6.678144563920796e-05)),(to_sfixed_a(0.009679693728685379)),(to_sfixed_a(9.233626769855618e-07)),(to_sfixed_a(0.0002811639569699764)),(to_sfixed_a(-4.5697179302806035e-05)),(to_sfixed_a(0.07892977446317673)),(to_sfixed_a(0.13906794786453247)),(to_sfixed_a(-0.04427460581064224)),(to_sfixed_a(-7.215669029392302e-06)),(to_sfixed_a(-0.29582974314689636)),(to_sfixed_a(-0.0009147184318862855)),(to_sfixed_a(5.903515557292849e-06)),(to_sfixed_a(-2.2367836209014058e-05)),(to_sfixed_a(0.00034630493610166013)),(to_sfixed_a(0.08833082765340805)),(to_sfixed_a(0.6035212278366089)),(to_sfixed_a(0.0011222029570490122)),(to_sfixed_a(-5.1455426728352904e-06)),(to_sfixed_a(0.002037087455391884)),(to_sfixed_a(-0.0045496211387217045)),(to_sfixed_a(-0.004655422177165747)),(to_sfixed_a(0.00010145437408937141)),(to_sfixed_a(-0.005423216614872217)),(to_sfixed_a(0.4907894730567932)),(to_sfixed_a(-0.05108022689819336)),(to_sfixed_a(-5.212277756072581e-07)),(to_sfixed_a(-0.005104289390146732)),(to_sfixed_a(0.0001160573010565713)),(to_sfixed_a(-0.00014547663158737123)),(to_sfixed_a(-0.00010993797332048416)),(to_sfixed_a(-0.002560919849202037)),(to_sfixed_a(0.002801071386784315)),(to_sfixed_a(0.008344834670424461)),(to_sfixed_a(3.9405473216902465e-05)),(to_sfixed_a(-0.5317007303237915)),(to_sfixed_a(4.963501851307228e-06)),(to_sfixed_a(0.4123334288597107)),(to_sfixed_a(-0.00010204499994870275)),(to_sfixed_a(-0.00010734271199908108)),(to_sfixed_a(-0.016894111409783363)),(to_sfixed_a(-0.006435609422624111)),(to_sfixed_a(-0.0015731947496533394)),(to_sfixed_a(-4.689085471909493e-05)),(to_sfixed_a(0.00020129079348407686)),(to_sfixed_a(-8.085524314083159e-06)),(to_sfixed_a(0.012401006184518337)),(to_sfixed_a(0.004380403086543083)),(to_sfixed_a(-0.0002475123037584126)),(to_sfixed_a(-0.0065841348841786385)),(to_sfixed_a(-0.0012371196644380689)),(to_sfixed_a(9.806311572901905e-05)),(to_sfixed_a(0.7140712141990662)),(to_sfixed_a(-0.005434155929833651)),(to_sfixed_a(0.00010687584290280938)),(to_sfixed_a(0.0008012035395950079)),(to_sfixed_a(0.03111514262855053)),(to_sfixed_a(-0.00014795918832533062)),(to_sfixed_a(7.228566391859204e-05)),(to_sfixed_a(-0.00011335244926158339)),(to_sfixed_a(-0.046672217547893524)),(to_sfixed_a(8.381630323128775e-05)),(to_sfixed_a(0.0003741762484423816)),(to_sfixed_a(-5.883842095499858e-05)),(to_sfixed_a(-0.00025253425701521337)),(to_sfixed_a(-2.654749187058769e-05)),(to_sfixed_a(-7.89841142250225e-05)),(to_sfixed_a(-1.3880198821425438e-06)),(to_sfixed_a(5.129895725985989e-07)),(to_sfixed_a(-0.00016569928266108036)),(to_sfixed_a(0.003954938612878323)),(to_sfixed_a(0.015673719346523285)),(to_sfixed_a(-3.574256334104575e-05)),(to_sfixed_a(-0.0020841544028371572)),(to_sfixed_a(0.0047883037477731705)),(to_sfixed_a(2.6666316443879623e-06)),(to_sfixed_a(0.00011205723421880975)),(to_sfixed_a(-6.963792111491784e-05)),(to_sfixed_a(4.501669536693953e-05)),(to_sfixed_a(-0.15665611624717712)),(to_sfixed_a(0.003302130149677396)),(to_sfixed_a(0.00011319720942992717)),(to_sfixed_a(-3.1486593798035756e-05)),(to_sfixed_a(8.010231249500066e-05)),(to_sfixed_a(-3.672088496387005e-06)),(to_sfixed_a(0.017666950821876526)),(to_sfixed_a(0.013764199800789356)),(to_sfixed_a(-0.00033412239281460643)),(to_sfixed_a(0.00015187029202934355)),(to_sfixed_a(-0.0006865494651719928)),(to_sfixed_a(1.0810868843691424e-05)),(to_sfixed_a(-0.00016676384257152677)),(to_sfixed_a(-0.00014876331260893494)),(to_sfixed_a(-0.00010668054164852947)),(to_sfixed_a(0.00010815532732522115)),(to_sfixed_a(-0.30016759037971497)),(to_sfixed_a(-0.005395551212131977)),(to_sfixed_a(0.00011638939758995548)),(to_sfixed_a(-0.0001296143454965204)),(to_sfixed_a(-0.00024743066751398146)),(to_sfixed_a(-3.1211522582452744e-05)),(to_sfixed_a(2.3235454136738554e-05)),(to_sfixed_a(-0.004324049223214388)),(to_sfixed_a(0.012354038655757904)),(to_sfixed_a(8.904952846933156e-05)),(to_sfixed_a(-2.9341812478378415e-05)),(to_sfixed_a(-0.3573648929595947)),(to_sfixed_a(-0.0006718853837810457)),(to_sfixed_a(0.0001438572653569281)),(to_sfixed_a(9.115582361118868e-05)),(to_sfixed_a(-4.677328252000734e-05)),(to_sfixed_a(7.506777183152735e-05)),(to_sfixed_a(-0.00042041816050186753)),(to_sfixed_a(-0.00030351357418112457)),(to_sfixed_a(-0.002663067076355219)),(to_sfixed_a(-0.00010109047434525564)),(to_sfixed_a(0.0013377359136939049)),(to_sfixed_a(-5.730174598284066e-05)),(to_sfixed_a(-0.0001664673036430031)),(to_sfixed_a(-0.0175054632127285)),(to_sfixed_a(-9.777760715223849e-05)),(to_sfixed_a(-8.488568710163236e-05)),(to_sfixed_a(0.006024069618433714)),(to_sfixed_a(0.00014315186126623303)),(to_sfixed_a(0.00011627688945736736)),(to_sfixed_a(0.015954365953803062)),(to_sfixed_a(1.9408364096307196e-05)),(to_sfixed_a(-0.0016391170211136341)),(to_sfixed_a(-0.00011736652231775224)),(to_sfixed_a(8.969110785983503e-05)),(to_sfixed_a(-0.00013085879618301988)),(to_sfixed_a(-1.0603165719658136e-05)),(to_sfixed_a(0.20659559965133667)),(to_sfixed_a(-0.004443921614438295)),(to_sfixed_a(9.018426499096677e-05)),(to_sfixed_a(-0.009470629505813122)),(to_sfixed_a(0.00010665693844202906)),(to_sfixed_a(0.003738190745934844)),(to_sfixed_a(0.0001082454837160185)),(to_sfixed_a(7.64656942919828e-05)),(to_sfixed_a(-0.004730915650725365)),(to_sfixed_a(-0.00607420364394784)),(to_sfixed_a(-0.004505305550992489)),(to_sfixed_a(0.0002518154797144234)),(to_sfixed_a(0.0014221828896552324)),(to_sfixed_a(-0.0008404154796153307)),(to_sfixed_a(-0.00036217260640114546)),(to_sfixed_a(0.2663962244987488)),(to_sfixed_a(-0.013333657756447792)),(to_sfixed_a(-0.44574761390686035)),(to_sfixed_a(-0.0012389017501845956)),(to_sfixed_a(-0.0025504152290523052)),(to_sfixed_a(-0.00019384526240173727)),(to_sfixed_a(6.10788119956851e-05)),(to_sfixed_a(-6.475578993558884e-05)),(to_sfixed_a(-7.834312418708578e-05)),(to_sfixed_a(-0.007156213745474815)),(to_sfixed_a(0.00132526527158916)),(to_sfixed_a(-0.004728080239146948)),(to_sfixed_a(-0.004059045575559139)),(to_sfixed_a(0.0043619475327432156)),(to_sfixed_a(3.6223780625732616e-05)),(to_sfixed_a(0.015912100672721863)),(to_sfixed_a(0.0016427116934210062)),(to_sfixed_a(0.00024585306528024375)),(to_sfixed_a(-0.24909371137619019)),(to_sfixed_a(0.00023725286882836372)),(to_sfixed_a(0.14074119925498962)),(to_sfixed_a(-0.002680707722902298)),(to_sfixed_a(0.000302967062452808)),(to_sfixed_a(5.71694690734148e-05)),(to_sfixed_a(-0.00010337230924051255)),(to_sfixed_a(-1.772039831848815e-05)),(to_sfixed_a(0.00010353900142945349)),(to_sfixed_a(0.00011990245548076928)),(to_sfixed_a(-0.0012903724564239383)),(to_sfixed_a(-0.003758067265152931)),(to_sfixed_a(-0.12996257841587067)),(to_sfixed_a(0.019016282632946968)),(to_sfixed_a(-0.004924679175019264)),(to_sfixed_a(0.17188963294029236)),(to_sfixed_a(-6.63165919831954e-05)),(to_sfixed_a(0.00015344578423537314)),(to_sfixed_a(7.60457623982802e-07)),(to_sfixed_a(-0.00015086746134329587)),(to_sfixed_a(-2.477153975632973e-05)),(to_sfixed_a(-0.00042621471220627427)),(to_sfixed_a(0.003471862291917205)),(to_sfixed_a(-0.05418219044804573)),(to_sfixed_a(1.703319685475435e-05)),(to_sfixed_a(-0.00023870433506090194)),(to_sfixed_a(0.0001460517814848572)),(to_sfixed_a(9.415802196599543e-05)),(to_sfixed_a(0.0006104860221967101)),(to_sfixed_a(0.001443564658984542)),(to_sfixed_a(-6.287623546086252e-05)),(to_sfixed_a(0.00011662197357509285)),(to_sfixed_a(-6.012823723722249e-05)),(to_sfixed_a(0.026686668395996094)),(to_sfixed_a(0.005485838744789362)),(to_sfixed_a(-0.00016798196884337813)),(to_sfixed_a(0.00015231080760713667)),(to_sfixed_a(-0.00011426019773352891)),(to_sfixed_a(-3.8106372812762856e-05)),(to_sfixed_a(0.008856835775077343)),(to_sfixed_a(0.40403634309768677)),(to_sfixed_a(-0.005423331633210182)),(to_sfixed_a(-3.897708666045219e-05)),(to_sfixed_a(-0.0035675298422574997)),(to_sfixed_a(0.000246217823587358)),(to_sfixed_a(-0.013423502445220947)),(to_sfixed_a(-6.162195495562628e-05)),(to_sfixed_a(0.0041090636514127254)),(to_sfixed_a(-0.00011613579408731312)),(to_sfixed_a(-0.018031107261776924)),(to_sfixed_a(-0.002734812907874584)),(to_sfixed_a(-0.001117622246965766)),(to_sfixed_a(0.3651728630065918)),(to_sfixed_a(-5.68139657843858e-05)),(to_sfixed_a(0.36364924907684326)),(to_sfixed_a(-0.0006786943413317204)),(to_sfixed_a(3.219767677364871e-05)),(to_sfixed_a(-0.0011445393320173025)),(to_sfixed_a(5.8444886235520244e-05)),(to_sfixed_a(5.270346446195617e-05)),(to_sfixed_a(0.009739469736814499)),(to_sfixed_a(-0.0011803850065916777)),(to_sfixed_a(-0.0004443828947842121)),(to_sfixed_a(-0.00028716985252685845)),(to_sfixed_a(0.0046288021840155125)),(to_sfixed_a(-0.00013461269554682076)),(to_sfixed_a(-0.0037480134051293135)),(to_sfixed_a(0.0002505416050553322)),(to_sfixed_a(7.034209556877613e-05)),(to_sfixed_a(-9.810255141928792e-05)),(to_sfixed_a(-0.04662545025348663)),(to_sfixed_a(4.0539438487030566e-05)),(to_sfixed_a(-6.854395905975252e-05)),(to_sfixed_a(-5.846258864039555e-05)),(to_sfixed_a(-0.005285106133669615)),(to_sfixed_a(0.31182920932769775)),(to_sfixed_a(-0.00010827968071680516)),(to_sfixed_a(-5.633105320157483e-05)),(to_sfixed_a(-1.6228230379056185e-05)),(to_sfixed_a(-0.00012101579341106117)),(to_sfixed_a(0.01705874316394329)),(to_sfixed_a(-0.007879482582211494)),(to_sfixed_a(-0.0026281101163476706)),(to_sfixed_a(0.003862250130623579)),(to_sfixed_a(-0.01144538912922144)),(to_sfixed_a(9.761461114976555e-07)),(to_sfixed_a(0.00014792928413953632)),(to_sfixed_a(-7.136352360248566e-05)),(to_sfixed_a(-0.0009848900372162461)),(to_sfixed_a(-0.0001701169239822775)),(to_sfixed_a(-7.054889283608645e-05)),(to_sfixed_a(-0.0025654996279627085)),(to_sfixed_a(-0.01694554276764393)),(to_sfixed_a(-1.0702548024710268e-05)),(to_sfixed_a(0.5326322913169861)),(to_sfixed_a(-0.0002747266844380647)),(to_sfixed_a(-0.006919840816408396)),(to_sfixed_a(-0.3272513151168823)),(to_sfixed_a(7.935440953588113e-05)),(to_sfixed_a(-0.0016631707549095154)),(to_sfixed_a(0.01305424328893423)),(to_sfixed_a(-0.0007479691412299871)),(to_sfixed_a(0.0002522203139960766)),(to_sfixed_a(0.004288596101105213)),(to_sfixed_a(0.4799380302429199)),(to_sfixed_a(-0.00016650294128339738)));

    constant weight_n2_40 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.029438402503728867)),(to_sfixed_a(0.3708868622779846)),(to_sfixed_a(0.23312516510486603)),(to_sfixed_a(5.804348620586097e-05)),(to_sfixed_a(0.13740137219429016)),(to_sfixed_a(2.9273134714458138e-05)),(to_sfixed_a(-0.00013003605999983847)),(to_sfixed_a(0.00027292472077533603)),(to_sfixed_a(0.00015389994950965047)),(to_sfixed_a(-0.00019253080245107412)),(to_sfixed_a(1.2129457900300622e-06)),(to_sfixed_a(-0.0034171033184975386)),(to_sfixed_a(-0.1389501541852951)),(to_sfixed_a(-0.00011454064224381)),(to_sfixed_a(-0.00010036141611635685)),(to_sfixed_a(0.00011633984104264528)),(to_sfixed_a(0.014395096339285374)),(to_sfixed_a(1.1692522093653679e-05)),(to_sfixed_a(0.011184087954461575)),(to_sfixed_a(-0.0011608753120526671)),(to_sfixed_a(0.0003018614661414176)),(to_sfixed_a(-0.00016705757298041135)),(to_sfixed_a(1.3477037100528833e-05)),(to_sfixed_a(-0.01374385878443718)),(to_sfixed_a(0.03870224207639694)),(to_sfixed_a(0.004068432841449976)),(to_sfixed_a(-4.397574230097234e-05)),(to_sfixed_a(3.9954444218892604e-05)),(to_sfixed_a(0.0005252882256172597)),(to_sfixed_a(3.1362156732939184e-05)),(to_sfixed_a(-0.0014120396226644516)),(to_sfixed_a(-0.00011757340689655393)),(to_sfixed_a(-0.012845329940319061)),(to_sfixed_a(-4.4606793380808085e-05)),(to_sfixed_a(-0.0002058235986623913)),(to_sfixed_a(-0.00015255746257025748)),(to_sfixed_a(0.004247007425874472)),(to_sfixed_a(-0.0033348065335303545)),(to_sfixed_a(0.004933226387947798)),(to_sfixed_a(-7.632119377376512e-05)),(to_sfixed_a(-0.12256857007741928)),(to_sfixed_a(0.1922432780265808)),(to_sfixed_a(0.00020044928533025086)),(to_sfixed_a(-0.00011321217607473955)),(to_sfixed_a(-0.3465253710746765)),(to_sfixed_a(-0.0014260096941143274)),(to_sfixed_a(0.4105011522769928)),(to_sfixed_a(0.0017747225938364863)),(to_sfixed_a(0.00018574143177829683)),(to_sfixed_a(-0.0008224545163102448)),(to_sfixed_a(0.0016850645188242197)),(to_sfixed_a(-0.00021264306269586086)),(to_sfixed_a(0.0002118283009622246)),(to_sfixed_a(1.2411146599333733e-05)),(to_sfixed_a(-0.01831742748618126)),(to_sfixed_a(0.3270929753780365)),(to_sfixed_a(-0.00014965074660722166)),(to_sfixed_a(-0.0020369826816022396)),(to_sfixed_a(-0.00010911629215115681)),(to_sfixed_a(0.00011742785864043981)),(to_sfixed_a(-2.5116052711382508e-05)),(to_sfixed_a(-0.00019213292398490012)),(to_sfixed_a(0.4186272919178009)),(to_sfixed_a(0.0018293448956683278)),(to_sfixed_a(4.889557749265805e-05)),(to_sfixed_a(0.41611671447753906)),(to_sfixed_a(-0.00014763032959308475)),(to_sfixed_a(-0.00126819615252316)),(to_sfixed_a(0.001127568306401372)),(to_sfixed_a(-1.0285099051543511e-05)),(to_sfixed_a(0.184289813041687)),(to_sfixed_a(-0.25239297747612)),(to_sfixed_a(0.23011663556098938)),(to_sfixed_a(-0.00016416139260400087)),(to_sfixed_a(7.115038170013577e-05)),(to_sfixed_a(-4.878368054050952e-05)),(to_sfixed_a(-0.3262423872947693)),(to_sfixed_a(-0.0008938178070820868)),(to_sfixed_a(-0.0002467230660840869)),(to_sfixed_a(0.009962612763047218)),(to_sfixed_a(-0.0008875172352418303)),(to_sfixed_a(6.574764120159671e-05)),(to_sfixed_a(0.2528136074542999)),(to_sfixed_a(0.0026117160450667143)),(to_sfixed_a(-7.304988685064018e-06)),(to_sfixed_a(-8.455348142888397e-05)),(to_sfixed_a(0.005903951823711395)),(to_sfixed_a(5.948677426204085e-07)),(to_sfixed_a(0.00023572078498546034)),(to_sfixed_a(-6.973029667278752e-05)),(to_sfixed_a(0.3358781337738037)),(to_sfixed_a(1.2745469575747848e-05)),(to_sfixed_a(0.002262710826471448)),(to_sfixed_a(0.0001542686513857916)),(to_sfixed_a(0.0003573825233615935)),(to_sfixed_a(0.0001688088959781453)),(to_sfixed_a(-2.520642738090828e-06)),(to_sfixed_a(0.00013079297787044197)),(to_sfixed_a(1.9832468751701526e-05)),(to_sfixed_a(-0.00016911856073420495)),(to_sfixed_a(-0.0067457701079547405)),(to_sfixed_a(-0.009090865030884743)),(to_sfixed_a(0.00018056451517622918)),(to_sfixed_a(-0.0013610536698251963)),(to_sfixed_a(0.0026714662089943886)),(to_sfixed_a(-5.315095040714368e-05)),(to_sfixed_a(-0.00019333376258146018)),(to_sfixed_a(-7.756045670248568e-05)),(to_sfixed_a(0.00010867534729186445)),(to_sfixed_a(-0.03129151090979576)),(to_sfixed_a(0.3542620837688446)),(to_sfixed_a(-1.8679718778003007e-05)),(to_sfixed_a(-0.0028779739513993263)),(to_sfixed_a(7.177163934102282e-05)),(to_sfixed_a(-0.0002202153264079243)),(to_sfixed_a(-0.1657683104276657)),(to_sfixed_a(-0.0057949949987232685)),(to_sfixed_a(-0.0044807856902480125)),(to_sfixed_a(4.498089037952013e-05)),(to_sfixed_a(-0.2178388088941574)),(to_sfixed_a(0.00016763228632044047)),(to_sfixed_a(0.000231029320275411)),(to_sfixed_a(0.00028540578205138445)),(to_sfixed_a(0.0001298672432312742)),(to_sfixed_a(-0.0002435945498291403)),(to_sfixed_a(-0.015225248411297798)),(to_sfixed_a(-0.0043251062743365765)),(to_sfixed_a(4.2561747250147164e-05)),(to_sfixed_a(0.0003816653334069997)),(to_sfixed_a(-0.00013531015429180115)),(to_sfixed_a(-0.00022607776918448508)),(to_sfixed_a(3.9092323277145624e-05)),(to_sfixed_a(0.0033344512339681387)),(to_sfixed_a(0.24379567801952362)),(to_sfixed_a(-5.4509262554347515e-05)),(to_sfixed_a(-8.538962720194831e-05)),(to_sfixed_a(0.031588055193424225)),(to_sfixed_a(0.00010720168938860297)),(to_sfixed_a(-0.00023574252554681152)),(to_sfixed_a(-0.00012017533299513161)),(to_sfixed_a(0.6035676002502441)),(to_sfixed_a(0.00012702334788627923)),(to_sfixed_a(-1.1541633284650743e-06)),(to_sfixed_a(3.8969232264207676e-05)),(to_sfixed_a(0.40858039259910583)),(to_sfixed_a(0.00019009647076018155)),(to_sfixed_a(-0.00707224290817976)),(to_sfixed_a(0.00013369059888646007)),(to_sfixed_a(0.00015591800911352038)),(to_sfixed_a(0.12974919378757477)),(to_sfixed_a(-0.00032282527536153793)),(to_sfixed_a(5.008940206607804e-06)),(to_sfixed_a(8.460514800390229e-05)),(to_sfixed_a(-6.732202018611133e-05)),(to_sfixed_a(0.00013671295891981572)),(to_sfixed_a(-0.002122262492775917)),(to_sfixed_a(0.0004213551292195916)),(to_sfixed_a(-0.00303790345788002)),(to_sfixed_a(-4.945584441884421e-05)),(to_sfixed_a(0.00011226684000575915)),(to_sfixed_a(-3.470056981313974e-05)),(to_sfixed_a(-6.502670294139534e-05)),(to_sfixed_a(0.011394323781132698)),(to_sfixed_a(0.29769060015678406)),(to_sfixed_a(-0.02728569693863392)),(to_sfixed_a(-0.5099737644195557)),(to_sfixed_a(9.061663877218962e-05)),(to_sfixed_a(-0.001067517208866775)),(to_sfixed_a(-0.00011212573008378968)),(to_sfixed_a(-5.742329085478559e-05)),(to_sfixed_a(-0.05819131061434746)),(to_sfixed_a(0.006382958497852087)),(to_sfixed_a(-0.0038335327990353107)),(to_sfixed_a(6.538725574500859e-05)),(to_sfixed_a(-0.40039315819740295)),(to_sfixed_a(-0.003125521820038557)),(to_sfixed_a(-0.00417762016877532)),(to_sfixed_a(0.00109548878390342)),(to_sfixed_a(0.26111772656440735)),(to_sfixed_a(0.2546682059764862)),(to_sfixed_a(-0.006879924330860376)),(to_sfixed_a(0.001823943923227489)),(to_sfixed_a(-0.00018279487267136574)),(to_sfixed_a(-0.00024180594482459128)),(to_sfixed_a(0.00010673694487195462)),(to_sfixed_a(-0.003585164900869131)),(to_sfixed_a(-0.01473757904022932)),(to_sfixed_a(-0.0005629068473353982)),(to_sfixed_a(0.22253210842609406)),(to_sfixed_a(-7.905382517492399e-06)),(to_sfixed_a(-0.017507413402199745)),(to_sfixed_a(-8.148031338350847e-05)),(to_sfixed_a(-0.006709700915962458)),(to_sfixed_a(9.811137715587392e-05)),(to_sfixed_a(-1.4968565665185452e-05)),(to_sfixed_a(0.002331262454390526)),(to_sfixed_a(-0.00016928199329413474)),(to_sfixed_a(-0.0060616969130933285)),(to_sfixed_a(0.22279101610183716)),(to_sfixed_a(6.176959141157568e-05)),(to_sfixed_a(-7.170950266299769e-05)),(to_sfixed_a(0.0001880540221463889)),(to_sfixed_a(9.027571650221944e-07)),(to_sfixed_a(-0.00015740575327072293)),(to_sfixed_a(0.00017388592823408544)),(to_sfixed_a(0.2524794936180115)),(to_sfixed_a(0.3583710789680481)),(to_sfixed_a(-0.000608637579716742)),(to_sfixed_a(-0.0012401939602568746)),(to_sfixed_a(-0.013692767359316349)),(to_sfixed_a(0.00015506541240029037)),(to_sfixed_a(0.00011871305468957871)),(to_sfixed_a(4.93209736305289e-05)),(to_sfixed_a(-0.00014678091974928975)),(to_sfixed_a(2.2667030862066895e-05)),(to_sfixed_a(0.00020858402422163635)),(to_sfixed_a(-0.007098960690200329)),(to_sfixed_a(-0.010791788809001446)),(to_sfixed_a(0.008774679154157639)),(to_sfixed_a(-3.870518412441015e-06)),(to_sfixed_a(3.293818008387461e-05)),(to_sfixed_a(-0.00019960432837251574)),(to_sfixed_a(-0.00021247110271360725)),(to_sfixed_a(5.407317075878382e-05)),(to_sfixed_a(-0.0041845859959721565)),(to_sfixed_a(-5.697896995116025e-06)),(to_sfixed_a(-1.4048302546143532e-05)),(to_sfixed_a(3.782528074225411e-05)),(to_sfixed_a(-0.36812716722488403)),(to_sfixed_a(0.38800597190856934)),(to_sfixed_a(0.1989699751138687)),(to_sfixed_a(-9.327041334472597e-05)),(to_sfixed_a(-2.9593065846711397e-06)),(to_sfixed_a(6.943016342120245e-05)),(to_sfixed_a(0.0004401108017191291)),(to_sfixed_a(-0.021147064864635468)),(to_sfixed_a(-0.29563120007514954)),(to_sfixed_a(7.152666512411088e-05)),(to_sfixed_a(8.489647007081658e-05)),(to_sfixed_a(0.0002897967351600528)),(to_sfixed_a(-0.03776749223470688)),(to_sfixed_a(7.524819375248626e-05)),(to_sfixed_a(0.22962161898612976)),(to_sfixed_a(0.00031584984390065074)),(to_sfixed_a(-0.005792318843305111)),(to_sfixed_a(-0.0015494741965085268)),(to_sfixed_a(0.01482983585447073)),(to_sfixed_a(-0.00013914049486629665)),(to_sfixed_a(0.00014880420349072665)),(to_sfixed_a(-0.0063341762870550156)),(to_sfixed_a(0.22914554178714752)),(to_sfixed_a(-0.00015704579709563404)),(to_sfixed_a(-0.0006751268520019948)),(to_sfixed_a(-0.00011560722487047315)),(to_sfixed_a(9.069346560863778e-05)),(to_sfixed_a(0.006725456099957228)),(to_sfixed_a(-0.0019738292321562767)),(to_sfixed_a(0.00018253465532325208)),(to_sfixed_a(-4.625194560503587e-05)),(to_sfixed_a(0.0003988310054410249)),(to_sfixed_a(-0.0001374330895487219)),(to_sfixed_a(0.0036041713319718838)),(to_sfixed_a(0.0003037671558558941)),(to_sfixed_a(-8.283546776510775e-06)),(to_sfixed_a(-0.00010309233039151877)),(to_sfixed_a(-0.41720616817474365)),(to_sfixed_a(0.00017609074711799622)),(to_sfixed_a(-1.7306883819401264e-06)),(to_sfixed_a(-0.00015209667617455125)),(to_sfixed_a(0.0018765690037980676)),(to_sfixed_a(-0.004277206026017666)),(to_sfixed_a(-3.5943230614066124e-07)),(to_sfixed_a(-1.8470709619577974e-05)),(to_sfixed_a(0.0001850746339187026)),(to_sfixed_a(0.0001463401858927682)),(to_sfixed_a(0.2517140805721283)),(to_sfixed_a(-0.18188415467739105)),(to_sfixed_a(-0.39217862486839294)),(to_sfixed_a(0.007515793666243553)),(to_sfixed_a(0.26636606454849243)),(to_sfixed_a(0.0001514446339569986)),(to_sfixed_a(8.376761979889125e-05)),(to_sfixed_a(-0.00015730458835605532)),(to_sfixed_a(0.20284684002399445)),(to_sfixed_a(6.0287911765044555e-05)),(to_sfixed_a(5.034533387515694e-06)),(to_sfixed_a(-0.002249437849968672)),(to_sfixed_a(-0.006194444373250008)),(to_sfixed_a(8.319050539284945e-05)),(to_sfixed_a(0.29370805621147156)),(to_sfixed_a(-0.00012745315325446427)),(to_sfixed_a(-0.5996347665786743)),(to_sfixed_a(0.0003774809592869133)),(to_sfixed_a(-0.00015611236449331045)),(to_sfixed_a(-0.004575884900987148)),(to_sfixed_a(-0.013667823746800423)),(to_sfixed_a(0.24867109954357147)),(to_sfixed_a(6.0676302382489666e-05)),(to_sfixed_a(-0.2614717185497284)),(to_sfixed_a(-0.0269466545432806)),(to_sfixed_a(-0.42474132776260376)));

    constant weight_n2_41 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.3807697892189026)),(to_sfixed_a(6.194716115714982e-05)),(to_sfixed_a(-0.00012353251804597676)),(to_sfixed_a(-1.6247446183115244e-05)),(to_sfixed_a(-0.00011914921924471855)),(to_sfixed_a(-0.00024748590658418834)),(to_sfixed_a(3.0634706490673125e-05)),(to_sfixed_a(5.602459714282304e-05)),(to_sfixed_a(-5.889611929887906e-05)),(to_sfixed_a(6.65973057039082e-05)),(to_sfixed_a(0.00018946111958939582)),(to_sfixed_a(-8.322124631376937e-05)),(to_sfixed_a(-2.9116952646290883e-05)),(to_sfixed_a(-0.0001163683264167048)),(to_sfixed_a(6.754390778951347e-05)),(to_sfixed_a(-1.5699384675826877e-05)),(to_sfixed_a(0.0001402752532158047)),(to_sfixed_a(-0.00011263557826168835)),(to_sfixed_a(-5.75225567445159e-06)),(to_sfixed_a(-7.697911496507004e-05)),(to_sfixed_a(-0.00018213674775324762)),(to_sfixed_a(-0.00011178894783370197)),(to_sfixed_a(-7.907191320555285e-05)),(to_sfixed_a(-8.349507697857916e-05)),(to_sfixed_a(0.00011949856707360595)),(to_sfixed_a(7.2962502599693835e-06)),(to_sfixed_a(-2.6417728804517537e-05)),(to_sfixed_a(-7.400979666272178e-05)),(to_sfixed_a(8.177013660315424e-05)),(to_sfixed_a(1.574158522998914e-05)),(to_sfixed_a(-4.538067878456786e-05)),(to_sfixed_a(-1.1296040611341596e-05)),(to_sfixed_a(-6.768778985133395e-05)),(to_sfixed_a(0.00013680517440661788)),(to_sfixed_a(-0.0001136425489676185)),(to_sfixed_a(0.00021452362125273794)),(to_sfixed_a(2.684121864149347e-05)),(to_sfixed_a(-2.7720303478417918e-05)),(to_sfixed_a(-0.00013019773177802563)),(to_sfixed_a(2.9837967304047197e-05)),(to_sfixed_a(1.2530465028248727e-05)),(to_sfixed_a(-4.6947541704867035e-05)),(to_sfixed_a(3.1842064345255494e-05)),(to_sfixed_a(-2.940031117759645e-05)),(to_sfixed_a(-1.2615124433068559e-05)),(to_sfixed_a(-2.9996830562595278e-05)),(to_sfixed_a(2.0342631614767015e-06)),(to_sfixed_a(8.608933421783149e-05)),(to_sfixed_a(1.5591664123348892e-05)),(to_sfixed_a(-2.535932435421273e-05)),(to_sfixed_a(2.8850918170064688e-06)),(to_sfixed_a(0.0002844023401848972)),(to_sfixed_a(-0.0001924818061525002)),(to_sfixed_a(-3.570373519323766e-05)),(to_sfixed_a(6.927482900209725e-06)),(to_sfixed_a(3.1965188100002706e-05)),(to_sfixed_a(2.3211272491607815e-05)),(to_sfixed_a(-5.8099685702472925e-06)),(to_sfixed_a(0.0001136036662501283)),(to_sfixed_a(0.00015743896074127406)),(to_sfixed_a(-0.0002354096359340474)),(to_sfixed_a(-0.00017954650684259832)),(to_sfixed_a(7.923637167550623e-05)),(to_sfixed_a(2.2089267076808028e-05)),(to_sfixed_a(-0.00011271436233073473)),(to_sfixed_a(-6.152880087029189e-05)),(to_sfixed_a(-7.271155482158065e-05)),(to_sfixed_a(-3.969802492065355e-05)),(to_sfixed_a(7.944807293824852e-05)),(to_sfixed_a(-9.8083201010013e-06)),(to_sfixed_a(-2.4019678676268086e-05)),(to_sfixed_a(0.00011172845552209765)),(to_sfixed_a(-0.00011871430615428835)),(to_sfixed_a(-6.782241689506918e-05)),(to_sfixed_a(4.6397370169870555e-05)),(to_sfixed_a(2.3914144549053162e-05)),(to_sfixed_a(5.8946494391420856e-05)),(to_sfixed_a(2.8483329515438527e-05)),(to_sfixed_a(0.0002014807250816375)),(to_sfixed_a(0.00021920895960647613)),(to_sfixed_a(-0.00023135743685998023)),(to_sfixed_a(0.00020171175128780305)),(to_sfixed_a(4.676809112424962e-05)),(to_sfixed_a(-0.00012191466521471739)),(to_sfixed_a(-0.00018583115888759494)),(to_sfixed_a(3.584422665880993e-05)),(to_sfixed_a(6.51638547424227e-05)),(to_sfixed_a(1.517155033070594e-05)),(to_sfixed_a(-1.142734254244715e-05)),(to_sfixed_a(-3.8271817174972966e-05)),(to_sfixed_a(9.389501792611554e-05)),(to_sfixed_a(0.00011396677291486412)),(to_sfixed_a(9.36853903112933e-05)),(to_sfixed_a(3.7346992030506954e-05)),(to_sfixed_a(-3.4903030609712005e-05)),(to_sfixed_a(1.7667865904513747e-05)),(to_sfixed_a(3.1312458304455504e-05)),(to_sfixed_a(-0.0001665608724579215)),(to_sfixed_a(-0.00017559982370585203)),(to_sfixed_a(-8.406132110394537e-06)),(to_sfixed_a(-0.00012270579463802278)),(to_sfixed_a(-0.00012613213039003313)),(to_sfixed_a(-8.559174602851272e-05)),(to_sfixed_a(-0.00012068638170603663)),(to_sfixed_a(0.00013542239321395755)),(to_sfixed_a(-1.5762430848553777e-05)),(to_sfixed_a(0.00014458045188803226)),(to_sfixed_a(8.06950411060825e-05)),(to_sfixed_a(0.00010060363274533302)),(to_sfixed_a(-0.00015143562632147223)),(to_sfixed_a(-2.440116077195853e-05)),(to_sfixed_a(-7.13221961632371e-05)),(to_sfixed_a(4.3062093027401716e-05)),(to_sfixed_a(0.0001146171271102503)),(to_sfixed_a(2.479749673511833e-05)),(to_sfixed_a(0.00013773696264252067)),(to_sfixed_a(-0.00016240938566625118)),(to_sfixed_a(0.00013780909648630768)),(to_sfixed_a(0.00021925933833699673)),(to_sfixed_a(-2.7555379347177222e-05)),(to_sfixed_a(1.8861312128137797e-05)),(to_sfixed_a(0.00017422655946575105)),(to_sfixed_a(0.00012037573469569907)),(to_sfixed_a(0.00022312902729026973)),(to_sfixed_a(-0.0002401791571173817)),(to_sfixed_a(-4.945868568029255e-05)),(to_sfixed_a(-9.254541510017589e-05)),(to_sfixed_a(-0.00028983154334127903)),(to_sfixed_a(-0.00020421970111783594)),(to_sfixed_a(6.636104080826044e-05)),(to_sfixed_a(-1.611042534932494e-05)),(to_sfixed_a(-3.53494833689183e-05)),(to_sfixed_a(-0.00012353579222690314)),(to_sfixed_a(1.8024822566076182e-05)),(to_sfixed_a(-0.0001187481902888976)),(to_sfixed_a(0.00013677489187102765)),(to_sfixed_a(-3.451652082731016e-05)),(to_sfixed_a(-2.9222865123301744e-05)),(to_sfixed_a(0.00012164349755039439)),(to_sfixed_a(-8.721969788894057e-05)),(to_sfixed_a(4.101514059584588e-05)),(to_sfixed_a(1.3224635040387511e-06)),(to_sfixed_a(-0.00022891111439093947)),(to_sfixed_a(-0.00012917305866722018)),(to_sfixed_a(0.00013194026541896164)),(to_sfixed_a(0.0002976452524308115)),(to_sfixed_a(0.00016240196418948472)),(to_sfixed_a(0.00020088521705474705)),(to_sfixed_a(0.00011589203495532274)),(to_sfixed_a(-3.318178642075509e-06)),(to_sfixed_a(-3.602400465751998e-05)),(to_sfixed_a(3.736716462299228e-05)),(to_sfixed_a(-0.00016916112508624792)),(to_sfixed_a(-0.0001418278698110953)),(to_sfixed_a(5.289461114443839e-06)),(to_sfixed_a(-3.312234184704721e-05)),(to_sfixed_a(0.0001709580683382228)),(to_sfixed_a(8.21671201265417e-05)),(to_sfixed_a(-8.747767424210906e-06)),(to_sfixed_a(0.00010807140643009916)),(to_sfixed_a(3.8572383346036077e-05)),(to_sfixed_a(-0.00028605456463992596)),(to_sfixed_a(1.695355967967771e-05)),(to_sfixed_a(-1.6102716472232714e-05)),(to_sfixed_a(-5.1480466936482117e-05)),(to_sfixed_a(3.58231773134321e-05)),(to_sfixed_a(-2.5583831302355975e-05)),(to_sfixed_a(8.021877147257328e-05)),(to_sfixed_a(-0.0002326493849977851)),(to_sfixed_a(8.310416887979954e-05)),(to_sfixed_a(0.14025498926639557)),(to_sfixed_a(4.403920320328325e-05)),(to_sfixed_a(-2.536516694817692e-05)),(to_sfixed_a(4.585628630593419e-06)),(to_sfixed_a(3.042053140234202e-05)),(to_sfixed_a(-0.0001304571924265474)),(to_sfixed_a(4.629560862667859e-06)),(to_sfixed_a(-0.00010887310781981796)),(to_sfixed_a(6.508597289212048e-05)),(to_sfixed_a(5.487192902364768e-05)),(to_sfixed_a(-0.00016074888117145747)),(to_sfixed_a(0.00012674054596573114)),(to_sfixed_a(-0.0001078133936971426)),(to_sfixed_a(-5.423745824373327e-05)),(to_sfixed_a(2.107306499965489e-06)),(to_sfixed_a(7.434649160131812e-05)),(to_sfixed_a(7.008311513345689e-06)),(to_sfixed_a(-2.253969978482928e-05)),(to_sfixed_a(-0.0001259276905329898)),(to_sfixed_a(0.00017530785407871008)),(to_sfixed_a(7.041694334475324e-05)),(to_sfixed_a(0.0002822483074851334)),(to_sfixed_a(0.00016363787290174514)),(to_sfixed_a(-8.424890256719664e-05)),(to_sfixed_a(0.00044957242789678276)),(to_sfixed_a(8.831637387629598e-06)),(to_sfixed_a(0.00011341266508679837)),(to_sfixed_a(-0.00019211355538573116)),(to_sfixed_a(0.00010584498522803187)),(to_sfixed_a(5.960897033219226e-05)),(to_sfixed_a(3.363885480212048e-05)),(to_sfixed_a(-1.1913689377252012e-06)),(to_sfixed_a(0.00010071460565086454)),(to_sfixed_a(5.494366632774472e-06)),(to_sfixed_a(-0.00020245296764187515)),(to_sfixed_a(3.2950338209047914e-05)),(to_sfixed_a(-0.00011677072325255722)),(to_sfixed_a(-6.148031388875097e-05)),(to_sfixed_a(-0.00017060125537682325)),(to_sfixed_a(-8.033588528633118e-05)),(to_sfixed_a(-2.009467061725445e-05)),(to_sfixed_a(0.00013548707647714764)),(to_sfixed_a(0.00015709282888565212)),(to_sfixed_a(-6.749120075255632e-06)),(to_sfixed_a(-0.00018452428048476577)),(to_sfixed_a(-4.11101063946262e-06)),(to_sfixed_a(-4.400488978717476e-05)),(to_sfixed_a(-1.471477298764512e-05)),(to_sfixed_a(-4.091859591426328e-05)),(to_sfixed_a(0.00016947016410995275)),(to_sfixed_a(6.151548586785793e-05)),(to_sfixed_a(0.0002444163546897471)),(to_sfixed_a(6.171679706312716e-05)),(to_sfixed_a(-5.3525291150435805e-06)),(to_sfixed_a(2.105567546095699e-05)),(to_sfixed_a(-2.780392242129892e-05)),(to_sfixed_a(0.00013754967949353158)),(to_sfixed_a(-8.380079816561192e-05)),(to_sfixed_a(6.96102506481111e-05)),(to_sfixed_a(1.4933259080862626e-05)),(to_sfixed_a(-0.12499641627073288)),(to_sfixed_a(0.00011576399265322834)),(to_sfixed_a(-0.0001576655195094645)),(to_sfixed_a(2.915321965701878e-05)),(to_sfixed_a(0.00022722748690284789)),(to_sfixed_a(-4.561919195111841e-05)),(to_sfixed_a(7.731076766503975e-05)),(to_sfixed_a(6.873526581330225e-05)),(to_sfixed_a(-5.0331578677287325e-05)),(to_sfixed_a(-3.3861317206174135e-05)),(to_sfixed_a(0.00018146642833016813)),(to_sfixed_a(-2.939363184850663e-05)),(to_sfixed_a(-5.721642082789913e-05)),(to_sfixed_a(-0.0001354472478851676)),(to_sfixed_a(6.172101711854339e-05)),(to_sfixed_a(-0.00012764424900524318)),(to_sfixed_a(-0.00015857318066991866)),(to_sfixed_a(2.7937938284594566e-05)),(to_sfixed_a(-0.00016971916193142533)),(to_sfixed_a(1.6537076589884236e-05)),(to_sfixed_a(-0.00016967469127848744)),(to_sfixed_a(0.0002970760688185692)),(to_sfixed_a(-2.6214747776975855e-05)),(to_sfixed_a(-0.0001297755225095898)),(to_sfixed_a(0.00023458871874026954)),(to_sfixed_a(-6.505561759695411e-05)),(to_sfixed_a(-6.675901386188343e-05)),(to_sfixed_a(-0.00022034818539395928)),(to_sfixed_a(-0.0001533290633233264)),(to_sfixed_a(0.00017938858945854008)),(to_sfixed_a(-0.00013085106911603361)),(to_sfixed_a(-0.00013756961561739445)),(to_sfixed_a(-7.45698343962431e-07)),(to_sfixed_a(9.605310333427042e-05)),(to_sfixed_a(-0.00016848048835527152)),(to_sfixed_a(4.075678589288145e-05)),(to_sfixed_a(3.639580972958356e-05)),(to_sfixed_a(-0.00021814453066326678)),(to_sfixed_a(3.3629825338721275e-05)),(to_sfixed_a(3.970947363995947e-05)),(to_sfixed_a(8.745562809053808e-06)),(to_sfixed_a(0.00019316165708005428)),(to_sfixed_a(-3.063051190110855e-05)),(to_sfixed_a(-0.00013038043107371777)),(to_sfixed_a(7.865978841437027e-05)),(to_sfixed_a(-2.8913091227877885e-05)),(to_sfixed_a(-9.892797970678657e-05)),(to_sfixed_a(6.380042032105848e-05)),(to_sfixed_a(-5.8193691074848175e-06)),(to_sfixed_a(8.39907443150878e-05)),(to_sfixed_a(0.00024039488926064223)),(to_sfixed_a(-0.00010654662037268281)),(to_sfixed_a(-1.598693779669702e-05)),(to_sfixed_a(1.8105471099261194e-05)),(to_sfixed_a(-6.028784264344722e-05)),(to_sfixed_a(6.309733726084232e-05)),(to_sfixed_a(-3.902643948094919e-05)),(to_sfixed_a(-9.71661793300882e-05)),(to_sfixed_a(0.00015602124040015042)),(to_sfixed_a(-2.3372704163193703e-06)),(to_sfixed_a(5.083900032332167e-05)),(to_sfixed_a(-7.594650378450751e-05)),(to_sfixed_a(8.92385869519785e-05)),(to_sfixed_a(2.4965826014522463e-05)),(to_sfixed_a(0.00017680699238553643)),(to_sfixed_a(-0.00010903101065196097)),(to_sfixed_a(4.9801270506577566e-05)),(to_sfixed_a(0.00024638924514874816)),(to_sfixed_a(-1.713083838694729e-05)),(to_sfixed_a(1.601031362952199e-05)),(to_sfixed_a(-5.953687650617212e-05)));

    constant weight_n2_42 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.33024075627326965)),(to_sfixed_a(0.0010981069644913077)),(to_sfixed_a(-0.001412191311828792)),(to_sfixed_a(-0.00024406301963608712)),(to_sfixed_a(-0.002205335069447756)),(to_sfixed_a(-2.4378565285587683e-05)),(to_sfixed_a(-0.0063086580485105515)),(to_sfixed_a(-0.00010011820995714515)),(to_sfixed_a(-0.0001891734718810767)),(to_sfixed_a(0.00018038001144304872)),(to_sfixed_a(-3.0436960514634848e-05)),(to_sfixed_a(0.0014813189627602696)),(to_sfixed_a(0.1809302568435669)),(to_sfixed_a(0.0022017396986484528)),(to_sfixed_a(0.00010503207158762962)),(to_sfixed_a(-0.0002378226927248761)),(to_sfixed_a(-0.0003758690145332366)),(to_sfixed_a(-3.7918063753750175e-05)),(to_sfixed_a(-0.00023630903160665184)),(to_sfixed_a(-0.0009790334152057767)),(to_sfixed_a(-5.747794784838334e-05)),(to_sfixed_a(0.00011650413216557354)),(to_sfixed_a(-6.687191489618272e-05)),(to_sfixed_a(-0.0027908661868423223)),(to_sfixed_a(-0.009775090962648392)),(to_sfixed_a(-0.0015053694369271398)),(to_sfixed_a(-8.831805462250486e-05)),(to_sfixed_a(-8.874628110788763e-05)),(to_sfixed_a(0.00017063895938917994)),(to_sfixed_a(-0.00024054931418504566)),(to_sfixed_a(-0.006478213705122471)),(to_sfixed_a(5.076704837847501e-05)),(to_sfixed_a(-0.0031796791590750217)),(to_sfixed_a(0.00011439079389674589)),(to_sfixed_a(0.00016306567704305053)),(to_sfixed_a(-3.8887374103069305e-06)),(to_sfixed_a(0.1600160300731659)),(to_sfixed_a(-0.10813070088624954)),(to_sfixed_a(-0.010484679602086544)),(to_sfixed_a(-2.6598936528898776e-06)),(to_sfixed_a(-0.14600211381912231)),(to_sfixed_a(-0.000702072458807379)),(to_sfixed_a(0.00013769780343864113)),(to_sfixed_a(0.00021166002261452377)),(to_sfixed_a(-0.000345804903190583)),(to_sfixed_a(0.00010098992061102763)),(to_sfixed_a(0.0009468364296481013)),(to_sfixed_a(-0.002741752890869975)),(to_sfixed_a(0.0001675860839895904)),(to_sfixed_a(-0.00214173411950469)),(to_sfixed_a(-0.3281281292438507)),(to_sfixed_a(-0.000650550180580467)),(to_sfixed_a(-2.177948772441596e-06)),(to_sfixed_a(-0.0012375748483464122)),(to_sfixed_a(-0.37219709157943726)),(to_sfixed_a(-0.011049623601138592)),(to_sfixed_a(0.00010587093129288405)),(to_sfixed_a(0.0018588671227917075)),(to_sfixed_a(-0.00024070042127277702)),(to_sfixed_a(0.0004232318024151027)),(to_sfixed_a(-0.0014589236816391349)),(to_sfixed_a(-0.0028510885313153267)),(to_sfixed_a(-9.631221473682672e-06)),(to_sfixed_a(-0.002785159507766366)),(to_sfixed_a(-3.223470048396848e-05)),(to_sfixed_a(-0.0009985044598579407)),(to_sfixed_a(9.532689000479877e-05)),(to_sfixed_a(-0.0950758159160614)),(to_sfixed_a(-0.004601822700351477)),(to_sfixed_a(6.139118340797722e-06)),(to_sfixed_a(0.0024446076713502407)),(to_sfixed_a(-0.00415465934202075)),(to_sfixed_a(6.751419277861714e-05)),(to_sfixed_a(-0.00011253349657636136)),(to_sfixed_a(0.0003200858482159674)),(to_sfixed_a(-9.171378042083234e-05)),(to_sfixed_a(-0.0004547313437797129)),(to_sfixed_a(-0.00417366623878479)),(to_sfixed_a(-1.465778041165322e-06)),(to_sfixed_a(0.004273109138011932)),(to_sfixed_a(0.0015858672559261322)),(to_sfixed_a(-6.557063898071647e-05)),(to_sfixed_a(-0.004590688273310661)),(to_sfixed_a(0.0010683551663532853)),(to_sfixed_a(-0.00010105570981977507)),(to_sfixed_a(-0.006173849105834961)),(to_sfixed_a(-0.0036167814396321774)),(to_sfixed_a(0.0016751711955294013)),(to_sfixed_a(3.0127186619210988e-05)),(to_sfixed_a(-2.7266709366813302e-05)),(to_sfixed_a(0.003924278542399406)),(to_sfixed_a(4.834886931348592e-05)),(to_sfixed_a(-0.0033958032727241516)),(to_sfixed_a(0.00020299162133596838)),(to_sfixed_a(-0.003944993484765291)),(to_sfixed_a(1.238364347955212e-05)),(to_sfixed_a(6.748773012077436e-05)),(to_sfixed_a(0.00017345647211186588)),(to_sfixed_a(-5.296968447510153e-05)),(to_sfixed_a(2.932195639004931e-05)),(to_sfixed_a(-0.0014561782591044903)),(to_sfixed_a(-0.0029754932038486004)),(to_sfixed_a(0.00029278313741087914)),(to_sfixed_a(-0.00618977565318346)),(to_sfixed_a(-0.003511545481160283)),(to_sfixed_a(-0.00019691625493578613)),(to_sfixed_a(-1.3989065337227657e-06)),(to_sfixed_a(2.278730971738696e-05)),(to_sfixed_a(-6.966909859329462e-05)),(to_sfixed_a(-0.0033627005759626627)),(to_sfixed_a(0.004313149489462376)),(to_sfixed_a(6.764999125152826e-05)),(to_sfixed_a(6.670189759461209e-05)),(to_sfixed_a(8.932022319640964e-05)),(to_sfixed_a(-0.00013913589646108449)),(to_sfixed_a(-0.008384318090975285)),(to_sfixed_a(0.00021023143199272454)),(to_sfixed_a(0.00021040583669673651)),(to_sfixed_a(-0.00018101933528669178)),(to_sfixed_a(-0.0006566905067302287)),(to_sfixed_a(-7.135100895538926e-05)),(to_sfixed_a(-6.538118032040074e-05)),(to_sfixed_a(-0.00013219841639511287)),(to_sfixed_a(-0.0002556189720053226)),(to_sfixed_a(1.4919467503204942e-05)),(to_sfixed_a(-0.0007308933418244123)),(to_sfixed_a(0.004964966792613268)),(to_sfixed_a(3.050832310691476e-05)),(to_sfixed_a(-0.0001741094165481627)),(to_sfixed_a(0.00015307344438042492)),(to_sfixed_a(-5.768996197730303e-05)),(to_sfixed_a(-6.466946797445416e-05)),(to_sfixed_a(-0.0012292537139728665)),(to_sfixed_a(0.0036999224685132504)),(to_sfixed_a(-0.0001994055201066658)),(to_sfixed_a(0.0001746859634295106)),(to_sfixed_a(-0.27287301421165466)),(to_sfixed_a(-7.170100434450433e-05)),(to_sfixed_a(1.5427656762767583e-05)),(to_sfixed_a(0.00019970825815107673)),(to_sfixed_a(0.002861375454813242)),(to_sfixed_a(-5.733182479161769e-05)),(to_sfixed_a(-3.693567123264074e-05)),(to_sfixed_a(5.45790717296768e-05)),(to_sfixed_a(-0.0008704972569830716)),(to_sfixed_a(0.00012175639858469367)),(to_sfixed_a(0.1932326704263687)),(to_sfixed_a(-2.3588039766764268e-05)),(to_sfixed_a(0.00011354642629157752)),(to_sfixed_a(0.0028120181523263454)),(to_sfixed_a(-0.0001175820580101572)),(to_sfixed_a(3.514922718750313e-05)),(to_sfixed_a(-0.10733254253864288)),(to_sfixed_a(3.065005148528144e-05)),(to_sfixed_a(0.000207088582101278)),(to_sfixed_a(0.0012367061572149396)),(to_sfixed_a(-1.715667895041406e-05)),(to_sfixed_a(-0.0006843769224360585)),(to_sfixed_a(3.588352046790533e-05)),(to_sfixed_a(-2.6048990548588336e-05)),(to_sfixed_a(-0.000104375125374645)),(to_sfixed_a(4.6390341594815254e-05)),(to_sfixed_a(0.006926513742655516)),(to_sfixed_a(0.0009558992460370064)),(to_sfixed_a(-0.002170740393921733)),(to_sfixed_a(0.0027831511106342077)),(to_sfixed_a(0.0002385443076491356)),(to_sfixed_a(-0.0033385809510946274)),(to_sfixed_a(0.0001869405823526904)),(to_sfixed_a(0.00012532452819868922)),(to_sfixed_a(-0.001669962308369577)),(to_sfixed_a(0.0002856240898836404)),(to_sfixed_a(1.0243005817756057e-05)),(to_sfixed_a(-0.00011909719614777714)),(to_sfixed_a(-0.00109389191493392)),(to_sfixed_a(-0.0006018953863531351)),(to_sfixed_a(-0.0021105362102389336)),(to_sfixed_a(-9.262458479497582e-05)),(to_sfixed_a(-0.0016940569039434195)),(to_sfixed_a(0.0007536670891568065)),(to_sfixed_a(-0.0010145928245037794)),(to_sfixed_a(-0.00019882808555848897)),(to_sfixed_a(7.18267256161198e-05)),(to_sfixed_a(0.0002403871767455712)),(to_sfixed_a(0.00017714317073114216)),(to_sfixed_a(-0.0002654880518093705)),(to_sfixed_a(-0.0008011558093130589)),(to_sfixed_a(-0.0012825271114706993)),(to_sfixed_a(0.0018658597255125642)),(to_sfixed_a(0.00043629464926198125)),(to_sfixed_a(-0.22913329303264618)),(to_sfixed_a(-5.081534618511796e-05)),(to_sfixed_a(-0.005796331912279129)),(to_sfixed_a(0.0001907732803374529)),(to_sfixed_a(4.0985600207932293e-05)),(to_sfixed_a(-0.000579319428652525)),(to_sfixed_a(6.836623651906848e-05)),(to_sfixed_a(-0.0022818087600171566)),(to_sfixed_a(-0.0035980287939310074)),(to_sfixed_a(0.00011382170487195253)),(to_sfixed_a(0.00041348530794493854)),(to_sfixed_a(4.426123632583767e-05)),(to_sfixed_a(1.4444085536524653e-05)),(to_sfixed_a(5.3394458518596366e-05)),(to_sfixed_a(-4.392248229123652e-05)),(to_sfixed_a(-0.0008666742942295969)),(to_sfixed_a(0.00309380772523582)),(to_sfixed_a(-0.00020544312428683043)),(to_sfixed_a(-0.0017838107887655497)),(to_sfixed_a(-0.0026403265073895454)),(to_sfixed_a(-0.0035780295729637146)),(to_sfixed_a(7.208655006252229e-09)),(to_sfixed_a(2.4775745259830728e-05)),(to_sfixed_a(-9.311700705438852e-05)),(to_sfixed_a(3.221970109734684e-05)),(to_sfixed_a(-1.9008431991096586e-05)),(to_sfixed_a(0.004109683446586132)),(to_sfixed_a(-0.0004643095307983458)),(to_sfixed_a(-0.27356910705566406)),(to_sfixed_a(1.057283952832222e-05)),(to_sfixed_a(-5.949266778770834e-06)),(to_sfixed_a(-5.695808067684993e-05)),(to_sfixed_a(3.082168404944241e-05)),(to_sfixed_a(0.000186545992619358)),(to_sfixed_a(-0.0006466592894867063)),(to_sfixed_a(-0.00014941726112738252)),(to_sfixed_a(-6.83319813106209e-05)),(to_sfixed_a(-0.00015347535372711718)),(to_sfixed_a(0.0023297439329326153)),(to_sfixed_a(-0.0025057303719222546)),(to_sfixed_a(-0.00024056457914412022)),(to_sfixed_a(-7.867375097703189e-05)),(to_sfixed_a(-8.837733912514523e-05)),(to_sfixed_a(-2.3066409994498827e-05)),(to_sfixed_a(0.0001854945730883628)),(to_sfixed_a(-0.0025395972188562155)),(to_sfixed_a(0.2266046404838562)),(to_sfixed_a(-0.00012944061018060893)),(to_sfixed_a(-0.0009011123911477625)),(to_sfixed_a(-0.0001005289814202115)),(to_sfixed_a(0.00016030148253776133)),(to_sfixed_a(0.00045202835462987423)),(to_sfixed_a(-0.001473442418500781)),(to_sfixed_a(0.00013016434968449175)),(to_sfixed_a(0.010372959077358246)),(to_sfixed_a(0.0025798336137086153)),(to_sfixed_a(-0.0009252472664229572)),(to_sfixed_a(-0.0009651270811446011)),(to_sfixed_a(-1.9387414795346558e-05)),(to_sfixed_a(-0.006456052418798208)),(to_sfixed_a(-0.000210518017411232)),(to_sfixed_a(-0.00015636722673662007)),(to_sfixed_a(0.0013735702959820628)),(to_sfixed_a(-0.00026823231019079685)),(to_sfixed_a(-0.0006007792544551194)),(to_sfixed_a(-0.009708949364721775)),(to_sfixed_a(-0.002807068871334195)),(to_sfixed_a(0.0004472954897210002)),(to_sfixed_a(-1.4553348592016846e-05)),(to_sfixed_a(-0.0016205162974074483)),(to_sfixed_a(5.030531610827893e-06)),(to_sfixed_a(0.002794686472043395)),(to_sfixed_a(-1.8244485545437783e-05)),(to_sfixed_a(-0.0012581886257976294)),(to_sfixed_a(-0.00013559543003793806)),(to_sfixed_a(-0.006790033541619778)),(to_sfixed_a(-0.00014855196059215814)),(to_sfixed_a(0.0001009884217637591)),(to_sfixed_a(-6.9249090302037075e-06)),(to_sfixed_a(0.1905476152896881)),(to_sfixed_a(-0.0031468947418034077)),(to_sfixed_a(7.578792428830639e-05)),(to_sfixed_a(-0.00021708215354010463)),(to_sfixed_a(0.00010374520206823945)),(to_sfixed_a(-0.00011696712317643687)),(to_sfixed_a(-0.006354296579957008)),(to_sfixed_a(-0.004811967723071575)),(to_sfixed_a(0.0007188867311924696)),(to_sfixed_a(0.1493416726589203)),(to_sfixed_a(0.0001387017546221614)),(to_sfixed_a(-1.945759868249297e-05)),(to_sfixed_a(-3.6960700526833534e-05)),(to_sfixed_a(-3.7323148717405275e-05)),(to_sfixed_a(-0.001441410044208169)),(to_sfixed_a(-5.7626733905635774e-05)),(to_sfixed_a(-9.104570926865563e-05)),(to_sfixed_a(0.0028215947095304728)),(to_sfixed_a(0.5466426014900208)),(to_sfixed_a(-1.4191318769007921e-05)),(to_sfixed_a(-0.0011401473311707377)),(to_sfixed_a(-0.00150221714284271)),(to_sfixed_a(-9.490589945926331e-06)),(to_sfixed_a(0.1985434889793396)),(to_sfixed_a(-0.00015608732064720243)),(to_sfixed_a(-0.004731619730591774)),(to_sfixed_a(0.002406272105872631)),(to_sfixed_a(-0.001185274450108409)),(to_sfixed_a(1.5274505130946636e-05)),(to_sfixed_a(0.0035502195823937654)),(to_sfixed_a(0.0010443812934681773)),(to_sfixed_a(-0.0060715083964169025)));

    constant weight_n2_43 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.1487203985452652)),(to_sfixed_a(-0.0029085788410156965)),(to_sfixed_a(0.3467563986778259)),(to_sfixed_a(6.435677642002702e-05)),(to_sfixed_a(0.004146211314946413)),(to_sfixed_a(0.000168586106155999)),(to_sfixed_a(-0.001485510845668614)),(to_sfixed_a(0.00026417814660817385)),(to_sfixed_a(0.00028963532531633973)),(to_sfixed_a(9.791876072995365e-05)),(to_sfixed_a(3.691673555294983e-05)),(to_sfixed_a(0.0015513418475165963)),(to_sfixed_a(-0.48807570338249207)),(to_sfixed_a(0.0021222559735178947)),(to_sfixed_a(5.792862066300586e-05)),(to_sfixed_a(9.159951150650159e-05)),(to_sfixed_a(0.17377996444702148)),(to_sfixed_a(-1.0901228961301968e-05)),(to_sfixed_a(0.2778453826904297)),(to_sfixed_a(-0.013497265055775642)),(to_sfixed_a(-8.453698683297262e-05)),(to_sfixed_a(-0.0002711321576498449)),(to_sfixed_a(0.00015699522919021547)),(to_sfixed_a(-0.001403974718414247)),(to_sfixed_a(-0.005567905958741903)),(to_sfixed_a(-0.0006141511257737875)),(to_sfixed_a(-0.000458134978543967)),(to_sfixed_a(0.0005940893897786736)),(to_sfixed_a(0.007012682501226664)),(to_sfixed_a(-4.6540211769752204e-05)),(to_sfixed_a(-0.03511752933263779)),(to_sfixed_a(0.00013144811964593828)),(to_sfixed_a(-0.009628979489207268)),(to_sfixed_a(1.2024756870232522e-06)),(to_sfixed_a(-4.13366942666471e-05)),(to_sfixed_a(4.020999767817557e-06)),(to_sfixed_a(-0.0005648054648190737)),(to_sfixed_a(-0.0020709766540676355)),(to_sfixed_a(0.011029301211237907)),(to_sfixed_a(-0.0001341810857411474)),(to_sfixed_a(0.4119277894496918)),(to_sfixed_a(0.20937605202198029)),(to_sfixed_a(0.0001224640873260796)),(to_sfixed_a(0.00012645476090256125)),(to_sfixed_a(0.00014246307546272874)),(to_sfixed_a(-0.2196088582277298)),(to_sfixed_a(0.3197697401046753)),(to_sfixed_a(0.6219861507415771)),(to_sfixed_a(-9.177959873341024e-05)),(to_sfixed_a(0.00399944419041276)),(to_sfixed_a(0.0980529636144638)),(to_sfixed_a(-0.0002223825140390545)),(to_sfixed_a(-0.00029294146224856377)),(to_sfixed_a(0.004312371835112572)),(to_sfixed_a(0.0012607991229742765)),(to_sfixed_a(-0.0016088407719507813)),(to_sfixed_a(-0.00023636895639356226)),(to_sfixed_a(-0.0007965476834215224)),(to_sfixed_a(3.6526813346426934e-05)),(to_sfixed_a(0.000200400419998914)),(to_sfixed_a(-0.01851540058851242)),(to_sfixed_a(0.0006121635087765753)),(to_sfixed_a(0.000507452292367816)),(to_sfixed_a(-0.4669477045536041)),(to_sfixed_a(-0.00026876968331635)),(to_sfixed_a(0.36476612091064453)),(to_sfixed_a(-1.0531981388339773e-05)),(to_sfixed_a(0.5098674297332764)),(to_sfixed_a(0.0004115033952984959)),(to_sfixed_a(-2.5119703423115425e-05)),(to_sfixed_a(-0.0031256284564733505)),(to_sfixed_a(-0.23627789318561554)),(to_sfixed_a(-0.21489623188972473)),(to_sfixed_a(-0.00015449429338332266)),(to_sfixed_a(0.0001500031939940527)),(to_sfixed_a(-7.190233009168878e-05)),(to_sfixed_a(-0.20550405979156494)),(to_sfixed_a(-0.001479440601542592)),(to_sfixed_a(3.0488041375065222e-05)),(to_sfixed_a(0.49701541662216187)),(to_sfixed_a(-0.0004659978440031409)),(to_sfixed_a(-0.00019347851048223674)),(to_sfixed_a(0.0013121376978233457)),(to_sfixed_a(-0.14377430081367493)),(to_sfixed_a(-9.244131797458977e-05)),(to_sfixed_a(5.031928594689816e-05)),(to_sfixed_a(-0.0010700846323743463)),(to_sfixed_a(0.004523417446762323)),(to_sfixed_a(6.417502299882472e-05)),(to_sfixed_a(0.0002370255097048357)),(to_sfixed_a(-0.001051601953804493)),(to_sfixed_a(0.0002700445184018463)),(to_sfixed_a(5.480338586494327e-06)),(to_sfixed_a(0.0004202217096462846)),(to_sfixed_a(-0.0021726302802562714)),(to_sfixed_a(-6.885520997457206e-05)),(to_sfixed_a(-6.448930071201175e-05)),(to_sfixed_a(1.847299608925823e-05)),(to_sfixed_a(-9.560221951687708e-05)),(to_sfixed_a(0.00014880491653457284)),(to_sfixed_a(0.00045354061876423657)),(to_sfixed_a(-0.0007804660126566887)),(to_sfixed_a(0.0001362904004054144)),(to_sfixed_a(-0.24150404334068298)),(to_sfixed_a(-0.27676859498023987)),(to_sfixed_a(0.0005810167640447617)),(to_sfixed_a(-0.00011321429337840527)),(to_sfixed_a(-1.1611223271756899e-06)),(to_sfixed_a(4.136960342293605e-05)),(to_sfixed_a(0.0003778286336455494)),(to_sfixed_a(-0.006971598137170076)),(to_sfixed_a(9.736220818012953e-06)),(to_sfixed_a(0.4240014851093292)),(to_sfixed_a(-0.00023651921947021037)),(to_sfixed_a(-0.00010827468213392422)),(to_sfixed_a(-0.0812031477689743)),(to_sfixed_a(-0.0024393093772232533)),(to_sfixed_a(0.000995442271232605)),(to_sfixed_a(-2.496343950042501e-05)),(to_sfixed_a(-0.001178950653411448)),(to_sfixed_a(2.000454333028756e-05)),(to_sfixed_a(-0.00013095236499793828)),(to_sfixed_a(0.0006254241452552378)),(to_sfixed_a(-0.00011726122465915978)),(to_sfixed_a(2.175063855247572e-05)),(to_sfixed_a(0.22737358510494232)),(to_sfixed_a(-0.0027096078265458345)),(to_sfixed_a(0.00029511755565181375)),(to_sfixed_a(-7.706972246523947e-05)),(to_sfixed_a(-3.7069694371894e-05)),(to_sfixed_a(-7.024359365459532e-05)),(to_sfixed_a(-1.4305616787169129e-05)),(to_sfixed_a(-0.0027378981467336416)),(to_sfixed_a(0.00025680821272544563)),(to_sfixed_a(-6.961397593840957e-05)),(to_sfixed_a(-2.699009928619489e-05)),(to_sfixed_a(0.3498561680316925)),(to_sfixed_a(0.3598153591156006)),(to_sfixed_a(0.00024202032363973558)),(to_sfixed_a(0.00020007468992844224)),(to_sfixed_a(0.35244220495224)),(to_sfixed_a(0.00023564440198242664)),(to_sfixed_a(5.7579774875193834e-05)),(to_sfixed_a(-5.585789040196687e-06)),(to_sfixed_a(-0.0025702607817947865)),(to_sfixed_a(-6.707017018925399e-05)),(to_sfixed_a(0.00020680180750787258)),(to_sfixed_a(-0.0001292597153224051)),(to_sfixed_a(-5.220333332545124e-05)),(to_sfixed_a(-0.0018766620196402073)),(to_sfixed_a(-9.002869774121791e-07)),(to_sfixed_a(-0.0001172911433968693)),(to_sfixed_a(-0.020400406792759895)),(to_sfixed_a(0.00045310985296964645)),(to_sfixed_a(0.00024245379609055817)),(to_sfixed_a(-0.39825379848480225)),(to_sfixed_a(-4.8513793444726616e-05)),(to_sfixed_a(0.0048086922615766525)),(to_sfixed_a(4.3091113184345886e-05)),(to_sfixed_a(-0.00028309368644841015)),(to_sfixed_a(6.177987233968452e-05)),(to_sfixed_a(-3.109373210463673e-05)),(to_sfixed_a(-0.006659075152128935)),(to_sfixed_a(-0.001276574213989079)),(to_sfixed_a(-0.033517781645059586)),(to_sfixed_a(-0.0008088427130132914)),(to_sfixed_a(0.0001481505751144141)),(to_sfixed_a(0.7030659317970276)),(to_sfixed_a(-7.086458208505064e-05)),(to_sfixed_a(-4.603634442901239e-05)),(to_sfixed_a(-4.900647036265582e-05)),(to_sfixed_a(-0.006256811786442995)),(to_sfixed_a(-0.002978693228214979)),(to_sfixed_a(-4.4825650547863916e-05)),(to_sfixed_a(0.39675000309944153)),(to_sfixed_a(-0.0018083363538607955)),(to_sfixed_a(0.09948424249887466)),(to_sfixed_a(0.3231375217437744)),(to_sfixed_a(0.0004892557044513524)),(to_sfixed_a(0.1274106353521347)),(to_sfixed_a(0.0012303013354539871)),(to_sfixed_a(0.1700485199689865)),(to_sfixed_a(0.00010490008571650833)),(to_sfixed_a(-7.701524009462446e-05)),(to_sfixed_a(0.00010227011080132797)),(to_sfixed_a(0.012432720512151718)),(to_sfixed_a(-0.015662480145692825)),(to_sfixed_a(0.004647143185138702)),(to_sfixed_a(-0.0009415022796019912)),(to_sfixed_a(-0.0015202021459117532)),(to_sfixed_a(-0.0017147529870271683)),(to_sfixed_a(-0.0002813769970089197)),(to_sfixed_a(0.4212338328361511)),(to_sfixed_a(0.0009916374692693353)),(to_sfixed_a(0.00018222807557322085)),(to_sfixed_a(0.0007808897644281387)),(to_sfixed_a(-6.824098818469793e-05)),(to_sfixed_a(-0.005964736919850111)),(to_sfixed_a(-0.001177978701889515)),(to_sfixed_a(-4.51933010481298e-05)),(to_sfixed_a(-0.00017758840112946928)),(to_sfixed_a(-0.00020501349354162812)),(to_sfixed_a(2.3427004634868354e-05)),(to_sfixed_a(6.031055090716109e-05)),(to_sfixed_a(0.00014800966891925782)),(to_sfixed_a(0.19623589515686035)),(to_sfixed_a(-0.002789827296510339)),(to_sfixed_a(0.14244942367076874)),(to_sfixed_a(7.883450598455966e-05)),(to_sfixed_a(0.0014181457227095962)),(to_sfixed_a(0.0033691562712192535)),(to_sfixed_a(1.959197106771171e-06)),(to_sfixed_a(-0.00011598174751270562)),(to_sfixed_a(-3.0216764571378008e-05)),(to_sfixed_a(2.002146720769815e-05)),(to_sfixed_a(-5.939014590694569e-05)),(to_sfixed_a(0.004499251954257488)),(to_sfixed_a(-0.0033159221056848764)),(to_sfixed_a(0.0020249129738658667)),(to_sfixed_a(1.7165708413813263e-05)),(to_sfixed_a(-0.00021980414749123156)),(to_sfixed_a(0.0002430482127238065)),(to_sfixed_a(-0.00011766879470087588)),(to_sfixed_a(0.0008781534852460027)),(to_sfixed_a(0.002065481850877404)),(to_sfixed_a(-0.0001145100177382119)),(to_sfixed_a(1.8380007531959563e-05)),(to_sfixed_a(4.432673449628055e-06)),(to_sfixed_a(-0.015171266160905361)),(to_sfixed_a(-0.000860820000525564)),(to_sfixed_a(0.2521263659000397)),(to_sfixed_a(-6.962964835111052e-05)),(to_sfixed_a(-0.00017211395606864244)),(to_sfixed_a(-0.00010170481982640922)),(to_sfixed_a(-0.0020283751655369997)),(to_sfixed_a(-0.0025023436173796654)),(to_sfixed_a(-0.006873671431094408)),(to_sfixed_a(0.00012713417527265847)),(to_sfixed_a(0.00015646246902178973)),(to_sfixed_a(-0.00028471992118284106)),(to_sfixed_a(-0.0048151277005672455)),(to_sfixed_a(-1.0584670235402882e-05)),(to_sfixed_a(0.010792168788611889)),(to_sfixed_a(0.00017355858290102333)),(to_sfixed_a(0.4009741246700287)),(to_sfixed_a(-0.002351614646613598)),(to_sfixed_a(0.00026514893397688866)),(to_sfixed_a(-0.0056333355605602264)),(to_sfixed_a(-1.7613820091355592e-07)),(to_sfixed_a(-0.008521178737282753)),(to_sfixed_a(0.00684881117194891)),(to_sfixed_a(-1.749761577229947e-05)),(to_sfixed_a(0.002061284612864256)),(to_sfixed_a(-9.801337000681087e-05)),(to_sfixed_a(0.0005426477291621268)),(to_sfixed_a(-0.0007916481117717922)),(to_sfixed_a(-0.0015740725211799145)),(to_sfixed_a(6.8432476837188e-05)),(to_sfixed_a(4.914507735520601e-05)),(to_sfixed_a(0.0019117306219413877)),(to_sfixed_a(-0.00015359089593403041)),(to_sfixed_a(0.004196206107735634)),(to_sfixed_a(-7.651936903130263e-05)),(to_sfixed_a(0.0007116791093721986)),(to_sfixed_a(2.3179753043223172e-05)),(to_sfixed_a(0.0006679671932943165)),(to_sfixed_a(8.743854414205998e-05)),(to_sfixed_a(7.68748577684164e-06)),(to_sfixed_a(7.11870234226808e-05)),(to_sfixed_a(-0.0005816928460262716)),(to_sfixed_a(0.0026615820825099945)),(to_sfixed_a(-0.00016902023344300687)),(to_sfixed_a(0.00016852928092703223)),(to_sfixed_a(0.00016967725241556764)),(to_sfixed_a(7.609504973515868e-05)),(to_sfixed_a(-0.004173845984041691)),(to_sfixed_a(0.446163535118103)),(to_sfixed_a(-0.00042854828643612564)),(to_sfixed_a(-0.013590446673333645)),(to_sfixed_a(-0.0025409776717424393)),(to_sfixed_a(3.8323218177538365e-05)),(to_sfixed_a(0.00029188813641667366)),(to_sfixed_a(-4.355644341558218e-05)),(to_sfixed_a(0.0006963365594856441)),(to_sfixed_a(3.794631629716605e-05)),(to_sfixed_a(-6.506985664600506e-05)),(to_sfixed_a(0.002059878082945943)),(to_sfixed_a(-0.7723646759986877)),(to_sfixed_a(1.113602047553286e-05)),(to_sfixed_a(-0.2208210527896881)),(to_sfixed_a(0.0003550209803506732)),(to_sfixed_a(-0.03396405279636383)),(to_sfixed_a(-0.010150429792702198)),(to_sfixed_a(-1.535149203846231e-05)),(to_sfixed_a(-0.010530155152082443)),(to_sfixed_a(0.33808523416519165)),(to_sfixed_a(0.008926312439143658)),(to_sfixed_a(3.905475023202598e-05)),(to_sfixed_a(-0.3858836889266968)),(to_sfixed_a(0.2122267782688141)),(to_sfixed_a(0.28012216091156006)));

    constant weight_n2_44 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.6011501550674438)),(to_sfixed_a(-0.5084386467933655)),(to_sfixed_a(-0.2359226793050766)),(to_sfixed_a(-3.933884727302939e-05)),(to_sfixed_a(-0.02490607462823391)),(to_sfixed_a(-2.3562148271594197e-05)),(to_sfixed_a(0.002435225760564208)),(to_sfixed_a(0.00012124293425586075)),(to_sfixed_a(-0.00011374062160030007)),(to_sfixed_a(0.00011643418110907078)),(to_sfixed_a(-0.00029343037749640644)),(to_sfixed_a(0.011759680695831776)),(to_sfixed_a(-0.01460241712629795)),(to_sfixed_a(0.062238287180662155)),(to_sfixed_a(3.732306504389271e-05)),(to_sfixed_a(-6.881384615553543e-05)),(to_sfixed_a(-0.016359075903892517)),(to_sfixed_a(-3.5311750252731144e-06)),(to_sfixed_a(-0.29623734951019287)),(to_sfixed_a(3.0486924515571445e-05)),(to_sfixed_a(0.00010645357542671263)),(to_sfixed_a(-4.753619577968493e-06)),(to_sfixed_a(-0.0012497048592194915)),(to_sfixed_a(-2.0098606910323724e-05)),(to_sfixed_a(0.4410634934902191)),(to_sfixed_a(0.007980716414749622)),(to_sfixed_a(-0.0001202055427711457)),(to_sfixed_a(-0.0017722249031066895)),(to_sfixed_a(-0.0033110177610069513)),(to_sfixed_a(0.0004516126064117998)),(to_sfixed_a(0.006370408460497856)),(to_sfixed_a(0.00038312163087539375)),(to_sfixed_a(0.001555274473503232)),(to_sfixed_a(0.00011498384992592037)),(to_sfixed_a(-0.00015533195983152837)),(to_sfixed_a(-9.147744276560843e-05)),(to_sfixed_a(-0.03561635687947273)),(to_sfixed_a(0.19048549234867096)),(to_sfixed_a(-0.004226257558912039)),(to_sfixed_a(-6.523995398310944e-05)),(to_sfixed_a(-0.00171829538885504)),(to_sfixed_a(-0.6394211649894714)),(to_sfixed_a(-8.55687540024519e-05)),(to_sfixed_a(-7.46329315006733e-05)),(to_sfixed_a(0.0001630703336559236)),(to_sfixed_a(-0.00452842004597187)),(to_sfixed_a(-0.6872386336326599)),(to_sfixed_a(-0.0011479324894025922)),(to_sfixed_a(4.619270112016238e-05)),(to_sfixed_a(0.003499767277389765)),(to_sfixed_a(-0.0075935791246593)),(to_sfixed_a(1.803341910999734e-05)),(to_sfixed_a(2.208063961006701e-05)),(to_sfixed_a(0.0011382605880498886)),(to_sfixed_a(0.008892347104847431)),(to_sfixed_a(0.23815196752548218)),(to_sfixed_a(-9.946330828825012e-05)),(to_sfixed_a(0.3189428448677063)),(to_sfixed_a(-0.00010816290887305513)),(to_sfixed_a(-3.1756128009874374e-05)),(to_sfixed_a(-0.0012871134094893932)),(to_sfixed_a(-0.000353459850884974)),(to_sfixed_a(0.12230633199214935)),(to_sfixed_a(-0.003480740124359727)),(to_sfixed_a(-4.619643732439727e-06)),(to_sfixed_a(0.00838871393352747)),(to_sfixed_a(0.0001150349125964567)),(to_sfixed_a(-0.12307195365428925)),(to_sfixed_a(0.0004897206090390682)),(to_sfixed_a(0.0001300251460634172)),(to_sfixed_a(0.00230032647959888)),(to_sfixed_a(0.005024376790970564)),(to_sfixed_a(-0.005435531493276358)),(to_sfixed_a(-0.00022951760911382735)),(to_sfixed_a(0.00044962228275835514)),(to_sfixed_a(1.0619072781992145e-05)),(to_sfixed_a(0.34937939047813416)),(to_sfixed_a(-0.007880130782723427)),(to_sfixed_a(-8.237402653321624e-07)),(to_sfixed_a(-0.6791402697563171)),(to_sfixed_a(-0.0018805130384862423)),(to_sfixed_a(3.821952850557864e-05)),(to_sfixed_a(-0.15226466953754425)),(to_sfixed_a(0.020127305760979652)),(to_sfixed_a(-0.0001016719252220355)),(to_sfixed_a(0.2073073536157608)),(to_sfixed_a(-0.006319072097539902)),(to_sfixed_a(0.0005170594668015838)),(to_sfixed_a(-1.466362300561741e-05)),(to_sfixed_a(6.0673351981677115e-05)),(to_sfixed_a(0.013360516168177128)),(to_sfixed_a(1.492553565185517e-06)),(to_sfixed_a(-0.001573925488628447)),(to_sfixed_a(-6.180333002703264e-05)),(to_sfixed_a(0.0006583862123079598)),(to_sfixed_a(-1.5072413589223288e-05)),(to_sfixed_a(-0.0002514371299184859)),(to_sfixed_a(-1.3090946595184505e-05)),(to_sfixed_a(-2.9522903787437826e-05)),(to_sfixed_a(0.0001291202788706869)),(to_sfixed_a(0.001876938040368259)),(to_sfixed_a(0.0028040683828294277)),(to_sfixed_a(6.958944140933454e-07)),(to_sfixed_a(0.0017900608945637941)),(to_sfixed_a(-0.18179234862327576)),(to_sfixed_a(4.630272451322526e-05)),(to_sfixed_a(0.0001990840391954407)),(to_sfixed_a(6.67073909426108e-05)),(to_sfixed_a(-0.0002647987275850028)),(to_sfixed_a(0.007440790068358183)),(to_sfixed_a(0.39657700061798096)),(to_sfixed_a(-0.00016759902064222842)),(to_sfixed_a(-0.3843412697315216)),(to_sfixed_a(0.00020573334768414497)),(to_sfixed_a(6.431753718061373e-05)),(to_sfixed_a(0.06814717501401901)),(to_sfixed_a(0.00010523635137360543)),(to_sfixed_a(0.0010121422819793224)),(to_sfixed_a(9.283973486162722e-05)),(to_sfixed_a(5.688726560038049e-06)),(to_sfixed_a(0.00014620166621170938)),(to_sfixed_a(-0.00011206661292817444)),(to_sfixed_a(-0.2720480263233185)),(to_sfixed_a(-0.000149753934238106)),(to_sfixed_a(1.2977507140021771e-06)),(to_sfixed_a(0.0064856200478971004)),(to_sfixed_a(0.004601308144629002)),(to_sfixed_a(1.3082441000733525e-05)),(to_sfixed_a(1.6929647244978696e-05)),(to_sfixed_a(0.0001134937338065356)),(to_sfixed_a(0.0001062298979377374)),(to_sfixed_a(2.2294989321380854e-06)),(to_sfixed_a(-0.0021274916362017393)),(to_sfixed_a(-0.031660474836826324)),(to_sfixed_a(-0.00015326541324611753)),(to_sfixed_a(-9.401427814736962e-05)),(to_sfixed_a(0.013737461529672146)),(to_sfixed_a(0.0024652283173054457)),(to_sfixed_a(0.0001553750626044348)),(to_sfixed_a(4.723740494227968e-05)),(to_sfixed_a(0.00016661763947922736)),(to_sfixed_a(-4.520990842138417e-05)),(to_sfixed_a(-0.0001963978575076908)),(to_sfixed_a(-4.237866960465908e-05)),(to_sfixed_a(-0.25632497668266296)),(to_sfixed_a(5.279892866383307e-05)),(to_sfixed_a(8.053703641053289e-05)),(to_sfixed_a(-0.00012698333011940122)),(to_sfixed_a(-0.0001508627610746771)),(to_sfixed_a(0.0033893603831529617)),(to_sfixed_a(3.123658098047599e-05)),(to_sfixed_a(-0.00014760592603124678)),(to_sfixed_a(0.0006677461205981672)),(to_sfixed_a(-6.350317562464625e-06)),(to_sfixed_a(5.689915269613266e-05)),(to_sfixed_a(0.23900353908538818)),(to_sfixed_a(2.1611558622680604e-05)),(to_sfixed_a(0.0033478448167443275)),(to_sfixed_a(0.00010778934665722772)),(to_sfixed_a(-6.367372407112271e-07)),(to_sfixed_a(-4.794525739271194e-05)),(to_sfixed_a(0.00016721492283977568)),(to_sfixed_a(-0.0019646508153527975)),(to_sfixed_a(0.0019512304570525885)),(to_sfixed_a(0.009127690456807613)),(to_sfixed_a(-0.0047969939187169075)),(to_sfixed_a(-7.169906166382134e-05)),(to_sfixed_a(-0.0009559452882967889)),(to_sfixed_a(-8.663279004395008e-06)),(to_sfixed_a(3.559797187335789e-05)),(to_sfixed_a(-0.05918155238032341)),(to_sfixed_a(0.26669415831565857)),(to_sfixed_a(0.0007713051163591444)),(to_sfixed_a(-0.00015077501302585006)),(to_sfixed_a(0.03018728829920292)),(to_sfixed_a(-0.00018662636284716427)),(to_sfixed_a(0.0031101536005735397)),(to_sfixed_a(0.01168828271329403)),(to_sfixed_a(0.0013539483770728111)),(to_sfixed_a(0.2904038429260254)),(to_sfixed_a(0.0007009030668996274)),(to_sfixed_a(-0.005256348289549351)),(to_sfixed_a(0.00010742879385361448)),(to_sfixed_a(4.59961338492576e-05)),(to_sfixed_a(1.0797048162203282e-06)),(to_sfixed_a(-0.00012935427366755903)),(to_sfixed_a(0.004408671986311674)),(to_sfixed_a(-0.0002705272054299712)),(to_sfixed_a(0.002347331028431654)),(to_sfixed_a(0.003972579725086689)),(to_sfixed_a(0.0024149215314537287)),(to_sfixed_a(-0.00011323828221065924)),(to_sfixed_a(-0.000322375213727355)),(to_sfixed_a(0.5259491801261902)),(to_sfixed_a(6.782356649637222e-06)),(to_sfixed_a(-0.010910495184361935)),(to_sfixed_a(-7.121037924662232e-05)),(to_sfixed_a(0.41466623544692993)),(to_sfixed_a(0.00433423463255167)),(to_sfixed_a(-0.00011374738096492365)),(to_sfixed_a(-3.1205054256133735e-06)),(to_sfixed_a(0.00015731426537968218)),(to_sfixed_a(1.2339995009824634e-05)),(to_sfixed_a(0.00016764143947511911)),(to_sfixed_a(-0.00010411131370346993)),(to_sfixed_a(0.0037110501434653997)),(to_sfixed_a(-0.42786189913749695)),(to_sfixed_a(-0.0903339609503746)),(to_sfixed_a(0.029375523328781128)),(to_sfixed_a(0.026684189215302467)),(to_sfixed_a(0.146108478307724)),(to_sfixed_a(1.337594585493207e-05)),(to_sfixed_a(-7.140538946259767e-05)),(to_sfixed_a(3.857155388686806e-05)),(to_sfixed_a(0.00024341090465895832)),(to_sfixed_a(-0.00019121075456496328)),(to_sfixed_a(0.23286154866218567)),(to_sfixed_a(0.020073292776942253)),(to_sfixed_a(0.00533608254045248)),(to_sfixed_a(0.00010807272337842733)),(to_sfixed_a(-4.5136075641494244e-05)),(to_sfixed_a(7.844355423003435e-07)),(to_sfixed_a(0.00012024734314763919)),(to_sfixed_a(-0.004881718661636114)),(to_sfixed_a(-0.28512677550315857)),(to_sfixed_a(2.4316956114489585e-05)),(to_sfixed_a(6.335030047921464e-05)),(to_sfixed_a(-6.808704347349703e-05)),(to_sfixed_a(-0.008550775237381458)),(to_sfixed_a(0.0018997048027813435)),(to_sfixed_a(-0.41743335127830505)),(to_sfixed_a(-0.00019268676987849176)),(to_sfixed_a(-3.140476837870665e-05)),(to_sfixed_a(5.659809539793059e-05)),(to_sfixed_a(0.0007627304876223207)),(to_sfixed_a(0.0002706774102989584)),(to_sfixed_a(0.005595676600933075)),(to_sfixed_a(0.00018280852236784995)),(to_sfixed_a(0.24158605933189392)),(to_sfixed_a(8.976461685961112e-05)),(to_sfixed_a(-0.5430245995521545)),(to_sfixed_a(-0.00021838920656591654)),(to_sfixed_a(-0.47016051411628723)),(to_sfixed_a(0.00013425221550278366)),(to_sfixed_a(-0.24094916880130768)),(to_sfixed_a(0.022004403173923492)),(to_sfixed_a(0.13331453502178192)),(to_sfixed_a(-0.4607459008693695)),(to_sfixed_a(0.00020498478261288255)),(to_sfixed_a(0.0031904312781989574)),(to_sfixed_a(-0.005045244935899973)),(to_sfixed_a(0.0001296460977755487)),(to_sfixed_a(-0.004313134588301182)),(to_sfixed_a(0.00011311795969959348)),(to_sfixed_a(-0.00018335260392632335)),(to_sfixed_a(-0.2899489402770996)),(to_sfixed_a(0.007833744399249554)),(to_sfixed_a(7.444975926773623e-05)),(to_sfixed_a(0.00037939357571303844)),(to_sfixed_a(0.005614979192614555)),(to_sfixed_a(-0.0001876412716228515)),(to_sfixed_a(7.671956700505689e-05)),(to_sfixed_a(2.1841173293069005e-05)),(to_sfixed_a(-5.070982297183946e-05)),(to_sfixed_a(-0.00010188711166847497)),(to_sfixed_a(0.34344199299812317)),(to_sfixed_a(-0.00011200486915186048)),(to_sfixed_a(-0.00017728247621562332)),(to_sfixed_a(-2.998085255967453e-05)),(to_sfixed_a(0.28720614314079285)),(to_sfixed_a(-0.2825104296207428)),(to_sfixed_a(-9.602250065654516e-05)),(to_sfixed_a(-2.931860217358917e-05)),(to_sfixed_a(5.165158654563129e-06)),(to_sfixed_a(5.805821274407208e-05)),(to_sfixed_a(-0.3400416672229767)),(to_sfixed_a(-0.014581064693629742)),(to_sfixed_a(0.3056868612766266)),(to_sfixed_a(0.4743273854255676)),(to_sfixed_a(-0.3150135278701782)),(to_sfixed_a(-0.00011595715477596968)),(to_sfixed_a(0.00032071833265945315)),(to_sfixed_a(-8.772968431003392e-05)),(to_sfixed_a(0.0005795059842057526)),(to_sfixed_a(1.535075716674328e-05)),(to_sfixed_a(4.309775249566883e-06)),(to_sfixed_a(0.0024983943440020084)),(to_sfixed_a(0.19846582412719727)),(to_sfixed_a(-0.00021707713312935084)),(to_sfixed_a(-0.3912844657897949)),(to_sfixed_a(0.005712066777050495)),(to_sfixed_a(0.009306092746555805)),(to_sfixed_a(0.000488003104692325)),(to_sfixed_a(-0.00010208963067270815)),(to_sfixed_a(0.021091146394610405)),(to_sfixed_a(-0.006283010356128216)),(to_sfixed_a(-0.00807157438248396)),(to_sfixed_a(-3.5312375985085964e-05)),(to_sfixed_a(0.19027197360992432)),(to_sfixed_a(-0.03364526852965355)),(to_sfixed_a(-0.0005592625238932669)));

    constant weight_n2_45 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.11818280816078186)),(to_sfixed_a(-0.0013038166798651218)),(to_sfixed_a(-0.004834326449781656)),(to_sfixed_a(-0.00011280480248387903)),(to_sfixed_a(-0.0006293238839134574)),(to_sfixed_a(-5.411478196037933e-05)),(to_sfixed_a(-0.01925460435450077)),(to_sfixed_a(1.6492762370035052e-05)),(to_sfixed_a(-4.670593625633046e-05)),(to_sfixed_a(-3.740319880307652e-05)),(to_sfixed_a(0.0003782060230150819)),(to_sfixed_a(-0.004942871164530516)),(to_sfixed_a(-0.0039819679223001)),(to_sfixed_a(0.29564738273620605)),(to_sfixed_a(-7.646431913599372e-05)),(to_sfixed_a(-4.74173721158877e-05)),(to_sfixed_a(0.0010526541154831648)),(to_sfixed_a(4.43633362010587e-05)),(to_sfixed_a(-0.35693788528442383)),(to_sfixed_a(0.10530120879411697)),(to_sfixed_a(0.0002464476856403053)),(to_sfixed_a(3.959426248911768e-05)),(to_sfixed_a(-7.737616397207603e-05)),(to_sfixed_a(-0.0022216413635760546)),(to_sfixed_a(-0.008816931396722794)),(to_sfixed_a(-0.5128848552703857)),(to_sfixed_a(0.00016587742720730603)),(to_sfixed_a(-7.04186677467078e-05)),(to_sfixed_a(-0.0019542076624929905)),(to_sfixed_a(5.729949043598026e-05)),(to_sfixed_a(-0.000987378298304975)),(to_sfixed_a(-9.95281880022958e-07)),(to_sfixed_a(0.291587233543396)),(to_sfixed_a(6.392288923962042e-05)),(to_sfixed_a(-0.00010781313176266849)),(to_sfixed_a(-0.00017241243040189147)),(to_sfixed_a(0.22381281852722168)),(to_sfixed_a(0.0003393166116438806)),(to_sfixed_a(-0.08060362935066223)),(to_sfixed_a(-6.571660924237221e-05)),(to_sfixed_a(-0.01335118617862463)),(to_sfixed_a(-0.006139141973108053)),(to_sfixed_a(-2.296115053468384e-05)),(to_sfixed_a(0.0001510970323579386)),(to_sfixed_a(-0.0009227970149368048)),(to_sfixed_a(0.48891741037368774)),(to_sfixed_a(0.008809893392026424)),(to_sfixed_a(0.0018681687070056796)),(to_sfixed_a(0.00041349715320393443)),(to_sfixed_a(-0.010268143378198147)),(to_sfixed_a(-0.16082504391670227)),(to_sfixed_a(-0.00010067808034364134)),(to_sfixed_a(4.71786770503968e-05)),(to_sfixed_a(-0.003536899806931615)),(to_sfixed_a(-0.0023073761258274317)),(to_sfixed_a(0.3411167562007904)),(to_sfixed_a(-0.00015590706607326865)),(to_sfixed_a(0.003886342281475663)),(to_sfixed_a(4.4452732254285365e-05)),(to_sfixed_a(0.00029373951838351786)),(to_sfixed_a(0.0008871892932802439)),(to_sfixed_a(0.00023205159232020378)),(to_sfixed_a(-2.08538185688667e-05)),(to_sfixed_a(-0.18287348747253418)),(to_sfixed_a(-0.00015231006545946002)),(to_sfixed_a(-8.368175622308627e-05)),(to_sfixed_a(0.0001162703410955146)),(to_sfixed_a(-0.004878444597125053)),(to_sfixed_a(0.007596383336931467)),(to_sfixed_a(-0.00010078707418870181)),(to_sfixed_a(-0.08817741274833679)),(to_sfixed_a(0.018764270469546318)),(to_sfixed_a(0.04705525189638138)),(to_sfixed_a(-4.832191189052537e-05)),(to_sfixed_a(-7.066693797241896e-05)),(to_sfixed_a(-1.869532570708543e-05)),(to_sfixed_a(0.0014380011707544327)),(to_sfixed_a(0.21062147617340088)),(to_sfixed_a(-0.00016639893874526024)),(to_sfixed_a(0.20559756457805634)),(to_sfixed_a(-0.001416739891283214)),(to_sfixed_a(-8.38537816889584e-05)),(to_sfixed_a(-0.005547000095248222)),(to_sfixed_a(-0.0020840733777731657)),(to_sfixed_a(-6.916416896274313e-05)),(to_sfixed_a(0.0016020371112972498)),(to_sfixed_a(0.1619851142168045)),(to_sfixed_a(-0.001969042466953397)),(to_sfixed_a(-6.0079535614931956e-05)),(to_sfixed_a(-6.313207995845005e-05)),(to_sfixed_a(0.011746710166335106)),(to_sfixed_a(0.00011453316255938262)),(to_sfixed_a(-8.999270357890055e-05)),(to_sfixed_a(-0.00021586506045423448)),(to_sfixed_a(-0.0013582648243755102)),(to_sfixed_a(0.00015109841478988528)),(to_sfixed_a(-6.158681208034977e-05)),(to_sfixed_a(-0.00020178747945465147)),(to_sfixed_a(-0.00010610454773996025)),(to_sfixed_a(6.145636143628508e-05)),(to_sfixed_a(0.2495703399181366)),(to_sfixed_a(0.0012185585219413042)),(to_sfixed_a(4.633697244571522e-06)),(to_sfixed_a(0.23453344404697418)),(to_sfixed_a(0.129976287484169)),(to_sfixed_a(0.0011960233096033335)),(to_sfixed_a(-9.315173520008102e-05)),(to_sfixed_a(-5.172316377866082e-05)),(to_sfixed_a(-0.00010244513396173716)),(to_sfixed_a(0.0011855850461870432)),(to_sfixed_a(-0.0006106624496169388)),(to_sfixed_a(-0.0001859617914306)),(to_sfixed_a(-0.004563146736472845)),(to_sfixed_a(0.0001612472115084529)),(to_sfixed_a(4.237094253767282e-05)),(to_sfixed_a(0.21986940503120422)),(to_sfixed_a(5.818644422106445e-05)),(to_sfixed_a(-0.006715106312185526)),(to_sfixed_a(8.415496995439753e-05)),(to_sfixed_a(0.3278736174106598)),(to_sfixed_a(-0.00028679397655650973)),(to_sfixed_a(-7.142525282688439e-05)),(to_sfixed_a(-0.4304850995540619)),(to_sfixed_a(0.00011747124517569318)),(to_sfixed_a(-5.888140731258318e-05)),(to_sfixed_a(-0.2658671438694)),(to_sfixed_a(-0.47942253947257996)),(to_sfixed_a(0.00016336685803253204)),(to_sfixed_a(0.00010494503658264875)),(to_sfixed_a(-4.477202310226858e-06)),(to_sfixed_a(-0.00018892424122896045)),(to_sfixed_a(-4.3170861317776144e-05)),(to_sfixed_a(0.000315213983412832)),(to_sfixed_a(-0.010809014551341534)),(to_sfixed_a(-0.00041871104622259736)),(to_sfixed_a(4.7475761675741524e-05)),(to_sfixed_a(-0.005990632344037294)),(to_sfixed_a(0.00023806867829989642)),(to_sfixed_a(-6.352181662805378e-05)),(to_sfixed_a(-7.174437632784247e-05)),(to_sfixed_a(-0.00012255598267074674)),(to_sfixed_a(6.12129078945145e-05)),(to_sfixed_a(0.000152383727254346)),(to_sfixed_a(-0.32105201482772827)),(to_sfixed_a(0.0018646626267582178)),(to_sfixed_a(6.472531822510064e-06)),(to_sfixed_a(0.0007793367258273065)),(to_sfixed_a(6.806074816267937e-05)),(to_sfixed_a(-2.420041710138321e-06)),(to_sfixed_a(0.0038080126978456974)),(to_sfixed_a(-5.8452213124837726e-05)),(to_sfixed_a(4.9423324526287615e-05)),(to_sfixed_a(0.0003357941750437021)),(to_sfixed_a(-9.849361958913505e-05)),(to_sfixed_a(2.290062911924906e-05)),(to_sfixed_a(0.13055235147476196)),(to_sfixed_a(0.00014766522508580238)),(to_sfixed_a(0.0008632222888991237)),(to_sfixed_a(-0.00018586491933092475)),(to_sfixed_a(-6.784546712879092e-05)),(to_sfixed_a(3.89518536394462e-05)),(to_sfixed_a(-9.883947495836765e-05)),(to_sfixed_a(-0.003833328140899539)),(to_sfixed_a(-0.0032476589549332857)),(to_sfixed_a(0.0020098660606890917)),(to_sfixed_a(-0.08569978177547455)),(to_sfixed_a(-0.0001290266664000228)),(to_sfixed_a(0.13551238179206848)),(to_sfixed_a(-6.967233639443293e-05)),(to_sfixed_a(0.00018982027540914714)),(to_sfixed_a(0.003712985198944807)),(to_sfixed_a(0.0014711474068462849)),(to_sfixed_a(-0.002971042413264513)),(to_sfixed_a(-3.190372444805689e-05)),(to_sfixed_a(0.007100480608642101)),(to_sfixed_a(0.00013246758317109197)),(to_sfixed_a(-0.23673057556152344)),(to_sfixed_a(0.002730662003159523)),(to_sfixed_a(0.34085744619369507)),(to_sfixed_a(-0.00294810114428401)),(to_sfixed_a(0.0006851834477856755)),(to_sfixed_a(0.0061001162976026535)),(to_sfixed_a(-0.00025645739515312016)),(to_sfixed_a(1.2524993508122861e-05)),(to_sfixed_a(5.559177225222811e-06)),(to_sfixed_a(-0.0024780158419162035)),(to_sfixed_a(-0.6672622561454773)),(to_sfixed_a(-0.0050354921258986)),(to_sfixed_a(-0.000701544398907572)),(to_sfixed_a(0.0010124810505658388)),(to_sfixed_a(-0.008479055017232895)),(to_sfixed_a(0.00046109588583931327)),(to_sfixed_a(-0.003460073843598366)),(to_sfixed_a(-0.00010408402886241674)),(to_sfixed_a(0.000282888620859012)),(to_sfixed_a(0.1309032440185547)),(to_sfixed_a(8.90491355676204e-05)),(to_sfixed_a(0.001978446962311864)),(to_sfixed_a(-0.2318652719259262)),(to_sfixed_a(-0.00021289548021741211)),(to_sfixed_a(-0.0001665326562942937)),(to_sfixed_a(6.52307498967275e-05)),(to_sfixed_a(3.56146483682096e-05)),(to_sfixed_a(-1.1982221622020006e-05)),(to_sfixed_a(5.680412868969142e-07)),(to_sfixed_a(-0.2104540765285492)),(to_sfixed_a(-0.004008103162050247)),(to_sfixed_a(-0.01923416368663311)),(to_sfixed_a(0.0014567531179636717)),(to_sfixed_a(0.0026247145142406225)),(to_sfixed_a(0.003088192315772176)),(to_sfixed_a(9.539422899251804e-05)),(to_sfixed_a(7.140845264075324e-05)),(to_sfixed_a(9.298442455474287e-05)),(to_sfixed_a(2.9792470741085708e-05)),(to_sfixed_a(1.8286678823642433e-05)),(to_sfixed_a(-0.0004670803318731487)),(to_sfixed_a(-0.004660366103053093)),(to_sfixed_a(0.003167166607454419)),(to_sfixed_a(-6.573605787707493e-06)),(to_sfixed_a(7.817296136636287e-05)),(to_sfixed_a(-6.75602350383997e-05)),(to_sfixed_a(2.657616278156638e-05)),(to_sfixed_a(-0.00508258817717433)),(to_sfixed_a(-0.0025913133285939693)),(to_sfixed_a(6.120166654000059e-05)),(to_sfixed_a(7.264126179507002e-05)),(to_sfixed_a(-3.4657827200135216e-05)),(to_sfixed_a(-0.6179602146148682)),(to_sfixed_a(0.5317504405975342)),(to_sfixed_a(-0.0009388932376168668)),(to_sfixed_a(-6.811208731960505e-05)),(to_sfixed_a(0.00020503689302131534)),(to_sfixed_a(-6.753468187525868e-05)),(to_sfixed_a(-0.37491753697395325)),(to_sfixed_a(0.3303464651107788)),(to_sfixed_a(-0.2555236220359802)),(to_sfixed_a(7.081230432959273e-05)),(to_sfixed_a(0.17825469374656677)),(to_sfixed_a(0.00029006306431256235)),(to_sfixed_a(-0.414975106716156)),(to_sfixed_a(-0.00019928408437408507)),(to_sfixed_a(0.23711548745632172)),(to_sfixed_a(-6.156692688819021e-05)),(to_sfixed_a(-0.20844592154026031)),(to_sfixed_a(0.004008050542324781)),(to_sfixed_a(0.004837299231439829)),(to_sfixed_a(0.00025821069721132517)),(to_sfixed_a(-1.7850878066383302e-05)),(to_sfixed_a(-0.0018075674306601286)),(to_sfixed_a(-0.0008769258856773376)),(to_sfixed_a(-0.00017090968322008848)),(to_sfixed_a(-0.006381602957844734)),(to_sfixed_a(0.00012694421457126737)),(to_sfixed_a(-0.0002935697848442942)),(to_sfixed_a(0.003606863785535097)),(to_sfixed_a(-0.008738130331039429)),(to_sfixed_a(-0.00011218790314160287)),(to_sfixed_a(-0.0001584486453793943)),(to_sfixed_a(7.311283843591809e-05)),(to_sfixed_a(0.00024803151609376073)),(to_sfixed_a(0.00035213999217376113)),(to_sfixed_a(-3.1010979000711814e-05)),(to_sfixed_a(0.0001401093031745404)),(to_sfixed_a(-0.00012691994197666645)),(to_sfixed_a(6.67861313559115e-05)),(to_sfixed_a(-6.657051562797278e-05)),(to_sfixed_a(0.0001141276370617561)),(to_sfixed_a(4.462647848413326e-05)),(to_sfixed_a(0.00196842267177999)),(to_sfixed_a(-0.004468111786991358)),(to_sfixed_a(-8.827639976516366e-05)),(to_sfixed_a(6.697280332446098e-05)),(to_sfixed_a(3.142231435049325e-07)),(to_sfixed_a(0.00026756033184938133)),(to_sfixed_a(0.0019651451148092747)),(to_sfixed_a(0.0019206214928999543)),(to_sfixed_a(0.21009540557861328)),(to_sfixed_a(0.005389922298491001)),(to_sfixed_a(-0.02262292243540287)),(to_sfixed_a(4.390021786093712e-06)),(to_sfixed_a(-0.00012967720977030694)),(to_sfixed_a(-5.623815377475694e-05)),(to_sfixed_a(-0.0025102419313043356)),(to_sfixed_a(0.00010397753794677556)),(to_sfixed_a(-2.6938985683955252e-05)),(to_sfixed_a(-0.005177405662834644)),(to_sfixed_a(0.001605871831998229)),(to_sfixed_a(8.822025847621262e-05)),(to_sfixed_a(-0.0009158133761957288)),(to_sfixed_a(0.0013220451073721051)),(to_sfixed_a(0.0007547604036517441)),(to_sfixed_a(0.36186957359313965)),(to_sfixed_a(0.00020367479010019451)),(to_sfixed_a(0.0004831702681258321)),(to_sfixed_a(0.0033188958186656237)),(to_sfixed_a(0.0016711672069504857)),(to_sfixed_a(0.00024232082068920135)),(to_sfixed_a(0.40176641941070557)),(to_sfixed_a(-0.006357159931212664)),(to_sfixed_a(-0.0010956055484712124)));

    constant weight_n2_46 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.29100531339645386)),(to_sfixed_a(-0.002723144832998514)),(to_sfixed_a(-0.0003011623921338469)),(to_sfixed_a(6.63755345158279e-05)),(to_sfixed_a(-0.006975517608225346)),(to_sfixed_a(-4.619266837835312e-05)),(to_sfixed_a(0.0005793426535092294)),(to_sfixed_a(-0.0001471949217375368)),(to_sfixed_a(-6.908199429744855e-05)),(to_sfixed_a(0.00010469370317878202)),(to_sfixed_a(0.00016836152644827962)),(to_sfixed_a(0.008360577747225761)),(to_sfixed_a(0.0001236082025570795)),(to_sfixed_a(0.0028468691743910313)),(to_sfixed_a(4.5255710574565455e-05)),(to_sfixed_a(0.00013344548642635345)),(to_sfixed_a(-0.0027980045415461063)),(to_sfixed_a(-0.00023159629199653864)),(to_sfixed_a(0.0012856345856562257)),(to_sfixed_a(-0.16746023297309875)),(to_sfixed_a(2.4051405489444733e-06)),(to_sfixed_a(0.0001299698487855494)),(to_sfixed_a(0.005187110044062138)),(to_sfixed_a(0.005795411765575409)),(to_sfixed_a(-0.006328332703560591)),(to_sfixed_a(0.006850182078778744)),(to_sfixed_a(-0.00031268454040400684)),(to_sfixed_a(2.737929389695637e-05)),(to_sfixed_a(0.00022148493735585362)),(to_sfixed_a(-7.4281851993873715e-06)),(to_sfixed_a(0.6049767136573792)),(to_sfixed_a(0.00019136090122628957)),(to_sfixed_a(-0.0009089091327041388)),(to_sfixed_a(0.00015393391367979348)),(to_sfixed_a(5.6783661420922726e-05)),(to_sfixed_a(2.95431527774781e-06)),(to_sfixed_a(-0.16270773112773895)),(to_sfixed_a(0.3752192556858063)),(to_sfixed_a(0.0016142267268151045)),(to_sfixed_a(-0.00012887064076494426)),(to_sfixed_a(0.011056727729737759)),(to_sfixed_a(0.006409918889403343)),(to_sfixed_a(1.850748958531767e-05)),(to_sfixed_a(0.00018218523473478854)),(to_sfixed_a(-0.004719426389783621)),(to_sfixed_a(-0.0003056564019061625)),(to_sfixed_a(-0.00166635075584054)),(to_sfixed_a(-0.002340503968298435)),(to_sfixed_a(0.00015911126683931798)),(to_sfixed_a(-0.0016449510585516691)),(to_sfixed_a(0.3653070330619812)),(to_sfixed_a(-0.0030877080280333757)),(to_sfixed_a(6.925790512468666e-05)),(to_sfixed_a(-0.4194648563861847)),(to_sfixed_a(0.014863580465316772)),(to_sfixed_a(-0.42424681782722473)),(to_sfixed_a(-5.071044142823666e-06)),(to_sfixed_a(0.0035947721917182207)),(to_sfixed_a(-0.0001340504240943119)),(to_sfixed_a(-0.00011329421249683946)),(to_sfixed_a(0.012806328013539314)),(to_sfixed_a(0.00724710151553154)),(to_sfixed_a(0.00012016540131298825)),(to_sfixed_a(0.4024008810520172)),(to_sfixed_a(1.784756750566885e-05)),(to_sfixed_a(-0.204468235373497)),(to_sfixed_a(-8.367547707166523e-05)),(to_sfixed_a(-0.036336954683065414)),(to_sfixed_a(-5.924295692238957e-05)),(to_sfixed_a(-2.7939866413362324e-05)),(to_sfixed_a(-0.06275945156812668)),(to_sfixed_a(-0.006936586927622557)),(to_sfixed_a(-0.0024676891043782234)),(to_sfixed_a(1.4561475836671889e-05)),(to_sfixed_a(-9.285857959184796e-05)),(to_sfixed_a(-4.2185638449154794e-05)),(to_sfixed_a(0.07125478982925415)),(to_sfixed_a(-0.01147963386029005)),(to_sfixed_a(-0.00011554003867786378)),(to_sfixed_a(0.016608862206339836)),(to_sfixed_a(-0.0009525521891191602)),(to_sfixed_a(-1.52934153447859e-05)),(to_sfixed_a(-0.10662005841732025)),(to_sfixed_a(-0.0035427215043455362)),(to_sfixed_a(0.00020169139315839857)),(to_sfixed_a(-0.00011948923201998696)),(to_sfixed_a(-0.00018548412481322885)),(to_sfixed_a(-8.365210305782966e-06)),(to_sfixed_a(-0.00037600757787004113)),(to_sfixed_a(-1.2466229236451909e-05)),(to_sfixed_a(-0.8507285714149475)),(to_sfixed_a(-0.00014822240336798131)),(to_sfixed_a(0.0001504191750427708)),(to_sfixed_a(1.1314208677504212e-05)),(to_sfixed_a(0.00549407210201025)),(to_sfixed_a(9.962379408534616e-06)),(to_sfixed_a(-0.00017427594866603613)),(to_sfixed_a(0.00015888584312051535)),(to_sfixed_a(-4.758105569635518e-05)),(to_sfixed_a(-1.2013570085400715e-06)),(to_sfixed_a(0.03322717547416687)),(to_sfixed_a(-0.0001497053453931585)),(to_sfixed_a(-1.999516098294407e-05)),(to_sfixed_a(0.21448910236358643)),(to_sfixed_a(-0.0022915720473974943)),(to_sfixed_a(0.3139897286891937)),(to_sfixed_a(0.00010327782365493476)),(to_sfixed_a(-3.238302451791242e-05)),(to_sfixed_a(0.0002636928402353078)),(to_sfixed_a(-0.0036099241115152836)),(to_sfixed_a(0.006327051669359207)),(to_sfixed_a(0.00012658353080041707)),(to_sfixed_a(-0.0043557183817029)),(to_sfixed_a(0.00011182680464116856)),(to_sfixed_a(4.046538379043341e-05)),(to_sfixed_a(-0.0027203222271054983)),(to_sfixed_a(0.0025316248647868633)),(to_sfixed_a(-0.00041190299089066684)),(to_sfixed_a(-0.00020804052473977208)),(to_sfixed_a(-0.002359686652198434)),(to_sfixed_a(-0.00026550376787781715)),(to_sfixed_a(6.092615512898192e-05)),(to_sfixed_a(0.00011161943257320672)),(to_sfixed_a(-6.723376282025129e-05)),(to_sfixed_a(9.218818013323471e-05)),(to_sfixed_a(0.0006324296118691564)),(to_sfixed_a(-0.0057097868993878365)),(to_sfixed_a(0.00023285247152671218)),(to_sfixed_a(3.209012720617466e-05)),(to_sfixed_a(-5.072351632406935e-05)),(to_sfixed_a(4.421470293891616e-05)),(to_sfixed_a(6.52357775834389e-05)),(to_sfixed_a(-0.00025774873211048543)),(to_sfixed_a(0.28407588601112366)),(to_sfixed_a(-0.0002641983446665108)),(to_sfixed_a(0.00022228527814149857)),(to_sfixed_a(0.0029072058387100697)),(to_sfixed_a(7.512423326261342e-05)),(to_sfixed_a(0.0001649431069381535)),(to_sfixed_a(0.00029595589148811996)),(to_sfixed_a(-0.37339815497398376)),(to_sfixed_a(-1.622956187929958e-05)),(to_sfixed_a(2.429058076813817e-05)),(to_sfixed_a(-0.000336633762344718)),(to_sfixed_a(-0.0008321244386024773)),(to_sfixed_a(0.0004610999603755772)),(to_sfixed_a(0.00124944350682199)),(to_sfixed_a(-0.0001643760479055345)),(to_sfixed_a(-0.00017937285883817822)),(to_sfixed_a(-0.0026597788091748953)),(to_sfixed_a(-0.0004445167141966522)),(to_sfixed_a(-8.184974285541102e-05)),(to_sfixed_a(0.26004406809806824)),(to_sfixed_a(0.00014589127385988832)),(to_sfixed_a(-0.0002506644232198596)),(to_sfixed_a(0.4104473888874054)),(to_sfixed_a(0.0002935619850177318)),(to_sfixed_a(0.1685391664505005)),(to_sfixed_a(8.216104470193386e-05)),(to_sfixed_a(-0.00017523960559628904)),(to_sfixed_a(6.075820783735253e-05)),(to_sfixed_a(-4.336061829235405e-05)),(to_sfixed_a(0.4543534517288208)),(to_sfixed_a(-0.10287604480981827)),(to_sfixed_a(0.033452633768320084)),(to_sfixed_a(0.5981802344322205)),(to_sfixed_a(-0.00024404327268712223)),(to_sfixed_a(1.959187284228392e-05)),(to_sfixed_a(-4.383530904306099e-05)),(to_sfixed_a(0.0001260380377061665)),(to_sfixed_a(0.00418707262724638)),(to_sfixed_a(0.0010517562041059136)),(to_sfixed_a(-0.000974050082731992)),(to_sfixed_a(-2.1087689674459398e-06)),(to_sfixed_a(0.004654897842556238)),(to_sfixed_a(-0.00032055351766757667)),(to_sfixed_a(-0.00046551611740142107)),(to_sfixed_a(0.5130948424339294)),(to_sfixed_a(-0.24661165475845337)),(to_sfixed_a(0.005553378723561764)),(to_sfixed_a(0.00025269004981964827)),(to_sfixed_a(-0.046560827642679214)),(to_sfixed_a(-0.0001683027803665027)),(to_sfixed_a(7.069003186188638e-05)),(to_sfixed_a(0.0004236674285493791)),(to_sfixed_a(0.008086401037871838)),(to_sfixed_a(0.2641581594944)),(to_sfixed_a(-0.161702960729599)),(to_sfixed_a(0.0038602007552981377)),(to_sfixed_a(0.36707931756973267)),(to_sfixed_a(-0.00010438838216941804)),(to_sfixed_a(-0.00015390968474093825)),(to_sfixed_a(0.035460419952869415)),(to_sfixed_a(0.0007566734566353261)),(to_sfixed_a(-0.00011376842303434387)),(to_sfixed_a(-0.004393777810037136)),(to_sfixed_a(-0.00012636801693588495)),(to_sfixed_a(0.2016240358352661)),(to_sfixed_a(-0.012874615378677845)),(to_sfixed_a(-1.4813209418207407e-05)),(to_sfixed_a(0.0002476298832334578)),(to_sfixed_a(-1.8392285710433498e-05)),(to_sfixed_a(-2.9694230761379004e-05)),(to_sfixed_a(-0.0002370034926570952)),(to_sfixed_a(4.435438313521445e-06)),(to_sfixed_a(0.0017456293571740389)),(to_sfixed_a(-0.127879798412323)),(to_sfixed_a(-0.2076028287410736)),(to_sfixed_a(0.01621408388018608)),(to_sfixed_a(-0.0005991060752421618)),(to_sfixed_a(-0.00012219294148962945)),(to_sfixed_a(0.00024274989846162498)),(to_sfixed_a(-7.665983139304444e-05)),(to_sfixed_a(-0.00018453187658451498)),(to_sfixed_a(-7.461522181984037e-05)),(to_sfixed_a(-7.11987740942277e-05)),(to_sfixed_a(-0.005158691667020321)),(to_sfixed_a(0.15387308597564697)),(to_sfixed_a(-0.13886044919490814)),(to_sfixed_a(6.21633225819096e-05)),(to_sfixed_a(0.00020468630827963352)),(to_sfixed_a(-7.852141425246373e-05)),(to_sfixed_a(-0.00024892244255170226)),(to_sfixed_a(0.001154493191279471)),(to_sfixed_a(-0.0037911420222371817)),(to_sfixed_a(6.608966941712424e-05)),(to_sfixed_a(6.529638631036505e-05)),(to_sfixed_a(-9.385003068018705e-07)),(to_sfixed_a(0.3200821876525879)),(to_sfixed_a(-0.2636938691139221)),(to_sfixed_a(-0.00035842976649291813)),(to_sfixed_a(0.00011671244283206761)),(to_sfixed_a(9.974234126275405e-05)),(to_sfixed_a(4.744111356558278e-05)),(to_sfixed_a(0.30035266280174255)),(to_sfixed_a(0.0063659329898655415)),(to_sfixed_a(0.011665833182632923)),(to_sfixed_a(0.00017479689267929643)),(to_sfixed_a(0.00016474726726301014)),(to_sfixed_a(0.00017080394900403917)),(to_sfixed_a(0.01796945370733738)),(to_sfixed_a(8.701699698576704e-05)),(to_sfixed_a(0.0003335624933242798)),(to_sfixed_a(-3.944485797546804e-06)),(to_sfixed_a(-0.0024530573282390833)),(to_sfixed_a(-0.0002291759301442653)),(to_sfixed_a(-0.13033781945705414)),(to_sfixed_a(-0.2645525336265564)),(to_sfixed_a(4.2527171899564564e-05)),(to_sfixed_a(-0.0014659998705610633)),(to_sfixed_a(0.00024665662203915417)),(to_sfixed_a(-0.00044638989493250847)),(to_sfixed_a(0.0001467389811296016)),(to_sfixed_a(2.0762268832186237e-05)),(to_sfixed_a(-0.0019354241667315364)),(to_sfixed_a(-0.0018794859061017632)),(to_sfixed_a(0.036639854311943054)),(to_sfixed_a(0.00010111099982168525)),(to_sfixed_a(7.17345392331481e-05)),(to_sfixed_a(0.00010042764915851876)),(to_sfixed_a(-0.0001693398371571675)),(to_sfixed_a(-0.001283678924664855)),(to_sfixed_a(7.859538163756952e-05)),(to_sfixed_a(8.835411790641956e-06)),(to_sfixed_a(-0.00010474491864442825)),(to_sfixed_a(0.05695132166147232)),(to_sfixed_a(-0.00018502341117709875)),(to_sfixed_a(8.020477253012359e-06)),(to_sfixed_a(2.360693906666711e-05)),(to_sfixed_a(-0.07058648020029068)),(to_sfixed_a(0.004686813335865736)),(to_sfixed_a(0.00023626491019967943)),(to_sfixed_a(6.231212319107726e-05)),(to_sfixed_a(7.019935583230108e-05)),(to_sfixed_a(0.000168251630384475)),(to_sfixed_a(0.017886318266391754)),(to_sfixed_a(0.24390269815921783)),(to_sfixed_a(0.29381895065307617)),(to_sfixed_a(-0.0003648450074251741)),(to_sfixed_a(0.0043732100166380405)),(to_sfixed_a(6.815665983594954e-05)),(to_sfixed_a(3.6771725717699155e-05)),(to_sfixed_a(-3.239980651414953e-05)),(to_sfixed_a(-0.0010488632833585143)),(to_sfixed_a(-3.816427488345653e-05)),(to_sfixed_a(-0.00014626866322942078)),(to_sfixed_a(-0.0007129278965294361)),(to_sfixed_a(0.0025336819235235453)),(to_sfixed_a(-5.7301760534755886e-05)),(to_sfixed_a(-0.029747983440756798)),(to_sfixed_a(0.0001723822351777926)),(to_sfixed_a(-0.0031888901721686125)),(to_sfixed_a(-0.5112093091011047)),(to_sfixed_a(-0.0002018249942921102)),(to_sfixed_a(-0.017639411613345146)),(to_sfixed_a(0.42751723527908325)),(to_sfixed_a(-0.1499665081501007)),(to_sfixed_a(-1.779975718818605e-06)),(to_sfixed_a(0.44539177417755127)),(to_sfixed_a(0.0004943907260894775)),(to_sfixed_a(0.4054794907569885)));

    constant weight_n2_47 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.3819226026535034)),(to_sfixed_a(0.00014152470976114273)),(to_sfixed_a(-0.0020625728648155928)),(to_sfixed_a(-7.243578875204548e-05)),(to_sfixed_a(-0.6002917289733887)),(to_sfixed_a(0.0001684638555161655)),(to_sfixed_a(0.09704626351594925)),(to_sfixed_a(-0.0001380286703351885)),(to_sfixed_a(1.5188161341939121e-06)),(to_sfixed_a(-8.677354344399646e-05)),(to_sfixed_a(-2.6272085960954428e-05)),(to_sfixed_a(0.002071739872917533)),(to_sfixed_a(0.00530533492565155)),(to_sfixed_a(-0.0013930010609328747)),(to_sfixed_a(-0.00011442331015132368)),(to_sfixed_a(0.0001459724153392017)),(to_sfixed_a(0.005047656130045652)),(to_sfixed_a(2.7657340979203582e-05)),(to_sfixed_a(0.004107220564037561)),(to_sfixed_a(-0.0005609930958598852)),(to_sfixed_a(-0.000301847408991307)),(to_sfixed_a(-0.00015742481627967209)),(to_sfixed_a(-0.0008601009612902999)),(to_sfixed_a(0.0006344971479848027)),(to_sfixed_a(0.29957273602485657)),(to_sfixed_a(-0.015737079083919525)),(to_sfixed_a(5.8066536439582705e-05)),(to_sfixed_a(3.548914537532255e-05)),(to_sfixed_a(0.00036056715180166066)),(to_sfixed_a(0.000104093698610086)),(to_sfixed_a(-0.34541401267051697)),(to_sfixed_a(6.338954699458554e-05)),(to_sfixed_a(0.01841946877539158)),(to_sfixed_a(-0.00016806001076474786)),(to_sfixed_a(3.240288788219914e-05)),(to_sfixed_a(-0.00014729709073435515)),(to_sfixed_a(0.37854471802711487)),(to_sfixed_a(-0.008921765722334385)),(to_sfixed_a(0.009520630352199078)),(to_sfixed_a(-0.00014962606655899435)),(to_sfixed_a(0.05496722832322121)),(to_sfixed_a(-0.0018448951886966825)),(to_sfixed_a(0.00045103931915946305)),(to_sfixed_a(6.942739128135145e-05)),(to_sfixed_a(0.0023826288525015116)),(to_sfixed_a(-0.2553250193595886)),(to_sfixed_a(0.0020495590288192034)),(to_sfixed_a(-0.000755783636122942)),(to_sfixed_a(0.00021629589900840074)),(to_sfixed_a(0.0021004467271268368)),(to_sfixed_a(0.0017594833625480533)),(to_sfixed_a(4.5013061026111245e-05)),(to_sfixed_a(-2.539590059313923e-05)),(to_sfixed_a(0.003532632952556014)),(to_sfixed_a(-0.22772030532360077)),(to_sfixed_a(0.0007900783093646169)),(to_sfixed_a(4.020195046905428e-05)),(to_sfixed_a(-0.020715754479169846)),(to_sfixed_a(-3.516109427437186e-05)),(to_sfixed_a(-0.00017358582408633083)),(to_sfixed_a(0.0001800484023988247)),(to_sfixed_a(-0.0016652164049446583)),(to_sfixed_a(-0.000184270873432979)),(to_sfixed_a(0.014756637625396252)),(to_sfixed_a(1.939140202011913e-05)),(to_sfixed_a(0.000855613499879837)),(to_sfixed_a(6.0264130297582597e-05)),(to_sfixed_a(-0.47292131185531616)),(to_sfixed_a(0.0045710098929703236)),(to_sfixed_a(0.000251673482125625)),(to_sfixed_a(0.012123754248023033)),(to_sfixed_a(0.004325964488089085)),(to_sfixed_a(0.0029713036492466927)),(to_sfixed_a(2.4371729523409158e-05)),(to_sfixed_a(-0.00017493439372628927)),(to_sfixed_a(-0.0001689687487669289)),(to_sfixed_a(0.1366082727909088)),(to_sfixed_a(0.004997251555323601)),(to_sfixed_a(-0.0001302915916312486)),(to_sfixed_a(-0.0027181857731193304)),(to_sfixed_a(0.0033408580347895622)),(to_sfixed_a(0.00015587439702358097)),(to_sfixed_a(-0.00021104683401063085)),(to_sfixed_a(-0.0038342310581356287)),(to_sfixed_a(-2.5460447432124056e-05)),(to_sfixed_a(0.0018682748777791858)),(to_sfixed_a(0.003022248623892665)),(to_sfixed_a(0.013704011216759682)),(to_sfixed_a(7.877540338085964e-05)),(to_sfixed_a(2.0559309632517397e-05)),(to_sfixed_a(-0.2618684470653534)),(to_sfixed_a(3.5375458537600935e-05)),(to_sfixed_a(0.0011558585101738572)),(to_sfixed_a(-8.00465713837184e-05)),(to_sfixed_a(-0.2221446931362152)),(to_sfixed_a(6.416478572646156e-05)),(to_sfixed_a(0.00031406874768435955)),(to_sfixed_a(0.00010221017873845994)),(to_sfixed_a(5.76642996747978e-05)),(to_sfixed_a(0.00015300011727958918)),(to_sfixed_a(0.0011162658920511603)),(to_sfixed_a(-0.0012936799321323633)),(to_sfixed_a(3.350935730850324e-05)),(to_sfixed_a(0.004485701210796833)),(to_sfixed_a(-0.000567088951356709)),(to_sfixed_a(-0.2647508680820465)),(to_sfixed_a(4.9239715735893697e-05)),(to_sfixed_a(4.848261596634984e-06)),(to_sfixed_a(7.090042345225811e-05)),(to_sfixed_a(0.007825701497495174)),(to_sfixed_a(0.009209498763084412)),(to_sfixed_a(-0.00013662301353178918)),(to_sfixed_a(-0.012086542323231697)),(to_sfixed_a(-6.449186184909195e-05)),(to_sfixed_a(-4.860905755776912e-05)),(to_sfixed_a(-0.02499077469110489)),(to_sfixed_a(0.003175707533955574)),(to_sfixed_a(0.00010568297875579447)),(to_sfixed_a(-7.131195161491632e-05)),(to_sfixed_a(0.004469454288482666)),(to_sfixed_a(9.83120480668731e-06)),(to_sfixed_a(-7.05847778590396e-05)),(to_sfixed_a(-0.019734730944037437)),(to_sfixed_a(0.00020029349252581596)),(to_sfixed_a(0.00012017529661534354)),(to_sfixed_a(0.009659882634878159)),(to_sfixed_a(0.24961313605308533)),(to_sfixed_a(-0.00015179663023445755)),(to_sfixed_a(3.436164843151346e-05)),(to_sfixed_a(-2.506781675037928e-05)),(to_sfixed_a(6.594053411390632e-05)),(to_sfixed_a(-6.881348235765472e-05)),(to_sfixed_a(-0.00020611472427845)),(to_sfixed_a(0.0059187444858253)),(to_sfixed_a(6.415629468392581e-05)),(to_sfixed_a(-5.55206133867614e-06)),(to_sfixed_a(-0.005498065613210201)),(to_sfixed_a(-0.24398966133594513)),(to_sfixed_a(-2.2095715394243598e-05)),(to_sfixed_a(5.858237273059785e-07)),(to_sfixed_a(-0.3657331168651581)),(to_sfixed_a(-4.35802576248534e-05)),(to_sfixed_a(-0.00031316454987972975)),(to_sfixed_a(-0.00012386984599288553)),(to_sfixed_a(-0.0012559995520859957)),(to_sfixed_a(-0.00013398914597928524)),(to_sfixed_a(-0.0007865680963732302)),(to_sfixed_a(6.295308412518352e-05)),(to_sfixed_a(5.264587525743991e-05)),(to_sfixed_a(0.0025695725344121456)),(to_sfixed_a(-4.992492904420942e-06)),(to_sfixed_a(0.00018032899242825806)),(to_sfixed_a(0.008636818267405033)),(to_sfixed_a(7.203831046354026e-06)),(to_sfixed_a(-0.00010078217746922746)),(to_sfixed_a(0.10078619420528412)),(to_sfixed_a(-1.6173376934602857e-05)),(to_sfixed_a(0.32716700434684753)),(to_sfixed_a(-4.164022175245918e-05)),(to_sfixed_a(0.00023262706235982478)),(to_sfixed_a(0.00011557650577742606)),(to_sfixed_a(0.00019460277690086514)),(to_sfixed_a(0.0026362952776253223)),(to_sfixed_a(0.003709173295646906)),(to_sfixed_a(0.25419121980667114)),(to_sfixed_a(0.34893640875816345)),(to_sfixed_a(-2.4807981390040368e-05)),(to_sfixed_a(-0.656957745552063)),(to_sfixed_a(7.81271155574359e-05)),(to_sfixed_a(0.00015922276361379772)),(to_sfixed_a(0.0042482600547373295)),(to_sfixed_a(-0.001056900480762124)),(to_sfixed_a(0.010860209353268147)),(to_sfixed_a(-5.751573189627379e-05)),(to_sfixed_a(0.05599258467555046)),(to_sfixed_a(0.002626137575134635)),(to_sfixed_a(-0.0013372490648180246)),(to_sfixed_a(-0.0006704666302539408)),(to_sfixed_a(-0.24640360474586487)),(to_sfixed_a(0.2999773621559143)),(to_sfixed_a(-0.0006433269591070712)),(to_sfixed_a(1.115284703701036e-05)),(to_sfixed_a(0.00011180752335349098)),(to_sfixed_a(2.226748620159924e-06)),(to_sfixed_a(-4.801556497113779e-05)),(to_sfixed_a(0.0005402277456596494)),(to_sfixed_a(0.2546735107898712)),(to_sfixed_a(-0.0011690679239109159)),(to_sfixed_a(0.0019313963130116463)),(to_sfixed_a(0.0030252868309617043)),(to_sfixed_a(0.005888015031814575)),(to_sfixed_a(-0.00011352464207448065)),(to_sfixed_a(-0.00044647487811744213)),(to_sfixed_a(0.002430162625387311)),(to_sfixed_a(4.8699192120693624e-05)),(to_sfixed_a(-0.27884340286254883)),(to_sfixed_a(-0.00014844922407064587)),(to_sfixed_a(0.2402818500995636)),(to_sfixed_a(-0.11025463789701462)),(to_sfixed_a(1.7770842532627285e-05)),(to_sfixed_a(-0.00019270549819339067)),(to_sfixed_a(-0.00011423085379647091)),(to_sfixed_a(-5.168813731870614e-05)),(to_sfixed_a(4.4444441300584e-05)),(to_sfixed_a(-5.5279968364629894e-05)),(to_sfixed_a(0.00016253971261903644)),(to_sfixed_a(0.40086236596107483)),(to_sfixed_a(0.0009251049486920238)),(to_sfixed_a(0.0011290523689240217)),(to_sfixed_a(0.36809781193733215)),(to_sfixed_a(0.0006917011924088001)),(to_sfixed_a(1.657813845667988e-05)),(to_sfixed_a(1.5256497135851532e-05)),(to_sfixed_a(6.013255551806651e-05)),(to_sfixed_a(-2.8911250410601497e-05)),(to_sfixed_a(-0.0001516241900390014)),(to_sfixed_a(0.004147510044276714)),(to_sfixed_a(0.005517643876373768)),(to_sfixed_a(-0.01044002827256918)),(to_sfixed_a(-0.00015040652942843735)),(to_sfixed_a(-0.00015263407840393484)),(to_sfixed_a(3.3514254027977586e-05)),(to_sfixed_a(0.00028674938948825)),(to_sfixed_a(-0.00012583677016664296)),(to_sfixed_a(0.18464641273021698)),(to_sfixed_a(6.353812932502478e-05)),(to_sfixed_a(-0.00044505810365080833)),(to_sfixed_a(-0.00019850001262966543)),(to_sfixed_a(-0.004546706099063158)),(to_sfixed_a(0.0004233169602230191)),(to_sfixed_a(-9.414897067472339e-05)),(to_sfixed_a(-0.00014721014304086566)),(to_sfixed_a(0.00018950695812236518)),(to_sfixed_a(0.00018842695862986147)),(to_sfixed_a(0.36230796575546265)),(to_sfixed_a(0.004265889059752226)),(to_sfixed_a(-0.005971348844468594)),(to_sfixed_a(-3.607925827964209e-05)),(to_sfixed_a(-0.0003035459667444229)),(to_sfixed_a(-3.026789090654347e-05)),(to_sfixed_a(0.3816165626049042)),(to_sfixed_a(-0.00021515584376174957)),(to_sfixed_a(0.0012046050978824496)),(to_sfixed_a(8.981299470178783e-05)),(to_sfixed_a(0.0005731640849262476)),(to_sfixed_a(0.008216185495257378)),(to_sfixed_a(0.043772224336862564)),(to_sfixed_a(-0.10518106073141098)),(to_sfixed_a(-5.44906833965797e-05)),(to_sfixed_a(0.007459825836122036)),(to_sfixed_a(-9.289942681789398e-05)),(to_sfixed_a(-2.4523782485630363e-05)),(to_sfixed_a(0.0020473182667046785)),(to_sfixed_a(0.0001683364826021716)),(to_sfixed_a(0.00199690368026495)),(to_sfixed_a(0.015458385460078716)),(to_sfixed_a(0.003614442888647318)),(to_sfixed_a(-7.285951869562268e-05)),(to_sfixed_a(9.824780136113986e-05)),(to_sfixed_a(0.0008138178964145482)),(to_sfixed_a(-2.6579538825899363e-05)),(to_sfixed_a(-0.25695890188217163)),(to_sfixed_a(0.00015543968765996397)),(to_sfixed_a(-4.309389987611212e-05)),(to_sfixed_a(-1.3512973964679986e-05)),(to_sfixed_a(0.00785174872726202)),(to_sfixed_a(0.00022942973009776324)),(to_sfixed_a(-1.298740244237706e-06)),(to_sfixed_a(-0.0003099634777754545)),(to_sfixed_a(0.5798467993736267)),(to_sfixed_a(0.006885869428515434)),(to_sfixed_a(-8.583505405113101e-05)),(to_sfixed_a(-1.3551936717703938e-05)),(to_sfixed_a(-6.577203748747706e-06)),(to_sfixed_a(-0.00010638288222253323)),(to_sfixed_a(0.007849717512726784)),(to_sfixed_a(-0.09460996836423874)),(to_sfixed_a(-0.0008969818591140211)),(to_sfixed_a(-7.091453881002963e-05)),(to_sfixed_a(0.3769439458847046)),(to_sfixed_a(1.1622756574070081e-05)),(to_sfixed_a(-3.192196163581684e-05)),(to_sfixed_a(-1.5947480278555304e-06)),(to_sfixed_a(-0.0008583071175962687)),(to_sfixed_a(-7.134603220038116e-05)),(to_sfixed_a(1.6958554624579847e-05)),(to_sfixed_a(0.007499853614717722)),(to_sfixed_a(0.0012674779864028096)),(to_sfixed_a(-5.4303163778968155e-06)),(to_sfixed_a(-0.02840440534055233)),(to_sfixed_a(-0.28307288885116577)),(to_sfixed_a(0.0028728204779326916)),(to_sfixed_a(0.006113190203905106)),(to_sfixed_a(-2.5583489332348108e-05)),(to_sfixed_a(0.1526748389005661)),(to_sfixed_a(0.0004959668149240315)),(to_sfixed_a(-0.0010756211122497916)),(to_sfixed_a(0.000149837345816195)),(to_sfixed_a(-0.005629445426166058)),(to_sfixed_a(-0.24706296622753143)),(to_sfixed_a(0.010300897993147373)));

    constant weight_n2_48 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.2917625904083252)),(to_sfixed_a(0.005466729402542114)),(to_sfixed_a(-0.0004054427263326943)),(to_sfixed_a(-0.00018971627287101)),(to_sfixed_a(-0.003861928591504693)),(to_sfixed_a(-0.00025065065710805357)),(to_sfixed_a(-0.01578875444829464)),(to_sfixed_a(-0.000286173599306494)),(to_sfixed_a(0.00021859639673493803)),(to_sfixed_a(1.9644692656584084e-05)),(to_sfixed_a(6.285553536145017e-05)),(to_sfixed_a(-0.3325853943824768)),(to_sfixed_a(-0.00018912123050540686)),(to_sfixed_a(-0.0006892221863381565)),(to_sfixed_a(-0.00029181837453506887)),(to_sfixed_a(9.95149093796499e-07)),(to_sfixed_a(0.00918243732303381)),(to_sfixed_a(6.929512892384082e-05)),(to_sfixed_a(0.0018661089707165956)),(to_sfixed_a(-0.0030642214696854353)),(to_sfixed_a(-6.102029510657303e-05)),(to_sfixed_a(-0.00021761965763289481)),(to_sfixed_a(-0.0022618176881223917)),(to_sfixed_a(-0.008857998996973038)),(to_sfixed_a(-0.0012869903584942222)),(to_sfixed_a(0.34700319170951843)),(to_sfixed_a(-0.00011563527368707582)),(to_sfixed_a(-0.005978688597679138)),(to_sfixed_a(-0.0021840219851583242)),(to_sfixed_a(6.366566231008619e-05)),(to_sfixed_a(0.10743030160665512)),(to_sfixed_a(-0.00010284699965268373)),(to_sfixed_a(-0.008735685609281063)),(to_sfixed_a(-0.00021183434000704437)),(to_sfixed_a(-0.00015717610949650407)),(to_sfixed_a(0.00027464033337309957)),(to_sfixed_a(0.018903015181422234)),(to_sfixed_a(-0.27286961674690247)),(to_sfixed_a(-0.0013274123193696141)),(to_sfixed_a(0.0003068673540838063)),(to_sfixed_a(-0.004686417523771524)),(to_sfixed_a(-0.002556051593273878)),(to_sfixed_a(0.00011315180745441467)),(to_sfixed_a(-0.00010434723662910983)),(to_sfixed_a(-0.002284580608829856)),(to_sfixed_a(0.4708244800567627)),(to_sfixed_a(0.0004702235455624759)),(to_sfixed_a(-0.011393816210329533)),(to_sfixed_a(-1.8305152480024844e-05)),(to_sfixed_a(-0.0015460319118574262)),(to_sfixed_a(0.00915388111025095)),(to_sfixed_a(0.005952494218945503)),(to_sfixed_a(5.7906559959519655e-05)),(to_sfixed_a(0.4245757460594177)),(to_sfixed_a(-0.008181551471352577)),(to_sfixed_a(-0.0007613579509779811)),(to_sfixed_a(5.117301770951599e-05)),(to_sfixed_a(-0.0007204572902992368)),(to_sfixed_a(-1.0364830814069137e-05)),(to_sfixed_a(-4.139351949561387e-05)),(to_sfixed_a(-2.9266506317071617e-05)),(to_sfixed_a(-0.003780063008889556)),(to_sfixed_a(-0.0014055707724764943)),(to_sfixed_a(-0.3004007041454315)),(to_sfixed_a(3.2329277019016445e-05)),(to_sfixed_a(0.6573424339294434)),(to_sfixed_a(6.502278847619891e-05)),(to_sfixed_a(-0.005203616339713335)),(to_sfixed_a(-0.00013803978799842298)),(to_sfixed_a(-6.803097494412214e-05)),(to_sfixed_a(0.2555074989795685)),(to_sfixed_a(0.0014212342211976647)),(to_sfixed_a(0.3114866316318512)),(to_sfixed_a(-4.684960003942251e-05)),(to_sfixed_a(-0.0001836252340581268)),(to_sfixed_a(-0.0001813927519833669)),(to_sfixed_a(-0.11268265545368195)),(to_sfixed_a(-0.0009430261561647058)),(to_sfixed_a(0.00011648600047919899)),(to_sfixed_a(-0.15531539916992188)),(to_sfixed_a(-0.00947259645909071)),(to_sfixed_a(-0.00011646667553577572)),(to_sfixed_a(0.000278201827313751)),(to_sfixed_a(0.0005112112266942859)),(to_sfixed_a(4.7319983423221856e-05)),(to_sfixed_a(0.005206046160310507)),(to_sfixed_a(-0.0002471369516570121)),(to_sfixed_a(-0.007516481447964907)),(to_sfixed_a(2.300393498444464e-05)),(to_sfixed_a(-0.00013689178740605712)),(to_sfixed_a(0.009325660765171051)),(to_sfixed_a(2.9450427973642945e-05)),(to_sfixed_a(0.38395261764526367)),(to_sfixed_a(-9.344980935566127e-05)),(to_sfixed_a(0.2725081741809845)),(to_sfixed_a(1.7717240552883595e-05)),(to_sfixed_a(0.0001508706045569852)),(to_sfixed_a(-3.72602189600002e-05)),(to_sfixed_a(-6.704388943035156e-05)),(to_sfixed_a(-0.0001354265696136281)),(to_sfixed_a(-0.012143361382186413)),(to_sfixed_a(-0.006730911787599325)),(to_sfixed_a(-0.00017875873891171068)),(to_sfixed_a(-0.008664869703352451)),(to_sfixed_a(0.2342786341905594)),(to_sfixed_a(-0.28146275877952576)),(to_sfixed_a(5.80874111619778e-05)),(to_sfixed_a(-9.340047836303711e-05)),(to_sfixed_a(-7.102829840732738e-05)),(to_sfixed_a(0.22315117716789246)),(to_sfixed_a(0.005215649493038654)),(to_sfixed_a(-0.0001206587694468908)),(to_sfixed_a(0.0016068682307377458)),(to_sfixed_a(-5.2463365136645734e-06)),(to_sfixed_a(1.8898965208791196e-05)),(to_sfixed_a(-0.009858550503849983)),(to_sfixed_a(-0.003934195730835199)),(to_sfixed_a(-0.0063340687192976475)),(to_sfixed_a(6.99699594406411e-05)),(to_sfixed_a(-0.0012717057252302766)),(to_sfixed_a(-6.503249460365623e-05)),(to_sfixed_a(-3.752380143851042e-05)),(to_sfixed_a(0.006771944463253021)),(to_sfixed_a(-5.389541911426932e-06)),(to_sfixed_a(4.424145299708471e-05)),(to_sfixed_a(0.012581096962094307)),(to_sfixed_a(0.008095627650618553)),(to_sfixed_a(2.8175831175758503e-05)),(to_sfixed_a(7.180790271377191e-05)),(to_sfixed_a(-0.00014740352344233543)),(to_sfixed_a(-0.0001495081523898989)),(to_sfixed_a(8.819538925308734e-05)),(to_sfixed_a(0.008928314782679081)),(to_sfixed_a(0.010748526081442833)),(to_sfixed_a(-1.62333162734285e-05)),(to_sfixed_a(0.0001509790017735213)),(to_sfixed_a(-0.6347106099128723)),(to_sfixed_a(0.00011698292655637488)),(to_sfixed_a(0.00010338866559322923)),(to_sfixed_a(-8.916727529140189e-05)),(to_sfixed_a(-0.0013007944216951728)),(to_sfixed_a(7.430691766785458e-05)),(to_sfixed_a(0.00013056042371317744)),(to_sfixed_a(-0.00013088577543385327)),(to_sfixed_a(0.005822279024869204)),(to_sfixed_a(-0.005695822648704052)),(to_sfixed_a(0.20628611743450165)),(to_sfixed_a(-0.00012912072998005897)),(to_sfixed_a(-2.5061501219170168e-05)),(to_sfixed_a(0.007425927557051182)),(to_sfixed_a(-4.392773553263396e-05)),(to_sfixed_a(6.507732905447483e-05)),(to_sfixed_a(-0.0018885063473135233)),(to_sfixed_a(0.00011582802835619077)),(to_sfixed_a(-7.141538662835956e-05)),(to_sfixed_a(-0.003557149786502123)),(to_sfixed_a(-0.0002658710000105202)),(to_sfixed_a(-0.007740972563624382)),(to_sfixed_a(0.024074682965874672)),(to_sfixed_a(8.046181028475985e-05)),(to_sfixed_a(6.07777874392923e-05)),(to_sfixed_a(9.044379112310708e-07)),(to_sfixed_a(0.03245604410767555)),(to_sfixed_a(0.3471267521381378)),(to_sfixed_a(0.26615381240844727)),(to_sfixed_a(-0.00604428444057703)),(to_sfixed_a(-0.00011814242316177115)),(to_sfixed_a(0.001696388004347682)),(to_sfixed_a(-0.0001292493980145082)),(to_sfixed_a(-0.00041332817636430264)),(to_sfixed_a(0.0004226278397254646)),(to_sfixed_a(0.006094690877944231)),(to_sfixed_a(-0.0025080100167542696)),(to_sfixed_a(0.00023747244267724454)),(to_sfixed_a(-0.5084218382835388)),(to_sfixed_a(0.00012756508658640087)),(to_sfixed_a(-0.010438453406095505)),(to_sfixed_a(-0.396009624004364)),(to_sfixed_a(0.29676496982574463)),(to_sfixed_a(0.0016333541134372354)),(to_sfixed_a(-0.0009604952065274119)),(to_sfixed_a(0.14857900142669678)),(to_sfixed_a(3.979577741120011e-06)),(to_sfixed_a(7.764116890029982e-05)),(to_sfixed_a(0.00011757787433452904)),(to_sfixed_a(0.42916926741600037)),(to_sfixed_a(0.012270299717783928)),(to_sfixed_a(0.350874125957489)),(to_sfixed_a(-7.532222662121058e-05)),(to_sfixed_a(0.007425223011523485)),(to_sfixed_a(-0.004902484826743603)),(to_sfixed_a(-4.157845978625119e-06)),(to_sfixed_a(-0.021320199593901634)),(to_sfixed_a(-0.01842365600168705)),(to_sfixed_a(5.584792234003544e-06)),(to_sfixed_a(0.41916748881340027)),(to_sfixed_a(-0.0001961169036803767)),(to_sfixed_a(0.0033255673479288816)),(to_sfixed_a(-0.008190292865037918)),(to_sfixed_a(-1.1732576240319759e-05)),(to_sfixed_a(-6.155224400572479e-05)),(to_sfixed_a(-0.00024448716430924833)),(to_sfixed_a(1.620875991648063e-06)),(to_sfixed_a(7.411121623590589e-05)),(to_sfixed_a(-0.0001128765579778701)),(to_sfixed_a(0.00035181306884624064)),(to_sfixed_a(-0.357642263174057)),(to_sfixed_a(0.02952299267053604)),(to_sfixed_a(-0.0014696733560413122)),(to_sfixed_a(-0.006918084807693958)),(to_sfixed_a(-0.0036380901001393795)),(to_sfixed_a(-5.7188102800864726e-05)),(to_sfixed_a(-2.473439963068813e-06)),(to_sfixed_a(2.3568856704514474e-05)),(to_sfixed_a(0.0001673468796070665)),(to_sfixed_a(-2.3377404431812465e-05)),(to_sfixed_a(0.009613551199436188)),(to_sfixed_a(0.0010866003576666117)),(to_sfixed_a(0.020122183486819267)),(to_sfixed_a(-0.00015222375805024058)),(to_sfixed_a(5.680557660525665e-05)),(to_sfixed_a(6.662858504569158e-05)),(to_sfixed_a(0.00015671004075556993)),(to_sfixed_a(0.3490750193595886)),(to_sfixed_a(0.4221835434436798)),(to_sfixed_a(-5.939260154264048e-05)),(to_sfixed_a(-0.0001562244287924841)),(to_sfixed_a(-7.509138958994299e-05)),(to_sfixed_a(-0.2720918357372284)),(to_sfixed_a(0.45267584919929504)),(to_sfixed_a(-0.0023130199406296015)),(to_sfixed_a(-0.0002896895457524806)),(to_sfixed_a(-3.075620043091476e-06)),(to_sfixed_a(-2.682596823433414e-05)),(to_sfixed_a(-0.008320844732224941)),(to_sfixed_a(0.007788887247443199)),(to_sfixed_a(-0.2675243020057678)),(to_sfixed_a(1.2236141628818586e-05)),(to_sfixed_a(0.003428908297792077)),(to_sfixed_a(-1.0100702638737857e-05)),(to_sfixed_a(0.00879389327019453)),(to_sfixed_a(-0.00017272811965085566)),(to_sfixed_a(-0.01062153372913599)),(to_sfixed_a(-8.717917080502957e-05)),(to_sfixed_a(-0.25055381655693054)),(to_sfixed_a(-0.00011220070155104622)),(to_sfixed_a(-0.01053667813539505)),(to_sfixed_a(0.00037792796501889825)),(to_sfixed_a(-0.00011261398321948946)),(to_sfixed_a(-0.40814444422721863)),(to_sfixed_a(-0.02465907298028469)),(to_sfixed_a(-3.704719347297214e-05)),(to_sfixed_a(-0.003081232775002718)),(to_sfixed_a(0.0003813485673163086)),(to_sfixed_a(-0.0001384462957503274)),(to_sfixed_a(0.0027668506372720003)),(to_sfixed_a(-0.21520468592643738)),(to_sfixed_a(0.00024334009503945708)),(to_sfixed_a(0.000168197468155995)),(to_sfixed_a(-0.00024546391796320677)),(to_sfixed_a(-0.00019863445777446032)),(to_sfixed_a(-0.00914948433637619)),(to_sfixed_a(-0.0002507773460820317)),(to_sfixed_a(-0.0004580671084113419)),(to_sfixed_a(-8.2532518717926e-05)),(to_sfixed_a(-0.011633610352873802)),(to_sfixed_a(0.0001475989120081067)),(to_sfixed_a(6.966076762182638e-05)),(to_sfixed_a(-0.00011517482926137745)),(to_sfixed_a(-0.007179551292210817)),(to_sfixed_a(-0.000399937795009464)),(to_sfixed_a(-2.025616413448006e-05)),(to_sfixed_a(0.0002905755245592445)),(to_sfixed_a(-0.00037855395930819213)),(to_sfixed_a(-6.800697883591056e-05)),(to_sfixed_a(0.001272597350180149)),(to_sfixed_a(-0.00314242672175169)),(to_sfixed_a(-0.5136958360671997)),(to_sfixed_a(0.31216099858283997)),(to_sfixed_a(0.0023534605279564857)),(to_sfixed_a(3.233598545193672e-05)),(to_sfixed_a(0.00029019612702541053)),(to_sfixed_a(-3.1469346140511334e-05)),(to_sfixed_a(-0.0013872203417122364)),(to_sfixed_a(-1.1403233656892553e-05)),(to_sfixed_a(0.00019791786326095462)),(to_sfixed_a(-0.005460056476294994)),(to_sfixed_a(0.012117237783968449)),(to_sfixed_a(6.797692913096398e-05)),(to_sfixed_a(-0.0007580571109429002)),(to_sfixed_a(-6.90455999574624e-05)),(to_sfixed_a(-0.0036173085682094097)),(to_sfixed_a(0.2096443623304367)),(to_sfixed_a(-7.65363365644589e-05)),(to_sfixed_a(0.0005861303652636707)),(to_sfixed_a(-0.21361476182937622)),(to_sfixed_a(-0.02234021946787834)),(to_sfixed_a(-6.945891072973609e-05)),(to_sfixed_a(-0.006762202829122543)),(to_sfixed_a(0.0015477604465559125)),(to_sfixed_a(-0.04515620321035385)));

    constant weight_n2_49 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.3593768775463104)),(to_sfixed_a(-0.0003307229490019381)),(to_sfixed_a(0.0011205546325072646)),(to_sfixed_a(3.2269308576360345e-06)),(to_sfixed_a(-0.3945358395576477)),(to_sfixed_a(6.363194552250206e-05)),(to_sfixed_a(0.00788792409002781)),(to_sfixed_a(5.957794201094657e-05)),(to_sfixed_a(-0.0002905106812249869)),(to_sfixed_a(-0.00016611705359537154)),(to_sfixed_a(-7.488924893550575e-05)),(to_sfixed_a(0.20332983136177063)),(to_sfixed_a(-0.0012242287630215287)),(to_sfixed_a(-0.0003289768937975168)),(to_sfixed_a(0.0001873207656899467)),(to_sfixed_a(0.0001675575040280819)),(to_sfixed_a(0.011706882156431675)),(to_sfixed_a(7.124892727006227e-05)),(to_sfixed_a(0.0012818868272006512)),(to_sfixed_a(-0.0024818407837301493)),(to_sfixed_a(-0.00015313908807002008)),(to_sfixed_a(-6.111527909524739e-05)),(to_sfixed_a(-0.0017547780880704522)),(to_sfixed_a(-0.0047223218716681)),(to_sfixed_a(-0.00010371285316068679)),(to_sfixed_a(0.0002225627686129883)),(to_sfixed_a(0.00016781926387920976)),(to_sfixed_a(0.0021231607533991337)),(to_sfixed_a(0.0004825158102903515)),(to_sfixed_a(-0.0001481351355323568)),(to_sfixed_a(0.003022381104528904)),(to_sfixed_a(-6.724359991494566e-05)),(to_sfixed_a(0.2119767814874649)),(to_sfixed_a(0.00023958869860507548)),(to_sfixed_a(4.288878699298948e-06)),(to_sfixed_a(8.481889381073415e-05)),(to_sfixed_a(-0.009878936223685741)),(to_sfixed_a(-0.08488615602254868)),(to_sfixed_a(0.002802174771204591)),(to_sfixed_a(-0.00018219355843029916)),(to_sfixed_a(0.003156391903758049)),(to_sfixed_a(-0.002616654383018613)),(to_sfixed_a(-0.0003046539204660803)),(to_sfixed_a(-0.0002216929424321279)),(to_sfixed_a(-0.16383235156536102)),(to_sfixed_a(0.014076541177928448)),(to_sfixed_a(0.0009325130376964808)),(to_sfixed_a(-0.11737975478172302)),(to_sfixed_a(0.00026130370679311454)),(to_sfixed_a(0.620796799659729)),(to_sfixed_a(-0.26731061935424805)),(to_sfixed_a(3.2572213967796415e-05)),(to_sfixed_a(7.197493687272072e-06)),(to_sfixed_a(-0.0011225119233131409)),(to_sfixed_a(-0.001092994469217956)),(to_sfixed_a(0.001946881297044456)),(to_sfixed_a(-0.0002201902971137315)),(to_sfixed_a(-0.0028002499602735043)),(to_sfixed_a(-0.000247381191002205)),(to_sfixed_a(0.00011533600627444685)),(to_sfixed_a(-0.00029323421767912805)),(to_sfixed_a(0.0002753061708062887)),(to_sfixed_a(-0.00013891459093429148)),(to_sfixed_a(0.010424613952636719)),(to_sfixed_a(0.00020335306180641055)),(to_sfixed_a(0.0017991196364164352)),(to_sfixed_a(3.946862125303596e-05)),(to_sfixed_a(-0.003228883957490325)),(to_sfixed_a(5.348475679056719e-05)),(to_sfixed_a(0.00010132571333087981)),(to_sfixed_a(-0.560573399066925)),(to_sfixed_a(0.04799720644950867)),(to_sfixed_a(-0.023135432973504066)),(to_sfixed_a(-6.541056791320443e-06)),(to_sfixed_a(-0.00017675358685664833)),(to_sfixed_a(-3.6232599086361006e-05)),(to_sfixed_a(-0.011866092681884766)),(to_sfixed_a(0.00015444849850609899)),(to_sfixed_a(1.2501717719715089e-05)),(to_sfixed_a(0.010818922892212868)),(to_sfixed_a(0.00011624019680311903)),(to_sfixed_a(-4.797431756742299e-06)),(to_sfixed_a(-0.011208727955818176)),(to_sfixed_a(0.007212251424789429)),(to_sfixed_a(0.00010223157005384564)),(to_sfixed_a(0.010713541880249977)),(to_sfixed_a(0.005773797631263733)),(to_sfixed_a(0.0035286799538880587)),(to_sfixed_a(-0.00011931764311157167)),(to_sfixed_a(6.225014658411965e-06)),(to_sfixed_a(0.0024011130444705486)),(to_sfixed_a(-3.953982377424836e-05)),(to_sfixed_a(0.004862206522375345)),(to_sfixed_a(1.0483243386261165e-05)),(to_sfixed_a(-0.00046853694948367774)),(to_sfixed_a(-6.508996739285067e-05)),(to_sfixed_a(0.0002050591865554452)),(to_sfixed_a(-7.026360981399193e-05)),(to_sfixed_a(1.138192237704061e-05)),(to_sfixed_a(-0.00015511178935412318)),(to_sfixed_a(-0.007831936702132225)),(to_sfixed_a(0.18223103880882263)),(to_sfixed_a(1.1744399671442807e-05)),(to_sfixed_a(-0.001414939877577126)),(to_sfixed_a(-0.017401179298758507)),(to_sfixed_a(-0.0004392522678244859)),(to_sfixed_a(0.00020183660672046244)),(to_sfixed_a(-8.910406904760748e-06)),(to_sfixed_a(-6.65349725750275e-05)),(to_sfixed_a(0.007917637005448341)),(to_sfixed_a(-0.01090956013649702)),(to_sfixed_a(-0.00016972066077869385)),(to_sfixed_a(0.031898003071546555)),(to_sfixed_a(1.7900412785820663e-05)),(to_sfixed_a(-4.322861786931753e-05)),(to_sfixed_a(-0.006386475171893835)),(to_sfixed_a(-0.005905963946133852)),(to_sfixed_a(0.00042682496132329106)),(to_sfixed_a(0.00017422337259631604)),(to_sfixed_a(-0.0006063145701773465)),(to_sfixed_a(-3.098975867033005e-07)),(to_sfixed_a(-9.776288061402738e-05)),(to_sfixed_a(-0.00288305152207613)),(to_sfixed_a(-6.896490231156349e-05)),(to_sfixed_a(-6.935887358849868e-05)),(to_sfixed_a(0.004527149256318808)),(to_sfixed_a(-0.47952800989151)),(to_sfixed_a(-8.79799627000466e-05)),(to_sfixed_a(0.00010468987602507696)),(to_sfixed_a(2.6267560315318406e-05)),(to_sfixed_a(0.00013055888121016324)),(to_sfixed_a(-0.0002371791924815625)),(to_sfixed_a(-0.002807374345138669)),(to_sfixed_a(-0.6331267356872559)),(to_sfixed_a(0.00016758800484240055)),(to_sfixed_a(0.00015256712504196912)),(to_sfixed_a(0.1995665282011032)),(to_sfixed_a(0.3745264410972595)),(to_sfixed_a(-2.840522938640788e-06)),(to_sfixed_a(-0.00010779986041598022)),(to_sfixed_a(0.005598567426204681)),(to_sfixed_a(0.0004195937071926892)),(to_sfixed_a(-0.00016606519056949764)),(to_sfixed_a(-8.996528049465269e-05)),(to_sfixed_a(0.0010649486212059855)),(to_sfixed_a(-0.0005352518055588007)),(to_sfixed_a(-0.000280361418845132)),(to_sfixed_a(0.00015061438898555934)),(to_sfixed_a(-5.9773705288534984e-05)),(to_sfixed_a(0.0013231333578005433)),(to_sfixed_a(8.436352800345048e-05)),(to_sfixed_a(8.518734102835879e-05)),(to_sfixed_a(-0.0068996865302324295)),(to_sfixed_a(8.555004023946822e-05)),(to_sfixed_a(-5.4422736866399646e-05)),(to_sfixed_a(0.003483860520645976)),(to_sfixed_a(0.00028874812414869666)),(to_sfixed_a(0.001515860902145505)),(to_sfixed_a(-9.967312507797033e-06)),(to_sfixed_a(7.250954513438046e-05)),(to_sfixed_a(0.00011599664867389947)),(to_sfixed_a(-7.804419146850705e-05)),(to_sfixed_a(-0.0025865540374070406)),(to_sfixed_a(0.005939437076449394)),(to_sfixed_a(-0.001243817969225347)),(to_sfixed_a(0.0031493394635617733)),(to_sfixed_a(0.00017189323261845857)),(to_sfixed_a(-0.3580264747142792)),(to_sfixed_a(2.361282895435579e-05)),(to_sfixed_a(-6.390372436726466e-05)),(to_sfixed_a(-0.35815683007240295)),(to_sfixed_a(0.001393222832120955)),(to_sfixed_a(0.006114307325333357)),(to_sfixed_a(-0.00017548564937897027)),(to_sfixed_a(0.2620520293712616)),(to_sfixed_a(-0.00016260994016192853)),(to_sfixed_a(0.19877572357654572)),(to_sfixed_a(0.00936782918870449)),(to_sfixed_a(-0.00017429063154850155)),(to_sfixed_a(-9.129435056820512e-06)),(to_sfixed_a(0.0010032592108473182)),(to_sfixed_a(-0.034209415316581726)),(to_sfixed_a(0.00013060911442153156)),(to_sfixed_a(-0.00017362157814204693)),(to_sfixed_a(0.0002446273574605584)),(to_sfixed_a(-0.0011810272699221969)),(to_sfixed_a(0.007133656181395054)),(to_sfixed_a(-0.0017969587352126837)),(to_sfixed_a(-0.0008342500077560544)),(to_sfixed_a(-0.5621764659881592)),(to_sfixed_a(-0.012718097306787968)),(to_sfixed_a(-0.00023022250388748944)),(to_sfixed_a(-0.008753887377679348)),(to_sfixed_a(0.0008211826789192855)),(to_sfixed_a(3.890343941748142e-05)),(to_sfixed_a(-0.010622699744999409)),(to_sfixed_a(0.00025099588674493134)),(to_sfixed_a(0.0014375537866726518)),(to_sfixed_a(0.3439231216907501)),(to_sfixed_a(-1.9851191609632224e-05)),(to_sfixed_a(-0.00011588264897000045)),(to_sfixed_a(0.0001658725377637893)),(to_sfixed_a(5.2710453019244596e-05)),(to_sfixed_a(7.066191028570756e-05)),(to_sfixed_a(-0.00012046004121657461)),(to_sfixed_a(0.0025139476638287306)),(to_sfixed_a(0.0019811848178505898)),(to_sfixed_a(0.3982621133327484)),(to_sfixed_a(0.24780461192131042)),(to_sfixed_a(0.32807260751724243)),(to_sfixed_a(-0.0030058224219828844)),(to_sfixed_a(-6.96259958203882e-05)),(to_sfixed_a(-2.9372058634180576e-06)),(to_sfixed_a(-7.033743895590305e-05)),(to_sfixed_a(-0.0001762132451403886)),(to_sfixed_a(-5.764816523878835e-05)),(to_sfixed_a(0.0036959671415388584)),(to_sfixed_a(0.002304127672687173)),(to_sfixed_a(0.20667818188667297)),(to_sfixed_a(-1.7738071619533002e-05)),(to_sfixed_a(-2.0547304302453995e-08)),(to_sfixed_a(-0.00010934439342236146)),(to_sfixed_a(-0.00015753789921291173)),(to_sfixed_a(0.00033841864205896854)),(to_sfixed_a(-0.11644736677408218)),(to_sfixed_a(1.8224796804133803e-05)),(to_sfixed_a(8.846462151268497e-05)),(to_sfixed_a(0.00027111946837976575)),(to_sfixed_a(0.0030158197041600943)),(to_sfixed_a(0.6173414587974548)),(to_sfixed_a(5.231564864516258e-05)),(to_sfixed_a(-7.195083162514493e-05)),(to_sfixed_a(0.00018514733528718352)),(to_sfixed_a(-1.1708267265930772e-05)),(to_sfixed_a(0.0061479355208575726)),(to_sfixed_a(-0.014893247745931149)),(to_sfixed_a(-0.27437615394592285)),(to_sfixed_a(4.960273508913815e-05)),(to_sfixed_a(0.000152075313962996)),(to_sfixed_a(-3.1299889087677e-05)),(to_sfixed_a(-0.28580597043037415)),(to_sfixed_a(-0.0002358811761951074)),(to_sfixed_a(0.0026010354049503803)),(to_sfixed_a(-8.546262688469142e-05)),(to_sfixed_a(-0.022299638018012047)),(to_sfixed_a(0.00537441112101078)),(to_sfixed_a(-0.0011386158876121044)),(to_sfixed_a(0.14763875305652618)),(to_sfixed_a(-0.0002850776072591543)),(to_sfixed_a(-0.21196751296520233)),(to_sfixed_a(0.0030432117637246847)),(to_sfixed_a(2.591172233223915e-05)),(to_sfixed_a(-0.0002930560440290719)),(to_sfixed_a(-0.0004447694809641689)),(to_sfixed_a(0.00030051852809265256)),(to_sfixed_a(0.48872050642967224)),(to_sfixed_a(0.2207014560699463)),(to_sfixed_a(0.00017536390805616975)),(to_sfixed_a(8.145820174831897e-05)),(to_sfixed_a(0.005223672837018967)),(to_sfixed_a(0.00013631265028379858)),(to_sfixed_a(0.0024318282958120108)),(to_sfixed_a(8.400483056902885e-05)),(to_sfixed_a(0.15881642699241638)),(to_sfixed_a(0.00013726107135880738)),(to_sfixed_a(0.00088644860079512)),(to_sfixed_a(4.335166158853099e-05)),(to_sfixed_a(-0.00018133049889001995)),(to_sfixed_a(0.00029532189364545047)),(to_sfixed_a(0.00894014723598957)),(to_sfixed_a(-0.2730468213558197)),(to_sfixed_a(8.988272747956216e-05)),(to_sfixed_a(0.00045971610234119)),(to_sfixed_a(2.719584881560877e-05)),(to_sfixed_a(5.9951107687084004e-05)),(to_sfixed_a(-0.0007279567653313279)),(to_sfixed_a(-0.002537144348025322)),(to_sfixed_a(-0.10944539308547974)),(to_sfixed_a(0.0371658056974411)),(to_sfixed_a(-0.0005133203230798244)),(to_sfixed_a(2.9685135814361274e-05)),(to_sfixed_a(-0.00020093933562748134)),(to_sfixed_a(2.0368835976114497e-05)),(to_sfixed_a(-0.0026565950829535723)),(to_sfixed_a(0.00029009004356339574)),(to_sfixed_a(9.923032484948635e-05)),(to_sfixed_a(0.00013755258987657726)),(to_sfixed_a(0.011737868189811707)),(to_sfixed_a(5.596955452347174e-05)),(to_sfixed_a(0.0002574846148490906)),(to_sfixed_a(-0.0051984284073114395)),(to_sfixed_a(0.0009568747482262552)),(to_sfixed_a(0.000541732064448297)),(to_sfixed_a(-7.83923824201338e-05)),(to_sfixed_a(0.2671334147453308)),(to_sfixed_a(4.161658580414951e-05)),(to_sfixed_a(0.003877856070175767)),(to_sfixed_a(-6.814872904215008e-05)),(to_sfixed_a(0.007052927743643522)),(to_sfixed_a(-0.02253410592675209)),(to_sfixed_a(0.012071073055267334)));

    constant weight_n2_50 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.03956938162446022)),(to_sfixed_a(-0.3169018030166626)),(to_sfixed_a(0.0009670755243860185)),(to_sfixed_a(-1.1858937796205282e-06)),(to_sfixed_a(0.017157215625047684)),(to_sfixed_a(0.00016822401084937155)),(to_sfixed_a(-0.02696909010410309)),(to_sfixed_a(-0.00017601906438358128)),(to_sfixed_a(8.49471689434722e-06)),(to_sfixed_a(-3.9448364987038076e-05)),(to_sfixed_a(7.232587813632563e-05)),(to_sfixed_a(0.01558738760650158)),(to_sfixed_a(-0.4903384745121002)),(to_sfixed_a(-0.0005730256671085954)),(to_sfixed_a(-9.879860590444878e-05)),(to_sfixed_a(-9.79842952801846e-05)),(to_sfixed_a(-0.0006949490052647889)),(to_sfixed_a(2.7642614440992475e-05)),(to_sfixed_a(-0.0073413727805018425)),(to_sfixed_a(-6.170067354105413e-05)),(to_sfixed_a(7.012393325567245e-05)),(to_sfixed_a(-5.69170260860119e-05)),(to_sfixed_a(0.00016196267097257078)),(to_sfixed_a(-0.0006777073722332716)),(to_sfixed_a(-0.00027845677686855197)),(to_sfixed_a(0.0006781991687603295)),(to_sfixed_a(0.00015096877177711576)),(to_sfixed_a(0.000546952651347965)),(to_sfixed_a(0.0005578225827775896)),(to_sfixed_a(4.127483407501131e-05)),(to_sfixed_a(-0.018559256568551064)),(to_sfixed_a(0.000104436170659028)),(to_sfixed_a(-0.0076686604879796505)),(to_sfixed_a(-5.745777161791921e-05)),(to_sfixed_a(1.3439981557894498e-05)),(to_sfixed_a(-0.00017805208335630596)),(to_sfixed_a(-0.34059780836105347)),(to_sfixed_a(0.24901796877384186)),(to_sfixed_a(0.006613234989345074)),(to_sfixed_a(-8.372122829314321e-05)),(to_sfixed_a(0.005632653832435608)),(to_sfixed_a(-0.0011814675526693463)),(to_sfixed_a(-1.0322673915652558e-06)),(to_sfixed_a(0.00010921909415628761)),(to_sfixed_a(-0.007659007329493761)),(to_sfixed_a(0.001492301351390779)),(to_sfixed_a(0.014268985949456692)),(to_sfixed_a(0.27698495984077454)),(to_sfixed_a(-6.444052269216627e-05)),(to_sfixed_a(0.001654129708185792)),(to_sfixed_a(-0.007193754892796278)),(to_sfixed_a(-0.0004602480912581086)),(to_sfixed_a(-1.9276987586636096e-05)),(to_sfixed_a(0.0013445564545691013)),(to_sfixed_a(-0.0002401743840891868)),(to_sfixed_a(0.00024941691663116217)),(to_sfixed_a(4.890243872068822e-07)),(to_sfixed_a(0.00044770928798243403)),(to_sfixed_a(0.0003062014002352953)),(to_sfixed_a(0.0001283212477574125)),(to_sfixed_a(-0.0005560726276598871)),(to_sfixed_a(-0.0003248946741223335)),(to_sfixed_a(0.00047251713112927973)),(to_sfixed_a(0.007891261018812656)),(to_sfixed_a(-0.00018353565246798098)),(to_sfixed_a(0.24205338954925537)),(to_sfixed_a(0.00011450536112533882)),(to_sfixed_a(0.303460031747818)),(to_sfixed_a(0.0005560955032706261)),(to_sfixed_a(0.0002881870314013213)),(to_sfixed_a(0.004039946477860212)),(to_sfixed_a(0.0028660830575972795)),(to_sfixed_a(0.0011596751864999533)),(to_sfixed_a(-6.90806336933747e-05)),(to_sfixed_a(0.00012904408504255116)),(to_sfixed_a(6.702124665025622e-05)),(to_sfixed_a(0.0019374657422304153)),(to_sfixed_a(-0.002781572286039591)),(to_sfixed_a(-2.1089217625558376e-06)),(to_sfixed_a(0.004941707942634821)),(to_sfixed_a(-9.841927385423332e-05)),(to_sfixed_a(-7.453963917214423e-05)),(to_sfixed_a(3.745290086953901e-05)),(to_sfixed_a(-0.443541556596756)),(to_sfixed_a(-0.00010468844266142696)),(to_sfixed_a(0.0007236718665808439)),(to_sfixed_a(-0.0047147804871201515)),(to_sfixed_a(-0.00013903211220167577)),(to_sfixed_a(0.00044544320553541183)),(to_sfixed_a(-0.00013637676602229476)),(to_sfixed_a(-0.009336929768323898)),(to_sfixed_a(4.887866089120507e-05)),(to_sfixed_a(0.00172870559617877)),(to_sfixed_a(-5.784626409877092e-06)),(to_sfixed_a(-0.005032431334257126)),(to_sfixed_a(0.13745594024658203)),(to_sfixed_a(-2.3296644940273836e-05)),(to_sfixed_a(2.7954942197538912e-05)),(to_sfixed_a(5.782274092780426e-05)),(to_sfixed_a(7.622933480888605e-05)),(to_sfixed_a(0.00045649291132576764)),(to_sfixed_a(-0.001157180406153202)),(to_sfixed_a(6.7112036049366e-05)),(to_sfixed_a(0.0024389722384512424)),(to_sfixed_a(0.007533828262239695)),(to_sfixed_a(0.00020702109031844884)),(to_sfixed_a(9.494615369476378e-07)),(to_sfixed_a(-6.288916483754292e-05)),(to_sfixed_a(0.00011207351053599268)),(to_sfixed_a(-0.012063104659318924)),(to_sfixed_a(-0.011362625285983086)),(to_sfixed_a(4.750759762828238e-05)),(to_sfixed_a(0.5183699727058411)),(to_sfixed_a(-0.00017808220582082868)),(to_sfixed_a(-0.00012964487541466951)),(to_sfixed_a(0.2202746570110321)),(to_sfixed_a(-0.0037554209120571613)),(to_sfixed_a(-7.058797200443223e-05)),(to_sfixed_a(-1.5077675925567746e-06)),(to_sfixed_a(0.00377066433429718)),(to_sfixed_a(5.633548062178306e-05)),(to_sfixed_a(0.0001214565199916251)),(to_sfixed_a(0.003034561639651656)),(to_sfixed_a(0.0001570989697938785)),(to_sfixed_a(-1.3010285329073668e-06)),(to_sfixed_a(0.2328515201807022)),(to_sfixed_a(-7.325431215576828e-05)),(to_sfixed_a(3.678610300994478e-05)),(to_sfixed_a(-8.531540515832603e-06)),(to_sfixed_a(6.923197361174971e-06)),(to_sfixed_a(0.00013294332893565297)),(to_sfixed_a(0.00017608472262509167)),(to_sfixed_a(4.617281229002401e-05)),(to_sfixed_a(-0.0010921533685177565)),(to_sfixed_a(-6.729621964041144e-05)),(to_sfixed_a(3.85728053515777e-05)),(to_sfixed_a(0.3941664695739746)),(to_sfixed_a(0.0011991815408691764)),(to_sfixed_a(0.00013303854211699218)),(to_sfixed_a(-0.00023685090127401054)),(to_sfixed_a(0.00010791392560349777)),(to_sfixed_a(-2.5094414013437927e-06)),(to_sfixed_a(3.316371294204146e-05)),(to_sfixed_a(1.0192095942329615e-05)),(to_sfixed_a(6.705775740556419e-05)),(to_sfixed_a(8.111324132187292e-05)),(to_sfixed_a(-0.00015408196486532688)),(to_sfixed_a(-3.0748375138500705e-05)),(to_sfixed_a(0.00010087353439303115)),(to_sfixed_a(0.0036171283572912216)),(to_sfixed_a(0.00010458067117724568)),(to_sfixed_a(7.06552091287449e-05)),(to_sfixed_a(-0.0035022138617932796)),(to_sfixed_a(-2.884220884880051e-05)),(to_sfixed_a(-4.506385448621586e-05)),(to_sfixed_a(-0.006247424520552158)),(to_sfixed_a(-2.2106512915343046e-05)),(to_sfixed_a(0.0012667503906413913)),(to_sfixed_a(5.0989452574867755e-05)),(to_sfixed_a(0.00010170145105803385)),(to_sfixed_a(8.926718874135986e-05)),(to_sfixed_a(0.0001299685100093484)),(to_sfixed_a(0.018544990569353104)),(to_sfixed_a(-0.07110114395618439)),(to_sfixed_a(-0.00993785634636879)),(to_sfixed_a(0.00037000825977884233)),(to_sfixed_a(-3.0512819648720324e-06)),(to_sfixed_a(-4.85373820993118e-05)),(to_sfixed_a(-0.00018796601216308773)),(to_sfixed_a(0.00011912449554074556)),(to_sfixed_a(-0.2815185487270355)),(to_sfixed_a(-0.00012254470493644476)),(to_sfixed_a(-1.217870885739103e-05)),(to_sfixed_a(0.00016513466835021973)),(to_sfixed_a(0.2892891466617584)),(to_sfixed_a(-0.0018045901088044047)),(to_sfixed_a(8.738896576687694e-05)),(to_sfixed_a(0.0006167658139020205)),(to_sfixed_a(0.2743300497531891)),(to_sfixed_a(-0.006327885203063488)),(to_sfixed_a(-0.0005531150964088738)),(to_sfixed_a(7.782589818816632e-05)),(to_sfixed_a(-3.784096406889148e-05)),(to_sfixed_a(0.00031453956034965813)),(to_sfixed_a(7.029091648291796e-05)),(to_sfixed_a(0.0012016710825264454)),(to_sfixed_a(0.00015853233344387263)),(to_sfixed_a(0.140494242310524)),(to_sfixed_a(3.192386793671176e-05)),(to_sfixed_a(2.21865157072898e-05)),(to_sfixed_a(-0.0002986053004860878)),(to_sfixed_a(-7.011587877059355e-05)),(to_sfixed_a(0.34850969910621643)),(to_sfixed_a(0.00043941469630226493)),(to_sfixed_a(-6.069015944376588e-05)),(to_sfixed_a(0.00017691077664494514)),(to_sfixed_a(-5.7261982874479145e-05)),(to_sfixed_a(-0.23307642340660095)),(to_sfixed_a(0.00033148148213513196)),(to_sfixed_a(-0.0004257207619957626)),(to_sfixed_a(-1.4574761735275388e-06)),(to_sfixed_a(0.0003218160127289593)),(to_sfixed_a(-2.466818841639906e-05)),(to_sfixed_a(6.911774835316464e-05)),(to_sfixed_a(6.14572927588597e-05)),(to_sfixed_a(-3.0284882086561993e-05)),(to_sfixed_a(-0.001720492378808558)),(to_sfixed_a(-0.00012340441753622144)),(to_sfixed_a(-0.012357104569673538)),(to_sfixed_a(0.0036642036866396666)),(to_sfixed_a(-0.0001590368920005858)),(to_sfixed_a(0.00023975274234544486)),(to_sfixed_a(0.00021694388124160469)),(to_sfixed_a(-2.8579597710631788e-05)),(to_sfixed_a(-1.4075558283366263e-05)),(to_sfixed_a(-4.285546310711652e-05)),(to_sfixed_a(-9.195946040563285e-05)),(to_sfixed_a(-0.010731350630521774)),(to_sfixed_a(0.0004092301242053509)),(to_sfixed_a(-0.00011389862629584968)),(to_sfixed_a(-0.00011461460235295817)),(to_sfixed_a(3.305007703602314e-05)),(to_sfixed_a(-1.3869983376935124e-05)),(to_sfixed_a(0.2999308109283447)),(to_sfixed_a(0.015171270817518234)),(to_sfixed_a(0.00012879370478913188)),(to_sfixed_a(-0.00020741349726449698)),(to_sfixed_a(-0.00020657562708947808)),(to_sfixed_a(-0.22124387323856354)),(to_sfixed_a(0.3897576332092285)),(to_sfixed_a(0.009684247896075249)),(to_sfixed_a(0.00011710124817909673)),(to_sfixed_a(2.5985185857280158e-05)),(to_sfixed_a(-3.170855052303523e-05)),(to_sfixed_a(-6.270752055570483e-05)),(to_sfixed_a(-0.0016651698388159275)),(to_sfixed_a(-0.256909042596817)),(to_sfixed_a(9.831647184910253e-05)),(to_sfixed_a(-0.00025425569037906826)),(to_sfixed_a(-0.0002767648547887802)),(to_sfixed_a(0.0002495837979950011)),(to_sfixed_a(-7.006420491961762e-05)),(to_sfixed_a(0.6178481578826904)),(to_sfixed_a(-1.8127320799976587e-05)),(to_sfixed_a(0.6660754084587097)),(to_sfixed_a(-0.0032193136867135763)),(to_sfixed_a(0.014318200759589672)),(to_sfixed_a(0.39877450466156006)),(to_sfixed_a(-1.6684338334016502e-05)),(to_sfixed_a(-0.25209012627601624)),(to_sfixed_a(7.263419684022665e-05)),(to_sfixed_a(-4.8264751967508346e-05)),(to_sfixed_a(-0.0009188160765916109)),(to_sfixed_a(1.789240923244506e-05)),(to_sfixed_a(0.00018971841200254858)),(to_sfixed_a(0.4390968084335327)),(to_sfixed_a(-0.0022757842671126127)),(to_sfixed_a(-1.1471096513560042e-05)),(to_sfixed_a(-9.807899914449081e-05)),(to_sfixed_a(-0.005630387458950281)),(to_sfixed_a(0.00010738411219790578)),(to_sfixed_a(0.0038581225089728832)),(to_sfixed_a(0.00023622480512131006)),(to_sfixed_a(0.2134837657213211)),(to_sfixed_a(7.545113476226106e-07)),(to_sfixed_a(-0.21543563902378082)),(to_sfixed_a(-0.00011543372238520533)),(to_sfixed_a(0.00010123100219061598)),(to_sfixed_a(-1.675952080404386e-05)),(to_sfixed_a(-0.04580208286643028)),(to_sfixed_a(0.0011417068308219314)),(to_sfixed_a(-7.852759154047817e-06)),(to_sfixed_a(0.00014867547724861652)),(to_sfixed_a(1.6325051547028124e-05)),(to_sfixed_a(-0.00013660872355103493)),(to_sfixed_a(0.4446163773536682)),(to_sfixed_a(0.0015152876731008291)),(to_sfixed_a(-0.0007866054656915367)),(to_sfixed_a(-0.43080973625183105)),(to_sfixed_a(0.0005781150539405644)),(to_sfixed_a(1.1055526556447148e-06)),(to_sfixed_a(-2.145526377717033e-05)),(to_sfixed_a(0.00014431524323299527)),(to_sfixed_a(0.00027728304849006236)),(to_sfixed_a(0.0002522446447983384)),(to_sfixed_a(-0.00011298068420728669)),(to_sfixed_a(0.0006560417823493481)),(to_sfixed_a(-0.3287794888019562)),(to_sfixed_a(0.00024908300838433206)),(to_sfixed_a(3.725448914337903e-05)),(to_sfixed_a(0.08770139515399933)),(to_sfixed_a(-0.010152912698686123)),(to_sfixed_a(0.003276925068348646)),(to_sfixed_a(-5.368207348510623e-05)),(to_sfixed_a(0.32438409328460693)),(to_sfixed_a(0.0003915834822691977)),(to_sfixed_a(0.0028620033990591764)),(to_sfixed_a(-7.745284528937191e-05)),(to_sfixed_a(-0.16278930008411407)),(to_sfixed_a(-0.010694578289985657)),(to_sfixed_a(0.0008979430422186852)));

    constant weight_n2_51 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.12365690618753433)),(to_sfixed_a(0.0014196953270584345)),(to_sfixed_a(-0.0036611100658774376)),(to_sfixed_a(-0.00030373010667972267)),(to_sfixed_a(0.006576417479664087)),(to_sfixed_a(-0.00023614108795300126)),(to_sfixed_a(-0.0014337345492094755)),(to_sfixed_a(-0.0001351881946902722)),(to_sfixed_a(-7.149855082388967e-05)),(to_sfixed_a(-0.00011720808106474578)),(to_sfixed_a(-0.00010338064021198079)),(to_sfixed_a(-0.5418473482131958)),(to_sfixed_a(0.0007535696495324373)),(to_sfixed_a(0.0028408134821802378)),(to_sfixed_a(0.00016838729789014906)),(to_sfixed_a(-5.895684807910584e-05)),(to_sfixed_a(0.3220156133174896)),(to_sfixed_a(-5.763376975664869e-05)),(to_sfixed_a(0.10932395607233047)),(to_sfixed_a(-0.015825532376766205)),(to_sfixed_a(0.0003144911315757781)),(to_sfixed_a(-0.00017781363567337394)),(to_sfixed_a(0.0002502668066881597)),(to_sfixed_a(-0.0019081616774201393)),(to_sfixed_a(-0.0023131188936531544)),(to_sfixed_a(0.3369392454624176)),(to_sfixed_a(0.00015518823056481779)),(to_sfixed_a(0.00016884898650459945)),(to_sfixed_a(0.36980581283569336)),(to_sfixed_a(-0.00028577528428286314)),(to_sfixed_a(-0.0012603213544934988)),(to_sfixed_a(0.00012804348079953343)),(to_sfixed_a(-0.001956716412678361)),(to_sfixed_a(3.226042099413462e-05)),(to_sfixed_a(0.00014937040396034718)),(to_sfixed_a(8.272600098280236e-05)),(to_sfixed_a(0.2507425844669342)),(to_sfixed_a(0.3038082420825958)),(to_sfixed_a(0.0031237704679369926)),(to_sfixed_a(-0.00020085403230041265)),(to_sfixed_a(-0.01873810403048992)),(to_sfixed_a(-0.01130695827305317)),(to_sfixed_a(-0.0001390089455526322)),(to_sfixed_a(-0.000142752323881723)),(to_sfixed_a(0.004586134105920792)),(to_sfixed_a(0.501054584980011)),(to_sfixed_a(0.0014423185493797064)),(to_sfixed_a(0.00723700225353241)),(to_sfixed_a(0.00023743341444060206)),(to_sfixed_a(-0.0008163654711097479)),(to_sfixed_a(0.4554823637008667)),(to_sfixed_a(0.0005966637982055545)),(to_sfixed_a(-0.00021874501544516534)),(to_sfixed_a(0.17350947856903076)),(to_sfixed_a(-0.003795844269916415)),(to_sfixed_a(-0.002537996042519808)),(to_sfixed_a(-0.00017430572188459337)),(to_sfixed_a(-0.004813395440578461)),(to_sfixed_a(2.954562660306692e-06)),(to_sfixed_a(-0.00017596119141671807)),(to_sfixed_a(0.007603376638144255)),(to_sfixed_a(-0.0024283549282699823)),(to_sfixed_a(0.0007446561940014362)),(to_sfixed_a(0.00445684976875782)),(to_sfixed_a(-9.86483137239702e-05)),(to_sfixed_a(0.3606870770454407)),(to_sfixed_a(-2.720265183597803e-05)),(to_sfixed_a(-0.0001068197307176888)),(to_sfixed_a(0.002212794730439782)),(to_sfixed_a(-0.00011635409464361146)),(to_sfixed_a(0.0006955131539143622)),(to_sfixed_a(0.025421833619475365)),(to_sfixed_a(0.02634432166814804)),(to_sfixed_a(-1.490165595896542e-05)),(to_sfixed_a(-7.733462553005666e-06)),(to_sfixed_a(-2.948539622593671e-05)),(to_sfixed_a(-0.7436113953590393)),(to_sfixed_a(0.14032739400863647)),(to_sfixed_a(4.360746606835164e-05)),(to_sfixed_a(-0.3224174678325653)),(to_sfixed_a(0.0032312232069671154)),(to_sfixed_a(-0.0002904599532485008)),(to_sfixed_a(0.004597383085638285)),(to_sfixed_a(-0.0015447826590389013)),(to_sfixed_a(-4.660659396904521e-05)),(to_sfixed_a(0.0007775748963467777)),(to_sfixed_a(0.2492436021566391)),(to_sfixed_a(-0.02208407036960125)),(to_sfixed_a(1.8776345314108767e-05)),(to_sfixed_a(6.211204890860245e-05)),(to_sfixed_a(0.008686878718435764)),(to_sfixed_a(4.764171899296343e-05)),(to_sfixed_a(0.23625318706035614)),(to_sfixed_a(-0.00012990995310246944)),(to_sfixed_a(0.2278350293636322)),(to_sfixed_a(9.459417196922004e-05)),(to_sfixed_a(9.343608689960092e-05)),(to_sfixed_a(9.047203639056534e-05)),(to_sfixed_a(3.913824912160635e-05)),(to_sfixed_a(0.00011317459575366229)),(to_sfixed_a(-0.004874371457844973)),(to_sfixed_a(-0.4139312505722046)),(to_sfixed_a(-0.00011654257104964927)),(to_sfixed_a(-0.011489407159388065)),(to_sfixed_a(0.013618230819702148)),(to_sfixed_a(-0.003836230840533972)),(to_sfixed_a(-0.00014948856551200151)),(to_sfixed_a(-1.9065480955759995e-05)),(to_sfixed_a(6.621998909395188e-05)),(to_sfixed_a(-0.0001495789474574849)),(to_sfixed_a(-0.002121181692928076)),(to_sfixed_a(6.981891056057066e-05)),(to_sfixed_a(0.24153442680835724)),(to_sfixed_a(8.561473805457354e-06)),(to_sfixed_a(1.4958932297304273e-05)),(to_sfixed_a(0.016114115715026855)),(to_sfixed_a(-0.005724216345697641)),(to_sfixed_a(1.1910171451745555e-05)),(to_sfixed_a(-2.9925347917014733e-05)),(to_sfixed_a(0.37609633803367615)),(to_sfixed_a(-0.00019966856052633375)),(to_sfixed_a(-0.00019347584748174995)),(to_sfixed_a(0.004924421198666096)),(to_sfixed_a(-3.543793718563393e-05)),(to_sfixed_a(0.00014821754302829504)),(to_sfixed_a(0.17307105660438538)),(to_sfixed_a(-0.399300754070282)),(to_sfixed_a(6.133028364274651e-05)),(to_sfixed_a(-4.336009078542702e-05)),(to_sfixed_a(0.0001666163734626025)),(to_sfixed_a(2.3836444597691298e-05)),(to_sfixed_a(7.97858665464446e-05)),(to_sfixed_a(0.0008161802543327212)),(to_sfixed_a(0.004176123533397913)),(to_sfixed_a(-7.458490290446207e-05)),(to_sfixed_a(0.00015380780678242445)),(to_sfixed_a(0.0019201108952984214)),(to_sfixed_a(0.0003916447749361396)),(to_sfixed_a(0.00016940383648034185)),(to_sfixed_a(0.0001138763691415079)),(to_sfixed_a(0.0017001208616420627)),(to_sfixed_a(-1.023900586005766e-05)),(to_sfixed_a(0.00037732013151980937)),(to_sfixed_a(2.6080986572196707e-05)),(to_sfixed_a(0.0002359657228225842)),(to_sfixed_a(-0.0001875523739727214)),(to_sfixed_a(0.0034468418452888727)),(to_sfixed_a(2.817958011291921e-05)),(to_sfixed_a(0.00030468276236206293)),(to_sfixed_a(-0.0058659459464251995)),(to_sfixed_a(1.9435930880717933e-05)),(to_sfixed_a(-0.00014860945520922542)),(to_sfixed_a(0.00035907927667722106)),(to_sfixed_a(0.0002066791639663279)),(to_sfixed_a(0.00020397845946718007)),(to_sfixed_a(-0.0278580691665411)),(to_sfixed_a(-0.00020514630887191743)),(to_sfixed_a(-0.0028417722787708044)),(to_sfixed_a(-0.00280912802554667)),(to_sfixed_a(-9.120158210862428e-07)),(to_sfixed_a(5.3289295465219766e-05)),(to_sfixed_a(-3.1588642741553485e-05)),(to_sfixed_a(-0.0026106438599526882)),(to_sfixed_a(0.015422857366502285)),(to_sfixed_a(-0.0108011020347476)),(to_sfixed_a(0.00043194054160267115)),(to_sfixed_a(0.0001786010543582961)),(to_sfixed_a(0.4128873646259308)),(to_sfixed_a(-6.914834375493228e-05)),(to_sfixed_a(0.00016825165948830545)),(to_sfixed_a(-0.20416121184825897)),(to_sfixed_a(-0.5183020234107971)),(to_sfixed_a(-0.26169002056121826)),(to_sfixed_a(-4.341599196777679e-05)),(to_sfixed_a(0.3102888762950897)),(to_sfixed_a(-0.3357275426387787)),(to_sfixed_a(-0.03730224072933197)),(to_sfixed_a(0.0006648239796049893)),(to_sfixed_a(-0.0026796269230544567)),(to_sfixed_a(0.3725053668022156)),(to_sfixed_a(0.0009054893744178116)),(to_sfixed_a(-0.0003296296636108309)),(to_sfixed_a(0.00013006202061660588)),(to_sfixed_a(-3.581927376217209e-05)),(to_sfixed_a(-0.00010403215128462762)),(to_sfixed_a(-0.0019687439780682325)),(to_sfixed_a(0.0033856912050396204)),(to_sfixed_a(0.0006940080784261227)),(to_sfixed_a(-0.004200170282274485)),(to_sfixed_a(-0.004118944983929396)),(to_sfixed_a(0.14197660982608795)),(to_sfixed_a(0.00014785431267227978)),(to_sfixed_a(-0.0015032000374048948)),(to_sfixed_a(0.010381458327174187)),(to_sfixed_a(0.00017593102529644966)),(to_sfixed_a(0.21108807623386383)),(to_sfixed_a(-2.662750193849206e-05)),(to_sfixed_a(-0.6857178807258606)),(to_sfixed_a(0.0015334765193983912)),(to_sfixed_a(-0.00011226487549720332)),(to_sfixed_a(0.00013664012658409774)),(to_sfixed_a(0.00011728639947250485)),(to_sfixed_a(-0.00015558101586066186)),(to_sfixed_a(8.917407831177115e-05)),(to_sfixed_a(-0.00023959571262821555)),(to_sfixed_a(0.0002691351983230561)),(to_sfixed_a(-0.0057817925699055195)),(to_sfixed_a(0.007851636968553066)),(to_sfixed_a(-0.3450562059879303)),(to_sfixed_a(-0.32350748777389526)),(to_sfixed_a(-0.19240841269493103)),(to_sfixed_a(-1.2463780876714736e-05)),(to_sfixed_a(-6.464503530878574e-05)),(to_sfixed_a(-0.00013714583474211395)),(to_sfixed_a(-5.419953595264815e-05)),(to_sfixed_a(-3.4790809877449647e-05)),(to_sfixed_a(0.34720379114151)),(to_sfixed_a(-0.011402374133467674)),(to_sfixed_a(0.03843117132782936)),(to_sfixed_a(6.561828922713175e-05)),(to_sfixed_a(-6.420569843612611e-05)),(to_sfixed_a(0.00016656582010909915)),(to_sfixed_a(-0.00042230478720739484)),(to_sfixed_a(0.00017942534759640694)),(to_sfixed_a(0.014343501068651676)),(to_sfixed_a(-1.2010539649054408e-05)),(to_sfixed_a(-5.686011718353257e-06)),(to_sfixed_a(-4.382913175504655e-06)),(to_sfixed_a(-0.19765068590641022)),(to_sfixed_a(-0.013686945661902428)),(to_sfixed_a(-0.012322073802351952)),(to_sfixed_a(0.00029044057009741664)),(to_sfixed_a(-2.9216898838058114e-05)),(to_sfixed_a(0.00011363464000169188)),(to_sfixed_a(-0.010382001288235188)),(to_sfixed_a(0.0007792434189468622)),(to_sfixed_a(-0.36086180806159973)),(to_sfixed_a(0.00011992107465630397)),(to_sfixed_a(0.002704498590901494)),(to_sfixed_a(-0.0002992756199091673)),(to_sfixed_a(0.027091586962342262)),(to_sfixed_a(-2.5228073354810476e-05)),(to_sfixed_a(0.0005790265277028084)),(to_sfixed_a(-6.416616815840825e-05)),(to_sfixed_a(0.08440110087394714)),(to_sfixed_a(0.0006622524233534932)),(to_sfixed_a(0.2419179528951645)),(to_sfixed_a(0.008980338461697102)),(to_sfixed_a(-0.00011202030873391777)),(to_sfixed_a(0.014900117181241512)),(to_sfixed_a(-0.010992970317602158)),(to_sfixed_a(-0.00010722665319917724)),(to_sfixed_a(0.37136325240135193)),(to_sfixed_a(0.00011278274178039283)),(to_sfixed_a(0.0005215186392888427)),(to_sfixed_a(0.015097185038030148)),(to_sfixed_a(-0.01049710437655449)),(to_sfixed_a(5.986283213132992e-06)),(to_sfixed_a(-0.0001749504590407014)),(to_sfixed_a(0.46787428855895996)),(to_sfixed_a(-0.00029296494903974235)),(to_sfixed_a(-0.0019585711415857077)),(to_sfixed_a(0.00011857652862090617)),(to_sfixed_a(0.0010287011973559856)),(to_sfixed_a(2.4680120986886322e-05)),(to_sfixed_a(0.0004595533828251064)),(to_sfixed_a(-7.405796350212768e-05)),(to_sfixed_a(-0.0002429768501315266)),(to_sfixed_a(0.00012967264046892524)),(to_sfixed_a(-0.6031407713890076)),(to_sfixed_a(0.0026783959474414587)),(to_sfixed_a(0.00017570311320014298)),(to_sfixed_a(-3.820491838268936e-05)),(to_sfixed_a(8.155846444424242e-05)),(to_sfixed_a(-0.0004248922341503203)),(to_sfixed_a(0.18246771395206451)),(to_sfixed_a(-0.18046315014362335)),(to_sfixed_a(-0.0010006690863519907)),(to_sfixed_a(-0.00914449617266655)),(to_sfixed_a(-0.00022202881518751383)),(to_sfixed_a(-6.529748497996479e-05)),(to_sfixed_a(2.1415151422843337e-05)),(to_sfixed_a(2.1076299162814394e-05)),(to_sfixed_a(-0.0010747292544692755)),(to_sfixed_a(-0.00011183533933945)),(to_sfixed_a(-0.0001808044034987688)),(to_sfixed_a(-0.005631266627460718)),(to_sfixed_a(-0.1370037943124771)),(to_sfixed_a(6.522091280203313e-05)),(to_sfixed_a(0.003239980898797512)),(to_sfixed_a(-0.00036870039184577763)),(to_sfixed_a(-0.00560429273173213)),(to_sfixed_a(0.004795054439455271)),(to_sfixed_a(-7.6376847573556e-05)),(to_sfixed_a(0.0012226466787979007)),(to_sfixed_a(-0.003501622239127755)),(to_sfixed_a(0.0008776720496825874)),(to_sfixed_a(-0.00018334358173888177)),(to_sfixed_a(-0.00828663632273674)),(to_sfixed_a(0.3121439218521118)),(to_sfixed_a(0.002371125156059861)));

    constant weight_n2_52 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.06524267792701721)),(to_sfixed_a(-0.003196715610101819)),(to_sfixed_a(-0.0010586980497464538)),(to_sfixed_a(-3.6969144275644794e-05)),(to_sfixed_a(3.7838355638086796e-05)),(to_sfixed_a(-6.740610842825845e-06)),(to_sfixed_a(0.010571543127298355)),(to_sfixed_a(0.00019402526959311217)),(to_sfixed_a(-0.00019361641898285598)),(to_sfixed_a(-0.0004508364072535187)),(to_sfixed_a(4.333368269726634e-05)),(to_sfixed_a(0.0008965543820522726)),(to_sfixed_a(0.0062926411628723145)),(to_sfixed_a(-0.0012392346980050206)),(to_sfixed_a(1.1894226190634072e-05)),(to_sfixed_a(2.8311995265539736e-05)),(to_sfixed_a(0.008337692357599735)),(to_sfixed_a(-1.508410059614107e-05)),(to_sfixed_a(-0.3618639409542084)),(to_sfixed_a(-0.002178631955757737)),(to_sfixed_a(6.634349119849503e-05)),(to_sfixed_a(0.00018228255794383585)),(to_sfixed_a(0.0009330885368399322)),(to_sfixed_a(-0.004091829061508179)),(to_sfixed_a(0.00804299395531416)),(to_sfixed_a(3.0983646865934134e-05)),(to_sfixed_a(0.00017567502800375223)),(to_sfixed_a(5.366408367990516e-05)),(to_sfixed_a(0.0008211329695768654)),(to_sfixed_a(0.0002926801680587232)),(to_sfixed_a(-0.0010798132279887795)),(to_sfixed_a(-0.0002857422223314643)),(to_sfixed_a(0.0013972235610708594)),(to_sfixed_a(0.00018903959426097572)),(to_sfixed_a(-7.122750685084611e-05)),(to_sfixed_a(-6.371863128151745e-05)),(to_sfixed_a(0.2080703228712082)),(to_sfixed_a(-0.008672905154526234)),(to_sfixed_a(0.16235283017158508)),(to_sfixed_a(4.522950257523917e-05)),(to_sfixed_a(-0.006476075854152441)),(to_sfixed_a(0.00043998996261507273)),(to_sfixed_a(-0.00013636886433232576)),(to_sfixed_a(0.00011214865662623197)),(to_sfixed_a(0.28899282217025757)),(to_sfixed_a(0.0063480194658041)),(to_sfixed_a(0.25488948822021484)),(to_sfixed_a(-0.505571186542511)),(to_sfixed_a(6.72978421789594e-06)),(to_sfixed_a(0.00011000739323208109)),(to_sfixed_a(0.0004884919035248458)),(to_sfixed_a(-0.0003136518644168973)),(to_sfixed_a(-9.192249126499519e-05)),(to_sfixed_a(-0.001026161015033722)),(to_sfixed_a(0.0077893552370369434)),(to_sfixed_a(-0.0011557149700820446)),(to_sfixed_a(-0.0002712909481488168)),(to_sfixed_a(0.001025608042255044)),(to_sfixed_a(0.00023771464475430548)),(to_sfixed_a(-3.9016042137518525e-05)),(to_sfixed_a(0.0005044706631451845)),(to_sfixed_a(0.00046347850002348423)),(to_sfixed_a(-0.00010462792124599218)),(to_sfixed_a(0.004641656298190355)),(to_sfixed_a(1.7384460079483688e-05)),(to_sfixed_a(-0.4623589813709259)),(to_sfixed_a(-7.754628313705325e-05)),(to_sfixed_a(-0.28927430510520935)),(to_sfixed_a(0.00030857627280056477)),(to_sfixed_a(0.00014065054710954428)),(to_sfixed_a(0.14056004583835602)),(to_sfixed_a(-0.013344754464924335)),(to_sfixed_a(0.0022738876286894083)),(to_sfixed_a(-1.2872202205471694e-05)),(to_sfixed_a(0.00045449897879734635)),(to_sfixed_a(0.00031502905767410994)),(to_sfixed_a(0.5096272230148315)),(to_sfixed_a(-0.005257018841803074)),(to_sfixed_a(-0.0001303316093981266)),(to_sfixed_a(0.6212862133979797)),(to_sfixed_a(0.002565076109021902)),(to_sfixed_a(-7.825481588952243e-05)),(to_sfixed_a(-0.00275541958399117)),(to_sfixed_a(-0.0027408646419644356)),(to_sfixed_a(0.00019678677199408412)),(to_sfixed_a(0.010619936510920525)),(to_sfixed_a(-0.002693610731512308)),(to_sfixed_a(0.35129985213279724)),(to_sfixed_a(2.9920156521257013e-06)),(to_sfixed_a(-6.03932530793827e-05)),(to_sfixed_a(0.0028498503379523754)),(to_sfixed_a(-4.594178972183727e-05)),(to_sfixed_a(0.004860149696469307)),(to_sfixed_a(-6.026432674843818e-05)),(to_sfixed_a(-0.0005698114982806146)),(to_sfixed_a(-6.013084203004837e-06)),(to_sfixed_a(1.0160372767131776e-05)),(to_sfixed_a(0.000215659718378447)),(to_sfixed_a(-6.349684554152191e-05)),(to_sfixed_a(-0.00025143491802737117)),(to_sfixed_a(-0.0033217105083167553)),(to_sfixed_a(-0.0027458257973194122)),(to_sfixed_a(0.00016770558431744576)),(to_sfixed_a(-0.0007641965639777482)),(to_sfixed_a(0.5861424803733826)),(to_sfixed_a(-0.0005067919264547527)),(to_sfixed_a(-8.551475912099704e-05)),(to_sfixed_a(3.801454295171425e-05)),(to_sfixed_a(7.321721932385117e-05)),(to_sfixed_a(0.0010362777393311262)),(to_sfixed_a(-0.39307326078414917)),(to_sfixed_a(-3.962579648941755e-05)),(to_sfixed_a(-0.28386572003364563)),(to_sfixed_a(8.589625940658152e-05)),(to_sfixed_a(1.6207166481763124e-05)),(to_sfixed_a(-0.00462455116212368)),(to_sfixed_a(0.4871586561203003)),(to_sfixed_a(0.08411522209644318)),(to_sfixed_a(-1.8265061953570694e-05)),(to_sfixed_a(-0.0003026441263500601)),(to_sfixed_a(-0.0004194549983367324)),(to_sfixed_a(0.00011642864410532638)),(to_sfixed_a(-0.4730064868927002)),(to_sfixed_a(-0.00011341294157318771)),(to_sfixed_a(1.2134805729147047e-06)),(to_sfixed_a(0.0032122046686708927)),(to_sfixed_a(-0.0032795441802591085)),(to_sfixed_a(-0.0001610197068657726)),(to_sfixed_a(0.0001888964034151286)),(to_sfixed_a(2.3127358872443438e-06)),(to_sfixed_a(0.00016814874834381044)),(to_sfixed_a(-4.461071512196213e-07)),(to_sfixed_a(-0.0022922453936189413)),(to_sfixed_a(0.0023858475033193827)),(to_sfixed_a(-6.51484660920687e-05)),(to_sfixed_a(-0.00010125673725269735)),(to_sfixed_a(0.006474669091403484)),(to_sfixed_a(1.8982689653057605e-05)),(to_sfixed_a(0.0002959890116471797)),(to_sfixed_a(0.00014959656982682645)),(to_sfixed_a(-0.5175394415855408)),(to_sfixed_a(-0.00017627204942982644)),(to_sfixed_a(3.68481851182878e-05)),(to_sfixed_a(1.0599937013466842e-05)),(to_sfixed_a(-0.0012550707906484604)),(to_sfixed_a(0.00017112278146669269)),(to_sfixed_a(0.0001954797189682722)),(to_sfixed_a(1.0591145837679505e-05)),(to_sfixed_a(0.00014897927758283913)),(to_sfixed_a(-0.0010192259214818478)),(to_sfixed_a(0.0002970771165564656)),(to_sfixed_a(3.0105351470410824e-05)),(to_sfixed_a(0.3090054988861084)),(to_sfixed_a(-6.500638846773654e-05)),(to_sfixed_a(3.3391730539733544e-05)),(to_sfixed_a(0.24666942656040192)),(to_sfixed_a(5.76349557377398e-05)),(to_sfixed_a(0.0013244114816188812)),(to_sfixed_a(-2.3121567210182548e-05)),(to_sfixed_a(-0.00026627880288287997)),(to_sfixed_a(2.5234065105905756e-05)),(to_sfixed_a(-0.00010531947191338986)),(to_sfixed_a(6.417452823370695e-05)),(to_sfixed_a(-0.00156799191609025)),(to_sfixed_a(0.0004285048053134233)),(to_sfixed_a(0.004543467424809933)),(to_sfixed_a(-4.0481972973793745e-07)),(to_sfixed_a(0.0007838192395865917)),(to_sfixed_a(9.563111962052062e-05)),(to_sfixed_a(-0.0001680606510490179)),(to_sfixed_a(0.012988310307264328)),(to_sfixed_a(-0.0035454609896987677)),(to_sfixed_a(0.003157511819154024)),(to_sfixed_a(-2.5050336262211204e-05)),(to_sfixed_a(0.06663773208856583)),(to_sfixed_a(0.0032496503554284573)),(to_sfixed_a(6.2017970776651055e-06)),(to_sfixed_a(0.0007582632824778557)),(to_sfixed_a(0.16723734140396118)),(to_sfixed_a(0.0036093576345592737)),(to_sfixed_a(-0.001878611627034843)),(to_sfixed_a(0.00010821786418091506)),(to_sfixed_a(-0.00011267293302807957)),(to_sfixed_a(0.00011645813356153667)),(to_sfixed_a(0.00013417478476185352)),(to_sfixed_a(0.0029662202578037977)),(to_sfixed_a(-0.22977565228939056)),(to_sfixed_a(-0.003066964680328965)),(to_sfixed_a(-0.0005092251230962574)),(to_sfixed_a(0.2415827065706253)),(to_sfixed_a(-0.0009645993704907596)),(to_sfixed_a(-0.0002204972697654739)),(to_sfixed_a(-0.2295711189508438)),(to_sfixed_a(0.0021165695507079363)),(to_sfixed_a(-3.230439324397594e-05)),(to_sfixed_a(0.0033667548559606075)),(to_sfixed_a(-2.4611355911474675e-05)),(to_sfixed_a(-0.002198603004217148)),(to_sfixed_a(0.01037590391933918)),(to_sfixed_a(-0.0001530372683191672)),(to_sfixed_a(-0.00031304676667787135)),(to_sfixed_a(0.00011924670252483338)),(to_sfixed_a(-0.0002431464963592589)),(to_sfixed_a(3.285666389274411e-05)),(to_sfixed_a(-0.00017987257160712034)),(to_sfixed_a(7.254523370647803e-05)),(to_sfixed_a(0.13738352060317993)),(to_sfixed_a(0.334106981754303)),(to_sfixed_a(-0.0014182263985276222)),(to_sfixed_a(0.21134017407894135)),(to_sfixed_a(-0.01579553820192814)),(to_sfixed_a(0.00013012628187425435)),(to_sfixed_a(4.5632419642060995e-05)),(to_sfixed_a(6.610910349991173e-05)),(to_sfixed_a(-0.00011026819265680388)),(to_sfixed_a(-0.00030962645541876554)),(to_sfixed_a(0.00023672338284086436)),(to_sfixed_a(0.003091333666816354)),(to_sfixed_a(-0.018713615834712982)),(to_sfixed_a(-8.952003554441035e-06)),(to_sfixed_a(0.0001685561437625438)),(to_sfixed_a(1.0051691788248718e-05)),(to_sfixed_a(0.00027293642051517963)),(to_sfixed_a(7.02047036611475e-05)),(to_sfixed_a(0.004019342828541994)),(to_sfixed_a(-0.0003125234507024288)),(to_sfixed_a(0.00013354937254916877)),(to_sfixed_a(-0.0002141204895451665)),(to_sfixed_a(0.46547070145606995)),(to_sfixed_a(0.0024059081915766)),(to_sfixed_a(-0.0063948193565011024)),(to_sfixed_a(0.00011688156519085169)),(to_sfixed_a(9.793560457183048e-05)),(to_sfixed_a(-0.00011675462883431464)),(to_sfixed_a(0.007465344853699207)),(to_sfixed_a(0.00021051152725704014)),(to_sfixed_a(-0.003613702952861786)),(to_sfixed_a(1.5492434613406658e-05)),(to_sfixed_a(-0.0017471647588536143)),(to_sfixed_a(-0.000290677446173504)),(to_sfixed_a(-0.002055530669167638)),(to_sfixed_a(0.0004474464221857488)),(to_sfixed_a(-0.0017342620994895697)),(to_sfixed_a(0.00013806117931380868)),(to_sfixed_a(-0.48472386598587036)),(to_sfixed_a(0.08400248736143112)),(to_sfixed_a(0.004237596411257982)),(to_sfixed_a(0.03863542526960373)),(to_sfixed_a(6.81709498167038e-05)),(to_sfixed_a(0.007116581313312054)),(to_sfixed_a(0.00034744635922834277)),(to_sfixed_a(6.958776793908328e-05)),(to_sfixed_a(-0.0005476415390148759)),(to_sfixed_a(-0.00012726374552585185)),(to_sfixed_a(-0.00010512817243579775)),(to_sfixed_a(0.0034233671613037586)),(to_sfixed_a(0.003176134079694748)),(to_sfixed_a(9.980978211387992e-05)),(to_sfixed_a(-3.605855454225093e-07)),(to_sfixed_a(0.007983623072504997)),(to_sfixed_a(-2.4916400434449315e-05)),(to_sfixed_a(-0.0029960437677800655)),(to_sfixed_a(0.00010131869930773973)),(to_sfixed_a(-0.0015536670107394457)),(to_sfixed_a(6.768250023014843e-05)),(to_sfixed_a(0.005735296290367842)),(to_sfixed_a(6.058676808606833e-05)),(to_sfixed_a(2.3363081709248945e-05)),(to_sfixed_a(-0.0004185524594504386)),(to_sfixed_a(0.0004496102046687156)),(to_sfixed_a(-0.004516643937677145)),(to_sfixed_a(4.935289325658232e-06)),(to_sfixed_a(0.0002683625789359212)),(to_sfixed_a(0.00018470489885658026)),(to_sfixed_a(-3.39573307428509e-05)),(to_sfixed_a(0.01121603511273861)),(to_sfixed_a(0.004109092056751251)),(to_sfixed_a(0.3914002478122711)),(to_sfixed_a(0.0015230963472276926)),(to_sfixed_a(-0.003788743633776903)),(to_sfixed_a(2.447152292006649e-05)),(to_sfixed_a(5.157825944479555e-05)),(to_sfixed_a(-0.00045229261741042137)),(to_sfixed_a(-0.0013821967877447605)),(to_sfixed_a(-7.582986290799454e-05)),(to_sfixed_a(0.0001569209125591442)),(to_sfixed_a(4.6846646000631154e-05)),(to_sfixed_a(-0.033372651785612106)),(to_sfixed_a(-3.846421168418601e-05)),(to_sfixed_a(0.4700663685798645)),(to_sfixed_a(-0.000998153118416667)),(to_sfixed_a(0.004093340132385492)),(to_sfixed_a(-0.002135914284735918)),(to_sfixed_a(0.00024161662440747023)),(to_sfixed_a(-0.0013908310793340206)),(to_sfixed_a(-0.00022156303748488426)),(to_sfixed_a(-0.0005622656317427754)),(to_sfixed_a(0.00013397051952779293)),(to_sfixed_a(0.4414817690849304)),(to_sfixed_a(-0.4473348557949066)),(to_sfixed_a(0.01756531558930874)));

    constant weight_n2_53 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.4088858366012573)),(to_sfixed_a(-0.004947203677147627)),(to_sfixed_a(0.0004935417091473937)),(to_sfixed_a(-9.485101327300072e-05)),(to_sfixed_a(-0.006575233768671751)),(to_sfixed_a(-3.621308133006096e-05)),(to_sfixed_a(-0.004966354463249445)),(to_sfixed_a(-0.00010723886953201145)),(to_sfixed_a(-7.827195076970384e-05)),(to_sfixed_a(-1.8505779735278338e-05)),(to_sfixed_a(0.0001492960873292759)),(to_sfixed_a(-0.0007033932488411665)),(to_sfixed_a(0.4187249541282654)),(to_sfixed_a(0.0037218634970486164)),(to_sfixed_a(-6.758278323104605e-05)),(to_sfixed_a(-0.00030093968962319195)),(to_sfixed_a(-0.0052515193819999695)),(to_sfixed_a(0.00030055874958634377)),(to_sfixed_a(-0.05585808679461479)),(to_sfixed_a(0.011934835463762283)),(to_sfixed_a(1.9813684048131108e-05)),(to_sfixed_a(7.059607014525682e-07)),(to_sfixed_a(3.4305812732782215e-05)),(to_sfixed_a(0.0009394004591740668)),(to_sfixed_a(-0.005678043235093355)),(to_sfixed_a(-0.004478564020246267)),(to_sfixed_a(-6.822565046604723e-05)),(to_sfixed_a(0.00018719019135460258)),(to_sfixed_a(-0.0008381491061300039)),(to_sfixed_a(0.00028941762866452336)),(to_sfixed_a(-0.6821476221084595)),(to_sfixed_a(-9.101413888856769e-05)),(to_sfixed_a(-0.005696902517229319)),(to_sfixed_a(1.4177596312947571e-05)),(to_sfixed_a(-4.591274773702025e-06)),(to_sfixed_a(0.00041712907841429114)),(to_sfixed_a(-0.006566837430000305)),(to_sfixed_a(-8.980801794677973e-06)),(to_sfixed_a(0.26679527759552)),(to_sfixed_a(7.414501305902377e-05)),(to_sfixed_a(-0.028671784326434135)),(to_sfixed_a(0.0025381906889379025)),(to_sfixed_a(-0.00010330394434276968)),(to_sfixed_a(-0.000406509090680629)),(to_sfixed_a(0.0002719741896726191)),(to_sfixed_a(-4.029223418910988e-05)),(to_sfixed_a(-0.31482163071632385)),(to_sfixed_a(-0.001647871918976307)),(to_sfixed_a(-9.385466546518728e-05)),(to_sfixed_a(-0.026063045486807823)),(to_sfixed_a(-0.002585784997791052)),(to_sfixed_a(-0.0006339988321997225)),(to_sfixed_a(0.00010995985940098763)),(to_sfixed_a(-0.000992374261841178)),(to_sfixed_a(-0.005346399731934071)),(to_sfixed_a(-0.015695830807089806)),(to_sfixed_a(-0.00015321196406148374)),(to_sfixed_a(0.000483682204503566)),(to_sfixed_a(1.1976033420069143e-05)),(to_sfixed_a(0.00010501734504941851)),(to_sfixed_a(-0.000516161322593689)),(to_sfixed_a(0.001497533405199647)),(to_sfixed_a(-0.0004670446505770087)),(to_sfixed_a(-0.001924623386003077)),(to_sfixed_a(3.7057758163427934e-05)),(to_sfixed_a(0.0007124810363166034)),(to_sfixed_a(-0.00020550757471937686)),(to_sfixed_a(0.0012635525781661272)),(to_sfixed_a(-0.006682675331830978)),(to_sfixed_a(2.6097990485141054e-05)),(to_sfixed_a(-0.012666876427829266)),(to_sfixed_a(-0.016628792509436607)),(to_sfixed_a(-0.02750157006084919)),(to_sfixed_a(-7.485543756047264e-05)),(to_sfixed_a(-3.086292781517841e-05)),(to_sfixed_a(-0.0001521184021839872)),(to_sfixed_a(-0.0022700554691255093)),(to_sfixed_a(-0.004170041531324387)),(to_sfixed_a(0.0002197600551880896)),(to_sfixed_a(-0.006109387613832951)),(to_sfixed_a(0.0025003980845212936)),(to_sfixed_a(5.512774805538356e-06)),(to_sfixed_a(-0.0025130249559879303)),(to_sfixed_a(-7.959073991514742e-05)),(to_sfixed_a(0.00028862213366664946)),(to_sfixed_a(-0.00041044646059162915)),(to_sfixed_a(0.0047336360439658165)),(to_sfixed_a(0.00014507495507132262)),(to_sfixed_a(-0.0001353810221189633)),(to_sfixed_a(0.00016749388305470347)),(to_sfixed_a(-0.0036415811628103256)),(to_sfixed_a(-2.637068973854184e-06)),(to_sfixed_a(0.00046161137288436294)),(to_sfixed_a(-0.00029255403205752373)),(to_sfixed_a(0.3330961763858795)),(to_sfixed_a(4.790692764800042e-05)),(to_sfixed_a(-9.265328844776377e-05)),(to_sfixed_a(-0.0003037467831745744)),(to_sfixed_a(9.195689926855266e-05)),(to_sfixed_a(-6.918392318766564e-05)),(to_sfixed_a(-0.00039547838969156146)),(to_sfixed_a(0.10721052438020706)),(to_sfixed_a(-0.0001279098796658218)),(to_sfixed_a(0.004436127375811338)),(to_sfixed_a(-0.027778886258602142)),(to_sfixed_a(-3.3023727155523375e-05)),(to_sfixed_a(0.00011610717774601653)),(to_sfixed_a(-0.00010348526848247275)),(to_sfixed_a(-0.00014810109860263765)),(to_sfixed_a(-0.0038648026529699564)),(to_sfixed_a(0.005010565277189016)),(to_sfixed_a(-2.3294192942557856e-05)),(to_sfixed_a(-0.004160770680755377)),(to_sfixed_a(-0.0002018586383201182)),(to_sfixed_a(-6.880451110191643e-05)),(to_sfixed_a(-0.0020960946567356586)),(to_sfixed_a(0.09868279099464417)),(to_sfixed_a(0.00019713136134669185)),(to_sfixed_a(-4.3793508666567504e-05)),(to_sfixed_a(0.0004796396242454648)),(to_sfixed_a(-1.4329198165796697e-05)),(to_sfixed_a(-0.00010432570707052946)),(to_sfixed_a(-0.00012406238238327205)),(to_sfixed_a(4.068003181600943e-05)),(to_sfixed_a(5.997602784191258e-05)),(to_sfixed_a(-0.0014700267929583788)),(to_sfixed_a(-0.000859788793604821)),(to_sfixed_a(-4.77068533655256e-06)),(to_sfixed_a(6.426605250453576e-05)),(to_sfixed_a(3.99789132643491e-05)),(to_sfixed_a(8.09076736913994e-05)),(to_sfixed_a(2.380781006650068e-05)),(to_sfixed_a(-0.003565294435247779)),(to_sfixed_a(-0.0039019123651087284)),(to_sfixed_a(5.877784133190289e-05)),(to_sfixed_a(-4.3573512812145054e-05)),(to_sfixed_a(-0.5116034150123596)),(to_sfixed_a(-0.0010218870593234897)),(to_sfixed_a(0.0002679739845916629)),(to_sfixed_a(-0.00017421290976926684)),(to_sfixed_a(-0.00010873240535147488)),(to_sfixed_a(6.627316906815395e-05)),(to_sfixed_a(3.5165568988304585e-05)),(to_sfixed_a(2.3724202037556097e-05)),(to_sfixed_a(-0.0009120692848227918)),(to_sfixed_a(-7.580621604574844e-05)),(to_sfixed_a(-0.00297724362462759)),(to_sfixed_a(-6.087208021199331e-05)),(to_sfixed_a(0.00023802007490303367)),(to_sfixed_a(-0.004245801828801632)),(to_sfixed_a(-4.574286504066549e-05)),(to_sfixed_a(-8.899785461835563e-05)),(to_sfixed_a(0.00014923645358067006)),(to_sfixed_a(-0.00011433252802817151)),(to_sfixed_a(-4.529874786385335e-05)),(to_sfixed_a(0.0003082775219809264)),(to_sfixed_a(-0.0001160846950369887)),(to_sfixed_a(0.006039824336767197)),(to_sfixed_a(1.0342278983443975e-05)),(to_sfixed_a(-0.00011315970914438367)),(to_sfixed_a(0.0003225863038096577)),(to_sfixed_a(-0.0001126554561778903)),(to_sfixed_a(0.24095579981803894)),(to_sfixed_a(-0.0032722419127821922)),(to_sfixed_a(-0.5173746347427368)),(to_sfixed_a(0.000757597095798701)),(to_sfixed_a(0.0001359243324259296)),(to_sfixed_a(-0.004073726013302803)),(to_sfixed_a(0.00041408787365071476)),(to_sfixed_a(-6.411383219528943e-05)),(to_sfixed_a(-0.012871021404862404)),(to_sfixed_a(-0.0065768808126449585)),(to_sfixed_a(-0.003191944444552064)),(to_sfixed_a(-1.2121137842768803e-05)),(to_sfixed_a(0.0017559684347361326)),(to_sfixed_a(1.2935936865687836e-05)),(to_sfixed_a(0.018618520349264145)),(to_sfixed_a(0.0006078844889998436)),(to_sfixed_a(0.0015466561308130622)),(to_sfixed_a(-0.4589572250843048)),(to_sfixed_a(-0.0004175754147581756)),(to_sfixed_a(-0.011704287491738796)),(to_sfixed_a(0.00013131108426023275)),(to_sfixed_a(-0.00025144542451016605)),(to_sfixed_a(0.0003839524579234421)),(to_sfixed_a(0.2885942757129669)),(to_sfixed_a(-0.009271778166294098)),(to_sfixed_a(-0.0019299436826258898)),(to_sfixed_a(0.0018088852521032095)),(to_sfixed_a(2.9451126465573907e-05)),(to_sfixed_a(0.016238674521446228)),(to_sfixed_a(3.731547622010112e-06)),(to_sfixed_a(0.004033894278109074)),(to_sfixed_a(-0.014113343320786953)),(to_sfixed_a(-6.86878920532763e-05)),(to_sfixed_a(-0.0061678760685026646)),(to_sfixed_a(-0.00011279356840532273)),(to_sfixed_a(-0.0003091417602263391)),(to_sfixed_a(-0.27661648392677307)),(to_sfixed_a(0.00012051505473209545)),(to_sfixed_a(-9.860342834144831e-05)),(to_sfixed_a(9.137656888924539e-07)),(to_sfixed_a(-8.793490269454196e-05)),(to_sfixed_a(0.0002895131183322519)),(to_sfixed_a(-0.00010148222645511851)),(to_sfixed_a(0.0001501519582234323)),(to_sfixed_a(-0.11915649473667145)),(to_sfixed_a(0.28040963411331177)),(to_sfixed_a(-0.0003907366772182286)),(to_sfixed_a(-0.0062302458100020885)),(to_sfixed_a(0.2338622510433197)),(to_sfixed_a(0.00024059318820945919)),(to_sfixed_a(-0.00010426182416267693)),(to_sfixed_a(-0.00020167554612271488)),(to_sfixed_a(0.00024009586195461452)),(to_sfixed_a(0.00019965152023360133)),(to_sfixed_a(0.002461434807628393)),(to_sfixed_a(0.0008991275681182742)),(to_sfixed_a(-0.027832036837935448)),(to_sfixed_a(-0.00027005749871023)),(to_sfixed_a(-0.0003210742142982781)),(to_sfixed_a(4.435126902535558e-05)),(to_sfixed_a(-2.6912122848443687e-05)),(to_sfixed_a(7.477428880520165e-06)),(to_sfixed_a(-0.4760521352291107)),(to_sfixed_a(-0.00018728349823504686)),(to_sfixed_a(-0.00011702307529048994)),(to_sfixed_a(-0.00010598699009278789)),(to_sfixed_a(0.0018373795319348574)),(to_sfixed_a(-0.7322578430175781)),(to_sfixed_a(-0.010178769007325172)),(to_sfixed_a(-0.00015112491382751614)),(to_sfixed_a(-0.0002900476101785898)),(to_sfixed_a(6.23675441602245e-05)),(to_sfixed_a(0.0009379533585160971)),(to_sfixed_a(0.011972315609455109)),(to_sfixed_a(0.001056350884027779)),(to_sfixed_a(-9.808994946070015e-05)),(to_sfixed_a(5.135536048328504e-05)),(to_sfixed_a(0.00021518944413401186)),(to_sfixed_a(-0.011264569126069546)),(to_sfixed_a(-0.00032332519185729325)),(to_sfixed_a(0.012832553125917912)),(to_sfixed_a(-0.0004208926111459732)),(to_sfixed_a(0.00872199796140194)),(to_sfixed_a(0.4394792318344116)),(to_sfixed_a(-0.026766043156385422)),(to_sfixed_a(-0.0010109452996402979)),(to_sfixed_a(0.0003033233806490898)),(to_sfixed_a(0.0005003963015042245)),(to_sfixed_a(0.0006975920405238867)),(to_sfixed_a(0.00013996662164572626)),(to_sfixed_a(0.0018679893109947443)),(to_sfixed_a(0.00021047733025625348)),(to_sfixed_a(0.00011101817653980106)),(to_sfixed_a(-0.011713827960193157)),(to_sfixed_a(0.005771535448729992)),(to_sfixed_a(-0.00014649283548351377)),(to_sfixed_a(-0.00010213694622507319)),(to_sfixed_a(-0.001019441056996584)),(to_sfixed_a(-0.0002183928736485541)),(to_sfixed_a(-0.0011778379557654262)),(to_sfixed_a(7.838886813260615e-05)),(to_sfixed_a(-0.0005235193530097604)),(to_sfixed_a(-7.687298057135195e-05)),(to_sfixed_a(-0.008315486833453178)),(to_sfixed_a(-0.00017279875464737415)),(to_sfixed_a(-0.0001823570637498051)),(to_sfixed_a(0.00022978548076935112)),(to_sfixed_a(-0.002996508264914155)),(to_sfixed_a(0.016265535727143288)),(to_sfixed_a(-3.038070644834079e-05)),(to_sfixed_a(-5.899804818909615e-05)),(to_sfixed_a(0.00010859256144613028)),(to_sfixed_a(-0.00017446934361942112)),(to_sfixed_a(-0.013859210535883904)),(to_sfixed_a(-0.0023187671322375536)),(to_sfixed_a(0.10515902191400528)),(to_sfixed_a(-0.07937967032194138)),(to_sfixed_a(-0.0015445258468389511)),(to_sfixed_a(-2.5365938199684024e-05)),(to_sfixed_a(-0.00012598828470800072)),(to_sfixed_a(-0.00021770074090454727)),(to_sfixed_a(0.010759834200143814)),(to_sfixed_a(5.95137826167047e-05)),(to_sfixed_a(0.00018602792988531291)),(to_sfixed_a(0.008615195751190186)),(to_sfixed_a(0.5055281519889832)),(to_sfixed_a(-0.00023740454344078898)),(to_sfixed_a(-0.0003631913859862834)),(to_sfixed_a(-0.00034761434653773904)),(to_sfixed_a(-0.004601949360221624)),(to_sfixed_a(-0.005516081117093563)),(to_sfixed_a(-0.00013460477930493653)),(to_sfixed_a(-0.0028206496499478817)),(to_sfixed_a(0.01478083711117506)),(to_sfixed_a(-0.0007870743284001946)),(to_sfixed_a(0.00023127731401473284)),(to_sfixed_a(0.3940190076828003)),(to_sfixed_a(0.0011837490601465106)),(to_sfixed_a(-0.003649928607046604)));

    constant weight_n2_54 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.19265209138393402)),(to_sfixed_a(-0.0024451296776533127)),(to_sfixed_a(0.003923745360225439)),(to_sfixed_a(-0.00041316793067380786)),(to_sfixed_a(0.29906901717185974)),(to_sfixed_a(-3.1827628845348954e-05)),(to_sfixed_a(-0.0043039945885539055)),(to_sfixed_a(2.3657030396861956e-05)),(to_sfixed_a(-6.685966218356043e-05)),(to_sfixed_a(-0.00011420845112297684)),(to_sfixed_a(-6.131101690698415e-05)),(to_sfixed_a(0.00023612652148585767)),(to_sfixed_a(-0.0011363074881955981)),(to_sfixed_a(0.004735007882118225)),(to_sfixed_a(-6.534100975841284e-05)),(to_sfixed_a(0.00024699399364180863)),(to_sfixed_a(-0.04392661154270172)),(to_sfixed_a(-2.4046385078690946e-06)),(to_sfixed_a(0.36482784152030945)),(to_sfixed_a(0.0011192351812496781)),(to_sfixed_a(2.684290666365996e-05)),(to_sfixed_a(-7.020728662610054e-05)),(to_sfixed_a(0.00044341228203848004)),(to_sfixed_a(0.007238556165248156)),(to_sfixed_a(-0.006661165971308947)),(to_sfixed_a(-0.004933822900056839)),(to_sfixed_a(3.772586569539271e-05)),(to_sfixed_a(0.0024262811057269573)),(to_sfixed_a(-1.2508753570728004e-05)),(to_sfixed_a(-4.6428467612713575e-06)),(to_sfixed_a(-0.10628621280193329)),(to_sfixed_a(3.4503966162446886e-05)),(to_sfixed_a(0.009337982162833214)),(to_sfixed_a(-3.0792169127380475e-05)),(to_sfixed_a(-1.0902149369940162e-06)),(to_sfixed_a(-3.943160845665261e-05)),(to_sfixed_a(-0.0005789247225038707)),(to_sfixed_a(0.004171160515397787)),(to_sfixed_a(0.0006029352080076933)),(to_sfixed_a(0.00017788067634683102)),(to_sfixed_a(0.010633337311446667)),(to_sfixed_a(0.005382264498621225)),(to_sfixed_a(-4.3100884795421734e-05)),(to_sfixed_a(1.820515899453312e-05)),(to_sfixed_a(-0.005636618006974459)),(to_sfixed_a(-0.002632878953590989)),(to_sfixed_a(-0.35644450783729553)),(to_sfixed_a(0.3572344481945038)),(to_sfixed_a(0.00011664917838061228)),(to_sfixed_a(-0.00373259955085814)),(to_sfixed_a(-0.007179485633969307)),(to_sfixed_a(-0.0002229191013611853)),(to_sfixed_a(-1.6311016224790365e-05)),(to_sfixed_a(0.0006633583689108491)),(to_sfixed_a(-0.007892664521932602)),(to_sfixed_a(-0.007347405422478914)),(to_sfixed_a(6.94787158863619e-05)),(to_sfixed_a(-0.00174221012275666)),(to_sfixed_a(-0.00019877144950442016)),(to_sfixed_a(7.896088209236041e-05)),(to_sfixed_a(-0.0014079053653404117)),(to_sfixed_a(2.7382471671444364e-05)),(to_sfixed_a(0.0006891007069498301)),(to_sfixed_a(0.23912765085697174)),(to_sfixed_a(0.00015542173059657216)),(to_sfixed_a(0.0014696716098114848)),(to_sfixed_a(-4.682575672632083e-05)),(to_sfixed_a(0.6113263368606567)),(to_sfixed_a(-0.0010677645914256573)),(to_sfixed_a(0.000117538555059582)),(to_sfixed_a(0.009211448021233082)),(to_sfixed_a(0.003272949019446969)),(to_sfixed_a(-0.0017706610960885882)),(to_sfixed_a(-6.289116572588682e-05)),(to_sfixed_a(2.6941634132526815e-05)),(to_sfixed_a(4.5286746171768755e-05)),(to_sfixed_a(-0.06965257227420807)),(to_sfixed_a(0.004299406427890062)),(to_sfixed_a(0.0003128224052488804)),(to_sfixed_a(0.004367210902273655)),(to_sfixed_a(-0.0029617154505103827)),(to_sfixed_a(-0.00014567148173227906)),(to_sfixed_a(0.00019334422540850937)),(to_sfixed_a(-0.002909279428422451)),(to_sfixed_a(0.00023866274568717927)),(to_sfixed_a(-0.0013363491743803024)),(to_sfixed_a(0.2680630087852478)),(to_sfixed_a(0.00012032382073812187)),(to_sfixed_a(0.00016499026969540864)),(to_sfixed_a(-2.3289991077035666e-05)),(to_sfixed_a(0.0025400256272405386)),(to_sfixed_a(-1.507924753241241e-05)),(to_sfixed_a(0.0006184803787618876)),(to_sfixed_a(-2.7061119908466935e-05)),(to_sfixed_a(0.01570981554687023)),(to_sfixed_a(-1.5965088095981628e-05)),(to_sfixed_a(0.00013353314716368914)),(to_sfixed_a(-0.00014875353372190148)),(to_sfixed_a(0.00032121999538503587)),(to_sfixed_a(-1.0128163921763189e-05)),(to_sfixed_a(-0.0018532575340941548)),(to_sfixed_a(0.008010899648070335)),(to_sfixed_a(-5.927229722146876e-05)),(to_sfixed_a(0.005185646470636129)),(to_sfixed_a(0.11408152431249619)),(to_sfixed_a(-0.003426586277782917)),(to_sfixed_a(4.1270752262789756e-05)),(to_sfixed_a(7.481418288080022e-05)),(to_sfixed_a(-0.00014923773414921016)),(to_sfixed_a(-0.00237478269264102)),(to_sfixed_a(-0.00028512769495137036)),(to_sfixed_a(-0.0002641452301759273)),(to_sfixed_a(0.5664883255958557)),(to_sfixed_a(0.0001802719198167324)),(to_sfixed_a(2.981346915476024e-05)),(to_sfixed_a(0.004619360901415348)),(to_sfixed_a(0.006920063868165016)),(to_sfixed_a(-0.0027636652812361717)),(to_sfixed_a(5.958581095910631e-05)),(to_sfixed_a(0.0035569374449551105)),(to_sfixed_a(-0.000168726866832003)),(to_sfixed_a(0.00010097583435708657)),(to_sfixed_a(0.005583855789154768)),(to_sfixed_a(-0.00017981103155761957)),(to_sfixed_a(0.00012911857629660517)),(to_sfixed_a(0.0014943428104743361)),(to_sfixed_a(-0.015547122806310654)),(to_sfixed_a(0.00018168363021686673)),(to_sfixed_a(3.175191523041576e-05)),(to_sfixed_a(6.944646884221584e-05)),(to_sfixed_a(0.00013528364070225507)),(to_sfixed_a(3.927743819076568e-05)),(to_sfixed_a(-0.25245222449302673)),(to_sfixed_a(0.009992532432079315)),(to_sfixed_a(-0.00013298835256136954)),(to_sfixed_a(0.00015203548537101597)),(to_sfixed_a(-0.007684173993766308)),(to_sfixed_a(0.0024394006468355656)),(to_sfixed_a(1.9002705812454224e-05)),(to_sfixed_a(-0.00018014652596320957)),(to_sfixed_a(0.008617526851594448)),(to_sfixed_a(-0.00010663471766747534)),(to_sfixed_a(-0.00022738731058780104)),(to_sfixed_a(0.00020424154354259372)),(to_sfixed_a(-0.37627625465393066)),(to_sfixed_a(0.002435401314869523)),(to_sfixed_a(0.00010591535829007626)),(to_sfixed_a(0.00010060802014777437)),(to_sfixed_a(0.00018371851183474064)),(to_sfixed_a(-0.009363939054310322)),(to_sfixed_a(9.506124479230493e-05)),(to_sfixed_a(2.6135443476960063e-05)),(to_sfixed_a(0.011311683803796768)),(to_sfixed_a(0.00022861592879053205)),(to_sfixed_a(9.817654790822417e-05)),(to_sfixed_a(0.006127969361841679)),(to_sfixed_a(-0.0004454055742826313)),(to_sfixed_a(0.0019426957005634904)),(to_sfixed_a(-5.654252163367346e-06)),(to_sfixed_a(-0.00010202421253779903)),(to_sfixed_a(7.908322004368529e-05)),(to_sfixed_a(0.0001543649414088577)),(to_sfixed_a(-0.006235712207853794)),(to_sfixed_a(-0.0006536625442095101)),(to_sfixed_a(-0.0001249477209057659)),(to_sfixed_a(0.0010575541527941823)),(to_sfixed_a(-0.000150279127410613)),(to_sfixed_a(0.3996768295764923)),(to_sfixed_a(-0.0002431934408377856)),(to_sfixed_a(2.3873075406299904e-05)),(to_sfixed_a(-0.024004502221941948)),(to_sfixed_a(-0.0023482725955545902)),(to_sfixed_a(-0.004630951676517725)),(to_sfixed_a(0.00011320706835249439)),(to_sfixed_a(-0.11940555274486542)),(to_sfixed_a(-0.0001545938866911456)),(to_sfixed_a(0.15578600764274597)),(to_sfixed_a(0.0026888656429946423)),(to_sfixed_a(-0.3240566551685333)),(to_sfixed_a(0.001676503918133676)),(to_sfixed_a(0.0005077699897810817)),(to_sfixed_a(0.15414422750473022)),(to_sfixed_a(3.7576392060145736e-05)),(to_sfixed_a(0.00012072196113876998)),(to_sfixed_a(0.0002024903369601816)),(to_sfixed_a(-0.007359403185546398)),(to_sfixed_a(-0.015915295109152794)),(to_sfixed_a(0.006830261088907719)),(to_sfixed_a(0.003424591151997447)),(to_sfixed_a(0.0027260873466730118)),(to_sfixed_a(0.009430446662008762)),(to_sfixed_a(-9.750466415425763e-05)),(to_sfixed_a(0.4044802188873291)),(to_sfixed_a(0.0034615446347743273)),(to_sfixed_a(0.00044831278501078486)),(to_sfixed_a(-0.04384544864296913)),(to_sfixed_a(-0.0002945760788861662)),(to_sfixed_a(0.003954180050641298)),(to_sfixed_a(-0.0016978479688987136)),(to_sfixed_a(-3.842415753751993e-05)),(to_sfixed_a(-0.00021862838184460998)),(to_sfixed_a(-8.551360224373639e-05)),(to_sfixed_a(-0.00017912720795720816)),(to_sfixed_a(0.00016771936498116702)),(to_sfixed_a(3.076387656619772e-05)),(to_sfixed_a(0.0007677776156924665)),(to_sfixed_a(-0.4026314914226532)),(to_sfixed_a(-0.2544156014919281)),(to_sfixed_a(0.003236297983676195)),(to_sfixed_a(0.006301191169768572)),(to_sfixed_a(0.005351838190108538)),(to_sfixed_a(-0.00011271486437181011)),(to_sfixed_a(6.917018617969006e-05)),(to_sfixed_a(-6.667439447483048e-05)),(to_sfixed_a(0.00014610822836402804)),(to_sfixed_a(0.00010866658703889698)),(to_sfixed_a(0.0032815607264637947)),(to_sfixed_a(0.0030302759259939194)),(to_sfixed_a(-0.2520693838596344)),(to_sfixed_a(-0.00015132504631765187)),(to_sfixed_a(0.00016726141620893031)),(to_sfixed_a(-8.833005267661065e-06)),(to_sfixed_a(7.606596045661718e-05)),(to_sfixed_a(0.003741135820746422)),(to_sfixed_a(0.21714021265506744)),(to_sfixed_a(-0.00015332602197304368)),(to_sfixed_a(-0.00028487585950642824)),(to_sfixed_a(-6.846408359706402e-05)),(to_sfixed_a(-0.20793041586875916)),(to_sfixed_a(-0.3436644375324249)),(to_sfixed_a(-0.05645216628909111)),(to_sfixed_a(-0.00010621469118632376)),(to_sfixed_a(-0.0001397782762069255)),(to_sfixed_a(2.4677367036929354e-05)),(to_sfixed_a(-0.0007760071312077343)),(to_sfixed_a(0.020283101126551628)),(to_sfixed_a(0.16872909665107727)),(to_sfixed_a(-0.0002398673095740378)),(to_sfixed_a(0.001192975090816617)),(to_sfixed_a(2.0523148123174906e-06)),(to_sfixed_a(-0.006466627586632967)),(to_sfixed_a(-0.00021796436340082437)),(to_sfixed_a(-0.16251790523529053)),(to_sfixed_a(0.00028655322967097163)),(to_sfixed_a(0.001850601751357317)),(to_sfixed_a(0.0016878076130524278)),(to_sfixed_a(-0.0047008320689201355)),(to_sfixed_a(0.00017599975399207324)),(to_sfixed_a(6.218752241693437e-05)),(to_sfixed_a(0.24027958512306213)),(to_sfixed_a(-0.01522605586796999)),(to_sfixed_a(3.1536579626845196e-05)),(to_sfixed_a(0.0003844103775918484)),(to_sfixed_a(-6.995955482125282e-05)),(to_sfixed_a(-0.23471280932426453)),(to_sfixed_a(-0.3275417387485504)),(to_sfixed_a(0.00024163616762962192)),(to_sfixed_a(0.00038356438744813204)),(to_sfixed_a(2.3118827812140808e-05)),(to_sfixed_a(0.3291756808757782)),(to_sfixed_a(2.439710806356743e-05)),(to_sfixed_a(-0.001047403085976839)),(to_sfixed_a(0.0001961074158316478)),(to_sfixed_a(0.0005217318539507687)),(to_sfixed_a(0.0002217428555013612)),(to_sfixed_a(-0.0026696152053773403)),(to_sfixed_a(-1.3174743799027056e-05)),(to_sfixed_a(0.0001502975937910378)),(to_sfixed_a(0.00027250187122263014)),(to_sfixed_a(-0.010361623018980026)),(to_sfixed_a(0.6415975689888)),(to_sfixed_a(-6.246305929380469e-06)),(to_sfixed_a(1.9910905393771827e-05)),(to_sfixed_a(-0.00041255546966567636)),(to_sfixed_a(-0.00010618048690957949)),(to_sfixed_a(-0.005215888377279043)),(to_sfixed_a(-0.010959464125335217)),(to_sfixed_a(-0.014006094075739384)),(to_sfixed_a(-0.16042840480804443)),(to_sfixed_a(0.0032113571651279926)),(to_sfixed_a(0.00018065868061967194)),(to_sfixed_a(-8.457628428004682e-05)),(to_sfixed_a(8.730260742595419e-05)),(to_sfixed_a(0.0005883525591343641)),(to_sfixed_a(0.00010715621465351433)),(to_sfixed_a(-2.914547803811729e-05)),(to_sfixed_a(0.0016446721274405718)),(to_sfixed_a(0.00943254865705967)),(to_sfixed_a(-0.000174654574948363)),(to_sfixed_a(-0.3059370815753937)),(to_sfixed_a(0.28472429513931274)),(to_sfixed_a(-0.025887440890073776)),(to_sfixed_a(-0.0026964701246470213)),(to_sfixed_a(1.7759863112587482e-05)),(to_sfixed_a(-0.002086765132844448)),(to_sfixed_a(0.2235173135995865)),(to_sfixed_a(-0.011543996632099152)),(to_sfixed_a(4.879791958956048e-05)),(to_sfixed_a(-0.001110417302697897)),(to_sfixed_a(0.4884578287601471)),(to_sfixed_a(-0.0062498170882463455)));

    constant weight_n2_55 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.6375442743301392)),(to_sfixed_a(0.0218668095767498)),(to_sfixed_a(0.00023334889556281269)),(to_sfixed_a(0.00011225510388612747)),(to_sfixed_a(-0.3786908686161041)),(to_sfixed_a(-2.3294272978091612e-05)),(to_sfixed_a(-0.0020237858407199383)),(to_sfixed_a(3.9337523048743606e-05)),(to_sfixed_a(-7.172998448368162e-05)),(to_sfixed_a(-0.00020078112720511854)),(to_sfixed_a(-7.862896018195897e-05)),(to_sfixed_a(9.811353811528534e-05)),(to_sfixed_a(0.002422645688056946)),(to_sfixed_a(0.004332392010837793)),(to_sfixed_a(7.355538400588557e-07)),(to_sfixed_a(6.498529546661302e-05)),(to_sfixed_a(0.0004343792097643018)),(to_sfixed_a(-0.00019956272444687784)),(to_sfixed_a(0.0051700701005756855)),(to_sfixed_a(0.0016764741158112884)),(to_sfixed_a(-0.00011669230298139155)),(to_sfixed_a(0.00011185904440935701)),(to_sfixed_a(-0.0033858646638691425)),(to_sfixed_a(0.0005834954208694398)),(to_sfixed_a(-0.0005424661794677377)),(to_sfixed_a(-0.3848251700401306)),(to_sfixed_a(-1.7138976545538753e-05)),(to_sfixed_a(-0.00013602094259113073)),(to_sfixed_a(-0.0003631303843576461)),(to_sfixed_a(-0.00024956819834187627)),(to_sfixed_a(-0.794856607913971)),(to_sfixed_a(-7.156326319091022e-05)),(to_sfixed_a(6.927950744284317e-05)),(to_sfixed_a(-7.083974196575582e-06)),(to_sfixed_a(0.00012599398905877024)),(to_sfixed_a(0.00022125169925857335)),(to_sfixed_a(0.019171474501490593)),(to_sfixed_a(0.016649845987558365)),(to_sfixed_a(0.0008667559595778584)),(to_sfixed_a(0.00013031861453782767)),(to_sfixed_a(0.2868000268936157)),(to_sfixed_a(0.003141046967357397)),(to_sfixed_a(3.944421769119799e-05)),(to_sfixed_a(2.1597275917883962e-05)),(to_sfixed_a(-0.00047892401926219463)),(to_sfixed_a(-0.42769110202789307)),(to_sfixed_a(-0.2748311460018158)),(to_sfixed_a(-0.0006289297598414123)),(to_sfixed_a(5.282504571368918e-05)),(to_sfixed_a(-0.00014655129052698612)),(to_sfixed_a(-0.0006128470413386822)),(to_sfixed_a(0.0004392365226522088)),(to_sfixed_a(-5.020730895921588e-06)),(to_sfixed_a(0.001824481994844973)),(to_sfixed_a(0.0056633418425917625)),(to_sfixed_a(-0.010420112870633602)),(to_sfixed_a(6.255839252844453e-05)),(to_sfixed_a(0.00013933845912106335)),(to_sfixed_a(4.6373104851227254e-05)),(to_sfixed_a(2.214945743617136e-05)),(to_sfixed_a(-0.017440464347600937)),(to_sfixed_a(-0.0036494790110737085)),(to_sfixed_a(-0.00037243723636493087)),(to_sfixed_a(-0.00019916502060368657)),(to_sfixed_a(-8.42090230435133e-05)),(to_sfixed_a(-0.0006961926119402051)),(to_sfixed_a(-0.00021726007980760187)),(to_sfixed_a(0.0033020530827343464)),(to_sfixed_a(-0.0036451020278036594)),(to_sfixed_a(-0.00011361001816112548)),(to_sfixed_a(0.019585145637392998)),(to_sfixed_a(0.0010596190113574266)),(to_sfixed_a(-0.000730629195459187)),(to_sfixed_a(-0.0002019875100813806)),(to_sfixed_a(0.00011272115807514638)),(to_sfixed_a(-7.006590021774173e-05)),(to_sfixed_a(-0.0014613235834985971)),(to_sfixed_a(-0.0006964525091461837)),(to_sfixed_a(-0.0003032372333109379)),(to_sfixed_a(0.004388227593153715)),(to_sfixed_a(0.0007621475961059332)),(to_sfixed_a(-0.0002048061287496239)),(to_sfixed_a(0.00047399982577189803)),(to_sfixed_a(0.016271190717816353)),(to_sfixed_a(-1.8697261111810803e-05)),(to_sfixed_a(-0.0019504472147673368)),(to_sfixed_a(0.00576007179915905)),(to_sfixed_a(0.00011156135587953031)),(to_sfixed_a(-0.00015253205492626876)),(to_sfixed_a(-0.00016924800002016127)),(to_sfixed_a(0.018636027351021767)),(to_sfixed_a(-1.1792901204898953e-05)),(to_sfixed_a(-0.0005746055976487696)),(to_sfixed_a(0.0001813699782360345)),(to_sfixed_a(-0.000598078069742769)),(to_sfixed_a(0.00011613142123678699)),(to_sfixed_a(-0.00018618624017108232)),(to_sfixed_a(-0.00014915474457666278)),(to_sfixed_a(-6.156010931590572e-05)),(to_sfixed_a(-0.00011649001680780202)),(to_sfixed_a(2.478017268003896e-05)),(to_sfixed_a(-0.0003454643883742392)),(to_sfixed_a(5.850879097124562e-05)),(to_sfixed_a(0.001377678825519979)),(to_sfixed_a(8.165922190528363e-05)),(to_sfixed_a(-0.001860063406638801)),(to_sfixed_a(0.00018997352162841707)),(to_sfixed_a(0.00014925276627764106)),(to_sfixed_a(4.344976332504302e-05)),(to_sfixed_a(0.0011003438849002123)),(to_sfixed_a(0.00288376584649086)),(to_sfixed_a(-0.0002385179395787418)),(to_sfixed_a(-0.004968124441802502)),(to_sfixed_a(6.848109478596598e-06)),(to_sfixed_a(9.336413495475426e-05)),(to_sfixed_a(0.02650080993771553)),(to_sfixed_a(-0.00010664550063665956)),(to_sfixed_a(0.00025638187071308494)),(to_sfixed_a(4.688296030508354e-05)),(to_sfixed_a(0.001413037651218474)),(to_sfixed_a(-9.639615745982155e-05)),(to_sfixed_a(5.8657125919125974e-05)),(to_sfixed_a(-0.00038039934588596225)),(to_sfixed_a(-0.00014684104826301336)),(to_sfixed_a(0.00010603482951410115)),(to_sfixed_a(-0.000497153087053448)),(to_sfixed_a(-0.03205152601003647)),(to_sfixed_a(-0.0003796694800257683)),(to_sfixed_a(0.00028607298736460507)),(to_sfixed_a(0.00016531416622456163)),(to_sfixed_a(2.4614122594357468e-05)),(to_sfixed_a(-1.0887852113228291e-06)),(to_sfixed_a(0.0005960009875707328)),(to_sfixed_a(0.009224362671375275)),(to_sfixed_a(-6.869681237731129e-05)),(to_sfixed_a(0.00011746047675842419)),(to_sfixed_a(0.3807581067085266)),(to_sfixed_a(-0.00011769912816816941)),(to_sfixed_a(-0.00017445559205953032)),(to_sfixed_a(0.0004107282729819417)),(to_sfixed_a(-0.0028092728462070227)),(to_sfixed_a(2.8750702767865732e-05)),(to_sfixed_a(-0.00044549640733748674)),(to_sfixed_a(-4.118573269806802e-05)),(to_sfixed_a(-0.00035049341386184096)),(to_sfixed_a(0.0003098673769272864)),(to_sfixed_a(-0.0010808466468006372)),(to_sfixed_a(-1.0403724445495754e-05)),(to_sfixed_a(-0.00016752797819208354)),(to_sfixed_a(2.6934467314276844e-05)),(to_sfixed_a(-0.00015142426127567887)),(to_sfixed_a(4.148656444158405e-05)),(to_sfixed_a(4.5217697334010154e-05)),(to_sfixed_a(-0.0002470139879733324)),(to_sfixed_a(-7.436554733430967e-05)),(to_sfixed_a(0.0024712327867746353)),(to_sfixed_a(-2.434523412375711e-05)),(to_sfixed_a(0.1712251901626587)),(to_sfixed_a(2.0771916751982644e-05)),(to_sfixed_a(0.00015173900465015322)),(to_sfixed_a(1.128315125242807e-05)),(to_sfixed_a(4.808196536032483e-05)),(to_sfixed_a(0.00043827539775520563)),(to_sfixed_a(0.00782693736255169)),(to_sfixed_a(-0.0007732242229394615)),(to_sfixed_a(-0.004031273070722818)),(to_sfixed_a(-5.719708133256063e-05)),(to_sfixed_a(-0.0005129611818119884)),(to_sfixed_a(3.5653069062391296e-05)),(to_sfixed_a(-0.00010853767889784649)),(to_sfixed_a(-0.2862425446510315)),(to_sfixed_a(-0.0016381720779463649)),(to_sfixed_a(0.0005492378259077668)),(to_sfixed_a(7.467404793715104e-05)),(to_sfixed_a(0.0004380311002023518)),(to_sfixed_a(0.0002109915076289326)),(to_sfixed_a(-2.1471025775099406e-06)),(to_sfixed_a(-0.001201302045956254)),(to_sfixed_a(-0.006771044805645943)),(to_sfixed_a(-0.4243778884410858)),(to_sfixed_a(0.0003706346615217626)),(to_sfixed_a(-0.15609623491764069)),(to_sfixed_a(0.00011939213436562568)),(to_sfixed_a(2.1775704226456583e-06)),(to_sfixed_a(-1.94706954061985e-05)),(to_sfixed_a(-0.0001631443010410294)),(to_sfixed_a(-0.014309004880487919)),(to_sfixed_a(0.0010759546421468258)),(to_sfixed_a(0.002079110126942396)),(to_sfixed_a(0.0061779264360666275)),(to_sfixed_a(0.009644805453717709)),(to_sfixed_a(0.0001921210205182433)),(to_sfixed_a(-0.0015930181834846735)),(to_sfixed_a(-0.0009200035128742456)),(to_sfixed_a(-0.00017573742661625147)),(to_sfixed_a(-0.2614574432373047)),(to_sfixed_a(-0.00020293291890993714)),(to_sfixed_a(-0.04133779555559158)),(to_sfixed_a(0.013244256377220154)),(to_sfixed_a(-0.00027107930509373546)),(to_sfixed_a(-0.00017230561934411526)),(to_sfixed_a(-0.00013849501556251198)),(to_sfixed_a(0.00011720314068952575)),(to_sfixed_a(-2.9426810215227306e-06)),(to_sfixed_a(-6.945656787138432e-05)),(to_sfixed_a(0.001374670653603971)),(to_sfixed_a(0.0013185052666813135)),(to_sfixed_a(0.2646830081939697)),(to_sfixed_a(0.2314033806324005)),(to_sfixed_a(0.17139476537704468)),(to_sfixed_a(-0.00063657684950158)),(to_sfixed_a(-0.00015186269592959434)),(to_sfixed_a(0.0002256013103760779)),(to_sfixed_a(5.2219926146790385e-05)),(to_sfixed_a(4.211542545817792e-06)),(to_sfixed_a(-0.00022209301823750138)),(to_sfixed_a(0.0016107199480757117)),(to_sfixed_a(-0.0008674405980855227)),(to_sfixed_a(-0.0006961406907066703)),(to_sfixed_a(-3.0499271815642715e-05)),(to_sfixed_a(9.5742943813093e-05)),(to_sfixed_a(-1.383785274811089e-06)),(to_sfixed_a(0.00015211620484478772)),(to_sfixed_a(-0.00020913974731229246)),(to_sfixed_a(0.013487178832292557)),(to_sfixed_a(-0.0001213081632158719)),(to_sfixed_a(0.00028079564799554646)),(to_sfixed_a(0.0002167748025385663)),(to_sfixed_a(0.17978547513484955)),(to_sfixed_a(-0.003055207198485732)),(to_sfixed_a(0.006449887994676828)),(to_sfixed_a(-5.715388397220522e-06)),(to_sfixed_a(1.52099528349936e-06)),(to_sfixed_a(-0.00016790836525615305)),(to_sfixed_a(0.0005492537748068571)),(to_sfixed_a(0.0001084784307749942)),(to_sfixed_a(0.004065864719450474)),(to_sfixed_a(0.00014571385690942407)),(to_sfixed_a(0.004683565814048052)),(to_sfixed_a(0.00021682424994651228)),(to_sfixed_a(0.0004322166496422142)),(to_sfixed_a(-5.870476161362603e-05)),(to_sfixed_a(-0.46028706431388855)),(to_sfixed_a(-0.00011551904754014686)),(to_sfixed_a(0.00273673958145082)),(to_sfixed_a(0.002007317030802369)),(to_sfixed_a(-0.37012314796447754)),(to_sfixed_a(-0.0003470456867944449)),(to_sfixed_a(-2.2267206077231094e-05)),(to_sfixed_a(0.0004676315584219992)),(to_sfixed_a(0.00039947443292476237)),(to_sfixed_a(7.025893137324601e-05)),(to_sfixed_a(0.002206140663474798)),(to_sfixed_a(-0.00023837503977119923)),(to_sfixed_a(-0.00012611686543095857)),(to_sfixed_a(-0.0019151533488184214)),(to_sfixed_a(-0.005063435062766075)),(to_sfixed_a(0.00015804263239260763)),(to_sfixed_a(-6.986955122556537e-05)),(to_sfixed_a(0.0015713567845523357)),(to_sfixed_a(-3.830311470665038e-06)),(to_sfixed_a(-0.0019735742826014757)),(to_sfixed_a(-0.00014997342077549547)),(to_sfixed_a(0.0004002661444246769)),(to_sfixed_a(2.9440183425322175e-05)),(to_sfixed_a(-0.0017231098609045148)),(to_sfixed_a(-5.636017885990441e-05)),(to_sfixed_a(-0.00010491137800272554)),(to_sfixed_a(4.425545921549201e-05)),(to_sfixed_a(0.0004494407039601356)),(to_sfixed_a(-0.009019692428410053)),(to_sfixed_a(0.0002905250294134021)),(to_sfixed_a(-0.00029984768480062485)),(to_sfixed_a(0.00014911213656887412)),(to_sfixed_a(0.00019968883134424686)),(to_sfixed_a(-0.3220239281654358)),(to_sfixed_a(0.0053365183994174)),(to_sfixed_a(-0.15329161286354065)),(to_sfixed_a(-0.00013445108197629452)),(to_sfixed_a(0.0015962414909154177)),(to_sfixed_a(8.903371053747833e-07)),(to_sfixed_a(-0.00011241246829740703)),(to_sfixed_a(6.591992860194296e-05)),(to_sfixed_a(0.003038890426978469)),(to_sfixed_a(2.7590212994255126e-06)),(to_sfixed_a(-4.494166205404326e-05)),(to_sfixed_a(0.0018179442267864943)),(to_sfixed_a(-0.0004918399499729276)),(to_sfixed_a(-0.0001558585063321516)),(to_sfixed_a(0.018527736887335777)),(to_sfixed_a(-0.00014037374057807028)),(to_sfixed_a(-0.00121692952234298)),(to_sfixed_a(0.16210557520389557)),(to_sfixed_a(0.00012123244960093871)),(to_sfixed_a(0.0005389657453633845)),(to_sfixed_a(-0.00020868569845333695)),(to_sfixed_a(-9.811996278585866e-06)),(to_sfixed_a(8.019960660021752e-05)),(to_sfixed_a(-0.004949295427650213)),(to_sfixed_a(0.0087415911257267)),(to_sfixed_a(0.00034518615575507283)));

    constant weight_n2_56 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.5289804339408875)),(to_sfixed_a(-0.5138644576072693)),(to_sfixed_a(-0.5799198150634766)),(to_sfixed_a(-6.550394755322486e-05)),(to_sfixed_a(0.21549652516841888)),(to_sfixed_a(-1.9261751731391996e-06)),(to_sfixed_a(0.3227634131908417)),(to_sfixed_a(-6.594440492335707e-05)),(to_sfixed_a(-0.0001305236219195649)),(to_sfixed_a(3.7485078792087734e-05)),(to_sfixed_a(-1.9257986423326656e-05)),(to_sfixed_a(0.0011932097841054201)),(to_sfixed_a(-0.006689231377094984)),(to_sfixed_a(0.0069667017087340355)),(to_sfixed_a(0.0001671957434155047)),(to_sfixed_a(6.228827260201797e-05)),(to_sfixed_a(0.05809149146080017)),(to_sfixed_a(-0.00018647988326847553)),(to_sfixed_a(0.15852071344852448)),(to_sfixed_a(0.004735034424811602)),(to_sfixed_a(-0.00018523455946706235)),(to_sfixed_a(0.00022454447753261775)),(to_sfixed_a(-0.001811683876439929)),(to_sfixed_a(0.00458682794123888)),(to_sfixed_a(-0.0015829490730538964)),(to_sfixed_a(0.0011474333005025983)),(to_sfixed_a(8.008049917407334e-06)),(to_sfixed_a(-0.0009482254972681403)),(to_sfixed_a(-0.0023867846466600895)),(to_sfixed_a(-0.00017448868311475962)),(to_sfixed_a(-0.0019305185414850712)),(to_sfixed_a(-0.00011804809037130326)),(to_sfixed_a(0.4566463828086853)),(to_sfixed_a(-8.457009244011715e-05)),(to_sfixed_a(4.636236553778872e-05)),(to_sfixed_a(-0.00011182806338183582)),(to_sfixed_a(-0.2840019762516022)),(to_sfixed_a(-0.03648076206445694)),(to_sfixed_a(-0.374925434589386)),(to_sfixed_a(-0.00018637775792740285)),(to_sfixed_a(-0.10996032506227493)),(to_sfixed_a(0.004782657139003277)),(to_sfixed_a(0.00016391607641708106)),(to_sfixed_a(-0.00010282434232067317)),(to_sfixed_a(-0.008233492262661457)),(to_sfixed_a(-0.3289485573768616)),(to_sfixed_a(-0.9611774682998657)),(to_sfixed_a(-0.006054259371012449)),(to_sfixed_a(0.00022586749400943518)),(to_sfixed_a(0.0027334284968674183)),(to_sfixed_a(-0.011129016056656837)),(to_sfixed_a(0.0001527152198832482)),(to_sfixed_a(-0.00018738521612249315)),(to_sfixed_a(0.001199220190756023)),(to_sfixed_a(0.00020691224199254066)),(to_sfixed_a(-0.0007035729358904064)),(to_sfixed_a(-0.00031664996640756726)),(to_sfixed_a(0.0016973491292446852)),(to_sfixed_a(-6.795018271077424e-05)),(to_sfixed_a(0.0001015970265143551)),(to_sfixed_a(-0.013224336318671703)),(to_sfixed_a(-0.001607157289981842)),(to_sfixed_a(-0.0011583863524720073)),(to_sfixed_a(-0.012782040983438492)),(to_sfixed_a(9.819441038416699e-05)),(to_sfixed_a(-0.34128108620643616)),(to_sfixed_a(-0.00017489047604613006)),(to_sfixed_a(0.1447744369506836)),(to_sfixed_a(-0.0021664765663444996)),(to_sfixed_a(2.6808149414137006e-05)),(to_sfixed_a(-0.1774817258119583)),(to_sfixed_a(-0.2578713297843933)),(to_sfixed_a(-0.005831554066389799)),(to_sfixed_a(-9.557980229146779e-05)),(to_sfixed_a(1.7346610547974706e-05)),(to_sfixed_a(4.579745655064471e-05)),(to_sfixed_a(-0.11019852012395859)),(to_sfixed_a(-0.0021854860242456198)),(to_sfixed_a(-3.035602276213467e-05)),(to_sfixed_a(-0.19165420532226562)),(to_sfixed_a(0.257725328207016)),(to_sfixed_a(0.00015069139772094786)),(to_sfixed_a(-0.30175355076789856)),(to_sfixed_a(2.577442501205951e-05)),(to_sfixed_a(5.425249401014298e-05)),(to_sfixed_a(-0.0011443514376878738)),(to_sfixed_a(0.009009172208607197)),(to_sfixed_a(8.987884211819619e-05)),(to_sfixed_a(3.656702028820291e-05)),(to_sfixed_a(3.8178128306753933e-05)),(to_sfixed_a(-0.03265003114938736)),(to_sfixed_a(2.5488676328677684e-05)),(to_sfixed_a(-0.2710712254047394)),(to_sfixed_a(4.49320359621197e-05)),(to_sfixed_a(-0.2131192535161972)),(to_sfixed_a(1.5866628018557094e-05)),(to_sfixed_a(-0.0001948637218447402)),(to_sfixed_a(0.00018609585822559893)),(to_sfixed_a(8.544159936718643e-05)),(to_sfixed_a(0.00011352711590006948)),(to_sfixed_a(0.0030040896963328123)),(to_sfixed_a(-0.0001222378050442785)),(to_sfixed_a(-0.00013690431660506874)),(to_sfixed_a(-0.002398653654381633)),(to_sfixed_a(-0.12544700503349304)),(to_sfixed_a(-0.0005524114822037518)),(to_sfixed_a(2.3372122086584568e-05)),(to_sfixed_a(-2.3360917111858726e-05)),(to_sfixed_a(-1.0483243386261165e-05)),(to_sfixed_a(-0.00014132105570752174)),(to_sfixed_a(0.525223433971405)),(to_sfixed_a(7.889760308898985e-05)),(to_sfixed_a(-0.3833804726600647)),(to_sfixed_a(0.00016933275037445128)),(to_sfixed_a(3.272480535088107e-05)),(to_sfixed_a(-0.005441182758659124)),(to_sfixed_a(0.0012602258939296007)),(to_sfixed_a(0.0010189099702984095)),(to_sfixed_a(-9.490233060205355e-05)),(to_sfixed_a(0.0021192680578678846)),(to_sfixed_a(7.148596341721714e-05)),(to_sfixed_a(0.00011740165064111352)),(to_sfixed_a(-0.0017957452218979597)),(to_sfixed_a(0.00014838544302619994)),(to_sfixed_a(5.7014927733689547e-05)),(to_sfixed_a(-0.17420659959316254)),(to_sfixed_a(0.28030070662498474)),(to_sfixed_a(-3.2263167668133974e-05)),(to_sfixed_a(-4.778581205755472e-05)),(to_sfixed_a(-0.0001686959294602275)),(to_sfixed_a(0.00015024565800558776)),(to_sfixed_a(-0.0002897733938880265)),(to_sfixed_a(0.00035936807398684323)),(to_sfixed_a(-0.001689300173893571)),(to_sfixed_a(4.6177061449270695e-05)),(to_sfixed_a(-0.00028899736935272813)),(to_sfixed_a(-0.06360068917274475)),(to_sfixed_a(-6.301906978478655e-05)),(to_sfixed_a(7.013219146756455e-05)),(to_sfixed_a(-0.00010142241808352992)),(to_sfixed_a(-0.0024104469921439886)),(to_sfixed_a(0.00015292323951143771)),(to_sfixed_a(4.923436790704727e-06)),(to_sfixed_a(3.262012614868581e-05)),(to_sfixed_a(-0.43227827548980713)),(to_sfixed_a(-4.891111166216433e-05)),(to_sfixed_a(0.22795230150222778)),(to_sfixed_a(-0.00014793231093790382)),(to_sfixed_a(-7.593294867547229e-05)),(to_sfixed_a(0.005937769077718258)),(to_sfixed_a(6.251037120819092e-05)),(to_sfixed_a(-0.00018185655062552541)),(to_sfixed_a(-0.26733964681625366)),(to_sfixed_a(0.00011275910219410434)),(to_sfixed_a(0.00024743235553614795)),(to_sfixed_a(-0.057798758149147034)),(to_sfixed_a(0.00018895234097726643)),(to_sfixed_a(0.13426634669303894)),(to_sfixed_a(-0.00012604201037902385)),(to_sfixed_a(-0.00019740559218917042)),(to_sfixed_a(-8.967712346930057e-06)),(to_sfixed_a(-0.00027033055084757507)),(to_sfixed_a(0.3438522219657898)),(to_sfixed_a(0.005360561888664961)),(to_sfixed_a(0.0029124044813215733)),(to_sfixed_a(-0.005422793794423342)),(to_sfixed_a(-0.00029868780984543264)),(to_sfixed_a(-0.003672835184261203)),(to_sfixed_a(1.4614270185120404e-05)),(to_sfixed_a(-3.1176023185253143e-07)),(to_sfixed_a(-0.0016974004684016109)),(to_sfixed_a(-0.02194170281291008)),(to_sfixed_a(-0.005102659575641155)),(to_sfixed_a(0.00013495099847204983)),(to_sfixed_a(0.32086315751075745)),(to_sfixed_a(-0.005803131964057684)),(to_sfixed_a(0.09355256706476212)),(to_sfixed_a(0.0005986502510495484)),(to_sfixed_a(-0.37758398056030273)),(to_sfixed_a(0.004551386926323175)),(to_sfixed_a(5.5684195103822276e-05)),(to_sfixed_a(0.27633926272392273)),(to_sfixed_a(-2.470986873959191e-05)),(to_sfixed_a(1.9751591025851667e-05)),(to_sfixed_a(-0.0001513328606961295)),(to_sfixed_a(-8.184561738744378e-05)),(to_sfixed_a(-0.002251480706036091)),(to_sfixed_a(0.0012941622408106923)),(to_sfixed_a(0.0019409263040870428)),(to_sfixed_a(0.00101340317633003)),(to_sfixed_a(0.010885123163461685)),(to_sfixed_a(0.0001905124372569844)),(to_sfixed_a(0.20447689294815063)),(to_sfixed_a(-0.004566481802612543)),(to_sfixed_a(0.00018709420692175627)),(to_sfixed_a(-0.007885191589593887)),(to_sfixed_a(0.0003795029188040644)),(to_sfixed_a(0.0005471163894981146)),(to_sfixed_a(-0.031325727701187134)),(to_sfixed_a(-0.00024212425341829658)),(to_sfixed_a(-0.00013699103146791458)),(to_sfixed_a(-0.0002374984323978424)),(to_sfixed_a(-3.901839954778552e-05)),(to_sfixed_a(3.6837074731010944e-05)),(to_sfixed_a(0.000249561300734058)),(to_sfixed_a(-0.00011183541209902614)),(to_sfixed_a(-0.530627965927124)),(to_sfixed_a(0.03102012164890766)),(to_sfixed_a(0.07567651569843292)),(to_sfixed_a(-0.0017746587982401252)),(to_sfixed_a(0.003677139524370432)),(to_sfixed_a(9.142291673924774e-06)),(to_sfixed_a(0.0004153571790084243)),(to_sfixed_a(-0.0001056143082678318)),(to_sfixed_a(6.70743320370093e-05)),(to_sfixed_a(-0.0002934057847596705)),(to_sfixed_a(0.0003096050932072103)),(to_sfixed_a(0.42162594199180603)),(to_sfixed_a(0.46486419439315796)),(to_sfixed_a(-0.00011566145985852927)),(to_sfixed_a(-0.00017197709530591965)),(to_sfixed_a(-3.0231101845856756e-05)),(to_sfixed_a(6.901482993271202e-05)),(to_sfixed_a(-0.0013510679127648473)),(to_sfixed_a(-0.28048425912857056)),(to_sfixed_a(5.69624244235456e-05)),(to_sfixed_a(0.00030670114210806787)),(to_sfixed_a(-0.00017565794405527413)),(to_sfixed_a(0.1824265718460083)),(to_sfixed_a(-0.01323789358139038)),(to_sfixed_a(-0.47221294045448303)),(to_sfixed_a(-2.760575443971902e-05)),(to_sfixed_a(0.0002354138414375484)),(to_sfixed_a(0.000156841502757743)),(to_sfixed_a(-1.1490490578580648e-05)),(to_sfixed_a(0.001995253609493375)),(to_sfixed_a(-0.021030070260167122)),(to_sfixed_a(-0.00011663547775242478)),(to_sfixed_a(8.336034079547971e-05)),(to_sfixed_a(-0.00019217398948967457)),(to_sfixed_a(-0.12155783921480179)),(to_sfixed_a(-0.00016730907373130322)),(to_sfixed_a(0.049622245132923126)),(to_sfixed_a(-0.00030271842842921615)),(to_sfixed_a(-0.0045157852582633495)),(to_sfixed_a(0.0009134444990195334)),(to_sfixed_a(-0.0038842891808599234)),(to_sfixed_a(-0.033985476940870285)),(to_sfixed_a(0.00011733404244296253)),(to_sfixed_a(-0.004230274818837643)),(to_sfixed_a(0.00954676978290081)),(to_sfixed_a(-0.00024554398260079324)),(to_sfixed_a(-0.29775750637054443)),(to_sfixed_a(0.00019066498498432338)),(to_sfixed_a(0.00019235454965382814)),(to_sfixed_a(-0.02167784795165062)),(to_sfixed_a(0.39405137300491333)),(to_sfixed_a(6.506333011202514e-05)),(to_sfixed_a(0.00016609836893621832)),(to_sfixed_a(0.003854539943858981)),(to_sfixed_a(8.265770156867802e-05)),(to_sfixed_a(0.058985017240047455)),(to_sfixed_a(-4.568522490444593e-05)),(to_sfixed_a(0.0002802588860504329)),(to_sfixed_a(-0.00011940315016545355)),(to_sfixed_a(0.1691126674413681)),(to_sfixed_a(-1.009533298201859e-05)),(to_sfixed_a(7.379871385637671e-05)),(to_sfixed_a(-6.525023491121829e-05)),(to_sfixed_a(0.06189161539077759)),(to_sfixed_a(0.4179679751396179)),(to_sfixed_a(2.3421798687195405e-05)),(to_sfixed_a(-0.0003157180326525122)),(to_sfixed_a(7.583475962746888e-06)),(to_sfixed_a(-0.00018515577539801598)),(to_sfixed_a(-0.0016792435199022293)),(to_sfixed_a(-0.004226052202284336)),(to_sfixed_a(0.002311921678483486)),(to_sfixed_a(-0.0015635265735909343)),(to_sfixed_a(0.0015422009164467454)),(to_sfixed_a(0.00012148384848842397)),(to_sfixed_a(-8.182003512047231e-06)),(to_sfixed_a(-4.373803676571697e-05)),(to_sfixed_a(0.005977093707770109)),(to_sfixed_a(-0.00011210267257411033)),(to_sfixed_a(7.574228220619261e-06)),(to_sfixed_a(0.00387611729092896)),(to_sfixed_a(0.001295586465857923)),(to_sfixed_a(5.939698894508183e-06)),(to_sfixed_a(-0.7230677008628845)),(to_sfixed_a(-0.00010848323290701956)),(to_sfixed_a(0.008107298985123634)),(to_sfixed_a(0.0007203692221082747)),(to_sfixed_a(-4.3500294850673527e-05)),(to_sfixed_a(-0.00046811820357106626)),(to_sfixed_a(-0.005665300879627466)),(to_sfixed_a(-0.00015179059118963778)),(to_sfixed_a(-1.0528525308473036e-05)),(to_sfixed_a(0.2854056656360626)),(to_sfixed_a(0.3930068910121918)),(to_sfixed_a(-0.021914692595601082)));

    constant weight_n2_57 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.5999822020530701)),(to_sfixed_a(0.003489825874567032)),(to_sfixed_a(-0.011854850687086582)),(to_sfixed_a(0.00015795149374753237)),(to_sfixed_a(-0.2448490858078003)),(to_sfixed_a(0.00020721078908536583)),(to_sfixed_a(0.0027183981146663427)),(to_sfixed_a(0.0001363138435408473)),(to_sfixed_a(0.00011304360668873414)),(to_sfixed_a(-0.00015205793897621334)),(to_sfixed_a(7.88498655310832e-05)),(to_sfixed_a(0.002171363215893507)),(to_sfixed_a(0.6434495449066162)),(to_sfixed_a(0.004792744759470224)),(to_sfixed_a(-0.00011414613982196897)),(to_sfixed_a(5.677336594089866e-05)),(to_sfixed_a(-0.2748972177505493)),(to_sfixed_a(0.00010590489546302706)),(to_sfixed_a(-0.22530202567577362)),(to_sfixed_a(0.22218674421310425)),(to_sfixed_a(-0.00018543584155850112)),(to_sfixed_a(6.353903154376894e-05)),(to_sfixed_a(-0.2652289867401123)),(to_sfixed_a(0.004246284253895283)),(to_sfixed_a(0.0070602488704025745)),(to_sfixed_a(-0.4218583106994629)),(to_sfixed_a(0.00020232470706105232)),(to_sfixed_a(0.0002284651855006814)),(to_sfixed_a(-0.004501113668084145)),(to_sfixed_a(3.0271883588284254e-05)),(to_sfixed_a(0.0007547001587226987)),(to_sfixed_a(-3.296589420642704e-05)),(to_sfixed_a(0.0006942905602045357)),(to_sfixed_a(-0.00011448224540799856)),(to_sfixed_a(-0.00028658195515163243)),(to_sfixed_a(-6.92267858539708e-05)),(to_sfixed_a(0.001411318895407021)),(to_sfixed_a(0.0047330730594694614)),(to_sfixed_a(0.0013382424367591739)),(to_sfixed_a(-0.00014637642016168684)),(to_sfixed_a(-0.04725959897041321)),(to_sfixed_a(0.014212590642273426)),(to_sfixed_a(-0.00020257275900803506)),(to_sfixed_a(-0.000256650906521827)),(to_sfixed_a(-0.001342406147159636)),(to_sfixed_a(-0.004366129171103239)),(to_sfixed_a(0.00034857267746701837)),(to_sfixed_a(-0.5686838626861572)),(to_sfixed_a(0.0002901041880249977)),(to_sfixed_a(0.11958303302526474)),(to_sfixed_a(-0.5409683585166931)),(to_sfixed_a(0.09741262346506119)),(to_sfixed_a(-0.00011764949886128306)),(to_sfixed_a(0.0004279840795788914)),(to_sfixed_a(0.007889258675277233)),(to_sfixed_a(-0.0024322711396962404)),(to_sfixed_a(-5.464607966132462e-07)),(to_sfixed_a(0.006661381106823683)),(to_sfixed_a(3.115608706139028e-06)),(to_sfixed_a(8.530073682777584e-05)),(to_sfixed_a(-0.0023222975432872772)),(to_sfixed_a(0.32147160172462463)),(to_sfixed_a(0.003781069302931428)),(to_sfixed_a(0.002483378630131483)),(to_sfixed_a(-0.00041799014434218407)),(to_sfixed_a(0.004316278733313084)),(to_sfixed_a(6.909741932759061e-05)),(to_sfixed_a(-0.558991551399231)),(to_sfixed_a(0.015463258139789104)),(to_sfixed_a(7.57470479584299e-05)),(to_sfixed_a(-0.1460350900888443)),(to_sfixed_a(-0.011818580329418182)),(to_sfixed_a(0.15725077688694)),(to_sfixed_a(-5.7962875871453434e-05)),(to_sfixed_a(0.00045132567174732685)),(to_sfixed_a(0.00021743786055594683)),(to_sfixed_a(0.004489127080887556)),(to_sfixed_a(-0.00391062255948782)),(to_sfixed_a(-6.0527498135343194e-05)),(to_sfixed_a(0.00016854408022481948)),(to_sfixed_a(0.001621092902496457)),(to_sfixed_a(-1.7252692487090826e-05)),(to_sfixed_a(0.0023302885238081217)),(to_sfixed_a(0.005700194276869297)),(to_sfixed_a(-0.00013658724492415786)),(to_sfixed_a(0.001180319464765489)),(to_sfixed_a(0.009312811307609081)),(to_sfixed_a(-7.706676115049049e-05)),(to_sfixed_a(2.300010237377137e-05)),(to_sfixed_a(2.295304147992283e-05)),(to_sfixed_a(0.00682409992441535)),(to_sfixed_a(0.00017262602341361344)),(to_sfixed_a(0.0004356609715614468)),(to_sfixed_a(0.00042131374357268214)),(to_sfixed_a(0.005705720279365778)),(to_sfixed_a(-2.9094899218762293e-05)),(to_sfixed_a(-0.0001149121526395902)),(to_sfixed_a(0.00041687930934131145)),(to_sfixed_a(0.0001065069081960246)),(to_sfixed_a(0.000244232447585091)),(to_sfixed_a(0.0026994459331035614)),(to_sfixed_a(0.31341752409935)),(to_sfixed_a(-3.950378595618531e-05)),(to_sfixed_a(-0.0005512955831363797)),(to_sfixed_a(0.003747569862753153)),(to_sfixed_a(-0.0002522955765016377)),(to_sfixed_a(0.0003137015155516565)),(to_sfixed_a(3.309329622425139e-05)),(to_sfixed_a(2.7792273613158613e-05)),(to_sfixed_a(0.00013834491255693138)),(to_sfixed_a(0.20883895456790924)),(to_sfixed_a(-0.00012684272951446474)),(to_sfixed_a(-0.7975652813911438)),(to_sfixed_a(2.3072119802236557e-05)),(to_sfixed_a(0.00011026275024050847)),(to_sfixed_a(0.008618823252618313)),(to_sfixed_a(0.24588324129581451)),(to_sfixed_a(0.0006957873702049255)),(to_sfixed_a(-9.078507719095796e-05)),(to_sfixed_a(0.02237575873732567)),(to_sfixed_a(5.0303795433137566e-05)),(to_sfixed_a(0.0001887841208372265)),(to_sfixed_a(-0.002434736816212535)),(to_sfixed_a(0.00012823572615161538)),(to_sfixed_a(-6.659870268777013e-05)),(to_sfixed_a(-0.2748298645019531)),(to_sfixed_a(0.00018020140123553574)),(to_sfixed_a(0.0002442648110445589)),(to_sfixed_a(-0.0002535140374675393)),(to_sfixed_a(1.4581710274796933e-05)),(to_sfixed_a(-6.274066981859505e-05)),(to_sfixed_a(0.00020758347818627954)),(to_sfixed_a(7.043882214929909e-05)),(to_sfixed_a(0.2385607361793518)),(to_sfixed_a(3.7173151213210076e-05)),(to_sfixed_a(0.00014955125516280532)),(to_sfixed_a(-0.00012504550977610052)),(to_sfixed_a(0.00010768361244117841)),(to_sfixed_a(-0.0002872769837267697)),(to_sfixed_a(-2.9872033337596804e-05)),(to_sfixed_a(-0.00355502194724977)),(to_sfixed_a(-0.00018081652524415404)),(to_sfixed_a(-4.262733273208141e-05)),(to_sfixed_a(4.073584568686783e-05)),(to_sfixed_a(0.0017271789256483316)),(to_sfixed_a(-0.00020884949481114745)),(to_sfixed_a(-0.0006666737026534975)),(to_sfixed_a(-2.070584741886705e-06)),(to_sfixed_a(-3.7650021113222465e-05)),(to_sfixed_a(0.0035103324335068464)),(to_sfixed_a(5.85465895710513e-05)),(to_sfixed_a(4.120522498851642e-05)),(to_sfixed_a(0.001822958467528224)),(to_sfixed_a(-0.00010659738472895697)),(to_sfixed_a(0.0002816463529597968)),(to_sfixed_a(0.33225512504577637)),(to_sfixed_a(-0.0001845939550548792)),(to_sfixed_a(0.37958914041519165)),(to_sfixed_a(0.0010178897064179182)),(to_sfixed_a(6.617672624997795e-05)),(to_sfixed_a(-7.660860137548298e-05)),(to_sfixed_a(-3.163859946653247e-05)),(to_sfixed_a(0.001704104244709015)),(to_sfixed_a(0.2967678904533386)),(to_sfixed_a(0.004568320699036121)),(to_sfixed_a(-0.004582920111715794)),(to_sfixed_a(-1.145264832302928e-06)),(to_sfixed_a(-0.2858983278274536)),(to_sfixed_a(0.00015075925330165774)),(to_sfixed_a(-4.969162546331063e-06)),(to_sfixed_a(0.005591315217316151)),(to_sfixed_a(0.00011927951709367335)),(to_sfixed_a(-0.0004807163786608726)),(to_sfixed_a(0.0002472737687639892)),(to_sfixed_a(-0.042254481464624405)),(to_sfixed_a(0.0003921141615137458)),(to_sfixed_a(0.007230826653540134)),(to_sfixed_a(0.0011069477768614888)),(to_sfixed_a(-0.005194749217480421)),(to_sfixed_a(0.0001333926775259897)),(to_sfixed_a(-0.00014880610979162157)),(to_sfixed_a(-0.0017263054614886642)),(to_sfixed_a(-1.1284679203527048e-05)),(to_sfixed_a(0.0002379492507316172)),(to_sfixed_a(-0.00011200044536963105)),(to_sfixed_a(0.0010854091960936785)),(to_sfixed_a(-0.265999972820282)),(to_sfixed_a(-0.0002677955199033022)),(to_sfixed_a(0.004160912707448006)),(to_sfixed_a(0.005186816677451134)),(to_sfixed_a(0.1986483335494995)),(to_sfixed_a(-3.419889253564179e-06)),(to_sfixed_a(-0.00032364617800340056)),(to_sfixed_a(0.21030941605567932)),(to_sfixed_a(-5.700226756744087e-05)),(to_sfixed_a(-0.35137858986854553)),(to_sfixed_a(-0.00011434721818659455)),(to_sfixed_a(-0.0015683415113016963)),(to_sfixed_a(0.007264238782227039)),(to_sfixed_a(0.0002303333894815296)),(to_sfixed_a(-0.00023054165649227798)),(to_sfixed_a(-1.0232797649223357e-05)),(to_sfixed_a(0.000193418629351072)),(to_sfixed_a(-6.808957550674677e-05)),(to_sfixed_a(0.00015707293641753495)),(to_sfixed_a(0.003189205192029476)),(to_sfixed_a(0.015560225583612919)),(to_sfixed_a(-0.0013135398039594293)),(to_sfixed_a(0.0017211779486387968)),(to_sfixed_a(0.0012963588815182447)),(to_sfixed_a(0.0039295325987041)),(to_sfixed_a(9.903006866807118e-05)),(to_sfixed_a(-0.00016823792248032987)),(to_sfixed_a(-0.0001005253943731077)),(to_sfixed_a(-2.9042585083516315e-05)),(to_sfixed_a(0.00024395823129452765)),(to_sfixed_a(0.005860599689185619)),(to_sfixed_a(0.003165467642247677)),(to_sfixed_a(0.47821328043937683)),(to_sfixed_a(-2.3062690161168575e-05)),(to_sfixed_a(2.6055662601720542e-05)),(to_sfixed_a(-0.00016852737462613732)),(to_sfixed_a(2.002027031267062e-06)),(to_sfixed_a(-0.00032243033638224006)),(to_sfixed_a(-0.05096219480037689)),(to_sfixed_a(0.00022744583839084953)),(to_sfixed_a(6.562324415426701e-06)),(to_sfixed_a(2.7941092412220314e-05)),(to_sfixed_a(0.3349202871322632)),(to_sfixed_a(0.0035337284207344055)),(to_sfixed_a(-0.0018631392158567905)),(to_sfixed_a(1.2345430150162429e-05)),(to_sfixed_a(-2.9859613277949393e-05)),(to_sfixed_a(0.000105326107586734)),(to_sfixed_a(0.0019244725117459893)),(to_sfixed_a(-0.0020382911898195744)),(to_sfixed_a(-0.15559230744838715)),(to_sfixed_a(3.6260546039557084e-05)),(to_sfixed_a(0.002659321529790759)),(to_sfixed_a(-5.81272215640638e-05)),(to_sfixed_a(0.015178359113633633)),(to_sfixed_a(-0.00020831817528232932)),(to_sfixed_a(0.3167724311351776)),(to_sfixed_a(0.00024803829728625715)),(to_sfixed_a(-0.26405468583106995)),(to_sfixed_a(0.005011842120438814)),(to_sfixed_a(-0.010821458883583546)),(to_sfixed_a(-0.3443559408187866)),(to_sfixed_a(-4.429678665474057e-05)),(to_sfixed_a(-6.0476784710772336e-05)),(to_sfixed_a(0.0068591502495110035)),(to_sfixed_a(9.466103074373677e-05)),(to_sfixed_a(0.1946732997894287)),(to_sfixed_a(1.8357277440372854e-05)),(to_sfixed_a(-0.0002650776004884392)),(to_sfixed_a(0.18382294476032257)),(to_sfixed_a(0.013261155225336552)),(to_sfixed_a(-0.00012838211841881275)),(to_sfixed_a(4.930492286803201e-05)),(to_sfixed_a(0.006176228169351816)),(to_sfixed_a(-0.00012683990644291043)),(to_sfixed_a(-0.00032868245034478605)),(to_sfixed_a(3.5765649954555556e-05)),(to_sfixed_a(-6.683587344014086e-06)),(to_sfixed_a(2.44125840254128e-06)),(to_sfixed_a(0.18654248118400574)),(to_sfixed_a(-6.897543789818883e-05)),(to_sfixed_a(0.000448276026872918)),(to_sfixed_a(2.4989894882310182e-05)),(to_sfixed_a(0.0024943421594798565)),(to_sfixed_a(-0.3206046223640442)),(to_sfixed_a(-0.0004109637229703367)),(to_sfixed_a(0.0001460413623135537)),(to_sfixed_a(-0.00031574463355354965)),(to_sfixed_a(6.470181688200682e-06)),(to_sfixed_a(0.00688279839232564)),(to_sfixed_a(0.009530765004456043)),(to_sfixed_a(0.0011303976643830538)),(to_sfixed_a(0.010154214687645435)),(to_sfixed_a(0.006980419158935547)),(to_sfixed_a(-0.00017599022248759866)),(to_sfixed_a(3.3630640245974064e-06)),(to_sfixed_a(-7.773296238156036e-05)),(to_sfixed_a(0.003452036762610078)),(to_sfixed_a(-6.80414741509594e-05)),(to_sfixed_a(8.65769834490493e-05)),(to_sfixed_a(0.0031903348863124847)),(to_sfixed_a(0.3773258924484253)),(to_sfixed_a(-0.00011691363761201501)),(to_sfixed_a(0.0005916432128287852)),(to_sfixed_a(0.0002447912411298603)),(to_sfixed_a(0.0034409796353429556)),(to_sfixed_a(0.006371443625539541)),(to_sfixed_a(-7.103103416739032e-05)),(to_sfixed_a(0.005142840091139078)),(to_sfixed_a(-0.009381517767906189)),(to_sfixed_a(0.0007546881679445505)),(to_sfixed_a(-6.172761641209945e-05)),(to_sfixed_a(0.4573090374469757)),(to_sfixed_a(-0.33910927176475525)),(to_sfixed_a(0.005178611259907484)));

    constant weight_n2_58 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.1754046082496643)),(to_sfixed_a(0.2729962170124054)),(to_sfixed_a(0.4129195213317871)),(to_sfixed_a(4.881851054960862e-05)),(to_sfixed_a(-0.0022533750161528587)),(to_sfixed_a(0.0002017488586716354)),(to_sfixed_a(-0.004210921004414558)),(to_sfixed_a(7.865719817345962e-05)),(to_sfixed_a(0.00023615082318428904)),(to_sfixed_a(7.166163413785398e-07)),(to_sfixed_a(-0.000119723379611969)),(to_sfixed_a(-0.008339956402778625)),(to_sfixed_a(0.003778050886467099)),(to_sfixed_a(0.00210491381585598)),(to_sfixed_a(7.083290256559849e-06)),(to_sfixed_a(-1.341786264674738e-05)),(to_sfixed_a(0.00967569462954998)),(to_sfixed_a(0.00011507173621794209)),(to_sfixed_a(0.004093446768820286)),(to_sfixed_a(0.0005084395525045693)),(to_sfixed_a(-0.00019693411013577133)),(to_sfixed_a(6.774781650165096e-05)),(to_sfixed_a(5.3027757530799136e-05)),(to_sfixed_a(0.004544689320027828)),(to_sfixed_a(0.005027380306273699)),(to_sfixed_a(0.0022495929151773453)),(to_sfixed_a(-3.576768722268753e-05)),(to_sfixed_a(-0.00010177730291616172)),(to_sfixed_a(-0.0005873679765500128)),(to_sfixed_a(1.0097955964738503e-06)),(to_sfixed_a(0.0015947401989251375)),(to_sfixed_a(-0.00010257153917336836)),(to_sfixed_a(0.0008828573627397418)),(to_sfixed_a(5.236714787315577e-05)),(to_sfixed_a(0.00012026139302179217)),(to_sfixed_a(-1.1781827197410166e-05)),(to_sfixed_a(0.007329908665269613)),(to_sfixed_a(-0.3278384208679199)),(to_sfixed_a(0.34471654891967773)),(to_sfixed_a(8.573185914428905e-05)),(to_sfixed_a(0.001552952453494072)),(to_sfixed_a(0.008813127875328064)),(to_sfixed_a(-2.9546003133873455e-05)),(to_sfixed_a(-0.0003741226391866803)),(to_sfixed_a(0.002780541777610779)),(to_sfixed_a(-0.0015766951255500317)),(to_sfixed_a(0.0005265463260002434)),(to_sfixed_a(-0.4883679151535034)),(to_sfixed_a(-1.1899886885657907e-05)),(to_sfixed_a(-0.014244724996387959)),(to_sfixed_a(-0.18539974093437195)),(to_sfixed_a(-0.0002740072086453438)),(to_sfixed_a(0.0003815765376202762)),(to_sfixed_a(0.0016764055471867323)),(to_sfixed_a(0.0006214859313331544)),(to_sfixed_a(0.07495802640914917)),(to_sfixed_a(0.00010805323836393654)),(to_sfixed_a(-0.011996733956038952)),(to_sfixed_a(-0.000232475736993365)),(to_sfixed_a(-1.6739795682951808e-05)),(to_sfixed_a(0.3117958605289459)),(to_sfixed_a(0.0016745670000091195)),(to_sfixed_a(8.390909351874143e-05)),(to_sfixed_a(0.011793486773967743)),(to_sfixed_a(-0.00010433950228616595)),(to_sfixed_a(0.17619982361793518)),(to_sfixed_a(0.00015035642718430609)),(to_sfixed_a(-0.30011874437332153)),(to_sfixed_a(-0.01171645987778902)),(to_sfixed_a(7.083329546730965e-05)),(to_sfixed_a(-0.006300320848822594)),(to_sfixed_a(-0.2199126034975052)),(to_sfixed_a(-0.02889963798224926)),(to_sfixed_a(0.0001556088827783242)),(to_sfixed_a(0.0003907921491190791)),(to_sfixed_a(-0.00011663060286082327)),(to_sfixed_a(-0.006172239314764738)),(to_sfixed_a(-0.15261822938919067)),(to_sfixed_a(-6.285133713390678e-05)),(to_sfixed_a(0.40687742829322815)),(to_sfixed_a(0.001298209186643362)),(to_sfixed_a(-4.9621405196376145e-05)),(to_sfixed_a(-0.0010559128131717443)),(to_sfixed_a(0.006506412290036678)),(to_sfixed_a(6.588226824533194e-06)),(to_sfixed_a(-0.3412136137485504)),(to_sfixed_a(0.0017446399433538318)),(to_sfixed_a(0.003631536616012454)),(to_sfixed_a(9.037675044964999e-05)),(to_sfixed_a(-0.00045143882744014263)),(to_sfixed_a(-0.0011259055463597178)),(to_sfixed_a(0.00015467000775970519)),(to_sfixed_a(-0.0030156681314110756)),(to_sfixed_a(2.2512071154778823e-05)),(to_sfixed_a(-0.004947743844240904)),(to_sfixed_a(0.00019867157971020788)),(to_sfixed_a(6.655769539065659e-05)),(to_sfixed_a(5.433757905848324e-06)),(to_sfixed_a(-3.1005460186861455e-05)),(to_sfixed_a(-0.0004495936445891857)),(to_sfixed_a(-0.5358709692955017)),(to_sfixed_a(0.0033219659235328436)),(to_sfixed_a(-6.878840213175863e-05)),(to_sfixed_a(0.01325293816626072)),(to_sfixed_a(0.15772461891174316)),(to_sfixed_a(0.0011082231067121029)),(to_sfixed_a(0.00022926318342797458)),(to_sfixed_a(-4.520497168414295e-05)),(to_sfixed_a(0.00010130461305379868)),(to_sfixed_a(0.012901552952826023)),(to_sfixed_a(-0.004295011050999165)),(to_sfixed_a(7.000282494118437e-05)),(to_sfixed_a(-0.0104218116030097)),(to_sfixed_a(-4.8325920943170786e-05)),(to_sfixed_a(-2.6633748348103836e-05)),(to_sfixed_a(-0.013569924049079418)),(to_sfixed_a(0.001985240960493684)),(to_sfixed_a(0.05874330550432205)),(to_sfixed_a(0.00014030672900844365)),(to_sfixed_a(-0.023961611092090607)),(to_sfixed_a(3.0368166335392743e-05)),(to_sfixed_a(3.0314564355649054e-05)),(to_sfixed_a(-0.014817122370004654)),(to_sfixed_a(-5.727593816118315e-05)),(to_sfixed_a(1.8232851289212704e-05)),(to_sfixed_a(0.002292126417160034)),(to_sfixed_a(-0.0015929697547107935)),(to_sfixed_a(0.00011814595927717164)),(to_sfixed_a(-0.00017568981274962425)),(to_sfixed_a(2.805798430927098e-06)),(to_sfixed_a(7.747279596515e-05)),(to_sfixed_a(-0.00011184746108483523)),(to_sfixed_a(0.0031850398518145084)),(to_sfixed_a(0.0029474031180143356)),(to_sfixed_a(0.00014905542775522918)),(to_sfixed_a(3.1449817470274866e-06)),(to_sfixed_a(-0.020244725048542023)),(to_sfixed_a(-0.00014373396697919816)),(to_sfixed_a(-6.86848652549088e-05)),(to_sfixed_a(0.00017373998707626015)),(to_sfixed_a(0.0029347592499107122)),(to_sfixed_a(0.00028736505191773176)),(to_sfixed_a(0.0002369616850046441)),(to_sfixed_a(-5.408970173448324e-05)),(to_sfixed_a(0.003055629087612033)),(to_sfixed_a(0.0006673862226307392)),(to_sfixed_a(-0.00553093571215868)),(to_sfixed_a(0.00017669133376330137)),(to_sfixed_a(0.00028246582951396704)),(to_sfixed_a(-0.0037886754143983126)),(to_sfixed_a(0.00019586477719713002)),(to_sfixed_a(0.00010211909102508798)),(to_sfixed_a(0.0010684425942599773)),(to_sfixed_a(7.966329576447606e-06)),(to_sfixed_a(5.857429641764611e-05)),(to_sfixed_a(0.008819449692964554)),(to_sfixed_a(3.5056000342592597e-06)),(to_sfixed_a(0.0036263691727072)),(to_sfixed_a(0.00010237906099064276)),(to_sfixed_a(-6.916929851286113e-05)),(to_sfixed_a(0.00018654789892025292)),(to_sfixed_a(7.70074111642316e-05)),(to_sfixed_a(-0.1989680677652359)),(to_sfixed_a(0.0027503317687660456)),(to_sfixed_a(0.007294125389307737)),(to_sfixed_a(0.009734703227877617)),(to_sfixed_a(5.7963239669334143e-05)),(to_sfixed_a(-0.005333642940968275)),(to_sfixed_a(0.00015359917597379535)),(to_sfixed_a(6.135564763098955e-05)),(to_sfixed_a(-0.027075989171862602)),(to_sfixed_a(0.001703679678030312)),(to_sfixed_a(0.004822855815291405)),(to_sfixed_a(5.0455018936190754e-05)),(to_sfixed_a(-0.005050355568528175)),(to_sfixed_a(0.0011441413080319762)),(to_sfixed_a(0.004213347565382719)),(to_sfixed_a(0.0016028555110096931)),(to_sfixed_a(0.3396948277950287)),(to_sfixed_a(-0.295746773481369)),(to_sfixed_a(-0.00022255536168813705)),(to_sfixed_a(8.737068128539249e-05)),(to_sfixed_a(0.00017650514200795442)),(to_sfixed_a(-0.0001898160990094766)),(to_sfixed_a(0.0001503660751041025)),(to_sfixed_a(-0.022175312042236328)),(to_sfixed_a(0.006137832999229431)),(to_sfixed_a(-0.002112775109708309)),(to_sfixed_a(0.001232309266924858)),(to_sfixed_a(7.733928214292973e-06)),(to_sfixed_a(0.006120261270552874)),(to_sfixed_a(-0.00019940256606787443)),(to_sfixed_a(-0.021875504404306412)),(to_sfixed_a(0.000877028563991189)),(to_sfixed_a(0.0001748425856931135)),(to_sfixed_a(-0.355633944272995)),(to_sfixed_a(-0.00011327808169880882)),(to_sfixed_a(0.004651596304029226)),(to_sfixed_a(0.7523541450500488)),(to_sfixed_a(-0.00013985713303554803)),(to_sfixed_a(2.3771863197907805e-06)),(to_sfixed_a(-1.2536256690509617e-06)),(to_sfixed_a(2.922771091107279e-05)),(to_sfixed_a(0.00023780157789587975)),(to_sfixed_a(0.00017170263163279742)),(to_sfixed_a(0.04934612661600113)),(to_sfixed_a(0.424211710691452)),(to_sfixed_a(0.3401870131492615)),(to_sfixed_a(0.2467341274023056)),(to_sfixed_a(0.17347505688667297)),(to_sfixed_a(-0.009861948899924755)),(to_sfixed_a(-7.794206612743437e-05)),(to_sfixed_a(-6.16660836385563e-05)),(to_sfixed_a(-2.406968269497156e-05)),(to_sfixed_a(7.69498510635458e-05)),(to_sfixed_a(-2.1881351131014526e-05)),(to_sfixed_a(-0.0030618684832006693)),(to_sfixed_a(0.0025483884382992983)),(to_sfixed_a(-0.007358202710747719)),(to_sfixed_a(7.681830174988136e-05)),(to_sfixed_a(2.7206602680962533e-05)),(to_sfixed_a(3.7583758967230096e-05)),(to_sfixed_a(-0.00010468839172972366)),(to_sfixed_a(0.00040401567821390927)),(to_sfixed_a(-0.0035960872191935778)),(to_sfixed_a(0.0002268899988848716)),(to_sfixed_a(-0.0002111121139023453)),(to_sfixed_a(0.00015761156100779772)),(to_sfixed_a(-0.0008784877136349678)),(to_sfixed_a(-0.01017099991440773)),(to_sfixed_a(-0.0005750394193455577)),(to_sfixed_a(-0.00012102589244022965)),(to_sfixed_a(-0.00028968683909624815)),(to_sfixed_a(-1.546118437545374e-05)),(to_sfixed_a(0.00834114383906126)),(to_sfixed_a(-0.011643868871033192)),(to_sfixed_a(0.23382675647735596)),(to_sfixed_a(-1.9471364794299006e-05)),(to_sfixed_a(-0.00016419099119957536)),(to_sfixed_a(9.430765203433111e-05)),(to_sfixed_a(-0.038545794785022736)),(to_sfixed_a(-0.0004129577719140798)),(to_sfixed_a(-0.03623685613274574)),(to_sfixed_a(-0.0001124707268900238)),(to_sfixed_a(-0.011277205310761929)),(to_sfixed_a(0.578146755695343)),(to_sfixed_a(0.007044672500342131)),(to_sfixed_a(0.14732244610786438)),(to_sfixed_a(1.0848936653928831e-05)),(to_sfixed_a(0.009147655218839645)),(to_sfixed_a(3.701238892972469e-05)),(to_sfixed_a(0.0002923869760707021)),(to_sfixed_a(0.0003150062693748623)),(to_sfixed_a(3.8578578823944554e-05)),(to_sfixed_a(-0.00011018490476999432)),(to_sfixed_a(-0.004418481141328812)),(to_sfixed_a(0.0048764050006866455)),(to_sfixed_a(6.794823275413364e-05)),(to_sfixed_a(-6.501466123154387e-05)),(to_sfixed_a(-0.1450587958097458)),(to_sfixed_a(0.0002790131256915629)),(to_sfixed_a(0.002445196034386754)),(to_sfixed_a(3.548167660483159e-05)),(to_sfixed_a(-0.0007507882546633482)),(to_sfixed_a(5.849760782439262e-05)),(to_sfixed_a(-0.035179171711206436)),(to_sfixed_a(-0.00020957767264917493)),(to_sfixed_a(7.475713937310502e-05)),(to_sfixed_a(0.00014607921184506267)),(to_sfixed_a(-0.000796228414401412)),(to_sfixed_a(-0.0044915927574038506)),(to_sfixed_a(1.7407852283213288e-05)),(to_sfixed_a(4.308909410610795e-06)),(to_sfixed_a(-3.363615178386681e-05)),(to_sfixed_a(3.285077400505543e-05)),(to_sfixed_a(-0.003200670937076211)),(to_sfixed_a(-0.0033400109969079494)),(to_sfixed_a(0.0024884610902518034)),(to_sfixed_a(0.3316771984100342)),(to_sfixed_a(0.2291480451822281)),(to_sfixed_a(3.996511804871261e-05)),(to_sfixed_a(-9.792856872081757e-05)),(to_sfixed_a(-6.980611942708492e-06)),(to_sfixed_a(-0.0002331181603949517)),(to_sfixed_a(0.00017506879521533847)),(to_sfixed_a(-7.142681715777144e-05)),(to_sfixed_a(0.0035557798109948635)),(to_sfixed_a(0.19634020328521729)),(to_sfixed_a(-0.00011442681716289371)),(to_sfixed_a(-0.00012974292621947825)),(to_sfixed_a(-0.0006543839117512107)),(to_sfixed_a(0.0038451075088232756)),(to_sfixed_a(0.14454534649848938)),(to_sfixed_a(-0.0001521065569249913)),(to_sfixed_a(-0.0032878092024475336)),(to_sfixed_a(-0.00224681687541306)),(to_sfixed_a(0.0013589265290647745)),(to_sfixed_a(7.874046423239633e-05)),(to_sfixed_a(-0.011809875257313251)),(to_sfixed_a(0.002477199537679553)),(to_sfixed_a(0.009882848709821701)));

    constant weight_n2_59 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.5780751705169678)),(to_sfixed_a(-0.0028316830284893513)),(to_sfixed_a(-0.35774853825569153)),(to_sfixed_a(-0.0002549403579905629)),(to_sfixed_a(-0.0038921525701880455)),(to_sfixed_a(1.3226126611698419e-05)),(to_sfixed_a(-0.0041079348884522915)),(to_sfixed_a(-0.00013754602696280926)),(to_sfixed_a(-8.264385542133823e-05)),(to_sfixed_a(4.452889697859064e-06)),(to_sfixed_a(-2.509209662093781e-05)),(to_sfixed_a(0.27895236015319824)),(to_sfixed_a(-0.012508331798017025)),(to_sfixed_a(0.28850629925727844)),(to_sfixed_a(-2.7632755518425256e-05)),(to_sfixed_a(0.0001788645749911666)),(to_sfixed_a(-0.12509246170520782)),(to_sfixed_a(0.00015528875519521534)),(to_sfixed_a(0.03754829242825508)),(to_sfixed_a(0.41144171357154846)),(to_sfixed_a(-0.00011269368405919522)),(to_sfixed_a(3.856948751490563e-06)),(to_sfixed_a(-0.0008652860415168107)),(to_sfixed_a(-0.0006229126593098044)),(to_sfixed_a(-0.006064211018383503)),(to_sfixed_a(-0.04844273254275322)),(to_sfixed_a(-2.0458510334719904e-05)),(to_sfixed_a(-0.0026152587961405516)),(to_sfixed_a(-0.005033798050135374)),(to_sfixed_a(-0.00015203229850158095)),(to_sfixed_a(-0.35080620646476746)),(to_sfixed_a(-6.254900654312223e-05)),(to_sfixed_a(-0.007128213066607714)),(to_sfixed_a(0.0001366143551422283)),(to_sfixed_a(-0.00012887318735010922)),(to_sfixed_a(0.00018043143791146576)),(to_sfixed_a(-0.08758246898651123)),(to_sfixed_a(0.016306664794683456)),(to_sfixed_a(0.0048318603076040745)),(to_sfixed_a(-8.411513408645988e-05)),(to_sfixed_a(0.004254782106727362)),(to_sfixed_a(0.004533151630312204)),(to_sfixed_a(0.0001131238677771762)),(to_sfixed_a(-6.408955960068852e-05)),(to_sfixed_a(-0.002043691463768482)),(to_sfixed_a(-0.3311269283294678)),(to_sfixed_a(-0.478998601436615)),(to_sfixed_a(-0.20976820588111877)),(to_sfixed_a(-0.00017728506645653397)),(to_sfixed_a(-0.000221485854126513)),(to_sfixed_a(-0.30358898639678955)),(to_sfixed_a(-0.0005897365626879036)),(to_sfixed_a(7.181008550105616e-05)),(to_sfixed_a(-0.00027180055622011423)),(to_sfixed_a(0.0012567879166454077)),(to_sfixed_a(-0.00711028603836894)),(to_sfixed_a(-0.000251743127591908)),(to_sfixed_a(0.016273144632577896)),(to_sfixed_a(-0.0001338272704742849)),(to_sfixed_a(-3.071907121920958e-05)),(to_sfixed_a(-0.0033287652768194675)),(to_sfixed_a(-0.0010011165868490934)),(to_sfixed_a(-0.0018192180432379246)),(to_sfixed_a(-0.0067109474912285805)),(to_sfixed_a(-6.396885146386921e-05)),(to_sfixed_a(2.6400746719446033e-05)),(to_sfixed_a(-0.00017611245857551694)),(to_sfixed_a(0.0004420778714120388)),(to_sfixed_a(-0.012763210572302341)),(to_sfixed_a(0.00011458187509560958)),(to_sfixed_a(-0.4870827794075012)),(to_sfixed_a(-0.3455829620361328)),(to_sfixed_a(-0.005499391350895166)),(to_sfixed_a(-5.61405613552779e-06)),(to_sfixed_a(-0.0001198167447000742)),(to_sfixed_a(9.894742106553167e-06)),(to_sfixed_a(-0.006598434876650572)),(to_sfixed_a(0.20677240192890167)),(to_sfixed_a(-4.009837721241638e-05)),(to_sfixed_a(-0.013306884095072746)),(to_sfixed_a(-0.0008814245229586959)),(to_sfixed_a(0.00011388817802071571)),(to_sfixed_a(-0.3890460133552551)),(to_sfixed_a(0.00025827856734395027)),(to_sfixed_a(2.0139857952017337e-05)),(to_sfixed_a(-0.26625657081604004)),(to_sfixed_a(-0.24685506522655487)),(to_sfixed_a(0.0006086267530918121)),(to_sfixed_a(-0.00027447205502539873)),(to_sfixed_a(2.978300108225085e-05)),(to_sfixed_a(-0.013019280508160591)),(to_sfixed_a(-5.662645708071068e-05)),(to_sfixed_a(-0.009616143070161343)),(to_sfixed_a(-9.929168300004676e-06)),(to_sfixed_a(0.0014171460643410683)),(to_sfixed_a(-4.1415871237404644e-05)),(to_sfixed_a(-0.00039300130447372794)),(to_sfixed_a(0.000290074065560475)),(to_sfixed_a(-0.00011983918375335634)),(to_sfixed_a(7.095497858244926e-05)),(to_sfixed_a(0.0009918429423123598)),(to_sfixed_a(-0.004978414159268141)),(to_sfixed_a(0.00015571006224490702)),(to_sfixed_a(0.2453383505344391)),(to_sfixed_a(-0.029190458357334137)),(to_sfixed_a(0.0008859592489898205)),(to_sfixed_a(0.000166371013619937)),(to_sfixed_a(-1.9934559531975538e-06)),(to_sfixed_a(-1.2464111932786182e-05)),(to_sfixed_a(-0.020767558366060257)),(to_sfixed_a(-0.00809774361550808)),(to_sfixed_a(0.00011228995572309941)),(to_sfixed_a(-0.2986426055431366)),(to_sfixed_a(-7.758937135804445e-05)),(to_sfixed_a(-0.00015039625577628613)),(to_sfixed_a(0.2503081262111664)),(to_sfixed_a(0.00041664947639219463)),(to_sfixed_a(-0.0005135885439813137)),(to_sfixed_a(0.0002076706732623279)),(to_sfixed_a(-0.24924317002296448)),(to_sfixed_a(-0.0003153050201945007)),(to_sfixed_a(0.00015330237511079758)),(to_sfixed_a(-0.0032955666538327932)),(to_sfixed_a(-0.00015028778580017388)),(to_sfixed_a(9.395467350259423e-05)),(to_sfixed_a(-6.106960063334554e-05)),(to_sfixed_a(-0.011900094337761402)),(to_sfixed_a(0.00018068419012706727)),(to_sfixed_a(-0.00010663162538548931)),(to_sfixed_a(0.00011858012294396758)),(to_sfixed_a(0.00012854972737841308)),(to_sfixed_a(-9.28579320316203e-05)),(to_sfixed_a(-0.31245237588882446)),(to_sfixed_a(-0.0006630672723986208)),(to_sfixed_a(0.00026544867432676256)),(to_sfixed_a(-0.00017654962721280754)),(to_sfixed_a(0.3140972852706909)),(to_sfixed_a(0.0015457989647984505)),(to_sfixed_a(-5.44582144357264e-06)),(to_sfixed_a(-0.0001079833455150947)),(to_sfixed_a(-0.00042987370397895575)),(to_sfixed_a(-0.00017830524302553385)),(to_sfixed_a(-9.874792158370838e-05)),(to_sfixed_a(0.00011532795906532556)),(to_sfixed_a(0.002182456897571683)),(to_sfixed_a(0.0003901589661836624)),(to_sfixed_a(-0.0013555039186030626)),(to_sfixed_a(-2.370115544181317e-05)),(to_sfixed_a(0.00038081983802840114)),(to_sfixed_a(0.0007314802496694028)),(to_sfixed_a(0.00010363315959693864)),(to_sfixed_a(-0.00039234530413523316)),(to_sfixed_a(-0.22332081198692322)),(to_sfixed_a(2.028832386713475e-05)),(to_sfixed_a(-2.843209949787706e-05)),(to_sfixed_a(0.0012175862211734056)),(to_sfixed_a(-0.00011345982784405351)),(to_sfixed_a(0.0005726132076233625)),(to_sfixed_a(6.2958897615317255e-06)),(to_sfixed_a(-3.046446363441646e-05)),(to_sfixed_a(-0.00011296285811113194)),(to_sfixed_a(-0.00024032809596974403)),(to_sfixed_a(-0.013166360557079315)),(to_sfixed_a(-0.000829123193398118)),(to_sfixed_a(-0.006261677946895361)),(to_sfixed_a(-0.0007648610044270754)),(to_sfixed_a(7.592898327857256e-07)),(to_sfixed_a(-0.0040346370078623295)),(to_sfixed_a(-3.6014491342939436e-05)),(to_sfixed_a(0.00026879680808633566)),(to_sfixed_a(-0.005367862526327372)),(to_sfixed_a(-0.0005303632351569831)),(to_sfixed_a(-0.008030645549297333)),(to_sfixed_a(-0.00011684249329846352)),(to_sfixed_a(0.30042845010757446)),(to_sfixed_a(-0.01170805748552084)),(to_sfixed_a(0.011292416602373123)),(to_sfixed_a(-0.018051812425255775)),(to_sfixed_a(0.0009242842788808048)),(to_sfixed_a(-0.18200050294399261)),(to_sfixed_a(-4.221560084261e-05)),(to_sfixed_a(-0.05306749418377876)),(to_sfixed_a(-4.376521974336356e-05)),(to_sfixed_a(-0.000249565695412457)),(to_sfixed_a(-0.00014883601397741586)),(to_sfixed_a(0.003226709086447954)),(to_sfixed_a(-0.03614204004406929)),(to_sfixed_a(-0.001914576510898769)),(to_sfixed_a(-0.0007016086019575596)),(to_sfixed_a(-0.0002922046696767211)),(to_sfixed_a(0.007821298204362392)),(to_sfixed_a(3.6676370655186474e-05)),(to_sfixed_a(-0.0020708038937300444)),(to_sfixed_a(-0.007187687326222658)),(to_sfixed_a(1.3417520676739514e-05)),(to_sfixed_a(-0.34654542803764343)),(to_sfixed_a(-0.00016278168186545372)),(to_sfixed_a(-0.02343306690454483)),(to_sfixed_a(0.6103612780570984)),(to_sfixed_a(3.586805541999638e-05)),(to_sfixed_a(-0.0002038459206232801)),(to_sfixed_a(-0.00015999538300093263)),(to_sfixed_a(1.3759010471403599e-05)),(to_sfixed_a(-6.64290419081226e-05)),(to_sfixed_a(0.00044686681940220296)),(to_sfixed_a(-0.00016270876221824437)),(to_sfixed_a(-0.332421213388443)),(to_sfixed_a(0.14022456109523773)),(to_sfixed_a(-0.021712714806199074)),(to_sfixed_a(0.0003064348711632192)),(to_sfixed_a(-0.00719647528603673)),(to_sfixed_a(-0.00022787446505390108)),(to_sfixed_a(0.000227299562538974)),(to_sfixed_a(0.00010758449207060039)),(to_sfixed_a(-3.696065687108785e-05)),(to_sfixed_a(-0.00015784241259098053)),(to_sfixed_a(-0.00014021116658113897)),(to_sfixed_a(0.5049706697463989)),(to_sfixed_a(-0.03166789561510086)),(to_sfixed_a(1.6853678971529007e-05)),(to_sfixed_a(-0.00010826317884493619)),(to_sfixed_a(-7.233220094349235e-05)),(to_sfixed_a(-7.4782437877729535e-06)),(to_sfixed_a(-0.004140161909162998)),(to_sfixed_a(-0.3906072974205017)),(to_sfixed_a(0.00016853261331561953)),(to_sfixed_a(0.00018225697567686439)),(to_sfixed_a(0.00015298623475246131)),(to_sfixed_a(-0.001886762329377234)),(to_sfixed_a(-0.00594426179304719)),(to_sfixed_a(-0.0010596744250506163)),(to_sfixed_a(0.00015506776981055737)),(to_sfixed_a(-3.386956814210862e-05)),(to_sfixed_a(2.027896698564291e-06)),(to_sfixed_a(-4.977284697815776e-05)),(to_sfixed_a(-0.0005311517743393779)),(to_sfixed_a(-0.017871828749775887)),(to_sfixed_a(8.192399400286376e-05)),(to_sfixed_a(4.528992576524615e-06)),(to_sfixed_a(-0.00018263846868649125)),(to_sfixed_a(-0.01583794318139553)),(to_sfixed_a(-0.00030561169842258096)),(to_sfixed_a(-0.0017578863771632314)),(to_sfixed_a(-0.00018827622989192605)),(to_sfixed_a(0.28387191891670227)),(to_sfixed_a(0.18463671207427979)),(to_sfixed_a(-0.014502786099910736)),(to_sfixed_a(-0.003491521580144763)),(to_sfixed_a(-0.0001691614743322134)),(to_sfixed_a(-0.0008978242985904217)),(to_sfixed_a(0.0019322169246152043)),(to_sfixed_a(-1.5197121683740988e-05)),(to_sfixed_a(-0.0027796670328825712)),(to_sfixed_a(0.00016681791748851538)),(to_sfixed_a(0.19797088205814362)),(to_sfixed_a(-0.027025045827031136)),(to_sfixed_a(0.012616906315088272)),(to_sfixed_a(-3.4392738598398864e-05)),(to_sfixed_a(0.00011000838276231661)),(to_sfixed_a(-0.002165663754567504)),(to_sfixed_a(-0.00013073479931335896)),(to_sfixed_a(0.36477771401405334)),(to_sfixed_a(8.322412031702697e-05)),(to_sfixed_a(-0.0008191175875253975)),(to_sfixed_a(0.00019980358774773777)),(to_sfixed_a(0.3353286385536194)),(to_sfixed_a(-2.8222581022419035e-05)),(to_sfixed_a(0.0001005678714136593)),(to_sfixed_a(-0.0001892993168439716)),(to_sfixed_a(0.36625272035598755)),(to_sfixed_a(-0.016768744215369225)),(to_sfixed_a(-0.00015507689386140555)),(to_sfixed_a(-0.0001347503566648811)),(to_sfixed_a(2.899768151110038e-05)),(to_sfixed_a(0.00010222555283689871)),(to_sfixed_a(-0.004954069387167692)),(to_sfixed_a(-0.0018847477622330189)),(to_sfixed_a(-0.0034945597872138023)),(to_sfixed_a(-0.03139685466885567)),(to_sfixed_a(-0.0017075322102755308)),(to_sfixed_a(0.00024945917539298534)),(to_sfixed_a(2.6922236429527402e-05)),(to_sfixed_a(6.431427755160257e-05)),(to_sfixed_a(0.008486342616379261)),(to_sfixed_a(-0.00010699634003685787)),(to_sfixed_a(6.12284493399784e-05)),(to_sfixed_a(0.004912794101983309)),(to_sfixed_a(-0.017528381198644638)),(to_sfixed_a(0.0001684495946392417)),(to_sfixed_a(-0.5816711187362671)),(to_sfixed_a(-0.0013356955023482442)),(to_sfixed_a(-0.012943804264068604)),(to_sfixed_a(0.15868757665157318)),(to_sfixed_a(-0.0001901494397316128)),(to_sfixed_a(0.1407289206981659)),(to_sfixed_a(-0.35395386815071106)),(to_sfixed_a(-0.0014203771715983748)),(to_sfixed_a(2.3683638573857024e-05)),(to_sfixed_a(-0.0034006324131041765)),(to_sfixed_a(-0.12147318571805954)),(to_sfixed_a(-0.008407779037952423)));

    constant weight_n2_60 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.13745366036891937)),(to_sfixed_a(-0.0016003098571673036)),(to_sfixed_a(-7.405151700368151e-05)),(to_sfixed_a(0.0001048251724569127)),(to_sfixed_a(0.0008823599200695753)),(to_sfixed_a(2.1691776055376977e-05)),(to_sfixed_a(0.01737716607749462)),(to_sfixed_a(-0.000207807999686338)),(to_sfixed_a(-1.5369732864201069e-06)),(to_sfixed_a(-0.00015454410458914936)),(to_sfixed_a(-4.4400017941370606e-05)),(to_sfixed_a(0.006219056900590658)),(to_sfixed_a(-0.001217240933328867)),(to_sfixed_a(-0.0026802904903888702)),(to_sfixed_a(-7.117990026017651e-05)),(to_sfixed_a(0.00029715962591581047)),(to_sfixed_a(0.008089917711913586)),(to_sfixed_a(-0.00013635613140650094)),(to_sfixed_a(-0.00362946349196136)),(to_sfixed_a(-0.00031002104515209794)),(to_sfixed_a(-0.0001530332228867337)),(to_sfixed_a(0.0004489057173486799)),(to_sfixed_a(0.002750806510448456)),(to_sfixed_a(-0.00026993604842573404)),(to_sfixed_a(0.014756325632333755)),(to_sfixed_a(-0.00022816486307419837)),(to_sfixed_a(-8.385948603972793e-05)),(to_sfixed_a(2.6039422664325684e-05)),(to_sfixed_a(-7.454799197148532e-05)),(to_sfixed_a(7.142445974750444e-05)),(to_sfixed_a(0.00533241406083107)),(to_sfixed_a(-6.006962212268263e-05)),(to_sfixed_a(0.006528765428811312)),(to_sfixed_a(1.801966573111713e-05)),(to_sfixed_a(-3.1029027013573796e-05)),(to_sfixed_a(5.40572582394816e-05)),(to_sfixed_a(-0.09788871556520462)),(to_sfixed_a(4.695986717706546e-05)),(to_sfixed_a(0.005058815702795982)),(to_sfixed_a(-3.248816938139498e-05)),(to_sfixed_a(0.013907663524150848)),(to_sfixed_a(-0.011939351446926594)),(to_sfixed_a(1.2124812201363966e-05)),(to_sfixed_a(-9.42931801546365e-05)),(to_sfixed_a(0.41771695017814636)),(to_sfixed_a(0.015717584639787674)),(to_sfixed_a(-0.0011807238915935159)),(to_sfixed_a(0.0002467166632413864)),(to_sfixed_a(0.00011530503979884088)),(to_sfixed_a(-8.760357741266489e-05)),(to_sfixed_a(0.003108266042545438)),(to_sfixed_a(0.0003154864825773984)),(to_sfixed_a(0.00029172273934818804)),(to_sfixed_a(-0.0008749798289500177)),(to_sfixed_a(0.03776738420128822)),(to_sfixed_a(0.21702785789966583)),(to_sfixed_a(-0.00019999899086542428)),(to_sfixed_a(0.020098760724067688)),(to_sfixed_a(3.1094925361685455e-05)),(to_sfixed_a(5.647664511343464e-05)),(to_sfixed_a(0.007768030744045973)),(to_sfixed_a(0.0059631322510540485)),(to_sfixed_a(-0.0012563277268782258)),(to_sfixed_a(-0.26948148012161255)),(to_sfixed_a(6.949857925064862e-05)),(to_sfixed_a(0.0014913579216226935)),(to_sfixed_a(-9.185952512780204e-05)),(to_sfixed_a(0.0001530604058643803)),(to_sfixed_a(0.021781668066978455)),(to_sfixed_a(0.0001908741978695616)),(to_sfixed_a(0.01787230186164379)),(to_sfixed_a(0.0013670905027538538)),(to_sfixed_a(0.0011127210455015302)),(to_sfixed_a(5.81460990360938e-05)),(to_sfixed_a(-7.134658517315984e-06)),(to_sfixed_a(7.155149069149047e-05)),(to_sfixed_a(0.3441690504550934)),(to_sfixed_a(-0.39119821786880493)),(to_sfixed_a(0.00011389315477572381)),(to_sfixed_a(0.3047318160533905)),(to_sfixed_a(0.010303240269422531)),(to_sfixed_a(1.493631862103939e-05)),(to_sfixed_a(-0.0015290938317775726)),(to_sfixed_a(2.160969415854197e-05)),(to_sfixed_a(-5.7209319493267685e-05)),(to_sfixed_a(0.008506587706506252)),(to_sfixed_a(-0.010982608422636986)),(to_sfixed_a(0.00010678725084289908)),(to_sfixed_a(7.263523002620786e-05)),(to_sfixed_a(-7.41111216484569e-05)),(to_sfixed_a(0.43935659527778625)),(to_sfixed_a(-0.00010365515481680632)),(to_sfixed_a(0.0154643589630723)),(to_sfixed_a(0.00011294118303339928)),(to_sfixed_a(0.00654170848429203)),(to_sfixed_a(-0.00015978349256329238)),(to_sfixed_a(-5.787326517747715e-05)),(to_sfixed_a(-7.090527651598677e-05)),(to_sfixed_a(-3.727236980921589e-05)),(to_sfixed_a(5.8297664509154856e-05)),(to_sfixed_a(0.0003047374193556607)),(to_sfixed_a(0.0048958128318190575)),(to_sfixed_a(5.672918632626534e-07)),(to_sfixed_a(-0.39812663197517395)),(to_sfixed_a(0.01122598722577095)),(to_sfixed_a(0.000999918789602816)),(to_sfixed_a(0.00010442910570418462)),(to_sfixed_a(6.327325536403805e-05)),(to_sfixed_a(2.6874236937146634e-05)),(to_sfixed_a(0.011346963234245777)),(to_sfixed_a(-0.25672900676727295)),(to_sfixed_a(-0.00014893378829583526)),(to_sfixed_a(-0.0005738551844842732)),(to_sfixed_a(-6.987839879002422e-05)),(to_sfixed_a(0.00010208362073171884)),(to_sfixed_a(-0.7474120259284973)),(to_sfixed_a(2.5875517167150974e-05)),(to_sfixed_a(0.011584097519516945)),(to_sfixed_a(2.7279238565824926e-05)),(to_sfixed_a(-0.0003757532685995102)),(to_sfixed_a(-6.342124834191054e-05)),(to_sfixed_a(-0.0001118493964895606)),(to_sfixed_a(0.006318606436252594)),(to_sfixed_a(3.2788258977234364e-05)),(to_sfixed_a(-0.00016613671323284507)),(to_sfixed_a(-0.351686030626297)),(to_sfixed_a(0.028372298926115036)),(to_sfixed_a(0.0002435502246953547)),(to_sfixed_a(-8.531605999451131e-07)),(to_sfixed_a(-9.438452980248258e-05)),(to_sfixed_a(0.0002955868258140981)),(to_sfixed_a(-0.00017557514365762472)),(to_sfixed_a(-0.0008888906450010836)),(to_sfixed_a(0.23663556575775146)),(to_sfixed_a(-0.00010415528959129006)),(to_sfixed_a(-6.483194010797888e-05)),(to_sfixed_a(0.07492532581090927)),(to_sfixed_a(0.0001716820988804102)),(to_sfixed_a(1.2295800843276083e-05)),(to_sfixed_a(-0.0002876909857150167)),(to_sfixed_a(0.006984231527894735)),(to_sfixed_a(0.00017491186736151576)),(to_sfixed_a(0.00031163261155597866)),(to_sfixed_a(4.723145684693009e-05)),(to_sfixed_a(0.0009942391188815236)),(to_sfixed_a(-2.5045665097422898e-08)),(to_sfixed_a(0.0007067238911986351)),(to_sfixed_a(-0.00011197332059964538)),(to_sfixed_a(-2.79650412267074e-05)),(to_sfixed_a(0.018720686435699463)),(to_sfixed_a(1.2310894817346707e-05)),(to_sfixed_a(3.691393067128956e-05)),(to_sfixed_a(-2.628024958539754e-06)),(to_sfixed_a(5.399268047767691e-05)),(to_sfixed_a(-1.8105944036506116e-05)),(to_sfixed_a(-0.33895012736320496)),(to_sfixed_a(-0.0002713938010856509)),(to_sfixed_a(0.009495649486780167)),(to_sfixed_a(1.1144999007228762e-05)),(to_sfixed_a(-7.635353540536016e-05)),(to_sfixed_a(0.00022882298799231648)),(to_sfixed_a(0.00025375105906277895)),(to_sfixed_a(0.001126241055317223)),(to_sfixed_a(-0.00012728996807709336)),(to_sfixed_a(0.004162808880209923)),(to_sfixed_a(0.0004984296392649412)),(to_sfixed_a(0.0002974200469907373)),(to_sfixed_a(0.0034900757018476725)),(to_sfixed_a(0.0001522386446595192)),(to_sfixed_a(-2.3409302229993045e-05)),(to_sfixed_a(-0.0005621819291263819)),(to_sfixed_a(0.014671994373202324)),(to_sfixed_a(-0.00010441498307045549)),(to_sfixed_a(0.00021567822841461748)),(to_sfixed_a(0.005358430556952953)),(to_sfixed_a(-0.11444837599992752)),(to_sfixed_a(0.003509087022393942)),(to_sfixed_a(0.23884007334709167)),(to_sfixed_a(-0.0011166651966050267)),(to_sfixed_a(-0.001851489651016891)),(to_sfixed_a(-0.0001455039600841701)),(to_sfixed_a(0.024311522021889687)),(to_sfixed_a(-8.433994662482291e-05)),(to_sfixed_a(-0.00015546957729384303)),(to_sfixed_a(5.8605975937098265e-05)),(to_sfixed_a(-7.99610570538789e-05)),(to_sfixed_a(-0.41301825642585754)),(to_sfixed_a(0.00045877715456299484)),(to_sfixed_a(-0.0014655994018539786)),(to_sfixed_a(-0.0064787063747644424)),(to_sfixed_a(-0.0038530060555785894)),(to_sfixed_a(-0.0002286417584400624)),(to_sfixed_a(0.00201806821860373)),(to_sfixed_a(0.008961498737335205)),(to_sfixed_a(-7.039285264909267e-05)),(to_sfixed_a(0.023449523374438286)),(to_sfixed_a(1.5818715837667696e-05)),(to_sfixed_a(0.0024140053428709507)),(to_sfixed_a(-0.0020991647616028786)),(to_sfixed_a(-1.0670992196537554e-06)),(to_sfixed_a(8.318581967614591e-05)),(to_sfixed_a(7.034548616502434e-05)),(to_sfixed_a(-1.1690899555105716e-05)),(to_sfixed_a(0.0001554307818878442)),(to_sfixed_a(-3.788489993894473e-05)),(to_sfixed_a(-0.002036679768934846)),(to_sfixed_a(-9.96551534626633e-06)),(to_sfixed_a(-0.0007560881786048412)),(to_sfixed_a(8.665402128826827e-05)),(to_sfixed_a(0.002348892390727997)),(to_sfixed_a(0.019567258656024933)),(to_sfixed_a(4.7299145080614835e-05)),(to_sfixed_a(6.644967652391642e-05)),(to_sfixed_a(-1.7342943465337157e-05)),(to_sfixed_a(-9.463978130952455e-06)),(to_sfixed_a(-0.0003155162266921252)),(to_sfixed_a(5.1164017349947244e-05)),(to_sfixed_a(0.0024367873556911945)),(to_sfixed_a(0.014558381401002407)),(to_sfixed_a(-7.10629319655709e-05)),(to_sfixed_a(8.741195779293776e-05)),(to_sfixed_a(0.00026757153682410717)),(to_sfixed_a(0.00029652711236849427)),(to_sfixed_a(-5.997479456709698e-05)),(to_sfixed_a(-0.0019447061931714416)),(to_sfixed_a(2.2743071895092726e-05)),(to_sfixed_a(-7.592374458909035e-06)),(to_sfixed_a(-0.00010569431469775736)),(to_sfixed_a(0.32092341780662537)),(to_sfixed_a(0.008075112476944923)),(to_sfixed_a(0.0005653110565617681)),(to_sfixed_a(0.00023810641141608357)),(to_sfixed_a(0.00018426644965074956)),(to_sfixed_a(-5.212862743064761e-05)),(to_sfixed_a(0.0057393331080675125)),(to_sfixed_a(0.005745162721723318)),(to_sfixed_a(0.006027999799698591)),(to_sfixed_a(-2.315541496500373e-05)),(to_sfixed_a(-0.0012024147436022758)),(to_sfixed_a(-0.00021434942027553916)),(to_sfixed_a(0.00012663302186410874)),(to_sfixed_a(1.5445417375303805e-05)),(to_sfixed_a(0.02143990993499756)),(to_sfixed_a(3.44429281540215e-06)),(to_sfixed_a(-0.4710310399532318)),(to_sfixed_a(-2.5120074496953748e-05)),(to_sfixed_a(0.014981313608586788)),(to_sfixed_a(0.004642740823328495)),(to_sfixed_a(6.435893737943843e-05)),(to_sfixed_a(0.01204997580498457)),(to_sfixed_a(0.008759581483900547)),(to_sfixed_a(-0.00015787765732966363)),(to_sfixed_a(-0.000571912620216608)),(to_sfixed_a(0.0001357157016173005)),(to_sfixed_a(-4.4562912080436945e-06)),(to_sfixed_a(0.0008409347501583397)),(to_sfixed_a(-0.0036866599693894386)),(to_sfixed_a(-0.00018574883870314807)),(to_sfixed_a(-1.6402060282416642e-05)),(to_sfixed_a(-0.013556195423007011)),(to_sfixed_a(6.1129750974942e-05)),(to_sfixed_a(-4.507879930315539e-05)),(to_sfixed_a(7.522612577304244e-07)),(to_sfixed_a(2.2443038687924854e-05)),(to_sfixed_a(0.00010162751277675852)),(to_sfixed_a(2.821587258949876e-05)),(to_sfixed_a(-0.00030785557464696467)),(to_sfixed_a(0.00016819355369079858)),(to_sfixed_a(3.8355505239451304e-05)),(to_sfixed_a(0.009181071072816849)),(to_sfixed_a(-0.0036656390875577927)),(to_sfixed_a(-0.00016768249042797834)),(to_sfixed_a(0.00023555940424557775)),(to_sfixed_a(2.8070935513824224e-05)),(to_sfixed_a(-6.986640801187605e-05)),(to_sfixed_a(-7.702635775785893e-05)),(to_sfixed_a(0.4941520094871521)),(to_sfixed_a(0.0020957530941814184)),(to_sfixed_a(0.012121566571295261)),(to_sfixed_a(-7.553604518761858e-05)),(to_sfixed_a(0.00017657523858360946)),(to_sfixed_a(8.018600783543661e-05)),(to_sfixed_a(2.972698894154746e-05)),(to_sfixed_a(2.164530087611638e-06)),(to_sfixed_a(-3.134476355626248e-05)),(to_sfixed_a(-5.181427695788443e-06)),(to_sfixed_a(7.025479135336354e-06)),(to_sfixed_a(-0.00021050682698842138)),(to_sfixed_a(7.048424595268443e-05)),(to_sfixed_a(5.0209833716508e-05)),(to_sfixed_a(-0.00010724109597504139)),(to_sfixed_a(0.013206413015723228)),(to_sfixed_a(0.046490129083395004)),(to_sfixed_a(2.6893161702901125e-05)),(to_sfixed_a(-0.0029900004155933857)),(to_sfixed_a(-2.479971772118006e-05)),(to_sfixed_a(0.009583322331309319)),(to_sfixed_a(0.0001740192819852382)),(to_sfixed_a(0.4725054204463959)),(to_sfixed_a(-0.39971134066581726)),(to_sfixed_a(0.0225245151668787)));

    constant weight_n2_61 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.0912046730518341)),(to_sfixed_a(0.0016352393431589007)),(to_sfixed_a(0.0007518390193581581)),(to_sfixed_a(3.0347699066624045e-05)),(to_sfixed_a(-0.0011621570447459817)),(to_sfixed_a(-0.00023923667322378606)),(to_sfixed_a(-0.0018575957510620356)),(to_sfixed_a(-0.000140962001751177)),(to_sfixed_a(0.00011276744771748781)),(to_sfixed_a(-0.00012891387450508773)),(to_sfixed_a(0.00012142954801674932)),(to_sfixed_a(0.201053649187088)),(to_sfixed_a(0.0036759250797331333)),(to_sfixed_a(0.0007499116472899914)),(to_sfixed_a(-6.70557637931779e-05)),(to_sfixed_a(-0.00011854979675263166)),(to_sfixed_a(-9.599282930139452e-05)),(to_sfixed_a(-9.611679706722498e-05)),(to_sfixed_a(0.0018662173533812165)),(to_sfixed_a(0.0018412641948089004)),(to_sfixed_a(8.876301581040025e-05)),(to_sfixed_a(0.00015102047473192215)),(to_sfixed_a(6.713548646075651e-05)),(to_sfixed_a(0.004201728384941816)),(to_sfixed_a(-0.00366231775842607)),(to_sfixed_a(-7.698861008975655e-05)),(to_sfixed_a(-1.079483627108857e-05)),(to_sfixed_a(4.751175583805889e-05)),(to_sfixed_a(-0.0003042881435249001)),(to_sfixed_a(-6.569728429894894e-05)),(to_sfixed_a(-0.0004433044232428074)),(to_sfixed_a(-0.0001013758301269263)),(to_sfixed_a(0.0046701314859092236)),(to_sfixed_a(-1.7277925508096814e-05)),(to_sfixed_a(-0.00024998554727062583)),(to_sfixed_a(-7.831271068425849e-05)),(to_sfixed_a(0.005684466101229191)),(to_sfixed_a(0.2308748960494995)),(to_sfixed_a(0.010911935940384865)),(to_sfixed_a(-0.00031342540751211345)),(to_sfixed_a(0.07834087312221527)),(to_sfixed_a(0.4451209604740143)),(to_sfixed_a(-2.4242686777142808e-05)),(to_sfixed_a(-7.720256689935923e-06)),(to_sfixed_a(0.00028386502526700497)),(to_sfixed_a(0.0018887275364249945)),(to_sfixed_a(3.107350130449049e-05)),(to_sfixed_a(0.00011728127719834447)),(to_sfixed_a(-0.00014429702423512936)),(to_sfixed_a(-0.0033271920401602983)),(to_sfixed_a(0.002425555605441332)),(to_sfixed_a(-6.98951625963673e-05)),(to_sfixed_a(-3.740331158041954e-05)),(to_sfixed_a(-0.00017720337200444192)),(to_sfixed_a(-0.003129074117168784)),(to_sfixed_a(-0.0007298529963009059)),(to_sfixed_a(-0.0001769961672835052)),(to_sfixed_a(-0.010649222880601883)),(to_sfixed_a(-0.0001307301572524011)),(to_sfixed_a(-1.5051300579216331e-05)),(to_sfixed_a(-0.0012077748542651534)),(to_sfixed_a(-0.0010460700141265988)),(to_sfixed_a(8.120272832456976e-05)),(to_sfixed_a(0.0023870922159403563)),(to_sfixed_a(-4.793488187715411e-06)),(to_sfixed_a(-1.5040851394587662e-05)),(to_sfixed_a(-9.423951269127429e-05)),(to_sfixed_a(0.3187798261642456)),(to_sfixed_a(-0.0014988607726991177)),(to_sfixed_a(0.00011088778410339728)),(to_sfixed_a(-0.0045640431344509125)),(to_sfixed_a(-0.5383875966072083)),(to_sfixed_a(0.0019570712465792894)),(to_sfixed_a(-0.00010913285950664431)),(to_sfixed_a(0.0001449501869501546)),(to_sfixed_a(-6.429362838389352e-05)),(to_sfixed_a(-0.2799631357192993)),(to_sfixed_a(0.0055057029239833355)),(to_sfixed_a(0.00022055752924643457)),(to_sfixed_a(0.006991230882704258)),(to_sfixed_a(-0.001514414674602449)),(to_sfixed_a(0.00018197987810708582)),(to_sfixed_a(0.009937075898051262)),(to_sfixed_a(-0.004432779271155596)),(to_sfixed_a(0.00018643496150616556)),(to_sfixed_a(0.0002903161512222141)),(to_sfixed_a(-0.002245516749098897)),(to_sfixed_a(-7.9877077951096e-05)),(to_sfixed_a(7.474009180441499e-07)),(to_sfixed_a(2.2227242880035192e-05)),(to_sfixed_a(-0.0018388634780421853)),(to_sfixed_a(-0.0001958551147254184)),(to_sfixed_a(0.0009724894189275801)),(to_sfixed_a(-7.03449040884152e-05)),(to_sfixed_a(-0.0016146646812558174)),(to_sfixed_a(2.2807318600825965e-05)),(to_sfixed_a(7.007254316704348e-05)),(to_sfixed_a(1.0709314665291458e-05)),(to_sfixed_a(0.0001974529295694083)),(to_sfixed_a(0.00020510998729150742)),(to_sfixed_a(0.005581803619861603)),(to_sfixed_a(0.007873745635151863)),(to_sfixed_a(-7.044474477879703e-05)),(to_sfixed_a(0.011987266130745411)),(to_sfixed_a(-0.3590428829193115)),(to_sfixed_a(0.0015946284402161837)),(to_sfixed_a(6.301799294305965e-05)),(to_sfixed_a(6.668638525297865e-05)),(to_sfixed_a(-4.408639142639004e-05)),(to_sfixed_a(-0.004258894827216864)),(to_sfixed_a(0.005359895993024111)),(to_sfixed_a(-0.0002297579194419086)),(to_sfixed_a(0.00046939431922510266)),(to_sfixed_a(0.00013667404709849507)),(to_sfixed_a(0.00010182222467847168)),(to_sfixed_a(-7.632034248672426e-05)),(to_sfixed_a(0.001283104531466961)),(to_sfixed_a(-5.412587051978335e-05)),(to_sfixed_a(-0.0002826607378665358)),(to_sfixed_a(0.2545223832130432)),(to_sfixed_a(-0.00015549507224932313)),(to_sfixed_a(3.0275172321125865e-05)),(to_sfixed_a(-0.00018941520829685032)),(to_sfixed_a(0.00028297858079895377)),(to_sfixed_a(-6.972550181671977e-07)),(to_sfixed_a(0.007374952081590891)),(to_sfixed_a(0.011379704810678959)),(to_sfixed_a(5.5787495512049645e-06)),(to_sfixed_a(-7.15527858119458e-06)),(to_sfixed_a(4.2822131945285946e-05)),(to_sfixed_a(-3.1162711820797995e-05)),(to_sfixed_a(6.70708977850154e-05)),(to_sfixed_a(-2.816114283632487e-05)),(to_sfixed_a(-0.002514092717319727)),(to_sfixed_a(0.00020155857782810926)),(to_sfixed_a(-1.9487306417431682e-06)),(to_sfixed_a(-0.003591802902519703)),(to_sfixed_a(-1.4068533346289769e-05)),(to_sfixed_a(-0.00020380222122184932)),(to_sfixed_a(0.00018242215446662158)),(to_sfixed_a(-0.0003227698616683483)),(to_sfixed_a(6.628797564189881e-05)),(to_sfixed_a(0.00020591313659679145)),(to_sfixed_a(-3.295938950031996e-05)),(to_sfixed_a(-7.976921915542334e-05)),(to_sfixed_a(-8.144844468915835e-05)),(to_sfixed_a(-0.00163773144595325)),(to_sfixed_a(-0.00011835178884211928)),(to_sfixed_a(-0.00019547012925613672)),(to_sfixed_a(-0.002168832579627633)),(to_sfixed_a(-0.0002891812182497233)),(to_sfixed_a(5.233897900325246e-05)),(to_sfixed_a(0.0001090177393052727)),(to_sfixed_a(0.00014625742915086448)),(to_sfixed_a(-0.00012721118400804698)),(to_sfixed_a(0.0024046902544796467)),(to_sfixed_a(-0.00044793004053644836)),(to_sfixed_a(0.003834249684587121)),(to_sfixed_a(0.03086959198117256)),(to_sfixed_a(-0.00013592703908216208)),(to_sfixed_a(-0.00014856294728815556)),(to_sfixed_a(0.0001079348148778081)),(to_sfixed_a(0.0007175551145337522)),(to_sfixed_a(-0.0016434246208518744)),(to_sfixed_a(-0.008176552131772041)),(to_sfixed_a(0.0007006992236711085)),(to_sfixed_a(7.079647912178189e-05)),(to_sfixed_a(-0.002320686588063836)),(to_sfixed_a(7.646785525139421e-05)),(to_sfixed_a(-0.0002667855005711317)),(to_sfixed_a(0.0026856190524995327)),(to_sfixed_a(0.0001829842512961477)),(to_sfixed_a(-0.0005243811174295843)),(to_sfixed_a(-6.682011007796973e-05)),(to_sfixed_a(0.0035367142409086227)),(to_sfixed_a(-0.0004581071261782199)),(to_sfixed_a(0.32216858863830566)),(to_sfixed_a(0.0007117476779967546)),(to_sfixed_a(0.006714111194014549)),(to_sfixed_a(-0.29172390699386597)),(to_sfixed_a(-0.00022206005814950913)),(to_sfixed_a(-0.03963810205459595)),(to_sfixed_a(0.00015252303273882717)),(to_sfixed_a(5.819246871396899e-05)),(to_sfixed_a(0.00011548969632713124)),(to_sfixed_a(-5.7207518693758175e-05)),(to_sfixed_a(0.0041214837692677975)),(to_sfixed_a(-0.0023609052877873182)),(to_sfixed_a(-0.0014682464534416795)),(to_sfixed_a(0.0002455135982017964)),(to_sfixed_a(0.0004031510034110397)),(to_sfixed_a(-1.912891457322985e-05)),(to_sfixed_a(0.4481872022151947)),(to_sfixed_a(0.001148595241829753)),(to_sfixed_a(6.929266237420961e-05)),(to_sfixed_a(-0.00015123152115847915)),(to_sfixed_a(0.00016719812992960215)),(to_sfixed_a(-0.12197653204202652)),(to_sfixed_a(-0.0004004209185950458)),(to_sfixed_a(0.00019832576799672097)),(to_sfixed_a(-4.99781162943691e-06)),(to_sfixed_a(-3.8793281419202685e-05)),(to_sfixed_a(0.00026871333830058575)),(to_sfixed_a(-6.112740811659023e-05)),(to_sfixed_a(0.00011535134399309754)),(to_sfixed_a(-0.00036457667010836303)),(to_sfixed_a(-0.003719981061294675)),(to_sfixed_a(0.006148098967969418)),(to_sfixed_a(-0.0012123011983931065)),(to_sfixed_a(-0.000982371042482555)),(to_sfixed_a(0.006171782035380602)),(to_sfixed_a(0.00015769785386510193)),(to_sfixed_a(0.00016744025924708694)),(to_sfixed_a(-9.80373442871496e-06)),(to_sfixed_a(-0.00027079437859356403)),(to_sfixed_a(0.0001365559292025864)),(to_sfixed_a(-0.0025117455516010523)),(to_sfixed_a(0.0001064608441083692)),(to_sfixed_a(-0.0017071387264877558)),(to_sfixed_a(-4.2992120143026114e-05)),(to_sfixed_a(0.00017877868958748877)),(to_sfixed_a(-1.4724231732543558e-05)),(to_sfixed_a(-0.0001689455530140549)),(to_sfixed_a(0.0008149972418323159)),(to_sfixed_a(-0.28269970417022705)),(to_sfixed_a(-1.0858930181711912e-06)),(to_sfixed_a(3.680640656966716e-05)),(to_sfixed_a(0.00015426866593770683)),(to_sfixed_a(-0.15636833012104034)),(to_sfixed_a(0.2697472870349884)),(to_sfixed_a(-0.3812439441680908)),(to_sfixed_a(-0.0001365135540254414)),(to_sfixed_a(2.8275553631829098e-05)),(to_sfixed_a(6.884002505103126e-05)),(to_sfixed_a(-0.0006313545163720846)),(to_sfixed_a(0.0006296219653449953)),(to_sfixed_a(0.0022298952098935843)),(to_sfixed_a(-7.772578101139516e-05)),(to_sfixed_a(-5.416309431893751e-05)),(to_sfixed_a(-0.00044377826270647347)),(to_sfixed_a(0.0001863956858869642)),(to_sfixed_a(-0.00014940713299438357)),(to_sfixed_a(-0.00043499493040144444)),(to_sfixed_a(-0.00024700560607016087)),(to_sfixed_a(-0.0022511817514896393)),(to_sfixed_a(-0.0027347698342055082)),(to_sfixed_a(-0.00039481359999626875)),(to_sfixed_a(0.24937626719474792)),(to_sfixed_a(8.949905168265104e-05)),(to_sfixed_a(-9.992389823310077e-05)),(to_sfixed_a(0.00022802843886893243)),(to_sfixed_a(-0.00010350051888963208)),(to_sfixed_a(-0.0022723174188286066)),(to_sfixed_a(0.00028650497552007437)),(to_sfixed_a(4.061315121361986e-05)),(to_sfixed_a(0.05966540053486824)),(to_sfixed_a(0.13127022981643677)),(to_sfixed_a(-0.00019329527276568115)),(to_sfixed_a(-9.727809811010957e-06)),(to_sfixed_a(0.00011491672921692953)),(to_sfixed_a(-6.787288293708116e-05)),(to_sfixed_a(0.48606300354003906)),(to_sfixed_a(-7.679538612137549e-06)),(to_sfixed_a(1.8752351024886593e-05)),(to_sfixed_a(0.0001482802035752684)),(to_sfixed_a(-0.001966190291568637)),(to_sfixed_a(-0.00011287411325611174)),(to_sfixed_a(4.2482388380449265e-06)),(to_sfixed_a(-0.00024303002282977104)),(to_sfixed_a(-0.16459518671035767)),(to_sfixed_a(0.023053260520100594)),(to_sfixed_a(5.529873305931687e-06)),(to_sfixed_a(0.00019960150530096143)),(to_sfixed_a(-9.354207577416673e-07)),(to_sfixed_a(0.00015457266999874264)),(to_sfixed_a(0.44235149025917053)),(to_sfixed_a(-0.004185643512755632)),(to_sfixed_a(-0.00014381793153006583)),(to_sfixed_a(-0.0051206923089921474)),(to_sfixed_a(-0.003882277524098754)),(to_sfixed_a(-2.3413565941154957e-05)),(to_sfixed_a(-4.688090120907873e-05)),(to_sfixed_a(-0.0001498337951488793)),(to_sfixed_a(0.0032025082036852837)),(to_sfixed_a(3.952439146814868e-05)),(to_sfixed_a(5.705835064873099e-06)),(to_sfixed_a(0.0021673578303307295)),(to_sfixed_a(0.009343262761831284)),(to_sfixed_a(4.533576429821551e-05)),(to_sfixed_a(-0.0003389034536667168)),(to_sfixed_a(-0.0012767721200361848)),(to_sfixed_a(-0.004026518203318119)),(to_sfixed_a(-0.23446473479270935)),(to_sfixed_a(0.00014892619219608605)),(to_sfixed_a(-0.002900456078350544)),(to_sfixed_a(0.013482406735420227)),(to_sfixed_a(-0.004238634370267391)),(to_sfixed_a(-2.3728494852548465e-05)),(to_sfixed_a(-0.29317381978034973)),(to_sfixed_a(0.31043344736099243)),(to_sfixed_a(0.2953740060329437)));

    constant weight_n2_62 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.3964781165122986)),(to_sfixed_a(0.0025567354168742895)),(to_sfixed_a(0.00397734809666872)),(to_sfixed_a(-6.677590135950595e-06)),(to_sfixed_a(-0.00034104904625564814)),(to_sfixed_a(0.00022643088595941663)),(to_sfixed_a(0.0003922799078281969)),(to_sfixed_a(-1.599938696017489e-05)),(to_sfixed_a(7.836327131371945e-05)),(to_sfixed_a(0.00017783153452910483)),(to_sfixed_a(-0.00016635858628433198)),(to_sfixed_a(-0.0034120227210223675)),(to_sfixed_a(-0.2512752115726471)),(to_sfixed_a(0.006874148268252611)),(to_sfixed_a(-0.00015212775906547904)),(to_sfixed_a(-7.81499402364716e-05)),(to_sfixed_a(0.1963854283094406)),(to_sfixed_a(-0.00011577548866625875)),(to_sfixed_a(0.008946167305111885)),(to_sfixed_a(0.00040100538171827793)),(to_sfixed_a(5.9908677940256894e-05)),(to_sfixed_a(-7.463966903742403e-05)),(to_sfixed_a(0.003395579755306244)),(to_sfixed_a(-0.0035757464356720448)),(to_sfixed_a(-0.006013742182403803)),(to_sfixed_a(0.012490684166550636)),(to_sfixed_a(0.00017258933803532273)),(to_sfixed_a(6.611109711229801e-05)),(to_sfixed_a(0.00381827331148088)),(to_sfixed_a(0.00016914220759645104)),(to_sfixed_a(0.0052720229141414165)),(to_sfixed_a(6.810465129092336e-05)),(to_sfixed_a(-0.003234399249777198)),(to_sfixed_a(0.0002510561898816377)),(to_sfixed_a(7.774170080665499e-05)),(to_sfixed_a(-2.5474364520050585e-05)),(to_sfixed_a(-0.0009246626286767423)),(to_sfixed_a(0.00040293988422490656)),(to_sfixed_a(0.002297856379300356)),(to_sfixed_a(0.0003119671600870788)),(to_sfixed_a(-0.13537874817848206)),(to_sfixed_a(0.3378683030605316)),(to_sfixed_a(7.144102710299194e-05)),(to_sfixed_a(3.0983719625510275e-06)),(to_sfixed_a(0.018958961591124535)),(to_sfixed_a(0.019779318943619728)),(to_sfixed_a(-0.0053034075535833836)),(to_sfixed_a(0.003959805238991976)),(to_sfixed_a(0.00011692135012708604)),(to_sfixed_a(-0.0002927431487478316)),(to_sfixed_a(0.012734227813780308)),(to_sfixed_a(0.00041531823808327317)),(to_sfixed_a(-0.00014327348617371172)),(to_sfixed_a(-0.002363271079957485)),(to_sfixed_a(0.008564437739551067)),(to_sfixed_a(0.3448896110057831)),(to_sfixed_a(0.00021364173153415322)),(to_sfixed_a(-0.02304897829890251)),(to_sfixed_a(3.4313219657633454e-05)),(to_sfixed_a(6.997189484536648e-05)),(to_sfixed_a(0.009396963752806187)),(to_sfixed_a(0.00748922023922205)),(to_sfixed_a(-5.596988557954319e-05)),(to_sfixed_a(0.0031307144090533257)),(to_sfixed_a(4.3820502469316125e-05)),(to_sfixed_a(0.5028066635131836)),(to_sfixed_a(0.00014971534255892038)),(to_sfixed_a(0.17682868242263794)),(to_sfixed_a(1.6909070836845785e-05)),(to_sfixed_a(-0.0001561164390295744)),(to_sfixed_a(-0.007670590188354254)),(to_sfixed_a(0.014892255887389183)),(to_sfixed_a(0.015157395973801613)),(to_sfixed_a(-4.008006362710148e-05)),(to_sfixed_a(0.00029323319904506207)),(to_sfixed_a(-8.283774513984099e-05)),(to_sfixed_a(-0.11988657712936401)),(to_sfixed_a(0.00036482553696259856)),(to_sfixed_a(-0.0001194247743114829)),(to_sfixed_a(-0.3028337359428406)),(to_sfixed_a(0.006509371101856232)),(to_sfixed_a(7.772824028506875e-05)),(to_sfixed_a(-0.0017360060010105371)),(to_sfixed_a(-0.004257506690919399)),(to_sfixed_a(-5.865204002475366e-05)),(to_sfixed_a(-0.0036008423194289207)),(to_sfixed_a(0.012260785326361656)),(to_sfixed_a(-0.00727984681725502)),(to_sfixed_a(0.0001498904312029481)),(to_sfixed_a(0.00021897633268963546)),(to_sfixed_a(0.0013129854341968894)),(to_sfixed_a(-0.00017007050337269902)),(to_sfixed_a(-0.00480251619592309)),(to_sfixed_a(-0.000113450747448951)),(to_sfixed_a(0.005450621247291565)),(to_sfixed_a(-0.00044164975406602025)),(to_sfixed_a(-0.000100561766885221)),(to_sfixed_a(-0.00016332075756508857)),(to_sfixed_a(-3.2786119845695794e-06)),(to_sfixed_a(1.7230740922968835e-06)),(to_sfixed_a(-0.004518113099038601)),(to_sfixed_a(0.002840417204424739)),(to_sfixed_a(-4.656852979678661e-06)),(to_sfixed_a(0.0052802604623138905)),(to_sfixed_a(-0.06560823321342468)),(to_sfixed_a(0.002433271612972021)),(to_sfixed_a(7.52951018512249e-06)),(to_sfixed_a(9.326783583674114e-06)),(to_sfixed_a(-0.00010635518265189603)),(to_sfixed_a(-0.029972923919558525)),(to_sfixed_a(-0.3664872944355011)),(to_sfixed_a(6.730109453201294e-05)),(to_sfixed_a(0.0033615368884056807)),(to_sfixed_a(0.0001482182851759717)),(to_sfixed_a(-7.006959640420973e-05)),(to_sfixed_a(0.0019192753825336695)),(to_sfixed_a(-0.0019057802855968475)),(to_sfixed_a(0.0008097145473584533)),(to_sfixed_a(0.00024602373014204204)),(to_sfixed_a(0.2765370011329651)),(to_sfixed_a(0.00011237048602197319)),(to_sfixed_a(0.0001554395566927269)),(to_sfixed_a(0.0007766406051814556)),(to_sfixed_a(-0.00013339624274522066)),(to_sfixed_a(-9.67967207543552e-06)),(to_sfixed_a(0.25341346859931946)),(to_sfixed_a(-0.1671902984380722)),(to_sfixed_a(5.0815287977457047e-08)),(to_sfixed_a(-2.206315184594132e-05)),(to_sfixed_a(-0.0001434302539564669)),(to_sfixed_a(2.815686457324773e-05)),(to_sfixed_a(0.0002483335556462407)),(to_sfixed_a(0.3783513903617859)),(to_sfixed_a(-0.0022664929274469614)),(to_sfixed_a(0.0003925490309484303)),(to_sfixed_a(-0.0001262879086425528)),(to_sfixed_a(0.022811854258179665)),(to_sfixed_a(0.0007860507466830313)),(to_sfixed_a(-0.0001515436451882124)),(to_sfixed_a(-0.00013556322664953768)),(to_sfixed_a(0.005082149989902973)),(to_sfixed_a(0.0002122127334587276)),(to_sfixed_a(-0.00016097357729449868)),(to_sfixed_a(-0.005297846160829067)),(to_sfixed_a(0.001074513653293252)),(to_sfixed_a(-9.390298509970307e-05)),(to_sfixed_a(-0.0021021340508013964)),(to_sfixed_a(0.00011505137081257999)),(to_sfixed_a(-8.475827053189278e-05)),(to_sfixed_a(-0.0019293945515528321)),(to_sfixed_a(1.0039657354354858e-05)),(to_sfixed_a(1.4237230061553419e-07)),(to_sfixed_a(-0.00037133932346478105)),(to_sfixed_a(8.535537199350074e-05)),(to_sfixed_a(5.734926526201889e-05)),(to_sfixed_a(-0.0012017188128083944)),(to_sfixed_a(-9.590288391336799e-05)),(to_sfixed_a(0.0013328870991244912)),(to_sfixed_a(4.002724017482251e-05)),(to_sfixed_a(-0.000180778035428375)),(to_sfixed_a(-6.697697972413152e-05)),(to_sfixed_a(-0.0002007479633903131)),(to_sfixed_a(-0.006342502776533365)),(to_sfixed_a(0.0025956197641789913)),(to_sfixed_a(-0.0052017406560480595)),(to_sfixed_a(-0.0025216725189238787)),(to_sfixed_a(-0.00011201507004443556)),(to_sfixed_a(0.2095952332019806)),(to_sfixed_a(5.975609383312985e-05)),(to_sfixed_a(0.00011631105007836595)),(to_sfixed_a(-0.000374576891772449)),(to_sfixed_a(-0.0019880691543221474)),(to_sfixed_a(0.0022679476533085108)),(to_sfixed_a(0.00016882896306924522)),(to_sfixed_a(-0.17263032495975494)),(to_sfixed_a(0.004625963978469372)),(to_sfixed_a(-0.5303172469139099)),(to_sfixed_a(0.32493454217910767)),(to_sfixed_a(-0.0038015181198716164)),(to_sfixed_a(0.7399805784225464)),(to_sfixed_a(0.0017386497929692268)),(to_sfixed_a(-0.023834852501749992)),(to_sfixed_a(-6.075343844713643e-05)),(to_sfixed_a(0.00018401199486106634)),(to_sfixed_a(-0.00016914785373955965)),(to_sfixed_a(0.004048920702189207)),(to_sfixed_a(0.25516071915626526)),(to_sfixed_a(-0.005309243220835924)),(to_sfixed_a(0.22872252762317657)),(to_sfixed_a(-0.016122911125421524)),(to_sfixed_a(-0.005380845628678799)),(to_sfixed_a(5.682814298779704e-05)),(to_sfixed_a(-0.009882871061563492)),(to_sfixed_a(0.007247674744576216)),(to_sfixed_a(2.9114409699104726e-05)),(to_sfixed_a(0.6054678559303284)),(to_sfixed_a(0.00017541449051350355)),(to_sfixed_a(-0.1298038214445114)),(to_sfixed_a(-0.0026464578695595264)),(to_sfixed_a(8.061361586442217e-05)),(to_sfixed_a(1.3831740943714976e-06)),(to_sfixed_a(0.00014851888408884406)),(to_sfixed_a(0.00021923180611338466)),(to_sfixed_a(-0.00011357721814420074)),(to_sfixed_a(0.0002749730774667114)),(to_sfixed_a(-0.002307344926521182)),(to_sfixed_a(-0.011634291149675846)),(to_sfixed_a(-0.5896345973014832)),(to_sfixed_a(4.3133608414791524e-05)),(to_sfixed_a(0.0032439481001347303)),(to_sfixed_a(-0.0023232512176036835)),(to_sfixed_a(1.2944990885443985e-05)),(to_sfixed_a(-0.00016659515677019954)),(to_sfixed_a(-0.00019214057829231024)),(to_sfixed_a(8.888619049685076e-07)),(to_sfixed_a(-7.113938772818074e-05)),(to_sfixed_a(-1.519000761618372e-05)),(to_sfixed_a(-0.0036297279875725508)),(to_sfixed_a(0.0017045049462467432)),(to_sfixed_a(-1.2080090527888387e-06)),(to_sfixed_a(0.00020811427384614944)),(to_sfixed_a(-0.00014658115105703473)),(to_sfixed_a(-0.0002276310115121305)),(to_sfixed_a(-0.006247712764889002)),(to_sfixed_a(-0.15681147575378418)),(to_sfixed_a(-7.094600005075336e-05)),(to_sfixed_a(-2.3169355699792504e-05)),(to_sfixed_a(-0.00018543517217040062)),(to_sfixed_a(0.0010267635807394981)),(to_sfixed_a(0.00944402813911438)),(to_sfixed_a(-0.0022781798616051674)),(to_sfixed_a(7.953053864184767e-05)),(to_sfixed_a(-0.00010137251229025424)),(to_sfixed_a(-0.00045984378084540367)),(to_sfixed_a(0.005853804759681225)),(to_sfixed_a(0.004706291016191244)),(to_sfixed_a(-0.5425775051116943)),(to_sfixed_a(-0.00025009637465700507)),(to_sfixed_a(-0.002113940427079797)),(to_sfixed_a(-2.8638794901780784e-05)),(to_sfixed_a(-0.008052659220993519)),(to_sfixed_a(-0.00011324059596518055)),(to_sfixed_a(0.09200646728277206)),(to_sfixed_a(-0.0001180529870907776)),(to_sfixed_a(0.014781991019845009)),(to_sfixed_a(0.005841435864567757)),(to_sfixed_a(0.5401577949523926)),(to_sfixed_a(-0.012109722942113876)),(to_sfixed_a(1.2472301023080945e-06)),(to_sfixed_a(0.12256282567977905)),(to_sfixed_a(-0.00015304436965379864)),(to_sfixed_a(7.028983236523345e-05)),(to_sfixed_a(0.00022231187904253602)),(to_sfixed_a(-0.000175075329025276)),(to_sfixed_a(9.718396904645488e-05)),(to_sfixed_a(0.008732874877750874)),(to_sfixed_a(-0.003353455103933811)),(to_sfixed_a(-5.8228892157785594e-05)),(to_sfixed_a(-0.0001486434048274532)),(to_sfixed_a(0.3540443480014801)),(to_sfixed_a(0.00024346262216567993)),(to_sfixed_a(-0.5227850079536438)),(to_sfixed_a(-0.0002039626706391573)),(to_sfixed_a(0.0004453863948583603)),(to_sfixed_a(-2.04151601792546e-05)),(to_sfixed_a(-0.0011198516003787518)),(to_sfixed_a(-0.00016583065735176206)),(to_sfixed_a(5.471920303534716e-07)),(to_sfixed_a(-1.401713234372437e-07)),(to_sfixed_a(-0.0007932125590741634)),(to_sfixed_a(0.000596114550717175)),(to_sfixed_a(-0.00014582497533410788)),(to_sfixed_a(5.838639481225982e-05)),(to_sfixed_a(0.0001489376008976251)),(to_sfixed_a(0.00016772988601587713)),(to_sfixed_a(-0.0045296913012862206)),(to_sfixed_a(0.009107621386647224)),(to_sfixed_a(0.21939769387245178)),(to_sfixed_a(-0.04226863384246826)),(to_sfixed_a(-0.0005000839591957629)),(to_sfixed_a(0.00010703925363486633)),(to_sfixed_a(0.000170580402482301)),(to_sfixed_a(-0.00015487706696148962)),(to_sfixed_a(0.0012797629460692406)),(to_sfixed_a(-6.642972584813833e-05)),(to_sfixed_a(0.00029726774664595723)),(to_sfixed_a(-0.16878639161586761)),(to_sfixed_a(0.008055517449975014)),(to_sfixed_a(3.947918594349176e-05)),(to_sfixed_a(-0.005813571624457836)),(to_sfixed_a(-0.021067151799798012)),(to_sfixed_a(0.0006443505990318954)),(to_sfixed_a(0.1994800865650177)),(to_sfixed_a(-2.048003261734266e-05)),(to_sfixed_a(-0.0038293912075459957)),(to_sfixed_a(0.0031945863738656044)),(to_sfixed_a(0.007954644970595837)),(to_sfixed_a(-6.893377576489002e-05)),(to_sfixed_a(-0.019076744094491005)),(to_sfixed_a(0.009930574335157871)),(to_sfixed_a(0.01214471273124218)));

    constant weight_n2_63 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.03792758285999298)),(to_sfixed_a(-0.26876991987228394)),(to_sfixed_a(-0.15874946117401123)),(to_sfixed_a(-0.00011300790356472135)),(to_sfixed_a(-0.001978490501642227)),(to_sfixed_a(3.837126132566482e-05)),(to_sfixed_a(0.0031313856597989798)),(to_sfixed_a(-0.00021812389604747295)),(to_sfixed_a(0.00016497616888955235)),(to_sfixed_a(7.706908218096942e-05)),(to_sfixed_a(-1.956777850864455e-07)),(to_sfixed_a(0.002506895223632455)),(to_sfixed_a(0.004170896951109171)),(to_sfixed_a(-0.0016922648064792156)),(to_sfixed_a(5.550937203224748e-06)),(to_sfixed_a(-0.00011810343858087435)),(to_sfixed_a(3.5651908547151834e-05)),(to_sfixed_a(7.180721149779856e-05)),(to_sfixed_a(-0.003004803555086255)),(to_sfixed_a(0.002416681731119752)),(to_sfixed_a(0.0001504092797404155)),(to_sfixed_a(0.00013376955757848918)),(to_sfixed_a(0.0017710445681586862)),(to_sfixed_a(0.0018817931413650513)),(to_sfixed_a(0.002914216835051775)),(to_sfixed_a(-3.170763739035465e-05)),(to_sfixed_a(-9.945491183316335e-05)),(to_sfixed_a(-0.00020654586842283607)),(to_sfixed_a(-0.0013364623300731182)),(to_sfixed_a(1.767536741681397e-05)),(to_sfixed_a(0.0020972085185348988)),(to_sfixed_a(0.00011622034071478993)),(to_sfixed_a(0.20472462475299835)),(to_sfixed_a(3.782966086873785e-05)),(to_sfixed_a(-0.0002459231182001531)),(to_sfixed_a(-0.00022138661006465554)),(to_sfixed_a(-0.3295843303203583)),(to_sfixed_a(-0.0012333635240793228)),(to_sfixed_a(0.00040484475903213024)),(to_sfixed_a(0.00017604778986424208)),(to_sfixed_a(0.004493482410907745)),(to_sfixed_a(-0.0018216350581496954)),(to_sfixed_a(1.7861908418126404e-05)),(to_sfixed_a(-3.491228198981844e-05)),(to_sfixed_a(0.00018173846183344722)),(to_sfixed_a(-0.00038284272886812687)),(to_sfixed_a(-0.16250482201576233)),(to_sfixed_a(-9.226157271768898e-05)),(to_sfixed_a(-0.00019465551304165274)),(to_sfixed_a(0.08667729049921036)),(to_sfixed_a(0.01661781221628189)),(to_sfixed_a(0.0005310210399329662)),(to_sfixed_a(-0.00023324944777414203)),(to_sfixed_a(-0.0031225483398884535)),(to_sfixed_a(0.0001456510362913832)),(to_sfixed_a(0.006297397892922163)),(to_sfixed_a(0.0002665205975063145)),(to_sfixed_a(0.010979007929563522)),(to_sfixed_a(-7.043856021482497e-05)),(to_sfixed_a(-0.00010582270624581724)),(to_sfixed_a(-0.0002770110440906137)),(to_sfixed_a(0.00449356297031045)),(to_sfixed_a(-0.000831166107673198)),(to_sfixed_a(3.3660424378467724e-05)),(to_sfixed_a(-4.580146196531132e-06)),(to_sfixed_a(0.001103140413761139)),(to_sfixed_a(-5.730547854909673e-05)),(to_sfixed_a(0.42025071382522583)),(to_sfixed_a(0.00524078868329525)),(to_sfixed_a(6.847808253951371e-05)),(to_sfixed_a(-0.1624099314212799)),(to_sfixed_a(0.0005721166962757707)),(to_sfixed_a(0.0012537436559796333)),(to_sfixed_a(3.7223901017569005e-05)),(to_sfixed_a(2.1761276002507657e-05)),(to_sfixed_a(0.00018278509378433228)),(to_sfixed_a(0.005986254196614027)),(to_sfixed_a(0.001906474120914936)),(to_sfixed_a(6.199852214194834e-05)),(to_sfixed_a(-0.009679058566689491)),(to_sfixed_a(0.0002503397117834538)),(to_sfixed_a(-8.561560389352962e-05)),(to_sfixed_a(-0.00330220814794302)),(to_sfixed_a(0.00010380722960690036)),(to_sfixed_a(-5.273250280879438e-06)),(to_sfixed_a(0.0013883971842005849)),(to_sfixed_a(0.006421985104680061)),(to_sfixed_a(0.0003213458985555917)),(to_sfixed_a(3.729107993422076e-05)),(to_sfixed_a(0.00016600577509962022)),(to_sfixed_a(0.0004414089780766517)),(to_sfixed_a(-5.7126773754134774e-05)),(to_sfixed_a(0.0006289619486778975)),(to_sfixed_a(0.00014006717537995428)),(to_sfixed_a(0.004001160617917776)),(to_sfixed_a(-2.9467977583408356e-05)),(to_sfixed_a(7.173894846346229e-05)),(to_sfixed_a(-7.1247253799811e-05)),(to_sfixed_a(-9.050132939592004e-05)),(to_sfixed_a(-1.1296302545815706e-05)),(to_sfixed_a(0.002188419457525015)),(to_sfixed_a(0.0010601709363982081)),(to_sfixed_a(-8.387837442569435e-05)),(to_sfixed_a(0.007229290436953306)),(to_sfixed_a(-0.29041680693626404)),(to_sfixed_a(0.0005831075832247734)),(to_sfixed_a(7.176223152782768e-05)),(to_sfixed_a(-0.0002739757183007896)),(to_sfixed_a(-6.880932778585702e-05)),(to_sfixed_a(0.0043458095751702785)),(to_sfixed_a(0.0016654765931889415)),(to_sfixed_a(0.00018953587277792394)),(to_sfixed_a(-0.00020614315872080624)),(to_sfixed_a(4.26650804001838e-05)),(to_sfixed_a(-4.5387667341856286e-05)),(to_sfixed_a(-0.001925838878378272)),(to_sfixed_a(-0.00021090780501253903)),(to_sfixed_a(0.0025472238194197416)),(to_sfixed_a(2.654443960636854e-06)),(to_sfixed_a(0.0011845971457660198)),(to_sfixed_a(-0.00017808123084250838)),(to_sfixed_a(-6.072673568269238e-05)),(to_sfixed_a(-0.0019879809115082026)),(to_sfixed_a(-7.935836038086563e-05)),(to_sfixed_a(8.073257049545646e-06)),(to_sfixed_a(0.006545563694089651)),(to_sfixed_a(0.003933336585760117)),(to_sfixed_a(0.00010552701860433444)),(to_sfixed_a(-0.00016643445997033268)),(to_sfixed_a(6.812354695284739e-05)),(to_sfixed_a(4.684982559410855e-05)),(to_sfixed_a(-0.00013517752813640982)),(to_sfixed_a(0.00031697319354861975)),(to_sfixed_a(-0.005167847964912653)),(to_sfixed_a(-0.0001813574490370229)),(to_sfixed_a(0.00010349987132940441)),(to_sfixed_a(0.006244776304811239)),(to_sfixed_a(0.0006512175896205008)),(to_sfixed_a(-6.729492451995611e-05)),(to_sfixed_a(7.935415487736464e-05)),(to_sfixed_a(-3.095805732300505e-05)),(to_sfixed_a(6.742827827110887e-05)),(to_sfixed_a(-0.0001973301696125418)),(to_sfixed_a(2.273278369102627e-06)),(to_sfixed_a(0.0025086253881454468)),(to_sfixed_a(0.0001361309114145115)),(to_sfixed_a(-0.0006463048048317432)),(to_sfixed_a(-6.696143100271001e-05)),(to_sfixed_a(-6.176450551720336e-05)),(to_sfixed_a(0.010648532770574093)),(to_sfixed_a(-6.513530388474464e-05)),(to_sfixed_a(-0.0002104148006765172)),(to_sfixed_a(-7.391256804112345e-05)),(to_sfixed_a(0.00010125700646312907)),(to_sfixed_a(7.891222048783675e-05)),(to_sfixed_a(0.24729643762111664)),(to_sfixed_a(-2.6131121558137238e-05)),(to_sfixed_a(0.007426534313708544)),(to_sfixed_a(4.764198820339516e-06)),(to_sfixed_a(-0.0002797903725877404)),(to_sfixed_a(-2.3735123249934986e-05)),(to_sfixed_a(-2.196443165303208e-05)),(to_sfixed_a(0.24247094988822937)),(to_sfixed_a(-9.426987526239827e-05)),(to_sfixed_a(0.0004764518525917083)),(to_sfixed_a(0.0008269259124062955)),(to_sfixed_a(-2.94740530080162e-05)),(to_sfixed_a(-0.0012499371077865362)),(to_sfixed_a(0.0001543681719340384)),(to_sfixed_a(5.838313518324867e-05)),(to_sfixed_a(0.0008307684329338372)),(to_sfixed_a(0.0025726796593517065)),(to_sfixed_a(0.0026701889000833035)),(to_sfixed_a(-0.00014876836212351918)),(to_sfixed_a(0.007816188968718052)),(to_sfixed_a(0.0005428103031590581)),(to_sfixed_a(0.004168905783444643)),(to_sfixed_a(0.15111559629440308)),(to_sfixed_a(-0.005557739641517401)),(to_sfixed_a(6.167087121866643e-05)),(to_sfixed_a(0.000287457718513906)),(to_sfixed_a(0.0174059197306633)),(to_sfixed_a(-3.603199729695916e-07)),(to_sfixed_a(6.0952392232138664e-05)),(to_sfixed_a(-0.00019990853616036475)),(to_sfixed_a(-0.0003446844930294901)),(to_sfixed_a(0.004859437700361013)),(to_sfixed_a(-0.0004883758374489844)),(to_sfixed_a(0.15238268673419952)),(to_sfixed_a(-0.00534841837361455)),(to_sfixed_a(-0.00022338939015753567)),(to_sfixed_a(-0.00030033523216843605)),(to_sfixed_a(0.07543322443962097)),(to_sfixed_a(-1.7641395970713347e-05)),(to_sfixed_a(-0.00015692262968514115)),(to_sfixed_a(0.0029381595086306334)),(to_sfixed_a(-0.00016184031846933067)),(to_sfixed_a(0.0037630556616932154)),(to_sfixed_a(-0.004723876714706421)),(to_sfixed_a(0.00030889728805050254)),(to_sfixed_a(-1.70044950209558e-05)),(to_sfixed_a(-6.639040657319129e-05)),(to_sfixed_a(1.3018448953516781e-05)),(to_sfixed_a(1.3647833839058876e-05)),(to_sfixed_a(2.822751412168145e-06)),(to_sfixed_a(-0.0020058348309248686)),(to_sfixed_a(-0.053688470274209976)),(to_sfixed_a(0.002504755975678563)),(to_sfixed_a(-0.00019016597070731223)),(to_sfixed_a(0.0025885605718940496)),(to_sfixed_a(0.01009355764836073)),(to_sfixed_a(0.00012893148232251406)),(to_sfixed_a(1.9665612853714265e-05)),(to_sfixed_a(-0.00015454919775947928)),(to_sfixed_a(-5.8500248997006565e-05)),(to_sfixed_a(0.00010539734648773447)),(to_sfixed_a(0.001089621800929308)),(to_sfixed_a(0.0014324388466775417)),(to_sfixed_a(0.007367252372205257)),(to_sfixed_a(0.00015541166067123413)),(to_sfixed_a(-0.0001511516165919602)),(to_sfixed_a(-0.0001930376747623086)),(to_sfixed_a(-0.00018338632071390748)),(to_sfixed_a(-0.000939849647693336)),(to_sfixed_a(-0.3553464114665985)),(to_sfixed_a(-0.00013683787256013602)),(to_sfixed_a(9.014271199703217e-06)),(to_sfixed_a(2.0281579054426402e-05)),(to_sfixed_a(-0.003831644309684634)),(to_sfixed_a(0.002947400324046612)),(to_sfixed_a(-0.3325175940990448)),(to_sfixed_a(-6.203028897289187e-05)),(to_sfixed_a(0.00010564114927547053)),(to_sfixed_a(-1.266312028747052e-05)),(to_sfixed_a(0.0002885445428546518)),(to_sfixed_a(0.2890062630176544)),(to_sfixed_a(-0.007706705015152693)),(to_sfixed_a(3.728092269739136e-05)),(to_sfixed_a(-0.0016525662504136562)),(to_sfixed_a(-1.5412369975820184e-06)),(to_sfixed_a(0.003675322514027357)),(to_sfixed_a(0.00011565773456823081)),(to_sfixed_a(0.0004159583477303386)),(to_sfixed_a(-0.00018668570555746555)),(to_sfixed_a(-0.0005387224373407662)),(to_sfixed_a(0.0023768434766680002)),(to_sfixed_a(0.004707151558250189)),(to_sfixed_a(-4.969693691236898e-05)),(to_sfixed_a(0.00029635129612870514)),(to_sfixed_a(0.0023750218097120523)),(to_sfixed_a(0.006988861598074436)),(to_sfixed_a(-9.101707837544382e-05)),(to_sfixed_a(5.959066766081378e-05)),(to_sfixed_a(5.811550363432616e-05)),(to_sfixed_a(-1.534070906927809e-05)),(to_sfixed_a(0.2860705554485321)),(to_sfixed_a(0.39915692806243896)),(to_sfixed_a(7.019265467533842e-05)),(to_sfixed_a(-4.236477252561599e-06)),(to_sfixed_a(-0.006404486950486898)),(to_sfixed_a(-0.00026304443599656224)),(to_sfixed_a(-0.0009486868511885405)),(to_sfixed_a(-1.0279145499225706e-05)),(to_sfixed_a(5.364037860999815e-05)),(to_sfixed_a(-0.00041985372081398964)),(to_sfixed_a(-1.4633835235144943e-05)),(to_sfixed_a(8.375493052881211e-06)),(to_sfixed_a(0.00021284091053530574)),(to_sfixed_a(4.765103221870959e-05)),(to_sfixed_a(0.00532059371471405)),(to_sfixed_a(-0.187758669257164)),(to_sfixed_a(6.333310011541471e-05)),(to_sfixed_a(0.00014138816914055496)),(to_sfixed_a(-6.400480924639851e-05)),(to_sfixed_a(-0.00014929073222447187)),(to_sfixed_a(-0.0019096223404631019)),(to_sfixed_a(-0.0056723845191299915)),(to_sfixed_a(0.0025179972872138023)),(to_sfixed_a(0.0029987080488353968)),(to_sfixed_a(-0.3069196939468384)),(to_sfixed_a(-0.00018594812718220055)),(to_sfixed_a(0.00015351340698543936)),(to_sfixed_a(-3.0099981813691556e-06)),(to_sfixed_a(0.0015788135351613164)),(to_sfixed_a(-0.00013541188673116267)),(to_sfixed_a(-4.6860441216267645e-06)),(to_sfixed_a(0.0028203721158206463)),(to_sfixed_a(0.0017494442872703075)),(to_sfixed_a(-0.00014540078700520098)),(to_sfixed_a(-0.3760404884815216)),(to_sfixed_a(-9.153752762358636e-05)),(to_sfixed_a(0.003633614396676421)),(to_sfixed_a(0.01682092621922493)),(to_sfixed_a(-9.997610322898254e-05)),(to_sfixed_a(-0.0009088970255106688)),(to_sfixed_a(-4.6421937440754846e-05)),(to_sfixed_a(-0.00029997900128364563)),(to_sfixed_a(0.00019717424584086984)),(to_sfixed_a(0.4588697850704193)),(to_sfixed_a(0.002980594988912344)),(to_sfixed_a(0.002214632695540786)));

    constant weight_n2_64 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.13560286164283752)),(to_sfixed_a(0.031668439507484436)),(to_sfixed_a(-0.4006825089454651)),(to_sfixed_a(0.0002270713885081932)),(to_sfixed_a(-0.004093949683010578)),(to_sfixed_a(-9.425348252989352e-07)),(to_sfixed_a(0.0028768451884388924)),(to_sfixed_a(-0.00018747174181044102)),(to_sfixed_a(-1.6852165572345257e-05)),(to_sfixed_a(-6.16033939877525e-05)),(to_sfixed_a(0.0001462748768972233)),(to_sfixed_a(-0.00029224593890830874)),(to_sfixed_a(0.004307041876018047)),(to_sfixed_a(-0.0005478317034430802)),(to_sfixed_a(0.0001619613030925393)),(to_sfixed_a(2.305445377714932e-06)),(to_sfixed_a(0.0005842173704877496)),(to_sfixed_a(6.276587373577058e-05)),(to_sfixed_a(-0.002679746365174651)),(to_sfixed_a(-0.00011602135782595724)),(to_sfixed_a(0.000227725860895589)),(to_sfixed_a(6.582727655768394e-05)),(to_sfixed_a(8.505125879310071e-05)),(to_sfixed_a(-0.00017750448023434728)),(to_sfixed_a(0.4031981825828552)),(to_sfixed_a(0.0031929968390613794)),(to_sfixed_a(0.00019926714594475925)),(to_sfixed_a(-5.7588982599554583e-05)),(to_sfixed_a(-0.00021096515411045402)),(to_sfixed_a(0.00020079873502254486)),(to_sfixed_a(0.3847103714942932)),(to_sfixed_a(-6.256654160097241e-06)),(to_sfixed_a(0.0014267824590206146)),(to_sfixed_a(1.922231967910193e-05)),(to_sfixed_a(-0.0002415027847746387)),(to_sfixed_a(-0.00017641051090322435)),(to_sfixed_a(-0.05263759568333626)),(to_sfixed_a(0.7052317261695862)),(to_sfixed_a(-0.24767880141735077)),(to_sfixed_a(-6.12335279583931e-05)),(to_sfixed_a(-0.0008849190198816359)),(to_sfixed_a(-0.00036759497015736997)),(to_sfixed_a(-6.134585419204086e-05)),(to_sfixed_a(4.938556230627e-06)),(to_sfixed_a(-0.002379519632086158)),(to_sfixed_a(0.4499166011810303)),(to_sfixed_a(-3.1046176445670426e-05)),(to_sfixed_a(-3.873130845022388e-05)),(to_sfixed_a(7.5836869655177e-06)),(to_sfixed_a(0.0008547752513550222)),(to_sfixed_a(0.000522713060490787)),(to_sfixed_a(6.44570536678657e-05)),(to_sfixed_a(-2.6775014703162014e-06)),(to_sfixed_a(-5.568181222770363e-07)),(to_sfixed_a(-0.00045618024887517095)),(to_sfixed_a(-0.027363071218132973)),(to_sfixed_a(1.5298675862140954e-05)),(to_sfixed_a(-0.004886792041361332)),(to_sfixed_a(7.442124478984624e-05)),(to_sfixed_a(0.00023636702098883688)),(to_sfixed_a(-0.4663046598434448)),(to_sfixed_a(-1.7774809748516418e-05)),(to_sfixed_a(-4.706444087787531e-05)),(to_sfixed_a(0.001778317498974502)),(to_sfixed_a(-4.5129745558369905e-06)),(to_sfixed_a(-0.1248612105846405)),(to_sfixed_a(0.00014080223627388477)),(to_sfixed_a(-0.00045829321607016027)),(to_sfixed_a(9.484343900112435e-05)),(to_sfixed_a(-7.151455793064088e-05)),(to_sfixed_a(0.0019681674893945456)),(to_sfixed_a(-0.0009444055613130331)),(to_sfixed_a(-9.989042155211791e-05)),(to_sfixed_a(2.3640342988073826e-05)),(to_sfixed_a(1.7347774701192975e-05)),(to_sfixed_a(-6.912174285389483e-06)),(to_sfixed_a(0.0014767531538382173)),(to_sfixed_a(0.2204631268978119)),(to_sfixed_a(5.8613994042389095e-05)),(to_sfixed_a(-0.00048598748981021345)),(to_sfixed_a(-0.0016008740058168769)),(to_sfixed_a(-0.00019909281400032341)),(to_sfixed_a(0.003247420070692897)),(to_sfixed_a(-0.007533102761954069)),(to_sfixed_a(-0.00016735019744373858)),(to_sfixed_a(0.3949466943740845)),(to_sfixed_a(-0.008008654229342937)),(to_sfixed_a(-0.0006073905387893319)),(to_sfixed_a(-2.771685103652999e-07)),(to_sfixed_a(-0.00020300140022300184)),(to_sfixed_a(-0.41105347871780396)),(to_sfixed_a(-8.608424832345918e-05)),(to_sfixed_a(0.3534521758556366)),(to_sfixed_a(0.0001489549467805773)),(to_sfixed_a(0.001846542814746499)),(to_sfixed_a(9.17065772227943e-05)),(to_sfixed_a(0.00014650961384177208)),(to_sfixed_a(-0.0001675028179306537)),(to_sfixed_a(3.193724842276424e-05)),(to_sfixed_a(0.00011202467430848628)),(to_sfixed_a(0.24983429908752441)),(to_sfixed_a(0.19721435010433197)),(to_sfixed_a(2.9729591915383935e-05)),(to_sfixed_a(-0.0002178964059567079)),(to_sfixed_a(0.00798804871737957)),(to_sfixed_a(-0.00015106437786016613)),(to_sfixed_a(-0.0001044178061420098)),(to_sfixed_a(0.00010673066572053358)),(to_sfixed_a(-0.00018792338960338384)),(to_sfixed_a(-0.0016496494645252824)),(to_sfixed_a(0.00723776500672102)),(to_sfixed_a(-0.00014909071614965796)),(to_sfixed_a(-3.641203511506319e-05)),(to_sfixed_a(7.076461042743176e-05)),(to_sfixed_a(5.777932528872043e-05)),(to_sfixed_a(0.0003888337523676455)),(to_sfixed_a(-0.0004327855131123215)),(to_sfixed_a(0.0001904835517052561)),(to_sfixed_a(-2.8098365874029696e-06)),(to_sfixed_a(0.14530372619628906)),(to_sfixed_a(-2.8115668101236224e-05)),(to_sfixed_a(-0.00019813215476460755)),(to_sfixed_a(-5.843104008818045e-05)),(to_sfixed_a(-0.0001785854110494256)),(to_sfixed_a(1.756608980940655e-05)),(to_sfixed_a(-0.15056893229484558)),(to_sfixed_a(-0.0016418768791481853)),(to_sfixed_a(-0.00019117558258585632)),(to_sfixed_a(-0.0002927092427853495)),(to_sfixed_a(0.00037758270627819)),(to_sfixed_a(0.0001181284460471943)),(to_sfixed_a(-0.0004456863389350474)),(to_sfixed_a(0.0022301976568996906)),(to_sfixed_a(-0.01817316561937332)),(to_sfixed_a(9.30262467591092e-06)),(to_sfixed_a(9.749017044669017e-05)),(to_sfixed_a(-0.0043825143948197365)),(to_sfixed_a(6.429240602301434e-05)),(to_sfixed_a(9.725859854370356e-06)),(to_sfixed_a(0.0001138309235102497)),(to_sfixed_a(-0.0002089870540658012)),(to_sfixed_a(-7.252964132931083e-05)),(to_sfixed_a(-0.00016900866467040032)),(to_sfixed_a(3.945691787521355e-05)),(to_sfixed_a(0.0007653482025489211)),(to_sfixed_a(-0.00011241218453506008)),(to_sfixed_a(0.00035501710954122245)),(to_sfixed_a(-4.4332045945338905e-07)),(to_sfixed_a(4.001241904916242e-05)),(to_sfixed_a(0.0005253205308690667)),(to_sfixed_a(-6.711453897878528e-05)),(to_sfixed_a(-0.00022942363284528255)),(to_sfixed_a(0.003059105249121785)),(to_sfixed_a(3.709815064212307e-05)),(to_sfixed_a(-0.00011578755220398307)),(to_sfixed_a(0.10869264602661133)),(to_sfixed_a(-0.0002292607823619619)),(to_sfixed_a(-0.002720697084441781)),(to_sfixed_a(-1.6972200683085248e-05)),(to_sfixed_a(-9.371413034386933e-05)),(to_sfixed_a(0.0004172809130977839)),(to_sfixed_a(-0.0001068624114850536)),(to_sfixed_a(0.4752846956253052)),(to_sfixed_a(-0.0803307518362999)),(to_sfixed_a(0.3576505184173584)),(to_sfixed_a(0.001344582880847156)),(to_sfixed_a(-0.00010364119953010231)),(to_sfixed_a(0.0007701233844272792)),(to_sfixed_a(-1.6323019735864364e-05)),(to_sfixed_a(0.0001167656882898882)),(to_sfixed_a(0.2054230123758316)),(to_sfixed_a(0.0002653352858033031)),(to_sfixed_a(0.0007252549985423684)),(to_sfixed_a(-1.3197437510825694e-05)),(to_sfixed_a(-0.0007022846257314086)),(to_sfixed_a(0.0007748507778160274)),(to_sfixed_a(0.001459105871617794)),(to_sfixed_a(0.27042585611343384)),(to_sfixed_a(-0.15624524652957916)),(to_sfixed_a(0.1418100893497467)),(to_sfixed_a(-6.39366771792993e-05)),(to_sfixed_a(0.004225455224514008)),(to_sfixed_a(5.745724047301337e-05)),(to_sfixed_a(-0.00024404824944213033)),(to_sfixed_a(-0.00023970955226104707)),(to_sfixed_a(-0.0006635623867623508)),(to_sfixed_a(0.007862295024096966)),(to_sfixed_a(-5.5763339332770556e-05)),(to_sfixed_a(-0.0002261977206217125)),(to_sfixed_a(0.0008812671876512468)),(to_sfixed_a(-0.0001960653462447226)),(to_sfixed_a(0.0003861271543428302)),(to_sfixed_a(0.00048791844164952636)),(to_sfixed_a(-0.0013167108409106731)),(to_sfixed_a(0.00011501460539875552)),(to_sfixed_a(-0.009891672059893608)),(to_sfixed_a(9.928048530127853e-05)),(to_sfixed_a(-0.00013122429663781077)),(to_sfixed_a(0.0035881015937775373)),(to_sfixed_a(6.901547749293968e-05)),(to_sfixed_a(-0.00011425757111283019)),(to_sfixed_a(0.00014744146028533578)),(to_sfixed_a(-0.00023516846704296768)),(to_sfixed_a(1.137666913564317e-06)),(to_sfixed_a(-4.7395213186973706e-05)),(to_sfixed_a(0.023284196853637695)),(to_sfixed_a(-0.0030271022114902735)),(to_sfixed_a(0.003450676565989852)),(to_sfixed_a(-0.2740180790424347)),(to_sfixed_a(-0.004290599375963211)),(to_sfixed_a(0.00127714267000556)),(to_sfixed_a(-1.8133141566067934e-06)),(to_sfixed_a(-0.00019167571736034006)),(to_sfixed_a(-2.667962689884007e-06)),(to_sfixed_a(-2.9311362595763057e-05)),(to_sfixed_a(-0.00018066824122797698)),(to_sfixed_a(-0.00169550406280905)),(to_sfixed_a(0.0003952966071665287)),(to_sfixed_a(-0.006299057509750128)),(to_sfixed_a(0.0003148661053273827)),(to_sfixed_a(1.7416139598935843e-05)),(to_sfixed_a(4.9636564654065296e-05)),(to_sfixed_a(6.278056389419362e-05)),(to_sfixed_a(-0.0005002682446502149)),(to_sfixed_a(0.06997241824865341)),(to_sfixed_a(-1.8014614397543482e-05)),(to_sfixed_a(-0.0002504762960597873)),(to_sfixed_a(-6.813888467149809e-05)),(to_sfixed_a(-0.002171281957998872)),(to_sfixed_a(0.2076970338821411)),(to_sfixed_a(0.0030814828351140022)),(to_sfixed_a(-6.864898023195565e-05)),(to_sfixed_a(6.323740672087297e-05)),(to_sfixed_a(-0.00011939689284190536)),(to_sfixed_a(0.002663961611688137)),(to_sfixed_a(-0.0005974891246296465)),(to_sfixed_a(-0.16182127594947815)),(to_sfixed_a(-0.0003101529146078974)),(to_sfixed_a(-0.00020074259373359382)),(to_sfixed_a(4.567147698253393e-06)),(to_sfixed_a(8.468073792755604e-05)),(to_sfixed_a(4.7493136662524194e-05)),(to_sfixed_a(-3.917526555596851e-05)),(to_sfixed_a(6.972204573685303e-05)),(to_sfixed_a(-6.727899017278105e-05)),(to_sfixed_a(-0.0008293448481708765)),(to_sfixed_a(0.2519491910934448)),(to_sfixed_a(0.0006228145211935043)),(to_sfixed_a(-7.103555253706872e-05)),(to_sfixed_a(0.3139457106590271)),(to_sfixed_a(0.0005132207297720015)),(to_sfixed_a(-0.0001032726067933254)),(to_sfixed_a(-0.0006292237085290253)),(to_sfixed_a(-2.9454946343321353e-05)),(to_sfixed_a(-2.6304311177227646e-05)),(to_sfixed_a(0.002678374294191599)),(to_sfixed_a(0.0027763687539845705)),(to_sfixed_a(-0.00020029456936754286)),(to_sfixed_a(-0.00020067585865035653)),(to_sfixed_a(-5.025685823056847e-07)),(to_sfixed_a(9.515234705759212e-05)),(to_sfixed_a(0.00013813888654112816)),(to_sfixed_a(0.0001302432647207752)),(to_sfixed_a(-8.571155922254547e-05)),(to_sfixed_a(5.692272679880261e-06)),(to_sfixed_a(0.001099891378544271)),(to_sfixed_a(3.843815647996962e-07)),(to_sfixed_a(8.559342677472159e-05)),(to_sfixed_a(-3.1466930522583425e-05)),(to_sfixed_a(-0.4840490520000458)),(to_sfixed_a(0.004806898534297943)),(to_sfixed_a(-7.144041592255235e-05)),(to_sfixed_a(4.528547287918627e-05)),(to_sfixed_a(-0.0001172009069705382)),(to_sfixed_a(6.788612517993897e-05)),(to_sfixed_a(0.004959996324032545)),(to_sfixed_a(0.000913107069209218)),(to_sfixed_a(-0.00019530230201780796)),(to_sfixed_a(-0.2827022671699524)),(to_sfixed_a(0.00064374681096524)),(to_sfixed_a(8.357070328202099e-06)),(to_sfixed_a(-0.0002873291668947786)),(to_sfixed_a(-6.624116213060915e-05)),(to_sfixed_a(9.489132935414091e-05)),(to_sfixed_a(-0.00010823797492776066)),(to_sfixed_a(-0.00011298054596409202)),(to_sfixed_a(0.0001505729742348194)),(to_sfixed_a(0.1461237072944641)),(to_sfixed_a(2.3471613531000912e-05)),(to_sfixed_a(-9.911393135553226e-05)),(to_sfixed_a(0.0006488108774647117)),(to_sfixed_a(0.00114907487295568)),(to_sfixed_a(-0.35179802775382996)),(to_sfixed_a(-2.634075644891709e-05)),(to_sfixed_a(0.0027064227033406496)),(to_sfixed_a(-0.38149553537368774)),(to_sfixed_a(-0.0017848036950454116)),(to_sfixed_a(-8.558069384889677e-05)),(to_sfixed_a(0.0009212970617227256)),(to_sfixed_a(0.014503605663776398)),(to_sfixed_a(0.0003713078622240573)));

    constant weight_n2_65 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.02419348619878292)),(to_sfixed_a(0.2644059658050537)),(to_sfixed_a(0.45517945289611816)),(to_sfixed_a(-0.00014924767310731113)),(to_sfixed_a(0.0018982948968186975)),(to_sfixed_a(-0.00011290119437035173)),(to_sfixed_a(0.007684969808906317)),(to_sfixed_a(1.3917015166953206e-06)),(to_sfixed_a(-6.73423201078549e-05)),(to_sfixed_a(-4.008215910289437e-06)),(to_sfixed_a(0.00030160180176608264)),(to_sfixed_a(-0.00310601107776165)),(to_sfixed_a(0.007823145017027855)),(to_sfixed_a(0.007074377965182066)),(to_sfixed_a(3.0502571462420747e-05)),(to_sfixed_a(0.00011608128261286765)),(to_sfixed_a(0.020298365503549576)),(to_sfixed_a(3.7569989217445254e-06)),(to_sfixed_a(-0.1906253546476364)),(to_sfixed_a(0.008235781453549862)),(to_sfixed_a(3.775360528379679e-05)),(to_sfixed_a(-0.00018280620861332864)),(to_sfixed_a(0.0015596951125189662)),(to_sfixed_a(0.3616219162940979)),(to_sfixed_a(0.007219282910227776)),(to_sfixed_a(0.0005985705065540969)),(to_sfixed_a(2.0560626580845565e-05)),(to_sfixed_a(-0.0013848096132278442)),(to_sfixed_a(0.00010523360106162727)),(to_sfixed_a(-1.3632845366373658e-05)),(to_sfixed_a(0.1512955278158188)),(to_sfixed_a(-0.0002370496658841148)),(to_sfixed_a(-0.00920606218278408)),(to_sfixed_a(8.993926167022437e-05)),(to_sfixed_a(0.00026494235498830676)),(to_sfixed_a(8.455090573988855e-05)),(to_sfixed_a(-0.010672718286514282)),(to_sfixed_a(-0.001736133941449225)),(to_sfixed_a(-0.17269881069660187)),(to_sfixed_a(-0.0001303462340729311)),(to_sfixed_a(0.013174718245863914)),(to_sfixed_a(0.03310484066605568)),(to_sfixed_a(-0.000107760148239322)),(to_sfixed_a(0.0002326963731320575)),(to_sfixed_a(0.03312670439481735)),(to_sfixed_a(-0.19975577294826508)),(to_sfixed_a(0.0006491929525509477)),(to_sfixed_a(0.010088139213621616)),(to_sfixed_a(0.00024279358331114054)),(to_sfixed_a(0.409753680229187)),(to_sfixed_a(0.0007864233339205384)),(to_sfixed_a(7.379155431408435e-05)),(to_sfixed_a(-4.441657802090049e-05)),(to_sfixed_a(-0.001314571825787425)),(to_sfixed_a(0.5087267160415649)),(to_sfixed_a(0.00032569500035606325)),(to_sfixed_a(-0.00024162551562767476)),(to_sfixed_a(0.04171251878142357)),(to_sfixed_a(1.7937109078047797e-06)),(to_sfixed_a(-0.00029821108910255134)),(to_sfixed_a(0.004322275519371033)),(to_sfixed_a(0.004893315024673939)),(to_sfixed_a(-0.0004591454635374248)),(to_sfixed_a(-0.0035729361698031425)),(to_sfixed_a(-0.00026216579135507345)),(to_sfixed_a(-0.4384821057319641)),(to_sfixed_a(-7.529921276727691e-05)),(to_sfixed_a(0.006097298115491867)),(to_sfixed_a(-0.0028091073036193848)),(to_sfixed_a(3.839243436232209e-05)),(to_sfixed_a(-0.9944912195205688)),(to_sfixed_a(-0.1102450042963028)),(to_sfixed_a(-0.3346887230873108)),(to_sfixed_a(-7.564904808532447e-05)),(to_sfixed_a(-1.1843185347970575e-05)),(to_sfixed_a(0.00044950353913009167)),(to_sfixed_a(-0.0018143029883503914)),(to_sfixed_a(0.0028642478864639997)),(to_sfixed_a(-0.00018655740132089704)),(to_sfixed_a(0.26152458786964417)),(to_sfixed_a(0.007726928219199181)),(to_sfixed_a(-3.0003349820617586e-05)),(to_sfixed_a(-0.003589688567444682)),(to_sfixed_a(0.004160259384661913)),(to_sfixed_a(3.679099609144032e-05)),(to_sfixed_a(0.0008299066103063524)),(to_sfixed_a(0.009239457547664642)),(to_sfixed_a(-0.00013902693171985447)),(to_sfixed_a(-0.0001686930627329275)),(to_sfixed_a(0.0003918416623491794)),(to_sfixed_a(0.32986167073249817)),(to_sfixed_a(-3.888584615197033e-06)),(to_sfixed_a(0.00875500962138176)),(to_sfixed_a(-0.0003161044733133167)),(to_sfixed_a(0.006959738675504923)),(to_sfixed_a(-7.741371518932283e-06)),(to_sfixed_a(0.00021793892665300518)),(to_sfixed_a(0.00010912014113273472)),(to_sfixed_a(-5.691176193067804e-05)),(to_sfixed_a(6.583382491953671e-05)),(to_sfixed_a(0.008515558205544949)),(to_sfixed_a(0.007652001921087503)),(to_sfixed_a(0.00011563238513190299)),(to_sfixed_a(0.017565779387950897)),(to_sfixed_a(0.006086112465709448)),(to_sfixed_a(0.007649134378880262)),(to_sfixed_a(0.00010922418005065992)),(to_sfixed_a(3.719756205100566e-05)),(to_sfixed_a(0.00012760046229232103)),(to_sfixed_a(0.007031908258795738)),(to_sfixed_a(0.007470931392163038)),(to_sfixed_a(-3.0200957553461194e-05)),(to_sfixed_a(0.0004339301958680153)),(to_sfixed_a(7.969041325850412e-05)),(to_sfixed_a(-0.0003011122753378004)),(to_sfixed_a(-0.1594850867986679)),(to_sfixed_a(0.003860385389998555)),(to_sfixed_a(0.0036192117258906364)),(to_sfixed_a(-0.00018071726663038135)),(to_sfixed_a(0.0034293984062969685)),(to_sfixed_a(-0.00013609291636385024)),(to_sfixed_a(5.004960257792845e-06)),(to_sfixed_a(0.0005505701992660761)),(to_sfixed_a(0.00013528249110095203)),(to_sfixed_a(0.00011293383431620896)),(to_sfixed_a(-0.5216110944747925)),(to_sfixed_a(0.027242032811045647)),(to_sfixed_a(-8.590222569182515e-05)),(to_sfixed_a(0.000300691113807261)),(to_sfixed_a(0.00011623678437899798)),(to_sfixed_a(0.00028769750497303903)),(to_sfixed_a(0.000290114403469488)),(to_sfixed_a(0.0009510965901426971)),(to_sfixed_a(-0.01860576681792736)),(to_sfixed_a(-0.00010395198478363454)),(to_sfixed_a(-0.00012859032722190022)),(to_sfixed_a(0.3522390127182007)),(to_sfixed_a(-0.003138905158266425)),(to_sfixed_a(0.00024373483029194176)),(to_sfixed_a(-0.00022006806102581322)),(to_sfixed_a(-0.002118667820468545)),(to_sfixed_a(0.00023727248481009156)),(to_sfixed_a(-9.597311145626009e-05)),(to_sfixed_a(0.4755669832229614)),(to_sfixed_a(0.24337010085582733)),(to_sfixed_a(0.19717863202095032)),(to_sfixed_a(-0.0018098182044923306)),(to_sfixed_a(6.78935248288326e-06)),(to_sfixed_a(3.699396984302439e-05)),(to_sfixed_a(0.0064136493019759655)),(to_sfixed_a(-5.625597987091169e-05)),(to_sfixed_a(1.7580241546966136e-06)),(to_sfixed_a(0.00066061329562217)),(to_sfixed_a(-2.565138856880367e-06)),(to_sfixed_a(-0.0001860566553659737)),(to_sfixed_a(-0.014134439639747143)),(to_sfixed_a(8.966483437689021e-05)),(to_sfixed_a(0.015310735441744328)),(to_sfixed_a(-0.00010332169767934829)),(to_sfixed_a(3.348422615090385e-05)),(to_sfixed_a(5.311179847922176e-06)),(to_sfixed_a(-3.8578451494686306e-05)),(to_sfixed_a(0.319335013628006)),(to_sfixed_a(0.00346489530056715)),(to_sfixed_a(0.0049974918365478516)),(to_sfixed_a(-0.0015056271804496646)),(to_sfixed_a(1.109373988583684e-05)),(to_sfixed_a(-0.00961316004395485)),(to_sfixed_a(-6.312462210189551e-05)),(to_sfixed_a(-0.0001306579215452075)),(to_sfixed_a(-0.0052419318817555904)),(to_sfixed_a(-0.00017149813356809318)),(to_sfixed_a(0.00497488584369421)),(to_sfixed_a(-2.9960610845591873e-05)),(to_sfixed_a(0.0035032941959798336)),(to_sfixed_a(0.0003366792807355523)),(to_sfixed_a(0.0023480765521526337)),(to_sfixed_a(-0.00013115935144014657)),(to_sfixed_a(0.007939069531857967)),(to_sfixed_a(0.00726043526083231)),(to_sfixed_a(-0.00022261192498262972)),(to_sfixed_a(-0.22715532779693604)),(to_sfixed_a(-0.000302697328152135)),(to_sfixed_a(-3.7059020542073995e-05)),(to_sfixed_a(-0.00020396422769408673)),(to_sfixed_a(-0.21149730682373047)),(to_sfixed_a(-0.48918795585632324)),(to_sfixed_a(-0.0019580742809921503)),(to_sfixed_a(-0.0010470820125192404)),(to_sfixed_a(-0.006106525659561157)),(to_sfixed_a(0.010899323038756847)),(to_sfixed_a(-2.5867366275633685e-05)),(to_sfixed_a(-0.2069995403289795)),(to_sfixed_a(0.0024881483986973763)),(to_sfixed_a(-0.00010557550558587536)),(to_sfixed_a(-0.329777330160141)),(to_sfixed_a(-0.00011354514572303742)),(to_sfixed_a(0.008449248038232327)),(to_sfixed_a(0.5030909776687622)),(to_sfixed_a(6.774053326807916e-05)),(to_sfixed_a(-0.00011622524471022189)),(to_sfixed_a(5.543469887925312e-05)),(to_sfixed_a(0.00017860250954981893)),(to_sfixed_a(-3.278259828221053e-05)),(to_sfixed_a(0.0002391243033343926)),(to_sfixed_a(0.15875208377838135)),(to_sfixed_a(0.0066507719457149506)),(to_sfixed_a(0.10725042223930359)),(to_sfixed_a(0.04989463835954666)),(to_sfixed_a(0.1073031947016716)),(to_sfixed_a(-0.12852059304714203)),(to_sfixed_a(-0.0001008486287901178)),(to_sfixed_a(5.335765308700502e-06)),(to_sfixed_a(3.7880672607570887e-06)),(to_sfixed_a(-0.00036873616045340896)),(to_sfixed_a(-0.0002203934418503195)),(to_sfixed_a(-0.0007842682534828782)),(to_sfixed_a(-0.0013872651616111398)),(to_sfixed_a(0.29676172137260437)),(to_sfixed_a(0.00011571998038562015)),(to_sfixed_a(-2.3673583200434223e-05)),(to_sfixed_a(-1.0352021490689367e-05)),(to_sfixed_a(8.521004929207265e-05)),(to_sfixed_a(-0.006053450051695108)),(to_sfixed_a(-0.530968189239502)),(to_sfixed_a(0.00015000553685240448)),(to_sfixed_a(-4.3995492887916043e-05)),(to_sfixed_a(-5.854664777871221e-06)),(to_sfixed_a(0.41107824444770813)),(to_sfixed_a(0.31842970848083496)),(to_sfixed_a(0.0004131795431021601)),(to_sfixed_a(0.00012868791236542165)),(to_sfixed_a(-1.1572912626434118e-05)),(to_sfixed_a(0.0001840031472966075)),(to_sfixed_a(0.009999768808484077)),(to_sfixed_a(-0.0021072274539619684)),(to_sfixed_a(-0.018902145326137543)),(to_sfixed_a(6.933573604328558e-05)),(to_sfixed_a(-0.0017275414429605007)),(to_sfixed_a(-0.00023553182836622)),(to_sfixed_a(0.005342049058526754)),(to_sfixed_a(0.0002619122969917953)),(to_sfixed_a(0.2916189134120941)),(to_sfixed_a(0.00016713391232769936)),(to_sfixed_a(-0.2820630371570587)),(to_sfixed_a(0.37202197313308716)),(to_sfixed_a(0.004823605064302683)),(to_sfixed_a(0.2541147470474243)),(to_sfixed_a(-5.74239093111828e-05)),(to_sfixed_a(0.013840219005942345)),(to_sfixed_a(0.025149976834654808)),(to_sfixed_a(-6.430577195715159e-05)),(to_sfixed_a(0.004120252560824156)),(to_sfixed_a(-4.538196662906557e-06)),(to_sfixed_a(6.330423639155924e-05)),(to_sfixed_a(-0.0011435498017817736)),(to_sfixed_a(0.2635750472545624)),(to_sfixed_a(-6.663668318651617e-05)),(to_sfixed_a(0.0004174144705757499)),(to_sfixed_a(0.0009293055045418441)),(to_sfixed_a(-0.00010443557403050363)),(to_sfixed_a(0.36336466670036316)),(to_sfixed_a(-8.452116162516177e-08)),(to_sfixed_a(-1.9840152162942104e-05)),(to_sfixed_a(-0.0001134836275014095)),(to_sfixed_a(0.006660341750830412)),(to_sfixed_a(0.0002317167673027143)),(to_sfixed_a(0.00024179357569664717)),(to_sfixed_a(0.0001936290500452742)),(to_sfixed_a(0.0024553542025387287)),(to_sfixed_a(-0.008790501393377781)),(to_sfixed_a(-0.0001674129016464576)),(to_sfixed_a(-0.0001792122784536332)),(to_sfixed_a(4.230349441058934e-05)),(to_sfixed_a(-0.00016738506383262575)),(to_sfixed_a(-0.0025849922094494104)),(to_sfixed_a(0.004856530111283064)),(to_sfixed_a(0.0016315599204972386)),(to_sfixed_a(0.23355485498905182)),(to_sfixed_a(0.002764349803328514)),(to_sfixed_a(6.199056224431843e-05)),(to_sfixed_a(0.00012815666559617966)),(to_sfixed_a(1.0806252248585224e-05)),(to_sfixed_a(0.008635650388896465)),(to_sfixed_a(0.00030333251925185323)),(to_sfixed_a(-1.4839890354778618e-05)),(to_sfixed_a(0.002140978118404746)),(to_sfixed_a(-0.00802409928292036)),(to_sfixed_a(-9.889910870697349e-05)),(to_sfixed_a(-1.747789792716503e-05)),(to_sfixed_a(0.003578060306608677)),(to_sfixed_a(0.0072498442605137825)),(to_sfixed_a(-0.0009428577614016831)),(to_sfixed_a(-0.00030798709485679865)),(to_sfixed_a(-0.002092055743560195)),(to_sfixed_a(0.00025549225392751396)),(to_sfixed_a(0.022641967982053757)),(to_sfixed_a(1.7651553207542747e-05)),(to_sfixed_a(0.0016876746667549014)),(to_sfixed_a(0.002624134300276637)),(to_sfixed_a(0.3692263960838318)));

    constant weight_n2_66 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.17055438458919525)),(to_sfixed_a(0.00010477962496224791)),(to_sfixed_a(0.0001844849466579035)),(to_sfixed_a(2.9138966056052595e-05)),(to_sfixed_a(0.0001652866485528648)),(to_sfixed_a(0.0001040961651597172)),(to_sfixed_a(-7.335772534133866e-05)),(to_sfixed_a(0.00044737086864188313)),(to_sfixed_a(7.165457645896822e-06)),(to_sfixed_a(0.00015751663886476308)),(to_sfixed_a(8.649483788758516e-06)),(to_sfixed_a(6.527705409098417e-05)),(to_sfixed_a(-4.541413363767788e-05)),(to_sfixed_a(0.00041109032463282347)),(to_sfixed_a(-0.00011414787877583876)),(to_sfixed_a(-2.1615363948512822e-05)),(to_sfixed_a(0.00022271972557064146)),(to_sfixed_a(-0.00015828940377105027)),(to_sfixed_a(0.000252982834354043)),(to_sfixed_a(6.922498869244009e-05)),(to_sfixed_a(-5.838979996042326e-05)),(to_sfixed_a(8.580250869272277e-05)),(to_sfixed_a(0.00013986359408590943)),(to_sfixed_a(0.0002793018938973546)),(to_sfixed_a(-7.160683162510395e-05)),(to_sfixed_a(-0.0001305319310631603)),(to_sfixed_a(0.00023812480503693223)),(to_sfixed_a(0.00014968356117606163)),(to_sfixed_a(-0.00010195114009547979)),(to_sfixed_a(-7.060374628053978e-05)),(to_sfixed_a(0.0001993879850488156)),(to_sfixed_a(-0.0002966249012388289)),(to_sfixed_a(-1.5336176147684455e-05)),(to_sfixed_a(-0.00041099078953266144)),(to_sfixed_a(0.0003776072117034346)),(to_sfixed_a(0.0001564388512633741)),(to_sfixed_a(-2.98367376672104e-05)),(to_sfixed_a(7.889913831604645e-05)),(to_sfixed_a(-8.639643783681095e-05)),(to_sfixed_a(0.0002193348773289472)),(to_sfixed_a(-0.0002209107915405184)),(to_sfixed_a(0.00015730716404505074)),(to_sfixed_a(-0.00016907989629544318)),(to_sfixed_a(5.352085281629115e-06)),(to_sfixed_a(1.7046782886609435e-05)),(to_sfixed_a(4.877030005445704e-05)),(to_sfixed_a(-4.337416248745285e-05)),(to_sfixed_a(-6.578141619684175e-05)),(to_sfixed_a(-0.0002170681400457397)),(to_sfixed_a(0.00015537533909082413)),(to_sfixed_a(4.5665205107070506e-05)),(to_sfixed_a(0.0002741919597610831)),(to_sfixed_a(0.0003049323568120599)),(to_sfixed_a(-5.773820885224268e-05)),(to_sfixed_a(-1.2217205949127674e-06)),(to_sfixed_a(7.991614256752655e-05)),(to_sfixed_a(-1.1926858860533684e-05)),(to_sfixed_a(-0.0002172531239921227)),(to_sfixed_a(3.971249680034816e-05)),(to_sfixed_a(-0.00011424170224927366)),(to_sfixed_a(-0.00019080484344158322)),(to_sfixed_a(-2.891496114898473e-05)),(to_sfixed_a(-3.076918073929846e-05)),(to_sfixed_a(-0.00037875340785831213)),(to_sfixed_a(8.230510866269469e-05)),(to_sfixed_a(5.1448434533085674e-05)),(to_sfixed_a(0.0002970660862047225)),(to_sfixed_a(0.00024192448472604156)),(to_sfixed_a(-9.784262510947883e-05)),(to_sfixed_a(-0.00014240659947972745)),(to_sfixed_a(-4.16113471146673e-06)),(to_sfixed_a(7.059339986881241e-05)),(to_sfixed_a(3.687491698656231e-07)),(to_sfixed_a(-0.0001136457285610959)),(to_sfixed_a(-5.850371962878853e-06)),(to_sfixed_a(-6.137811578810215e-05)),(to_sfixed_a(0.00015943715698085725)),(to_sfixed_a(3.310990723548457e-05)),(to_sfixed_a(8.66283371578902e-05)),(to_sfixed_a(5.964328011032194e-05)),(to_sfixed_a(0.00041391560807824135)),(to_sfixed_a(6.431622023228556e-05)),(to_sfixed_a(-7.063017983455211e-05)),(to_sfixed_a(-4.080160579178482e-06)),(to_sfixed_a(-0.00014192222442943603)),(to_sfixed_a(-0.00028007946093566716)),(to_sfixed_a(0.000306333793560043)),(to_sfixed_a(1.8751306924968958e-06)),(to_sfixed_a(-1.1209220247110352e-05)),(to_sfixed_a(-2.282725108671002e-05)),(to_sfixed_a(-0.00018858778639696538)),(to_sfixed_a(-1.0888905308092944e-05)),(to_sfixed_a(-0.0001765812048688531)),(to_sfixed_a(0.00016570906154811382)),(to_sfixed_a(0.00010320820729248226)),(to_sfixed_a(-0.0001130359378294088)),(to_sfixed_a(0.00013737489643972367)),(to_sfixed_a(-0.00010701817518565804)),(to_sfixed_a(0.00023769179824739695)),(to_sfixed_a(6.111571565270424e-05)),(to_sfixed_a(-0.00016799740842543542)),(to_sfixed_a(-0.0001016385795082897)),(to_sfixed_a(3.78317927243188e-05)),(to_sfixed_a(0.00020387755648698658)),(to_sfixed_a(6.778151873731986e-05)),(to_sfixed_a(-0.00023650257207918912)),(to_sfixed_a(0.00011295151489321142)),(to_sfixed_a(-8.456901559839025e-05)),(to_sfixed_a(6.0215410485398024e-05)),(to_sfixed_a(0.00027023901930078864)),(to_sfixed_a(-0.0003796291712205857)),(to_sfixed_a(0.0001566567225381732)),(to_sfixed_a(6.48364657536149e-05)),(to_sfixed_a(-0.0004475715395528823)),(to_sfixed_a(-0.0004511058214120567)),(to_sfixed_a(1.834895374486223e-05)),(to_sfixed_a(-2.2591266315430403e-06)),(to_sfixed_a(-5.8312863984610885e-05)),(to_sfixed_a(6.259114161366597e-05)),(to_sfixed_a(-6.820631824666634e-05)),(to_sfixed_a(-7.875292067183182e-05)),(to_sfixed_a(-3.531946276780218e-05)),(to_sfixed_a(-0.00011610927322180942)),(to_sfixed_a(-6.274945189943537e-05)),(to_sfixed_a(-6.827813922427595e-05)),(to_sfixed_a(3.6579524021362886e-05)),(to_sfixed_a(0.00023497849178966135)),(to_sfixed_a(0.00018426190945319831)),(to_sfixed_a(-0.00011207375791855156)),(to_sfixed_a(-8.708775567356497e-08)),(to_sfixed_a(9.343784768134356e-08)),(to_sfixed_a(-1.2574739230331033e-05)),(to_sfixed_a(-0.00015473528765141964)),(to_sfixed_a(-0.00030482670990750194)),(to_sfixed_a(-3.11750773107633e-06)),(to_sfixed_a(-5.039482130086981e-05)),(to_sfixed_a(4.60985247627832e-05)),(to_sfixed_a(0.0002869424642995)),(to_sfixed_a(5.6812270486261696e-05)),(to_sfixed_a(0.00024388672318309546)),(to_sfixed_a(-0.00015927344793453813)),(to_sfixed_a(-4.509113568929024e-05)),(to_sfixed_a(0.00011393496242817491)),(to_sfixed_a(-0.0003821327700279653)),(to_sfixed_a(-0.0002214340347563848)),(to_sfixed_a(2.375073017901741e-05)),(to_sfixed_a(9.487002535024658e-05)),(to_sfixed_a(-7.102621748344973e-05)),(to_sfixed_a(-0.00019268014875706285)),(to_sfixed_a(-0.0001843368954723701)),(to_sfixed_a(-5.7136581744998693e-05)),(to_sfixed_a(-5.706944648409262e-05)),(to_sfixed_a(-1.0536734407651238e-05)),(to_sfixed_a(-0.00020436802878975868)),(to_sfixed_a(0.00011676319991238415)),(to_sfixed_a(-4.3833948438987136e-05)),(to_sfixed_a(-3.3117845305241644e-05)),(to_sfixed_a(-0.0002507091558072716)),(to_sfixed_a(0.00013708836922887713)),(to_sfixed_a(-5.821811646455899e-05)),(to_sfixed_a(-0.00019875170255545527)),(to_sfixed_a(-0.0001329329825239256)),(to_sfixed_a(-0.00018101930618286133)),(to_sfixed_a(0.0003132063720840961)),(to_sfixed_a(-4.604662171914242e-05)),(to_sfixed_a(-0.00024098341236822307)),(to_sfixed_a(5.079348193248734e-05)),(to_sfixed_a(-0.00013731957005802542)),(to_sfixed_a(6.945956556592137e-05)),(to_sfixed_a(0.00024660181952640414)),(to_sfixed_a(-0.00030511562363244593)),(to_sfixed_a(-6.873606616863981e-05)),(to_sfixed_a(6.508601654786617e-05)),(to_sfixed_a(5.1742972573265433e-08)),(to_sfixed_a(4.290704964660108e-07)),(to_sfixed_a(3.2759409805294126e-05)),(to_sfixed_a(0.00021998226293362677)),(to_sfixed_a(-2.305013913428411e-05)),(to_sfixed_a(-0.0002923218999058008)),(to_sfixed_a(-2.284030051669106e-05)),(to_sfixed_a(-0.00013672737986780703)),(to_sfixed_a(-6.245528493309394e-05)),(to_sfixed_a(-0.00010864966316148639)),(to_sfixed_a(6.267438584472984e-05)),(to_sfixed_a(-0.00019124700338579714)),(to_sfixed_a(1.956555206561461e-05)),(to_sfixed_a(-6.967002991586924e-05)),(to_sfixed_a(-0.00024766867863945663)),(to_sfixed_a(0.0001580747775733471)),(to_sfixed_a(7.780094165354967e-06)),(to_sfixed_a(-7.544511754531413e-05)),(to_sfixed_a(4.714121678262018e-05)),(to_sfixed_a(0.00038511023740284145)),(to_sfixed_a(0.00015178814646787941)),(to_sfixed_a(3.584354999475181e-06)),(to_sfixed_a(0.0002150968211935833)),(to_sfixed_a(-1.5684054233133793e-07)),(to_sfixed_a(-0.000129492866108194)),(to_sfixed_a(-0.00030545939807780087)),(to_sfixed_a(-0.00017466314602643251)),(to_sfixed_a(0.00011192054080311209)),(to_sfixed_a(2.198667061747983e-07)),(to_sfixed_a(5.980227069812827e-05)),(to_sfixed_a(-0.00029030669247731566)),(to_sfixed_a(-0.00016707685426808894)),(to_sfixed_a(7.43759810575284e-05)),(to_sfixed_a(-0.00029460040968842804)),(to_sfixed_a(-6.0251310060266405e-05)),(to_sfixed_a(0.0001689615601208061)),(to_sfixed_a(6.401113932952285e-05)),(to_sfixed_a(0.00011298392928438261)),(to_sfixed_a(-2.184387994930148e-06)),(to_sfixed_a(0.0001270273351110518)),(to_sfixed_a(-5.5841559515101835e-05)),(to_sfixed_a(1.0325617040507495e-05)),(to_sfixed_a(-0.0001668372133281082)),(to_sfixed_a(-1.528080611024052e-05)),(to_sfixed_a(-0.00010777503484860063)),(to_sfixed_a(-3.5184348234906793e-06)),(to_sfixed_a(-0.0003005088656209409)),(to_sfixed_a(-0.0002756146132014692)),(to_sfixed_a(-0.0002980824501719326)),(to_sfixed_a(4.7457935579586774e-05)),(to_sfixed_a(-0.00011427610297687352)),(to_sfixed_a(2.9258430004119873e-05)),(to_sfixed_a(0.00011884467676281929)),(to_sfixed_a(0.00013241672422736883)),(to_sfixed_a(0.00012840703129768372)),(to_sfixed_a(-0.00010377381113357842)),(to_sfixed_a(-0.00020298815798014402)),(to_sfixed_a(-3.9388047298416495e-05)),(to_sfixed_a(0.0001679689739830792)),(to_sfixed_a(0.0001584849233040586)),(to_sfixed_a(-0.00016665158909745514)),(to_sfixed_a(0.00017060444224625826)),(to_sfixed_a(-1.0789372026920319e-06)),(to_sfixed_a(5.5720047384966165e-05)),(to_sfixed_a(4.1895429603755474e-05)),(to_sfixed_a(1.787279143172782e-05)),(to_sfixed_a(-2.2146634364617057e-05)),(to_sfixed_a(-1.1390955478418618e-05)),(to_sfixed_a(-0.00014822956291027367)),(to_sfixed_a(0.0001686706964392215)),(to_sfixed_a(-0.00016133402823470533)),(to_sfixed_a(-8.109891496133059e-07)),(to_sfixed_a(-2.4030716303968802e-05)),(to_sfixed_a(7.144617848098278e-05)),(to_sfixed_a(2.317547841812484e-05)),(to_sfixed_a(-0.00015654046728741378)),(to_sfixed_a(7.342911703744903e-05)),(to_sfixed_a(0.00016250165936071426)),(to_sfixed_a(-5.188251088839024e-05)),(to_sfixed_a(-0.00011641602031886578)),(to_sfixed_a(3.263326652813703e-05)),(to_sfixed_a(0.00010028201359091327)),(to_sfixed_a(0.00022905250079929829)),(to_sfixed_a(0.00011268363596173003)),(to_sfixed_a(0.00014951961929909885)),(to_sfixed_a(-2.320075873285532e-05)),(to_sfixed_a(-7.95236264821142e-05)),(to_sfixed_a(-8.910530596040189e-05)),(to_sfixed_a(-0.0002453152264934033)),(to_sfixed_a(3.5582655982580036e-05)),(to_sfixed_a(0.0001647969038458541)),(to_sfixed_a(-0.00011893654300365597)),(to_sfixed_a(0.00021457027469296008)),(to_sfixed_a(0.0001899976487038657)),(to_sfixed_a(-8.948370668804273e-05)),(to_sfixed_a(0.00044479206553660333)),(to_sfixed_a(3.878996358253062e-05)),(to_sfixed_a(0.00012230062566231936)),(to_sfixed_a(4.864639777224511e-06)),(to_sfixed_a(0.00030027629691176116)),(to_sfixed_a(-9.123874770011753e-05)),(to_sfixed_a(6.636149191763252e-05)),(to_sfixed_a(-1.9972749214502983e-05)),(to_sfixed_a(-0.00011681742034852505)),(to_sfixed_a(-1.1650387023109943e-05)),(to_sfixed_a(-0.00012722982501145452)),(to_sfixed_a(0.0002928077010437846)),(to_sfixed_a(-0.0001661409914959222)),(to_sfixed_a(0.00015738379443064332)),(to_sfixed_a(-6.262330862227827e-05)),(to_sfixed_a(7.069025014061481e-05)),(to_sfixed_a(-6.766855221940205e-05)),(to_sfixed_a(-0.00015166381490416825)),(to_sfixed_a(-0.00014561551506631076)),(to_sfixed_a(2.5144880055449903e-05)),(to_sfixed_a(4.4800595787819475e-05)),(to_sfixed_a(2.5625500711612403e-05)),(to_sfixed_a(4.314687248552218e-05)),(to_sfixed_a(0.00015623973740730435)),(to_sfixed_a(3.294059570180252e-05)),(to_sfixed_a(-0.0002573792007751763)),(to_sfixed_a(-0.00010565005504759029)),(to_sfixed_a(-0.00012957362923771143)),(to_sfixed_a(-6.462071905843914e-05)),(to_sfixed_a(-0.00014723515778314322)),(to_sfixed_a(-0.00013050198322162032)),(to_sfixed_a(-5.107604374643415e-05)),(to_sfixed_a(-0.000187645127880387)));

    constant weight_n2_67 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.018768737092614174)),(to_sfixed_a(0.0058620041236281395)),(to_sfixed_a(-0.227173313498497)),(to_sfixed_a(-6.900053995195776e-05)),(to_sfixed_a(-0.00317795155569911)),(to_sfixed_a(0.00042391757597215474)),(to_sfixed_a(-0.0036912139039486647)),(to_sfixed_a(6.928792572580278e-06)),(to_sfixed_a(1.083263850887306e-05)),(to_sfixed_a(6.528032827191055e-05)),(to_sfixed_a(9.393460641149431e-05)),(to_sfixed_a(-0.0004958901554346085)),(to_sfixed_a(0.000287980365101248)),(to_sfixed_a(-0.0032456570770591497)),(to_sfixed_a(-1.740917650749907e-05)),(to_sfixed_a(-0.0002392241731286049)),(to_sfixed_a(0.20012317597866058)),(to_sfixed_a(-0.0002915227669291198)),(to_sfixed_a(0.1623273491859436)),(to_sfixed_a(-0.0013095058966428041)),(to_sfixed_a(0.00023845906252972782)),(to_sfixed_a(0.0002515811356715858)),(to_sfixed_a(0.0006912383250892162)),(to_sfixed_a(0.00040838008862920105)),(to_sfixed_a(-0.008771664462983608)),(to_sfixed_a(0.3378383219242096)),(to_sfixed_a(0.00010985043627442792)),(to_sfixed_a(0.000679382064845413)),(to_sfixed_a(5.5437954870285466e-05)),(to_sfixed_a(-0.00011588783672777936)),(to_sfixed_a(0.12771232426166534)),(to_sfixed_a(0.00010579702939139679)),(to_sfixed_a(0.010240352712571621)),(to_sfixed_a(-2.5067958631552756e-05)),(to_sfixed_a(-0.00012764048005919904)),(to_sfixed_a(-0.00018466226174496114)),(to_sfixed_a(0.23937951028347015)),(to_sfixed_a(0.016132568940520287)),(to_sfixed_a(0.0009732822072692215)),(to_sfixed_a(0.00015533748955931515)),(to_sfixed_a(-0.15930438041687012)),(to_sfixed_a(-0.0010877971071749926)),(to_sfixed_a(-0.0001812674745451659)),(to_sfixed_a(-9.989844329538755e-06)),(to_sfixed_a(-0.000449911633040756)),(to_sfixed_a(0.16452158987522125)),(to_sfixed_a(-0.0012349422322586179)),(to_sfixed_a(-0.006116847507655621)),(to_sfixed_a(-0.00018330762395635247)),(to_sfixed_a(-0.24620378017425537)),(to_sfixed_a(-0.0002888780436478555)),(to_sfixed_a(-0.0005964648444205523)),(to_sfixed_a(-4.039478881168179e-06)),(to_sfixed_a(-0.0012793107889592648)),(to_sfixed_a(-0.0020491264294832945)),(to_sfixed_a(-0.002696490380913019)),(to_sfixed_a(-0.00031028533703647554)),(to_sfixed_a(-0.3670267164707184)),(to_sfixed_a(0.00010002800263464451)),(to_sfixed_a(-4.403836283017881e-05)),(to_sfixed_a(0.00439379783347249)),(to_sfixed_a(0.13677643239498138)),(to_sfixed_a(0.0006268125725910068)),(to_sfixed_a(0.3648611903190613)),(to_sfixed_a(4.173125489614904e-07)),(to_sfixed_a(0.000177523004822433)),(to_sfixed_a(9.408795449417084e-07)),(to_sfixed_a(-0.27671903371810913)),(to_sfixed_a(-0.462368369102478)),(to_sfixed_a(0.0003043293545488268)),(to_sfixed_a(0.0028758139815181494)),(to_sfixed_a(-0.008726630359888077)),(to_sfixed_a(-0.0041144536808133125)),(to_sfixed_a(0.00010967137495754287)),(to_sfixed_a(1.9409133528824896e-05)),(to_sfixed_a(1.0951385775115341e-05)),(to_sfixed_a(-0.0007228718022815883)),(to_sfixed_a(-0.0010571556631475687)),(to_sfixed_a(0.00010669017501641065)),(to_sfixed_a(0.0066507053561508656)),(to_sfixed_a(-0.005592638161033392)),(to_sfixed_a(-0.00018368710880167782)),(to_sfixed_a(-0.001390698365867138)),(to_sfixed_a(0.4239853620529175)),(to_sfixed_a(-5.62022250960581e-05)),(to_sfixed_a(-0.008232778869569302)),(to_sfixed_a(-9.710356971481815e-05)),(to_sfixed_a(0.0004650001064874232)),(to_sfixed_a(-1.9495208107400686e-05)),(to_sfixed_a(-7.484428351745009e-06)),(to_sfixed_a(-0.08286137133836746)),(to_sfixed_a(-0.00011751792044378817)),(to_sfixed_a(-0.004626184701919556)),(to_sfixed_a(-6.845211464678869e-05)),(to_sfixed_a(0.0007734441314823925)),(to_sfixed_a(0.00010958432540064678)),(to_sfixed_a(2.9713744879700243e-05)),(to_sfixed_a(-2.6326692022848874e-05)),(to_sfixed_a(0.00018347047443967313)),(to_sfixed_a(5.861031240783632e-06)),(to_sfixed_a(-0.0026126601733267307)),(to_sfixed_a(-0.0008031127508729696)),(to_sfixed_a(0.00012812591739930212)),(to_sfixed_a(0.009328910149633884)),(to_sfixed_a(0.08458968251943588)),(to_sfixed_a(-0.003599474672228098)),(to_sfixed_a(-0.00011165507748955861)),(to_sfixed_a(6.818637484684587e-05)),(to_sfixed_a(0.00011206404451513663)),(to_sfixed_a(-0.003050764324143529)),(to_sfixed_a(-0.002831777324900031)),(to_sfixed_a(0.0004503463860601187)),(to_sfixed_a(0.32786351442337036)),(to_sfixed_a(-3.720878157764673e-05)),(to_sfixed_a(7.245377491926774e-05)),(to_sfixed_a(0.0052751884795725346)),(to_sfixed_a(0.006492132321000099)),(to_sfixed_a(-0.0014073867350816727)),(to_sfixed_a(1.804545900085941e-05)),(to_sfixed_a(0.005792503245174885)),(to_sfixed_a(0.00013714280794374645)),(to_sfixed_a(7.056893809931353e-05)),(to_sfixed_a(-0.0009197630570270121)),(to_sfixed_a(6.689805741189048e-05)),(to_sfixed_a(3.0060677090659738e-05)),(to_sfixed_a(0.0002334045566385612)),(to_sfixed_a(0.0029755043797194958)),(to_sfixed_a(-0.00011443662515375763)),(to_sfixed_a(-0.00017922029655892402)),(to_sfixed_a(-3.451141674304381e-05)),(to_sfixed_a(5.240253813099116e-06)),(to_sfixed_a(1.1635671398835257e-05)),(to_sfixed_a(0.006957840174436569)),(to_sfixed_a(0.0003602424985729158)),(to_sfixed_a(0.00014806445688009262)),(to_sfixed_a(-4.6472523536067456e-05)),(to_sfixed_a(-0.458223432302475)),(to_sfixed_a(-0.3803183138370514)),(to_sfixed_a(1.9296070604468696e-05)),(to_sfixed_a(0.00026963657001033425)),(to_sfixed_a(0.008564909920096397)),(to_sfixed_a(0.00010774573456728831)),(to_sfixed_a(-0.00014598631241824478)),(to_sfixed_a(0.0001165691064670682)),(to_sfixed_a(0.0011223435867577791)),(to_sfixed_a(0.0002373642782913521)),(to_sfixed_a(-0.0020731198601424694)),(to_sfixed_a(0.00015752892068121582)),(to_sfixed_a(-6.478876457549632e-06)),(to_sfixed_a(0.005163389258086681)),(to_sfixed_a(0.00016699508705642074)),(to_sfixed_a(-8.806315599940717e-05)),(to_sfixed_a(0.011429434642195702)),(to_sfixed_a(-0.00016546309052500874)),(to_sfixed_a(-4.110993177164346e-05)),(to_sfixed_a(0.007498462684452534)),(to_sfixed_a(6.397676770575345e-07)),(to_sfixed_a(-0.0023738353047519922)),(to_sfixed_a(-4.19962962041609e-05)),(to_sfixed_a(-6.075177589082159e-05)),(to_sfixed_a(-1.8156017176806927e-05)),(to_sfixed_a(-9.03757827472873e-05)),(to_sfixed_a(0.0011313938302919269)),(to_sfixed_a(-0.004690167959779501)),(to_sfixed_a(0.0020852016750723124)),(to_sfixed_a(0.23665757477283478)),(to_sfixed_a(4.727357008960098e-05)),(to_sfixed_a(-0.5525032877922058)),(to_sfixed_a(-6.172920984681696e-05)),(to_sfixed_a(5.658692680299282e-05)),(to_sfixed_a(0.150405615568161)),(to_sfixed_a(0.24778710305690765)),(to_sfixed_a(-0.0003680000372696668)),(to_sfixed_a(-2.5255143555114046e-05)),(to_sfixed_a(-0.427401065826416)),(to_sfixed_a(-0.00045930349733680487)),(to_sfixed_a(-0.0011339980410411954)),(to_sfixed_a(-0.0004067165427841246)),(to_sfixed_a(-0.06889329850673676)),(to_sfixed_a(-0.0026817063335329294)),(to_sfixed_a(-0.0024067938793450594)),(to_sfixed_a(0.01626516878604889)),(to_sfixed_a(-0.00032168274628929794)),(to_sfixed_a(0.0001791691465768963)),(to_sfixed_a(0.00011275420547463)),(to_sfixed_a(-0.010120815597474575)),(to_sfixed_a(0.22734999656677246)),(to_sfixed_a(-0.001195372431538999)),(to_sfixed_a(0.000691224355250597)),(to_sfixed_a(-0.0015214710729196668)),(to_sfixed_a(0.00010116385237779468)),(to_sfixed_a(-0.0002766994875855744)),(to_sfixed_a(0.23881906270980835)),(to_sfixed_a(-0.1908724009990692)),(to_sfixed_a(-8.81175947142765e-06)),(to_sfixed_a(0.0002039847313426435)),(to_sfixed_a(1.049692218657583e-05)),(to_sfixed_a(0.31171637773513794)),(to_sfixed_a(-0.019968457520008087)),(to_sfixed_a(-2.619758015498519e-05)),(to_sfixed_a(-4.496147812460549e-05)),(to_sfixed_a(1.173109922092408e-05)),(to_sfixed_a(-0.00018684726092033088)),(to_sfixed_a(0.0001147485600085929)),(to_sfixed_a(0.000105122038803529)),(to_sfixed_a(0.001255081151612103)),(to_sfixed_a(0.0001478111371397972)),(to_sfixed_a(-0.5737327933311462)),(to_sfixed_a(-0.36816269159317017)),(to_sfixed_a(-0.301445335149765)),(to_sfixed_a(-0.0022047844249755144)),(to_sfixed_a(-0.00015352238551713526)),(to_sfixed_a(0.00013568345457315445)),(to_sfixed_a(-1.2001401046290994e-06)),(to_sfixed_a(1.9103805243503302e-05)),(to_sfixed_a(0.00032566607114858925)),(to_sfixed_a(0.0023720215540379286)),(to_sfixed_a(0.002284080721437931)),(to_sfixed_a(-0.36676743626594543)),(to_sfixed_a(-6.508986552944407e-05)),(to_sfixed_a(-5.4159496357897297e-05)),(to_sfixed_a(-0.0002278934116475284)),(to_sfixed_a(-1.0754763934528455e-05)),(to_sfixed_a(0.001654263585805893)),(to_sfixed_a(0.3930896818637848)),(to_sfixed_a(0.00015821527631487697)),(to_sfixed_a(-3.2336381991626695e-05)),(to_sfixed_a(3.3956759580178186e-05)),(to_sfixed_a(0.29969656467437744)),(to_sfixed_a(-0.2960550785064697)),(to_sfixed_a(0.0011665369383990765)),(to_sfixed_a(2.1014129742980003e-06)),(to_sfixed_a(-4.969180736225098e-06)),(to_sfixed_a(-0.00011439326772233471)),(to_sfixed_a(-0.00043596926843747497)),(to_sfixed_a(0.02151252143085003)),(to_sfixed_a(-9.280195081373677e-05)),(to_sfixed_a(6.106216460466385e-05)),(to_sfixed_a(9.17181750992313e-05)),(to_sfixed_a(-1.414847793057561e-05)),(to_sfixed_a(0.39249569177627563)),(to_sfixed_a(8.060159598244354e-05)),(to_sfixed_a(0.003424422349780798)),(to_sfixed_a(-1.0742478480096906e-05)),(to_sfixed_a(-0.007304946891963482)),(to_sfixed_a(-0.00013417258742265403)),(to_sfixed_a(0.0557694211602211)),(to_sfixed_a(0.0004613028431776911)),(to_sfixed_a(-0.00018168975657317787)),(to_sfixed_a(0.0034267345909029245)),(to_sfixed_a(-0.012925758957862854)),(to_sfixed_a(-0.00023651070659980178)),(to_sfixed_a(-5.2467617933871225e-05)),(to_sfixed_a(5.87801041547209e-05)),(to_sfixed_a(0.005437040701508522)),(to_sfixed_a(0.0015131820691749454)),(to_sfixed_a(-0.009910853579640388)),(to_sfixed_a(-6.552260310854763e-05)),(to_sfixed_a(0.00014914826897438616)),(to_sfixed_a(-0.0026597394607961178)),(to_sfixed_a(3.193523662048392e-05)),(to_sfixed_a(-0.0017283596098423004)),(to_sfixed_a(-5.80345731577836e-05)),(to_sfixed_a(-0.0013711097417399287)),(to_sfixed_a(0.00023740969481877983)),(to_sfixed_a(-0.010636309161782265)),(to_sfixed_a(2.523025978007354e-05)),(to_sfixed_a(-6.654839671682566e-05)),(to_sfixed_a(0.00017360845231451094)),(to_sfixed_a(0.002521627815440297)),(to_sfixed_a(-0.003365106415003538)),(to_sfixed_a(6.678879435639828e-05)),(to_sfixed_a(0.00024421184207312763)),(to_sfixed_a(-0.00024367606965824962)),(to_sfixed_a(6.327367736957967e-05)),(to_sfixed_a(0.00925865676254034)),(to_sfixed_a(-0.008807804435491562)),(to_sfixed_a(-0.0007052121218293905)),(to_sfixed_a(-0.007165734656155109)),(to_sfixed_a(0.0011518375249579549)),(to_sfixed_a(4.578045627567917e-05)),(to_sfixed_a(-0.0003088662924710661)),(to_sfixed_a(6.253930041566491e-05)),(to_sfixed_a(0.018904242664575577)),(to_sfixed_a(-0.00027576505090110004)),(to_sfixed_a(2.5555487809469923e-05)),(to_sfixed_a(-0.061293620616197586)),(to_sfixed_a(0.17152734100818634)),(to_sfixed_a(0.0001055059110512957)),(to_sfixed_a(-0.0006138097960501909)),(to_sfixed_a(-0.0005928806494921446)),(to_sfixed_a(0.3051016330718994)),(to_sfixed_a(-0.1436815708875656)),(to_sfixed_a(-0.00015216306201182306)),(to_sfixed_a(-0.002074396936222911)),(to_sfixed_a(0.0014482589904218912)),(to_sfixed_a(-0.012983767315745354)),(to_sfixed_a(3.039046350750141e-05)),(to_sfixed_a(-0.00192259659525007)),(to_sfixed_a(0.0005963699659332633)),(to_sfixed_a(-0.0027946163900196552)));

    constant weight_n2_68 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.16064637899398804)),(to_sfixed_a(0.0003749360330402851)),(to_sfixed_a(0.001825879793614149)),(to_sfixed_a(0.0001622883282834664)),(to_sfixed_a(-0.0003264980623498559)),(to_sfixed_a(5.0764378102030605e-05)),(to_sfixed_a(0.004762684460729361)),(to_sfixed_a(4.6398810809478164e-05)),(to_sfixed_a(-0.00010095354082295671)),(to_sfixed_a(0.00018737393838819116)),(to_sfixed_a(0.00015055114636197686)),(to_sfixed_a(0.005672133527696133)),(to_sfixed_a(6.019206921337172e-06)),(to_sfixed_a(-0.011985759250819683)),(to_sfixed_a(6.336237129289657e-05)),(to_sfixed_a(-0.0002199753507738933)),(to_sfixed_a(0.0030711479485034943)),(to_sfixed_a(6.54981704428792e-05)),(to_sfixed_a(-0.3827626705169678)),(to_sfixed_a(0.00017348365508951247)),(to_sfixed_a(0.00010649923206074163)),(to_sfixed_a(-0.00028234237106516957)),(to_sfixed_a(-9.800177213037387e-05)),(to_sfixed_a(2.4279026547446847e-05)),(to_sfixed_a(-0.018995316699147224)),(to_sfixed_a(0.00023926369613036513)),(to_sfixed_a(0.00026968930615112185)),(to_sfixed_a(-0.00041184856672771275)),(to_sfixed_a(0.0004773661494255066)),(to_sfixed_a(0.00015051671653054655)),(to_sfixed_a(0.003107902593910694)),(to_sfixed_a(6.25846951152198e-05)),(to_sfixed_a(0.003739945823326707)),(to_sfixed_a(0.00014810920401941985)),(to_sfixed_a(0.0001347191573586315)),(to_sfixed_a(6.298976950347424e-05)),(to_sfixed_a(-0.029479756951332092)),(to_sfixed_a(0.0006471263477578759)),(to_sfixed_a(0.010911926627159119)),(to_sfixed_a(-2.109894558088854e-05)),(to_sfixed_a(0.002326009562239051)),(to_sfixed_a(-0.010753149166703224)),(to_sfixed_a(-0.00015646680549252778)),(to_sfixed_a(-9.753467747941613e-05)),(to_sfixed_a(0.009141982533037663)),(to_sfixed_a(0.014823938719928265)),(to_sfixed_a(0.0010550011647865176)),(to_sfixed_a(0.0070382533594965935)),(to_sfixed_a(6.794153887312859e-05)),(to_sfixed_a(-0.00045626884093508124)),(to_sfixed_a(-0.0045704604126513)),(to_sfixed_a(0.0006186259561218321)),(to_sfixed_a(-0.00015327607979997993)),(to_sfixed_a(-0.0011914529604837298)),(to_sfixed_a(0.0044516162015497684)),(to_sfixed_a(0.0015913434326648712)),(to_sfixed_a(-0.0001544467086205259)),(to_sfixed_a(0.014528443105518818)),(to_sfixed_a(-0.00022374774562194943)),(to_sfixed_a(0.00017442082753404975)),(to_sfixed_a(0.00786147452890873)),(to_sfixed_a(0.0012621720088645816)),(to_sfixed_a(-0.0006961353938095272)),(to_sfixed_a(0.005751060787588358)),(to_sfixed_a(5.608690116787329e-05)),(to_sfixed_a(0.0008212840184569359)),(to_sfixed_a(-0.00016876182053238153)),(to_sfixed_a(-0.0011210101656615734)),(to_sfixed_a(0.007510931696742773)),(to_sfixed_a(-1.2549542589113116e-05)),(to_sfixed_a(0.010363386943936348)),(to_sfixed_a(0.014261444099247456)),(to_sfixed_a(0.001460682600736618)),(to_sfixed_a(0.000126411541714333)),(to_sfixed_a(-9.622928337194026e-05)),(to_sfixed_a(-0.0002863455156330019)),(to_sfixed_a(0.011394539847970009)),(to_sfixed_a(0.005002275109291077)),(to_sfixed_a(-6.599484186153859e-05)),(to_sfixed_a(0.0009872500086203218)),(to_sfixed_a(0.008817227557301521)),(to_sfixed_a(9.154609870165586e-07)),(to_sfixed_a(0.28597214818000793)),(to_sfixed_a(-0.009399449452757835)),(to_sfixed_a(-1.4350674973684363e-05)),(to_sfixed_a(0.0005616131238639355)),(to_sfixed_a(-0.005110196303576231)),(to_sfixed_a(0.00015263208479154855)),(to_sfixed_a(-0.0001546737621538341)),(to_sfixed_a(-0.00015149317914620042)),(to_sfixed_a(0.010897470638155937)),(to_sfixed_a(-0.00010003217903431505)),(to_sfixed_a(0.009514815174043179)),(to_sfixed_a(-0.00029321512556634843)),(to_sfixed_a(0.0029083574190735817)),(to_sfixed_a(-0.0004180604009889066)),(to_sfixed_a(-1.386128133162856e-06)),(to_sfixed_a(-0.0002470386680215597)),(to_sfixed_a(0.00010753805690910667)),(to_sfixed_a(-6.898125138832256e-05)),(to_sfixed_a(0.00014885740529280156)),(to_sfixed_a(0.006159014999866486)),(to_sfixed_a(0.00016872193373274058)),(to_sfixed_a(0.00707531813532114)),(to_sfixed_a(0.009208261966705322)),(to_sfixed_a(0.00033649595570750535)),(to_sfixed_a(5.839435107191093e-05)),(to_sfixed_a(-9.836880781222135e-05)),(to_sfixed_a(0.00016712755314074457)),(to_sfixed_a(0.005739902146160603)),(to_sfixed_a(0.003027903148904443)),(to_sfixed_a(-0.00011624998296611011)),(to_sfixed_a(0.004954407457262278)),(to_sfixed_a(-0.00019048296962864697)),(to_sfixed_a(7.102305971784517e-05)),(to_sfixed_a(0.0009190295822918415)),(to_sfixed_a(1.4923782146070153e-05)),(to_sfixed_a(0.004878317005932331)),(to_sfixed_a(0.000420364027377218)),(to_sfixed_a(0.004739203490316868)),(to_sfixed_a(0.00011617783457040787)),(to_sfixed_a(-9.426493488717824e-05)),(to_sfixed_a(0.007433649152517319)),(to_sfixed_a(8.987673936644569e-05)),(to_sfixed_a(-0.00017350452253594995)),(to_sfixed_a(-0.20775461196899414)),(to_sfixed_a(-0.0011052609188482165)),(to_sfixed_a(-0.00019454091670922935)),(to_sfixed_a(0.00018176648882217705)),(to_sfixed_a(-0.00010922276123892516)),(to_sfixed_a(-7.99732151790522e-05)),(to_sfixed_a(-0.00020037118520122021)),(to_sfixed_a(-0.0008372088195756078)),(to_sfixed_a(0.004976935219019651)),(to_sfixed_a(-0.00015251357399392873)),(to_sfixed_a(-0.00011637775605777279)),(to_sfixed_a(0.025956040248274803)),(to_sfixed_a(0.0011276907753199339)),(to_sfixed_a(5.6966331612784415e-05)),(to_sfixed_a(-6.844159361207858e-05)),(to_sfixed_a(0.002953980816528201)),(to_sfixed_a(-4.480571078602225e-06)),(to_sfixed_a(5.888981104362756e-05)),(to_sfixed_a(3.973461571149528e-05)),(to_sfixed_a(0.0009322295081801713)),(to_sfixed_a(-3.121140252915211e-05)),(to_sfixed_a(-0.00014312288840301335)),(to_sfixed_a(-1.6037294699344784e-05)),(to_sfixed_a(-0.00023799158225301653)),(to_sfixed_a(0.010166153311729431)),(to_sfixed_a(-0.00012839461851399392)),(to_sfixed_a(-0.00020572844368871301)),(to_sfixed_a(-4.624690336640924e-05)),(to_sfixed_a(3.845013998216018e-05)),(to_sfixed_a(7.968211866682395e-05)),(to_sfixed_a(0.010313517414033413)),(to_sfixed_a(3.647806806839071e-05)),(to_sfixed_a(0.0012508210493251681)),(to_sfixed_a(-0.0001812463451642543)),(to_sfixed_a(0.00018072778766509145)),(to_sfixed_a(0.0001785702770575881)),(to_sfixed_a(3.7369332858361304e-05)),(to_sfixed_a(-0.0007709618657827377)),(to_sfixed_a(0.00036074797390028834)),(to_sfixed_a(-0.001852886052802205)),(to_sfixed_a(-0.00013293520896695554)),(to_sfixed_a(-0.00015333712508436292)),(to_sfixed_a(0.0040413811802864075)),(to_sfixed_a(0.00020041759125888348)),(to_sfixed_a(3.147995812469162e-05)),(to_sfixed_a(-7.614486094098538e-06)),(to_sfixed_a(0.0048147342167794704)),(to_sfixed_a(-0.00010034300794359297)),(to_sfixed_a(0.00010284571908414364)),(to_sfixed_a(0.007763995323330164)),(to_sfixed_a(2.7853853680426255e-05)),(to_sfixed_a(-0.0004349040682427585)),(to_sfixed_a(0.00191610271576792)),(to_sfixed_a(0.001177057740278542)),(to_sfixed_a(0.009230240248143673)),(to_sfixed_a(0.0002735318266786635)),(to_sfixed_a(0.01794537715613842)),(to_sfixed_a(1.8358456145506352e-05)),(to_sfixed_a(0.00024367248988710344)),(to_sfixed_a(3.226862463634461e-05)),(to_sfixed_a(-0.00011901515972567722)),(to_sfixed_a(-0.4760810136795044)),(to_sfixed_a(-0.004511741921305656)),(to_sfixed_a(-0.0071580917574465275)),(to_sfixed_a(-0.009025738574564457)),(to_sfixed_a(-0.007505423855036497)),(to_sfixed_a(-0.00032316124998033047)),(to_sfixed_a(0.005627342499792576)),(to_sfixed_a(0.0074307881295681)),(to_sfixed_a(0.00023593484365846962)),(to_sfixed_a(-0.00036198936868458986)),(to_sfixed_a(-4.086362605448812e-05)),(to_sfixed_a(0.0012052258243784308)),(to_sfixed_a(-0.009807627648115158)),(to_sfixed_a(-0.00010224025027127936)),(to_sfixed_a(1.741227606544271e-07)),(to_sfixed_a(4.225148586556315e-06)),(to_sfixed_a(6.184908124851063e-05)),(to_sfixed_a(0.00015316359349526465)),(to_sfixed_a(0.00017424763063900173)),(to_sfixed_a(-0.0031826950144022703)),(to_sfixed_a(0.00033270561834797263)),(to_sfixed_a(9.85413498710841e-05)),(to_sfixed_a(0.0006688915891572833)),(to_sfixed_a(0.008959806524217129)),(to_sfixed_a(0.007119388319551945)),(to_sfixed_a(-2.4550521629862487e-05)),(to_sfixed_a(2.9228722269181162e-05)),(to_sfixed_a(0.00017391619621776044)),(to_sfixed_a(2.4254273739643395e-05)),(to_sfixed_a(-3.0333438189700246e-05)),(to_sfixed_a(-0.0001485609682276845)),(to_sfixed_a(-0.001755259814672172)),(to_sfixed_a(-0.011425376869738102)),(to_sfixed_a(-4.904113302472979e-05)),(to_sfixed_a(-0.00011663367331493646)),(to_sfixed_a(-7.983700197655708e-05)),(to_sfixed_a(-6.971739639993757e-05)),(to_sfixed_a(0.00010038880282081664)),(to_sfixed_a(0.0074869245290756226)),(to_sfixed_a(2.3975644580787048e-05)),(to_sfixed_a(-6.767128070350736e-05)),(to_sfixed_a(8.300868648802862e-05)),(to_sfixed_a(0.004034625366330147)),(to_sfixed_a(-2.1414962247945368e-08)),(to_sfixed_a(-0.0012100182939320803)),(to_sfixed_a(-4.199970135232434e-06)),(to_sfixed_a(6.816095992689952e-05)),(to_sfixed_a(-7.171102333813906e-05)),(to_sfixed_a(0.0017924611456692219)),(to_sfixed_a(0.0038653675001114607)),(to_sfixed_a(0.010893930681049824)),(to_sfixed_a(-0.00010149664740310982)),(to_sfixed_a(-0.0028673307970166206)),(to_sfixed_a(0.00019413346308283508)),(to_sfixed_a(7.11124885128811e-05)),(to_sfixed_a(0.00014180794823914766)),(to_sfixed_a(0.0009720881935209036)),(to_sfixed_a(-0.00017392158042639494)),(to_sfixed_a(-0.16973675787448883)),(to_sfixed_a(7.835878932382911e-07)),(to_sfixed_a(0.015403573401272297)),(to_sfixed_a(0.30594363808631897)),(to_sfixed_a(0.00019537133630365133)),(to_sfixed_a(0.016639403998851776)),(to_sfixed_a(0.0012278123758733273)),(to_sfixed_a(9.718994260765612e-05)),(to_sfixed_a(-0.00017375044990330935)),(to_sfixed_a(-0.0002238908491563052)),(to_sfixed_a(-4.747927960124798e-05)),(to_sfixed_a(0.013876613229513168)),(to_sfixed_a(-0.016404641792178154)),(to_sfixed_a(-0.0001288278290303424)),(to_sfixed_a(0.00020488556765485555)),(to_sfixed_a(0.0007138578221201897)),(to_sfixed_a(-1.1280979379080236e-05)),(to_sfixed_a(0.0024742495734244585)),(to_sfixed_a(0.00025200884556397796)),(to_sfixed_a(-6.095442586229183e-05)),(to_sfixed_a(0.00028794220997951925)),(to_sfixed_a(2.5021814508363605e-05)),(to_sfixed_a(0.00016067101387307048)),(to_sfixed_a(-0.0001767520880093798)),(to_sfixed_a(-7.356443529715762e-05)),(to_sfixed_a(0.004488943610340357)),(to_sfixed_a(-0.027806589379906654)),(to_sfixed_a(-8.499543037032709e-05)),(to_sfixed_a(5.2531337132677436e-05)),(to_sfixed_a(0.00010460095654707402)),(to_sfixed_a(-3.085161733906716e-05)),(to_sfixed_a(-2.279003820149228e-05)),(to_sfixed_a(-0.0015590903349220753)),(to_sfixed_a(0.003911648411303759)),(to_sfixed_a(0.5053724646568298)),(to_sfixed_a(0.0003488787333481014)),(to_sfixed_a(7.097366324160248e-05)),(to_sfixed_a(3.670441219583154e-05)),(to_sfixed_a(5.6084973039105535e-06)),(to_sfixed_a(0.0004099197976756841)),(to_sfixed_a(-7.567898865090683e-05)),(to_sfixed_a(-0.00016375046106986701)),(to_sfixed_a(4.294576501706615e-05)),(to_sfixed_a(-7.870485569583252e-05)),(to_sfixed_a(0.0001294638786930591)),(to_sfixed_a(-0.00015927347703836858)),(to_sfixed_a(0.00016439642058685422)),(to_sfixed_a(0.005024057812988758)),(to_sfixed_a(-0.002167119411751628)),(to_sfixed_a(-2.8934096917510033e-05)),(to_sfixed_a(-6.664253305643797e-05)),(to_sfixed_a(-0.00027566711651161313)),(to_sfixed_a(0.00881236232817173)),(to_sfixed_a(-5.955873348284513e-06)),(to_sfixed_a(0.19042128324508667)),(to_sfixed_a(-0.0007368900114670396)),(to_sfixed_a(0.013094470836222172)));

    constant weight_n2_69 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.021321171894669533)),(to_sfixed_a(-0.14693978428840637)),(to_sfixed_a(-0.00017683768237475306)),(to_sfixed_a(2.6687979698181152e-05)),(to_sfixed_a(-0.00899468082934618)),(to_sfixed_a(1.1107928003184497e-05)),(to_sfixed_a(-0.004909760318696499)),(to_sfixed_a(-0.00018481114238966256)),(to_sfixed_a(-0.00011655554408207536)),(to_sfixed_a(-0.00018524061306379735)),(to_sfixed_a(-0.00027129618683829904)),(to_sfixed_a(-0.001160788699053228)),(to_sfixed_a(0.4418184757232666)),(to_sfixed_a(-0.000644522428046912)),(to_sfixed_a(-9.169264376396313e-05)),(to_sfixed_a(0.00016088075062725693)),(to_sfixed_a(-0.0016573728062212467)),(to_sfixed_a(-3.75605741282925e-05)),(to_sfixed_a(-0.02361091412603855)),(to_sfixed_a(0.006462139077484608)),(to_sfixed_a(0.00028424206539057195)),(to_sfixed_a(0.00010056810424430296)),(to_sfixed_a(4.4664222514256835e-05)),(to_sfixed_a(-0.031077664345502853)),(to_sfixed_a(-0.00348193128593266)),(to_sfixed_a(-0.25353705883026123)),(to_sfixed_a(7.125127740437165e-05)),(to_sfixed_a(-0.00035630696220323443)),(to_sfixed_a(-0.010627849027514458)),(to_sfixed_a(-0.00014127408212516457)),(to_sfixed_a(-0.012657544575631618)),(to_sfixed_a(-1.824661740101874e-05)),(to_sfixed_a(-0.004664760548621416)),(to_sfixed_a(4.093674215255305e-05)),(to_sfixed_a(-3.2555952202528715e-05)),(to_sfixed_a(-0.00015475120744667947)),(to_sfixed_a(0.2399594485759735)),(to_sfixed_a(0.2193586528301239)),(to_sfixed_a(0.017668591812253)),(to_sfixed_a(1.4207078493200243e-05)),(to_sfixed_a(-0.014935004524886608)),(to_sfixed_a(-0.0002097111864713952)),(to_sfixed_a(0.00011257143341936171)),(to_sfixed_a(9.392313950229436e-05)),(to_sfixed_a(-0.00484379893168807)),(to_sfixed_a(0.5779188275337219)),(to_sfixed_a(0.0003918232978321612)),(to_sfixed_a(-0.0158085934817791)),(to_sfixed_a(-0.00018618347530718893)),(to_sfixed_a(-0.008930515497922897)),(to_sfixed_a(-0.0015058285789564252)),(to_sfixed_a(-0.001242010504938662)),(to_sfixed_a(-0.00011334721784805879)),(to_sfixed_a(-0.0010571860475465655)),(to_sfixed_a(-0.005856611765921116)),(to_sfixed_a(0.0012146258959546685)),(to_sfixed_a(-0.00011313670256640762)),(to_sfixed_a(-0.0021179248578846455)),(to_sfixed_a(2.3957734811119735e-05)),(to_sfixed_a(-6.93409820087254e-05)),(to_sfixed_a(-0.0004102906968910247)),(to_sfixed_a(-0.0021112910471856594)),(to_sfixed_a(0.00026897696079686284)),(to_sfixed_a(0.020233934745192528)),(to_sfixed_a(3.158633626298979e-05)),(to_sfixed_a(0.0011945331934839487)),(to_sfixed_a(-1.9840030290652066e-05)),(to_sfixed_a(-0.3942195177078247)),(to_sfixed_a(5.585350299952552e-05)),(to_sfixed_a(-0.00028590759029611945)),(to_sfixed_a(0.10388283431529999)),(to_sfixed_a(0.009617749601602554)),(to_sfixed_a(0.22312018275260925)),(to_sfixed_a(-0.00011646775237750262)),(to_sfixed_a(-1.8044291209662333e-05)),(to_sfixed_a(-6.957250298000872e-05)),(to_sfixed_a(-0.00011268626258242875)),(to_sfixed_a(-0.0008428136352449656)),(to_sfixed_a(6.873243546579033e-05)),(to_sfixed_a(0.0005597688141278923)),(to_sfixed_a(0.00019968478591181338)),(to_sfixed_a(7.609630847582594e-05)),(to_sfixed_a(-0.0007978520588949323)),(to_sfixed_a(-0.00224841246381402)),(to_sfixed_a(0.0001160158499260433)),(to_sfixed_a(-0.0028527688700705767)),(to_sfixed_a(0.0025510459672659636)),(to_sfixed_a(-0.0003273199254181236)),(to_sfixed_a(0.00024527229834347963)),(to_sfixed_a(-0.0001156005819211714)),(to_sfixed_a(0.00109367654658854)),(to_sfixed_a(-0.00016106276598293334)),(to_sfixed_a(0.0018998893210664392)),(to_sfixed_a(3.69735062122345e-05)),(to_sfixed_a(0.0006207820260897279)),(to_sfixed_a(9.827988833421841e-06)),(to_sfixed_a(-0.00018044511671178043)),(to_sfixed_a(-0.00017472250328864902)),(to_sfixed_a(0.00024348945589736104)),(to_sfixed_a(1.63383774633985e-05)),(to_sfixed_a(-0.000858538318425417)),(to_sfixed_a(-2.9585222364403307e-05)),(to_sfixed_a(-7.313209789572284e-05)),(to_sfixed_a(0.24363937973976135)),(to_sfixed_a(-0.0008436902426183224)),(to_sfixed_a(-0.00629581930115819)),(to_sfixed_a(7.174238271545619e-05)),(to_sfixed_a(4.0366241591982543e-05)),(to_sfixed_a(-3.6885830922983587e-07)),(to_sfixed_a(-0.006341917905956507)),(to_sfixed_a(-0.024244019761681557)),(to_sfixed_a(0.00011637808347586542)),(to_sfixed_a(-0.002422436373308301)),(to_sfixed_a(6.790892803110182e-05)),(to_sfixed_a(1.6773723473306745e-05)),(to_sfixed_a(0.003965658601373434)),(to_sfixed_a(0.002516786102205515)),(to_sfixed_a(-0.0010885512456297874)),(to_sfixed_a(5.35885410499759e-05)),(to_sfixed_a(0.3114193081855774)),(to_sfixed_a(1.424683432560414e-05)),(to_sfixed_a(-0.00023686198983341455)),(to_sfixed_a(-6.8458124587778e-05)),(to_sfixed_a(2.9391812859103084e-05)),(to_sfixed_a(-8.454931958112866e-05)),(to_sfixed_a(-0.0033818779047578573)),(to_sfixed_a(-0.00011497173545649275)),(to_sfixed_a(0.00021946057677268982)),(to_sfixed_a(-8.641235763207078e-05)),(to_sfixed_a(-4.6600052883150056e-05)),(to_sfixed_a(-8.498500392306596e-07)),(to_sfixed_a(0.000109880231320858)),(to_sfixed_a(-0.00031180543010123074)),(to_sfixed_a(-0.0002973020018544048)),(to_sfixed_a(-0.00011398311471566558)),(to_sfixed_a(-0.0002088695764541626)),(to_sfixed_a(-0.3733576238155365)),(to_sfixed_a(0.0001893416338134557)),(to_sfixed_a(0.0002230534446425736)),(to_sfixed_a(7.148533768486232e-05)),(to_sfixed_a(0.0065423110499978065)),(to_sfixed_a(1.1358170013409108e-06)),(to_sfixed_a(-1.2570104445330799e-05)),(to_sfixed_a(2.965495514217764e-05)),(to_sfixed_a(1.7365109670208767e-06)),(to_sfixed_a(4.5210705138742924e-05)),(to_sfixed_a(0.00021674024173989892)),(to_sfixed_a(9.330517059424892e-05)),(to_sfixed_a(-5.9013393183704466e-05)),(to_sfixed_a(-0.0007077567861415446)),(to_sfixed_a(0.00016725290333852172)),(to_sfixed_a(6.424127786885947e-05)),(to_sfixed_a(0.007699521724134684)),(to_sfixed_a(-0.0001161227046395652)),(to_sfixed_a(6.721311365254223e-05)),(to_sfixed_a(0.12236358225345612)),(to_sfixed_a(-0.0002184732147725299)),(to_sfixed_a(-0.003238525241613388)),(to_sfixed_a(-7.517401172663085e-07)),(to_sfixed_a(-6.764347926946357e-05)),(to_sfixed_a(-9.288742148783058e-07)),(to_sfixed_a(1.094288018066436e-05)),(to_sfixed_a(0.0011287418892607093)),(to_sfixed_a(-0.20754949748516083)),(to_sfixed_a(-0.21784470975399017)),(to_sfixed_a(0.0001040396819007583)),(to_sfixed_a(-0.0003220912185497582)),(to_sfixed_a(0.007210101000964642)),(to_sfixed_a(0.00020535651128739119)),(to_sfixed_a(0.00016820483142510056)),(to_sfixed_a(0.35602429509162903)),(to_sfixed_a(2.9536106012528762e-05)),(to_sfixed_a(-0.001600240240804851)),(to_sfixed_a(-0.00012026209878968075)),(to_sfixed_a(-0.16024059057235718)),(to_sfixed_a(0.00029895181069150567)),(to_sfixed_a(0.00017355740419588983)),(to_sfixed_a(-0.0007079612114466727)),(to_sfixed_a(0.00157740933354944)),(to_sfixed_a(0.014084932394325733)),(to_sfixed_a(-0.002052305731922388)),(to_sfixed_a(-0.0067093889228999615)),(to_sfixed_a(0.0002368500136071816)),(to_sfixed_a(-0.00018398121756035835)),(to_sfixed_a(-0.00011916588118765503)),(to_sfixed_a(0.32120540738105774)),(to_sfixed_a(-0.0015599472681060433)),(to_sfixed_a(-0.00145675556268543)),(to_sfixed_a(1.7379097698722035e-06)),(to_sfixed_a(-2.4825703803799115e-05)),(to_sfixed_a(-0.00014778428885620087)),(to_sfixed_a(-7.444896618835628e-05)),(to_sfixed_a(-0.0012845637975260615)),(to_sfixed_a(0.0007664794684387743)),(to_sfixed_a(0.0003037798742298037)),(to_sfixed_a(0.28756675124168396)),(to_sfixed_a(0.00018772849580273032)),(to_sfixed_a(0.0013604048872366548)),(to_sfixed_a(-0.3017311990261078)),(to_sfixed_a(0.00011260727478656918)),(to_sfixed_a(4.433834692463279e-05)),(to_sfixed_a(0.00017953114002011716)),(to_sfixed_a(0.0003104271017946303)),(to_sfixed_a(0.00013405721983872354)),(to_sfixed_a(1.4409182767849416e-05)),(to_sfixed_a(0.00033254866139031947)),(to_sfixed_a(9.71224217209965e-05)),(to_sfixed_a(0.022053292021155357)),(to_sfixed_a(-0.0005830125301145017)),(to_sfixed_a(-0.006818877533078194)),(to_sfixed_a(0.002465815283358097)),(to_sfixed_a(1.6309386410284787e-06)),(to_sfixed_a(-0.0001925388933159411)),(to_sfixed_a(-0.00017535853839945048)),(to_sfixed_a(4.3520434701349586e-05)),(to_sfixed_a(-0.0001062787341652438)),(to_sfixed_a(-0.00021988118533045053)),(to_sfixed_a(0.0006063461187295616)),(to_sfixed_a(-0.3453019857406616)),(to_sfixed_a(2.1414016373455524e-06)),(to_sfixed_a(-7.110602018656209e-05)),(to_sfixed_a(7.075116445776075e-05)),(to_sfixed_a(-0.00023655107361264527)),(to_sfixed_a(-0.0005035484791733325)),(to_sfixed_a(-0.0031780756544321775)),(to_sfixed_a(-3.447139170020819e-05)),(to_sfixed_a(-0.00017842126544564962)),(to_sfixed_a(0.00021781670511700213)),(to_sfixed_a(-0.009535192511975765)),(to_sfixed_a(0.0007438617176376283)),(to_sfixed_a(-0.24426764249801636)),(to_sfixed_a(0.000278186023933813)),(to_sfixed_a(0.00012133138079661876)),(to_sfixed_a(-0.00012933154357597232)),(to_sfixed_a(0.00011214765254408121)),(to_sfixed_a(0.0046376753598451614)),(to_sfixed_a(0.010552474297583103)),(to_sfixed_a(-7.100836228346452e-05)),(to_sfixed_a(1.8931677914224565e-06)),(to_sfixed_a(0.00041812710696831346)),(to_sfixed_a(-0.0008914015488699079)),(to_sfixed_a(2.227618097094819e-05)),(to_sfixed_a(0.22294364869594574)),(to_sfixed_a(6.818499969085678e-05)),(to_sfixed_a(-0.02812284417450428)),(to_sfixed_a(0.007921939715743065)),(to_sfixed_a(-0.0048731472343206406)),(to_sfixed_a(-0.008659053593873978)),(to_sfixed_a(0.00020516868971753865)),(to_sfixed_a(6.186299287946895e-05)),(to_sfixed_a(-0.009632382541894913)),(to_sfixed_a(0.00014619450666941702)),(to_sfixed_a(-0.0016208022134378552)),(to_sfixed_a(4.8197667638305575e-05)),(to_sfixed_a(0.0002629375958349556)),(to_sfixed_a(-0.007330566179007292)),(to_sfixed_a(-0.0006030381773598492)),(to_sfixed_a(0.00041433892329223454)),(to_sfixed_a(-0.0001522109523648396)),(to_sfixed_a(-0.002188921207562089)),(to_sfixed_a(-0.00010675600788090378)),(to_sfixed_a(-8.808130951365456e-05)),(to_sfixed_a(0.00020579741976689547)),(to_sfixed_a(-0.0007780923042446375)),(to_sfixed_a(-0.00029318209271878004)),(to_sfixed_a(-0.007182282395660877)),(to_sfixed_a(-3.1947012757882476e-05)),(to_sfixed_a(-1.9440496544120833e-05)),(to_sfixed_a(6.264105468289927e-05)),(to_sfixed_a(-0.0061963279731571674)),(to_sfixed_a(-0.19843249022960663)),(to_sfixed_a(0.0001556806528242305)),(to_sfixed_a(-0.00016068978584371507)),(to_sfixed_a(0.00019090935529675335)),(to_sfixed_a(1.744591281749308e-05)),(to_sfixed_a(0.0002778297639451921)),(to_sfixed_a(-0.6230766773223877)),(to_sfixed_a(-0.0018166692461818457)),(to_sfixed_a(-0.27525612711906433)),(to_sfixed_a(-0.24353472888469696)),(to_sfixed_a(-4.708046617452055e-06)),(to_sfixed_a(-0.00012806773884221911)),(to_sfixed_a(1.2330157915130258e-05)),(to_sfixed_a(0.18741653859615326)),(to_sfixed_a(2.1040370484115556e-05)),(to_sfixed_a(-3.3590848033782095e-05)),(to_sfixed_a(1.4101424312684685e-06)),(to_sfixed_a(0.32596156001091003)),(to_sfixed_a(5.998130654916167e-05)),(to_sfixed_a(-0.00027201228658668697)),(to_sfixed_a(-0.0004350020899437368)),(to_sfixed_a(-0.007174456957727671)),(to_sfixed_a(0.011269956827163696)),(to_sfixed_a(0.00013643709826283157)),(to_sfixed_a(-0.0024213874712586403)),(to_sfixed_a(-0.002912824507802725)),(to_sfixed_a(-0.008908920921385288)),(to_sfixed_a(4.830060061067343e-05)),(to_sfixed_a(0.2800523042678833)),(to_sfixed_a(-0.6981225609779358)),(to_sfixed_a(0.2881714999675751)));

    constant weight_n2_70 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.34269073605537415)),(to_sfixed_a(-0.0007191718323156238)),(to_sfixed_a(0.39375051856040955)),(to_sfixed_a(-0.00011540178093127906)),(to_sfixed_a(0.23756751418113708)),(to_sfixed_a(-3.126348019577563e-06)),(to_sfixed_a(-0.021273192018270493)),(to_sfixed_a(-0.00022982692462392151)),(to_sfixed_a(9.838573168963194e-05)),(to_sfixed_a(0.00013080482312943786)),(to_sfixed_a(-2.0966679585399106e-05)),(to_sfixed_a(0.02417881414294243)),(to_sfixed_a(-0.0011501837288960814)),(to_sfixed_a(0.00015619114856235683)),(to_sfixed_a(-0.00026577687822282314)),(to_sfixed_a(-0.0001287904306082055)),(to_sfixed_a(0.0008404466207139194)),(to_sfixed_a(-1.9151921151205897e-06)),(to_sfixed_a(0.0046765487641096115)),(to_sfixed_a(0.0004895463353022933)),(to_sfixed_a(0.00012989020615350455)),(to_sfixed_a(-6.12010044278577e-05)),(to_sfixed_a(0.0002705795341171324)),(to_sfixed_a(-0.0038950988091528416)),(to_sfixed_a(0.0029610414057970047)),(to_sfixed_a(-0.0008278583409264684)),(to_sfixed_a(8.609191718278453e-05)),(to_sfixed_a(0.3252953588962555)),(to_sfixed_a(-0.00012370060721877962)),(to_sfixed_a(0.0002921409031841904)),(to_sfixed_a(-0.008608772419393063)),(to_sfixed_a(0.00010353947436669841)),(to_sfixed_a(-0.0077471486292779446)),(to_sfixed_a(7.087890116963536e-05)),(to_sfixed_a(-4.349699156591669e-05)),(to_sfixed_a(0.00022025787620805204)),(to_sfixed_a(-4.189410537946969e-05)),(to_sfixed_a(0.1480139195919037)),(to_sfixed_a(0.006113127339631319)),(to_sfixed_a(0.00025212031323462725)),(to_sfixed_a(-0.007499277591705322)),(to_sfixed_a(0.0013910492416471243)),(to_sfixed_a(1.7580394342076033e-05)),(to_sfixed_a(0.00013219595712143928)),(to_sfixed_a(-0.0070934114046394825)),(to_sfixed_a(-0.0010863144416362047)),(to_sfixed_a(0.003316994523629546)),(to_sfixed_a(0.48437365889549255)),(to_sfixed_a(-0.0002738577895797789)),(to_sfixed_a(0.000982443685643375)),(to_sfixed_a(-0.0064498018473386765)),(to_sfixed_a(0.0002011200413107872)),(to_sfixed_a(0.00012950606469530612)),(to_sfixed_a(0.0035928545985370874)),(to_sfixed_a(-0.0001993637706618756)),(to_sfixed_a(-0.002613473916426301)),(to_sfixed_a(0.00015418145630974323)),(to_sfixed_a(0.00027829522150568664)),(to_sfixed_a(0.0003024021571036428)),(to_sfixed_a(0.00010708154877647758)),(to_sfixed_a(0.0007829134119674563)),(to_sfixed_a(0.0007188101299107075)),(to_sfixed_a(0.0018918371060863137)),(to_sfixed_a(-0.3021858036518097)),(to_sfixed_a(8.941579289967194e-05)),(to_sfixed_a(0.00010957672930089757)),(to_sfixed_a(1.1557829566299915e-05)),(to_sfixed_a(0.0008506863377988338)),(to_sfixed_a(0.00045877060620114207)),(to_sfixed_a(0.00030381526448763907)),(to_sfixed_a(-0.003256535157561302)),(to_sfixed_a(0.001614508219063282)),(to_sfixed_a(-0.010251765139400959)),(to_sfixed_a(-0.00020505257998593152)),(to_sfixed_a(-0.0001492229785071686)),(to_sfixed_a(0.00010521236981730908)),(to_sfixed_a(0.02881285920739174)),(to_sfixed_a(0.00017075422510970384)),(to_sfixed_a(0.00013660980039276183)),(to_sfixed_a(0.08181974291801453)),(to_sfixed_a(-0.006335774436593056)),(to_sfixed_a(2.1010986529290676e-05)),(to_sfixed_a(0.00028585444670170546)),(to_sfixed_a(-0.1614745408296585)),(to_sfixed_a(-0.00012791490007657558)),(to_sfixed_a(-0.016595367342233658)),(to_sfixed_a(0.024753984063863754)),(to_sfixed_a(0.002404274418950081)),(to_sfixed_a(-0.00018011500651482493)),(to_sfixed_a(2.0526211301330477e-05)),(to_sfixed_a(-0.00012628702097572386)),(to_sfixed_a(-1.1237661965424195e-06)),(to_sfixed_a(0.00279080867767334)),(to_sfixed_a(0.00011676781286951154)),(to_sfixed_a(0.001219684723764658)),(to_sfixed_a(-6.020941509632394e-05)),(to_sfixed_a(-1.6161444364115596e-05)),(to_sfixed_a(0.00023673813848290592)),(to_sfixed_a(-0.0001517074415460229)),(to_sfixed_a(-0.00012538168812170625)),(to_sfixed_a(0.0008614328107796609)),(to_sfixed_a(-0.004475634545087814)),(to_sfixed_a(7.639623072464019e-05)),(to_sfixed_a(-0.006267184857279062)),(to_sfixed_a(-0.003668963210657239)),(to_sfixed_a(0.0012945614289492369)),(to_sfixed_a(-0.00016837345901876688)),(to_sfixed_a(6.124261562945321e-05)),(to_sfixed_a(-0.0003763873246498406)),(to_sfixed_a(-0.011928740888834)),(to_sfixed_a(-0.8674494624137878)),(to_sfixed_a(-8.955210068961605e-05)),(to_sfixed_a(0.3003241717815399)),(to_sfixed_a(-0.00016861918265931308)),(to_sfixed_a(-0.00022286936291493475)),(to_sfixed_a(-0.01083375047892332)),(to_sfixed_a(-0.00010021701746154577)),(to_sfixed_a(-0.30392807722091675)),(to_sfixed_a(-7.41479016141966e-05)),(to_sfixed_a(-0.008185047656297684)),(to_sfixed_a(0.00010506785474717617)),(to_sfixed_a(0.00017502595437690616)),(to_sfixed_a(0.0017555771628394723)),(to_sfixed_a(-3.061799725401215e-05)),(to_sfixed_a(-0.00029863585950806737)),(to_sfixed_a(-0.00675848638638854)),(to_sfixed_a(-0.0021336690988391638)),(to_sfixed_a(-8.382396481465548e-05)),(to_sfixed_a(0.0002158928255084902)),(to_sfixed_a(-0.0001519562501925975)),(to_sfixed_a(0.0001498773053754121)),(to_sfixed_a(-0.00012076528219040483)),(to_sfixed_a(0.0016245378646999598)),(to_sfixed_a(0.005538858938962221)),(to_sfixed_a(-2.2763477318221703e-05)),(to_sfixed_a(-1.0907897376455367e-06)),(to_sfixed_a(0.001443674205802381)),(to_sfixed_a(0.00017371689318679273)),(to_sfixed_a(6.62858656141907e-05)),(to_sfixed_a(-0.00020033417968079448)),(to_sfixed_a(-3.342776471981779e-05)),(to_sfixed_a(7.28662998881191e-05)),(to_sfixed_a(-1.8807841115631163e-05)),(to_sfixed_a(6.542788469232619e-05)),(to_sfixed_a(-7.295540126506239e-05)),(to_sfixed_a(-0.0011158070992678404)),(to_sfixed_a(-4.28723797085695e-06)),(to_sfixed_a(-0.00017455563647672534)),(to_sfixed_a(9.295774361817166e-06)),(to_sfixed_a(0.0021641310304403305)),(to_sfixed_a(0.00017855141777545214)),(to_sfixed_a(-1.241968129761517e-05)),(to_sfixed_a(0.0002135721588274464)),(to_sfixed_a(3.0274488381110132e-05)),(to_sfixed_a(-0.00023533799685537815)),(to_sfixed_a(0.012665975838899612)),(to_sfixed_a(-0.00014291155093815178)),(to_sfixed_a(0.001867438666522503)),(to_sfixed_a(6.873661186546087e-05)),(to_sfixed_a(-6.356541416607797e-05)),(to_sfixed_a(-0.00012135522410972044)),(to_sfixed_a(5.665874050464481e-05)),(to_sfixed_a(0.013729309663176537)),(to_sfixed_a(1.651020284043625e-05)),(to_sfixed_a(0.00019316771067678928)),(to_sfixed_a(-0.0029125583823770285)),(to_sfixed_a(-0.00029928318690508604)),(to_sfixed_a(0.3992876410484314)),(to_sfixed_a(-8.154565148288384e-05)),(to_sfixed_a(0.0001369442616123706)),(to_sfixed_a(-9.962219337467104e-06)),(to_sfixed_a(8.772595901973546e-05)),(to_sfixed_a(-0.0017476006178185344)),(to_sfixed_a(-6.53843380860053e-05)),(to_sfixed_a(-0.0021567856892943382)),(to_sfixed_a(0.0004443901707418263)),(to_sfixed_a(0.17709538340568542)),(to_sfixed_a(-0.0031524954829365015)),(to_sfixed_a(0.4728798270225525)),(to_sfixed_a(-0.002211229410022497)),(to_sfixed_a(0.0004493730375543237)),(to_sfixed_a(-0.011341563425958157)),(to_sfixed_a(-3.322505654068664e-05)),(to_sfixed_a(2.9131952032912523e-05)),(to_sfixed_a(-0.00010158627992495894)),(to_sfixed_a(0.0005469830939546227)),(to_sfixed_a(0.0008253557025454938)),(to_sfixed_a(-0.00011334288137732074)),(to_sfixed_a(-4.13102243328467e-05)),(to_sfixed_a(0.00024271823349408805)),(to_sfixed_a(-0.0025737506803125143)),(to_sfixed_a(5.0803944759536535e-05)),(to_sfixed_a(0.016813049092888832)),(to_sfixed_a(-0.0024772952310740948)),(to_sfixed_a(7.688580808462575e-05)),(to_sfixed_a(-0.002639466430991888)),(to_sfixed_a(6.937790021765977e-05)),(to_sfixed_a(-0.009486607275903225)),(to_sfixed_a(0.0029262586031109095)),(to_sfixed_a(-6.543667404912412e-05)),(to_sfixed_a(4.7721750888740644e-05)),(to_sfixed_a(6.521263276226819e-05)),(to_sfixed_a(-0.0002512557548470795)),(to_sfixed_a(-0.00010548443242441863)),(to_sfixed_a(3.5969598684459925e-05)),(to_sfixed_a(2.480918374203611e-05)),(to_sfixed_a(-0.0013706450117751956)),(to_sfixed_a(0.0014561109710484743)),(to_sfixed_a(-0.01799551583826542)),(to_sfixed_a(-0.0003724727139342576)),(to_sfixed_a(0.009762070141732693)),(to_sfixed_a(6.402867438737303e-05)),(to_sfixed_a(-4.5957705879118294e-05)),(to_sfixed_a(-0.00012822328426409513)),(to_sfixed_a(3.0434090149356052e-05)),(to_sfixed_a(-1.3153476174920797e-07)),(to_sfixed_a(-0.0040665664710104465)),(to_sfixed_a(-0.0014675735728815198)),(to_sfixed_a(0.0015895761316642165)),(to_sfixed_a(-0.0004156621580477804)),(to_sfixed_a(4.66024357592687e-06)),(to_sfixed_a(3.780067345360294e-05)),(to_sfixed_a(0.0001528523425804451)),(to_sfixed_a(0.0019912279676645994)),(to_sfixed_a(0.11738590896129608)),(to_sfixed_a(9.579915058566257e-05)),(to_sfixed_a(0.00023590459022670984)),(to_sfixed_a(0.00010451434354763478)),(to_sfixed_a(0.002617449266836047)),(to_sfixed_a(0.00026190740754827857)),(to_sfixed_a(0.006161988712847233)),(to_sfixed_a(8.609460201114416e-05)),(to_sfixed_a(3.732943150680512e-05)),(to_sfixed_a(6.492192187579349e-05)),(to_sfixed_a(-0.007851975969970226)),(to_sfixed_a(-0.0029545314610004425)),(to_sfixed_a(-0.005906716920435429)),(to_sfixed_a(-0.00015332559996750206)),(to_sfixed_a(5.431383033283055e-05)),(to_sfixed_a(0.0002546661999076605)),(to_sfixed_a(-0.0001084171308320947)),(to_sfixed_a(6.93602196406573e-05)),(to_sfixed_a(0.002716262824833393)),(to_sfixed_a(-0.00010856729932129383)),(to_sfixed_a(0.13480333983898163)),(to_sfixed_a(-0.0028155252803117037)),(to_sfixed_a(-0.005931801162660122)),(to_sfixed_a(0.17352642118930817)),(to_sfixed_a(-0.00018243142403662205)),(to_sfixed_a(-0.0013707856414839625)),(to_sfixed_a(-0.00020620744908228517)),(to_sfixed_a(7.764052134007215e-05)),(to_sfixed_a(-0.00019665008585434407)),(to_sfixed_a(-0.00012873552623204887)),(to_sfixed_a(0.00014720215403940529)),(to_sfixed_a(-0.008926333859562874)),(to_sfixed_a(-0.0011754067381843925)),(to_sfixed_a(0.0001117853753385134)),(to_sfixed_a(-0.0001769974041962996)),(to_sfixed_a(-0.003098869463428855)),(to_sfixed_a(2.0248990040272474e-06)),(to_sfixed_a(0.0004858853935729712)),(to_sfixed_a(0.000135816095280461)),(to_sfixed_a(0.0006275451160036027)),(to_sfixed_a(1.6318932466674596e-05)),(to_sfixed_a(-0.016707731410861015)),(to_sfixed_a(4.4500731746666133e-05)),(to_sfixed_a(-0.00017471081810072064)),(to_sfixed_a(5.777863407274708e-05)),(to_sfixed_a(-0.001578143797814846)),(to_sfixed_a(0.000347000895999372)),(to_sfixed_a(-0.00030569176306016743)),(to_sfixed_a(-0.00020600849529728293)),(to_sfixed_a(-3.501421451801434e-05)),(to_sfixed_a(-6.413558730855584e-05)),(to_sfixed_a(-8.460076787741855e-05)),(to_sfixed_a(0.18951156735420227)),(to_sfixed_a(-0.003880937583744526)),(to_sfixed_a(-0.019570695236325264)),(to_sfixed_a(0.0013028536923229694)),(to_sfixed_a(7.691193604841828e-05)),(to_sfixed_a(0.00011693441774696112)),(to_sfixed_a(1.8381309928372502e-05)),(to_sfixed_a(0.0004842568887397647)),(to_sfixed_a(-0.00045020144898444414)),(to_sfixed_a(0.00013515834871213883)),(to_sfixed_a(-0.0006472887471318245)),(to_sfixed_a(9.753649646881968e-05)),(to_sfixed_a(9.27170185605064e-05)),(to_sfixed_a(-0.00017129132174886763)),(to_sfixed_a(0.00025379389990121126)),(to_sfixed_a(-0.006359782535582781)),(to_sfixed_a(0.0012239476200193167)),(to_sfixed_a(0.00011381784861441702)),(to_sfixed_a(0.0003993733262177557)),(to_sfixed_a(0.11588577181100845)),(to_sfixed_a(0.00037589360726997256)),(to_sfixed_a(-0.00030777600477449596)),(to_sfixed_a(0.00206114468164742)),(to_sfixed_a(0.003237253287807107)),(to_sfixed_a(-0.00356938224285841)));

    constant weight_n2_71 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.10557638853788376)),(to_sfixed_a(0.15839596092700958)),(to_sfixed_a(-0.0010266228346154094)),(to_sfixed_a(0.0001826184889068827)),(to_sfixed_a(0.011846152134239674)),(to_sfixed_a(2.235391002614051e-05)),(to_sfixed_a(0.00046447766362689435)),(to_sfixed_a(-6.527664663735777e-05)),(to_sfixed_a(-0.00018075318075716496)),(to_sfixed_a(0.00017661036690697074)),(to_sfixed_a(-1.8189854017691687e-05)),(to_sfixed_a(-0.0010779683943837881)),(to_sfixed_a(0.4129253923892975)),(to_sfixed_a(-0.0004913541488349438)),(to_sfixed_a(0.00017400231445208192)),(to_sfixed_a(0.00013687075988855213)),(to_sfixed_a(0.0041869585402309895)),(to_sfixed_a(0.0001672374055488035)),(to_sfixed_a(-0.2357560694217682)),(to_sfixed_a(-0.0007023952202871442)),(to_sfixed_a(6.509765808004886e-05)),(to_sfixed_a(-1.8991457181982696e-05)),(to_sfixed_a(3.55995653080754e-05)),(to_sfixed_a(0.0002517353859730065)),(to_sfixed_a(0.0007252019713632762)),(to_sfixed_a(0.0009591178386472166)),(to_sfixed_a(0.0004220609553158283)),(to_sfixed_a(5.323192453943193e-05)),(to_sfixed_a(0.0002874083293136209)),(to_sfixed_a(2.3335396690526977e-05)),(to_sfixed_a(-0.0007262712460942566)),(to_sfixed_a(0.00041790155228227377)),(to_sfixed_a(0.0021434780210256577)),(to_sfixed_a(0.00020406272960826755)),(to_sfixed_a(0.00010591211321298033)),(to_sfixed_a(-7.772224489599466e-05)),(to_sfixed_a(0.110618457198143)),(to_sfixed_a(0.004268005955964327)),(to_sfixed_a(0.21304459869861603)),(to_sfixed_a(-0.00019889470422640443)),(to_sfixed_a(-0.004265645518898964)),(to_sfixed_a(0.0013420562027022243)),(to_sfixed_a(-0.00022488817921839654)),(to_sfixed_a(0.0001535859191790223)),(to_sfixed_a(-0.0007649053004570305)),(to_sfixed_a(0.39660680294036865)),(to_sfixed_a(0.0008633121615275741)),(to_sfixed_a(-0.4374648928642273)),(to_sfixed_a(-0.0001590804458828643)),(to_sfixed_a(-0.0012106436770409346)),(to_sfixed_a(-0.1818958967924118)),(to_sfixed_a(-0.0005386081757023931)),(to_sfixed_a(-4.29321953561157e-05)),(to_sfixed_a(0.0013094197493046522)),(to_sfixed_a(0.0018531633540987968)),(to_sfixed_a(-0.0009893454844132066)),(to_sfixed_a(-3.667139753815718e-05)),(to_sfixed_a(-0.0001279425050597638)),(to_sfixed_a(2.521665010135621e-05)),(to_sfixed_a(-0.00010597660730127245)),(to_sfixed_a(-0.000569372670724988)),(to_sfixed_a(-0.0019042430212721229)),(to_sfixed_a(0.00027569083613343537)),(to_sfixed_a(0.004264465533196926)),(to_sfixed_a(0.00019299877749290317)),(to_sfixed_a(0.0019308694172650576)),(to_sfixed_a(5.725960363633931e-06)),(to_sfixed_a(-0.4598816931247711)),(to_sfixed_a(-0.0004877836909145117)),(to_sfixed_a(-3.807854955084622e-05)),(to_sfixed_a(-0.001152743585407734)),(to_sfixed_a(-0.0016893285792320967)),(to_sfixed_a(-0.01672513410449028)),(to_sfixed_a(0.00021750091400463134)),(to_sfixed_a(-0.00018008542247116566)),(to_sfixed_a(1.5005483874119818e-05)),(to_sfixed_a(-0.0006168583640828729)),(to_sfixed_a(-2.3646149202249944e-05)),(to_sfixed_a(0.00024770392337813973)),(to_sfixed_a(0.007285716477781534)),(to_sfixed_a(-0.00020604341989383101)),(to_sfixed_a(3.0042474463698454e-05)),(to_sfixed_a(0.00034576281905174255)),(to_sfixed_a(0.009586403146386147)),(to_sfixed_a(-0.00014932401245459914)),(to_sfixed_a(0.0010604115668684244)),(to_sfixed_a(-0.00981347169727087)),(to_sfixed_a(5.209031223785132e-05)),(to_sfixed_a(-0.00012669115676544607)),(to_sfixed_a(7.393702253466472e-05)),(to_sfixed_a(0.0008862162940204144)),(to_sfixed_a(0.00028826232301071286)),(to_sfixed_a(-3.6099452700000256e-05)),(to_sfixed_a(0.0001133381447289139)),(to_sfixed_a(0.21878692507743835)),(to_sfixed_a(-4.963911487720907e-05)),(to_sfixed_a(-0.0003133390564471483)),(to_sfixed_a(0.0004144567355979234)),(to_sfixed_a(0.00010875429870793596)),(to_sfixed_a(1.082509697880596e-06)),(to_sfixed_a(-0.00030498357955366373)),(to_sfixed_a(-0.0002884953864850104)),(to_sfixed_a(-8.028392039705068e-05)),(to_sfixed_a(-2.7598600354394875e-05)),(to_sfixed_a(0.003028406063094735)),(to_sfixed_a(-9.605495870346203e-05)),(to_sfixed_a(7.010546687524766e-05)),(to_sfixed_a(6.404898158507422e-07)),(to_sfixed_a(0.000304173183394596)),(to_sfixed_a(0.00038408415275625885)),(to_sfixed_a(0.003222930710762739)),(to_sfixed_a(0.00023605399474035949)),(to_sfixed_a(-4.7427674871869385e-05)),(to_sfixed_a(-0.00011576660472201183)),(to_sfixed_a(-0.00020160069107078016)),(to_sfixed_a(0.003201617393642664)),(to_sfixed_a(0.0005625698831863701)),(to_sfixed_a(-0.00011797060869866982)),(to_sfixed_a(6.65256375214085e-05)),(to_sfixed_a(0.03223053365945816)),(to_sfixed_a(-5.366692857933231e-05)),(to_sfixed_a(6.523980118799955e-05)),(to_sfixed_a(0.00020219816360622644)),(to_sfixed_a(-8.45128670334816e-06)),(to_sfixed_a(7.383958291029558e-05)),(to_sfixed_a(0.0011855058837682009)),(to_sfixed_a(0.004449437838047743)),(to_sfixed_a(7.107491546776146e-05)),(to_sfixed_a(-0.0001948393473867327)),(to_sfixed_a(-0.0004586017457768321)),(to_sfixed_a(0.0002964164305012673)),(to_sfixed_a(-3.846293839160353e-05)),(to_sfixed_a(-0.0017170370556414127)),(to_sfixed_a(0.00865844450891018)),(to_sfixed_a(0.0002914378419518471)),(to_sfixed_a(1.4121906133368611e-07)),(to_sfixed_a(-0.23753072321414948)),(to_sfixed_a(0.0006011469522491097)),(to_sfixed_a(-2.3070093448041007e-05)),(to_sfixed_a(0.00012272717140149325)),(to_sfixed_a(0.0009916587732732296)),(to_sfixed_a(-0.00021943078900221735)),(to_sfixed_a(-0.0002403043763479218)),(to_sfixed_a(1.1980290764768142e-05)),(to_sfixed_a(-0.00045876012882217765)),(to_sfixed_a(-3.9039106923155487e-05)),(to_sfixed_a(-0.00011804982204921544)),(to_sfixed_a(-0.00010781749006127939)),(to_sfixed_a(-0.00044904660899192095)),(to_sfixed_a(0.0035403689835220575)),(to_sfixed_a(-0.0002945244195871055)),(to_sfixed_a(0.00019603371038101614)),(to_sfixed_a(0.005584534257650375)),(to_sfixed_a(-5.66349845030345e-05)),(to_sfixed_a(8.741274359636009e-05)),(to_sfixed_a(0.110594242811203)),(to_sfixed_a(-0.00013174483319744468)),(to_sfixed_a(-3.120761539321393e-05)),(to_sfixed_a(-4.1296323615824804e-05)),(to_sfixed_a(2.725647937040776e-05)),(to_sfixed_a(-6.884454342070967e-05)),(to_sfixed_a(0.00018789850582834333)),(to_sfixed_a(0.011079560965299606)),(to_sfixed_a(-0.0002737566828727722)),(to_sfixed_a(0.002615602919831872)),(to_sfixed_a(0.003029188374057412)),(to_sfixed_a(-0.0001067468838300556)),(to_sfixed_a(-0.21946598589420319)),(to_sfixed_a(0.000239882298046723)),(to_sfixed_a(-0.00015284294204320759)),(to_sfixed_a(0.00010577149805612862)),(to_sfixed_a(0.0021484943572431803)),(to_sfixed_a(0.0017071921611204743)),(to_sfixed_a(4.424805229064077e-05)),(to_sfixed_a(0.0033017368987202644)),(to_sfixed_a(0.0003378767869435251)),(to_sfixed_a(-0.0009182203793898225)),(to_sfixed_a(0.0008465484715998173)),(to_sfixed_a(0.030966462567448616)),(to_sfixed_a(-0.0001663801376707852)),(to_sfixed_a(-0.001495556440204382)),(to_sfixed_a(0.008268150500953197)),(to_sfixed_a(-5.678509478457272e-05)),(to_sfixed_a(4.5736393076367676e-05)),(to_sfixed_a(-0.00011263163469266146)),(to_sfixed_a(-0.000549072865396738)),(to_sfixed_a(0.001315227011218667)),(to_sfixed_a(-0.0009180563502013683)),(to_sfixed_a(3.65300802513957e-05)),(to_sfixed_a(0.00011240683670621365)),(to_sfixed_a(-2.5928588001988828e-05)),(to_sfixed_a(6.920780288055539e-05)),(to_sfixed_a(0.004534376319497824)),(to_sfixed_a(0.0004116272903047502)),(to_sfixed_a(-0.00015998497838154435)),(to_sfixed_a(0.006424945313483477)),(to_sfixed_a(0.0001370281825074926)),(to_sfixed_a(0.3297640085220337)),(to_sfixed_a(0.00429786229506135)),(to_sfixed_a(-1.211209746543318e-05)),(to_sfixed_a(0.0002186103374697268)),(to_sfixed_a(-5.9093727031722665e-06)),(to_sfixed_a(-2.8493115678429604e-05)),(to_sfixed_a(-0.00024217639293055981)),(to_sfixed_a(-0.00022197648650035262)),(to_sfixed_a(0.0025895971339195967)),(to_sfixed_a(0.23448817431926727)),(to_sfixed_a(0.30315855145454407)),(to_sfixed_a(-0.029194099828600883)),(to_sfixed_a(-0.0017125641461461782)),(to_sfixed_a(0.001983123831450939)),(to_sfixed_a(-5.5561045883223414e-05)),(to_sfixed_a(3.8135884096845984e-05)),(to_sfixed_a(7.122757961042225e-05)),(to_sfixed_a(-0.00013621035031974316)),(to_sfixed_a(0.00013868248788639903)),(to_sfixed_a(0.00014557907707057893)),(to_sfixed_a(0.0016149289440363646)),(to_sfixed_a(-0.0003510660899337381)),(to_sfixed_a(-6.274646875681356e-05)),(to_sfixed_a(5.7602301239967346e-05)),(to_sfixed_a(-9.061252058017999e-06)),(to_sfixed_a(5.6996403145603836e-05)),(to_sfixed_a(0.29087215662002563)),(to_sfixed_a(0.37924614548683167)),(to_sfixed_a(-0.0001919036149047315)),(to_sfixed_a(4.115277261007577e-05)),(to_sfixed_a(0.00019520011846907437)),(to_sfixed_a(0.0015124842757359147)),(to_sfixed_a(0.22960177063941956)),(to_sfixed_a(-0.0025891170371323824)),(to_sfixed_a(-8.620700100436807e-07)),(to_sfixed_a(-0.0002174425608245656)),(to_sfixed_a(0.0002881533873733133)),(to_sfixed_a(0.0029819600749760866)),(to_sfixed_a(-0.00041278719436377287)),(to_sfixed_a(0.010216306895017624)),(to_sfixed_a(0.00015657389303669333)),(to_sfixed_a(-0.00011678635200951248)),(to_sfixed_a(0.00014345849922392517)),(to_sfixed_a(0.000686502200551331)),(to_sfixed_a(-0.0002843828115146607)),(to_sfixed_a(-0.016351943835616112)),(to_sfixed_a(-0.00014233925321605057)),(to_sfixed_a(-0.36457425355911255)),(to_sfixed_a(-0.00033745390828698874)),(to_sfixed_a(0.0006165255908854306)),(to_sfixed_a(0.0009415795793756843)),(to_sfixed_a(-0.0001443721994291991)),(to_sfixed_a(0.0008666125941090286)),(to_sfixed_a(0.00018274672038387507)),(to_sfixed_a(0.0004110482113901526)),(to_sfixed_a(-0.00047333622933365405)),(to_sfixed_a(-0.0001474725577281788)),(to_sfixed_a(-0.00045588024659082294)),(to_sfixed_a(0.008566346019506454)),(to_sfixed_a(-0.0016668590251356363)),(to_sfixed_a(8.884555427357554e-06)),(to_sfixed_a(-6.980048055993393e-05)),(to_sfixed_a(0.009630112908780575)),(to_sfixed_a(5.7128963817376643e-05)),(to_sfixed_a(-0.0016044043004512787)),(to_sfixed_a(-0.00011412890307838097)),(to_sfixed_a(-0.0011577238328754902)),(to_sfixed_a(0.00019109167624264956)),(to_sfixed_a(0.005949580576270819)),(to_sfixed_a(2.5905887014232576e-05)),(to_sfixed_a(0.00015572598204016685)),(to_sfixed_a(1.013074506772682e-05)),(to_sfixed_a(0.0009208493283949792)),(to_sfixed_a(0.003981187008321285)),(to_sfixed_a(-0.00017205390031449497)),(to_sfixed_a(2.9486101993825287e-05)),(to_sfixed_a(-4.435762093635276e-06)),(to_sfixed_a(9.860369027592242e-05)),(to_sfixed_a(0.0053454916924238205)),(to_sfixed_a(-0.20170927047729492)),(to_sfixed_a(0.0007554280455224216)),(to_sfixed_a(0.0027386248111724854)),(to_sfixed_a(-0.0023781706113368273)),(to_sfixed_a(-3.738316081580706e-05)),(to_sfixed_a(7.934014138299972e-05)),(to_sfixed_a(-0.0004455870948731899)),(to_sfixed_a(-0.0011660639429464936)),(to_sfixed_a(-6.763963028788567e-05)),(to_sfixed_a(0.00030140415765345097)),(to_sfixed_a(-0.0002386566047789529)),(to_sfixed_a(0.5089545845985413)),(to_sfixed_a(0.00010062688670586795)),(to_sfixed_a(0.3045128583908081)),(to_sfixed_a(-0.0005052300402894616)),(to_sfixed_a(0.0030574235133826733)),(to_sfixed_a(0.007432727143168449)),(to_sfixed_a(-0.00018235872266814113)),(to_sfixed_a(0.21668507158756256)),(to_sfixed_a(0.00011014474875992164)),(to_sfixed_a(-0.0005572510999627411)),(to_sfixed_a(-5.789388524135575e-05)),(to_sfixed_a(0.002471936633810401)),(to_sfixed_a(-0.40058261156082153)),(to_sfixed_a(0.0032409951090812683)));

    constant weight_n2_72 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.03376784920692444)),(to_sfixed_a(0.32538902759552)),(to_sfixed_a(0.18471331894397736)),(to_sfixed_a(0.00021240323258098215)),(to_sfixed_a(-0.007667138706892729)),(to_sfixed_a(-0.00023684589541517198)),(to_sfixed_a(-0.0022543154191225767)),(to_sfixed_a(-5.456844519358128e-06)),(to_sfixed_a(0.00011470923345768824)),(to_sfixed_a(-0.00014937650121282786)),(to_sfixed_a(-1.028574479278177e-05)),(to_sfixed_a(-0.014584130607545376)),(to_sfixed_a(-0.002899260027334094)),(to_sfixed_a(-0.00013960438081994653)),(to_sfixed_a(-7.838382589397952e-05)),(to_sfixed_a(-0.0002002236433327198)),(to_sfixed_a(0.0013737054541707039)),(to_sfixed_a(6.588229007320479e-05)),(to_sfixed_a(0.005088410340249538)),(to_sfixed_a(0.0015656366012990475)),(to_sfixed_a(-0.0001275358663406223)),(to_sfixed_a(-2.8695849323412403e-05)),(to_sfixed_a(8.280493784695864e-05)),(to_sfixed_a(0.006659494247287512)),(to_sfixed_a(-0.006207022815942764)),(to_sfixed_a(-0.001302359509281814)),(to_sfixed_a(-0.00018169675604440272)),(to_sfixed_a(0.0006071508396416903)),(to_sfixed_a(0.0003465065383352339)),(to_sfixed_a(-4.625648580258712e-05)),(to_sfixed_a(-0.001004425110295415)),(to_sfixed_a(-6.821005081292242e-05)),(to_sfixed_a(0.005009246990084648)),(to_sfixed_a(-0.00010085711983265355)),(to_sfixed_a(-0.00011833137250505388)),(to_sfixed_a(-2.964909072034061e-06)),(to_sfixed_a(0.20528879761695862)),(to_sfixed_a(0.01849181391298771)),(to_sfixed_a(-0.02470952272415161)),(to_sfixed_a(-0.00018360874673817307)),(to_sfixed_a(0.0009625709499232471)),(to_sfixed_a(6.0960395785514265e-05)),(to_sfixed_a(4.717505362350494e-06)),(to_sfixed_a(0.00022161102970130742)),(to_sfixed_a(-0.013788055628538132)),(to_sfixed_a(-0.013553480617702007)),(to_sfixed_a(0.000682633079122752)),(to_sfixed_a(-0.005704923532903194)),(to_sfixed_a(4.98828012496233e-06)),(to_sfixed_a(-0.005146434996277094)),(to_sfixed_a(-0.0015767294680699706)),(to_sfixed_a(-5.316847818903625e-06)),(to_sfixed_a(1.056285691447556e-05)),(to_sfixed_a(5.200070881983265e-05)),(to_sfixed_a(-0.01570403389632702)),(to_sfixed_a(0.0030505747999995947)),(to_sfixed_a(0.00014883668336551636)),(to_sfixed_a(-0.016481716185808182)),(to_sfixed_a(3.804365042014979e-05)),(to_sfixed_a(-0.00015551589604001492)),(to_sfixed_a(-0.011400808580219746)),(to_sfixed_a(-0.0021891717333346605)),(to_sfixed_a(-0.0009370885672979057)),(to_sfixed_a(0.35442158579826355)),(to_sfixed_a(7.080085924826562e-05)),(to_sfixed_a(-0.001984243281185627)),(to_sfixed_a(-0.00019504287047311664)),(to_sfixed_a(0.04931700602173805)),(to_sfixed_a(-0.0002252942358609289)),(to_sfixed_a(-5.650187813444063e-05)),(to_sfixed_a(0.01429660338908434)),(to_sfixed_a(0.0012267460115253925)),(to_sfixed_a(0.005359850358217955)),(to_sfixed_a(-0.00013401043543126434)),(to_sfixed_a(-0.00023328234965447336)),(to_sfixed_a(-7.049127452773973e-05)),(to_sfixed_a(-0.4162960946559906)),(to_sfixed_a(0.3607979118824005)),(to_sfixed_a(1.275792601518333e-05)),(to_sfixed_a(0.012742401100695133)),(to_sfixed_a(-0.009831557981669903)),(to_sfixed_a(-1.954461185960099e-05)),(to_sfixed_a(0.46651700139045715)),(to_sfixed_a(-0.001840225886553526)),(to_sfixed_a(-0.00010087640839628875)),(to_sfixed_a(0.00748463673517108)),(to_sfixed_a(-0.0008422020473517478)),(to_sfixed_a(0.0017779483459889889)),(to_sfixed_a(0.0002516638778615743)),(to_sfixed_a(7.048206316540018e-05)),(to_sfixed_a(-0.012686043977737427)),(to_sfixed_a(-3.6072760849492624e-05)),(to_sfixed_a(-0.005971561186015606)),(to_sfixed_a(-2.9334798455238342e-05)),(to_sfixed_a(0.04501976817846298)),(to_sfixed_a(2.5265639123972505e-05)),(to_sfixed_a(0.0001489425776526332)),(to_sfixed_a(-4.733716923510656e-05)),(to_sfixed_a(-7.110301521606743e-05)),(to_sfixed_a(0.00020008068531751633)),(to_sfixed_a(-0.002676416886970401)),(to_sfixed_a(0.002941317390650511)),(to_sfixed_a(0.0002116963005391881)),(to_sfixed_a(0.001082350267097354)),(to_sfixed_a(0.0005763547378592193)),(to_sfixed_a(-0.002542453818023205)),(to_sfixed_a(4.3090403778478503e-07)),(to_sfixed_a(-4.916290345136076e-05)),(to_sfixed_a(-0.0001513720053480938)),(to_sfixed_a(0.0028540324419736862)),(to_sfixed_a(0.002386373933404684)),(to_sfixed_a(-0.000319607846904546)),(to_sfixed_a(0.37697333097457886)),(to_sfixed_a(0.00015029881615191698)),(to_sfixed_a(-1.2877731933258474e-05)),(to_sfixed_a(0.0028496405575424433)),(to_sfixed_a(0.008970912545919418)),(to_sfixed_a(-0.003338045673444867)),(to_sfixed_a(-1.422091736458242e-05)),(to_sfixed_a(0.0003703833499457687)),(to_sfixed_a(-0.00014413168537430465)),(to_sfixed_a(-0.0002943685685750097)),(to_sfixed_a(0.40639981627464294)),(to_sfixed_a(-4.245017407811247e-05)),(to_sfixed_a(0.0001557570940349251)),(to_sfixed_a(-0.0022270865738391876)),(to_sfixed_a(-0.0037113858852535486)),(to_sfixed_a(0.0002612223324831575)),(to_sfixed_a(-0.0003123139322269708)),(to_sfixed_a(-6.342925189528614e-07)),(to_sfixed_a(-2.986927211168222e-05)),(to_sfixed_a(8.610928489360958e-06)),(to_sfixed_a(-7.211350020952523e-05)),(to_sfixed_a(-0.005209416151046753)),(to_sfixed_a(0.0002849109878297895)),(to_sfixed_a(0.00011642474419204518)),(to_sfixed_a(-0.016492819413542747)),(to_sfixed_a(-0.0002066157612716779)),(to_sfixed_a(-0.00014835043111816049)),(to_sfixed_a(1.3800148735754192e-05)),(to_sfixed_a(0.22839486598968506)),(to_sfixed_a(5.6085809774231166e-06)),(to_sfixed_a(-0.0002986521867569536)),(to_sfixed_a(0.004328875336796045)),(to_sfixed_a(-0.0028962513897567987)),(to_sfixed_a(0.004348854534327984)),(to_sfixed_a(-0.0015904189785942435)),(to_sfixed_a(0.00011237481521675363)),(to_sfixed_a(-0.00023734082060400397)),(to_sfixed_a(-0.00895608589053154)),(to_sfixed_a(-2.3381522623822093e-05)),(to_sfixed_a(0.00015440437709912658)),(to_sfixed_a(0.00784937385469675)),(to_sfixed_a(-4.461963544599712e-05)),(to_sfixed_a(-1.1212196113774553e-06)),(to_sfixed_a(-0.0024108721408993006)),(to_sfixed_a(-0.00041593058267608285)),(to_sfixed_a(-3.248808206990361e-05)),(to_sfixed_a(-0.00017748857499100268)),(to_sfixed_a(3.222384111722931e-05)),(to_sfixed_a(4.020577762275934e-06)),(to_sfixed_a(0.000247310585109517)),(to_sfixed_a(0.007273424416780472)),(to_sfixed_a(-0.0027948827482759953)),(to_sfixed_a(-0.0033552993554621935)),(to_sfixed_a(0.008694066666066647)),(to_sfixed_a(-0.00015441939467564225)),(to_sfixed_a(0.004764455370604992)),(to_sfixed_a(-0.0002439470263198018)),(to_sfixed_a(5.878355295863003e-07)),(to_sfixed_a(-0.011097948998212814)),(to_sfixed_a(-0.0002446948201395571)),(to_sfixed_a(-0.0023420609068125486)),(to_sfixed_a(2.7107831556349993e-05)),(to_sfixed_a(-0.2745296061038971)),(to_sfixed_a(-0.001384971896186471)),(to_sfixed_a(-0.00013684443547390401)),(to_sfixed_a(-0.002347630448639393)),(to_sfixed_a(0.008565523661673069)),(to_sfixed_a(-0.011674159206449986)),(to_sfixed_a(-0.0009445277391932905)),(to_sfixed_a(0.016578763723373413)),(to_sfixed_a(5.732747376896441e-05)),(to_sfixed_a(3.592365828808397e-05)),(to_sfixed_a(0.0001562477700645104)),(to_sfixed_a(-0.004594453610479832)),(to_sfixed_a(-0.005342586897313595)),(to_sfixed_a(0.006145352963358164)),(to_sfixed_a(-0.00030340757803060114)),(to_sfixed_a(-0.0005844865227118134)),(to_sfixed_a(0.007851775735616684)),(to_sfixed_a(-0.00013718963600695133)),(to_sfixed_a(-9.394971129950136e-05)),(to_sfixed_a(0.0016544387908652425)),(to_sfixed_a(2.868819865398109e-05)),(to_sfixed_a(0.011148128658533096)),(to_sfixed_a(0.00012713903561234474)),(to_sfixed_a(-0.30756473541259766)),(to_sfixed_a(-0.008377481251955032)),(to_sfixed_a(0.0001272635709028691)),(to_sfixed_a(0.0001531880407128483)),(to_sfixed_a(-0.00010326967458240688)),(to_sfixed_a(3.37259225489106e-05)),(to_sfixed_a(-1.566046557854861e-05)),(to_sfixed_a(0.00014649747754447162)),(to_sfixed_a(0.24774612486362457)),(to_sfixed_a(-0.0029052505269646645)),(to_sfixed_a(0.0016813846305012703)),(to_sfixed_a(-0.0009635672904551029)),(to_sfixed_a(-0.0012586787343025208)),(to_sfixed_a(0.003979164641350508)),(to_sfixed_a(-4.31919761467725e-06)),(to_sfixed_a(-5.644520570058376e-06)),(to_sfixed_a(-0.00010985838162014261)),(to_sfixed_a(-0.0001989408629015088)),(to_sfixed_a(-0.00014311181439552456)),(to_sfixed_a(-0.0004660828853957355)),(to_sfixed_a(0.00031343073351308703)),(to_sfixed_a(-0.001167083391919732)),(to_sfixed_a(-2.9743478080490604e-05)),(to_sfixed_a(6.240999209694564e-05)),(to_sfixed_a(-2.953000512206927e-05)),(to_sfixed_a(-0.00013689174375031143)),(to_sfixed_a(0.29063206911087036)),(to_sfixed_a(-0.005492720752954483)),(to_sfixed_a(7.633803761564195e-06)),(to_sfixed_a(-0.00016808792133815587)),(to_sfixed_a(-0.00015444440941791981)),(to_sfixed_a(-0.34061485528945923)),(to_sfixed_a(-0.0003168111725244671)),(to_sfixed_a(-0.002585489070042968)),(to_sfixed_a(0.0002879348467104137)),(to_sfixed_a(-0.0001913346495712176)),(to_sfixed_a(6.584259972441941e-05)),(to_sfixed_a(-0.0014377186307683587)),(to_sfixed_a(0.010609699413180351)),(to_sfixed_a(0.0028094439767301083)),(to_sfixed_a(-9.645873797126114e-05)),(to_sfixed_a(-0.005981996189802885)),(to_sfixed_a(0.00027098413556814194)),(to_sfixed_a(-0.009963431395590305)),(to_sfixed_a(0.0001914385356940329)),(to_sfixed_a(0.0032617757096886635)),(to_sfixed_a(-8.102157153189182e-06)),(to_sfixed_a(0.004454857669770718)),(to_sfixed_a(-0.0008365956600755453)),(to_sfixed_a(-0.31951746344566345)),(to_sfixed_a(0.5260167717933655)),(to_sfixed_a(3.1081526685738936e-05)),(to_sfixed_a(-0.015524414367973804)),(to_sfixed_a(-0.019921978935599327)),(to_sfixed_a(-3.551200279616751e-05)),(to_sfixed_a(-0.0010279510170221329)),(to_sfixed_a(-0.00020408135605975986)),(to_sfixed_a(0.0002164213510695845)),(to_sfixed_a(0.17884740233421326)),(to_sfixed_a(-0.0027659954503178596)),(to_sfixed_a(9.835488890530542e-05)),(to_sfixed_a(0.00022727533360011876)),(to_sfixed_a(0.000718997442163527)),(to_sfixed_a(-0.00023782970674801618)),(to_sfixed_a(0.3570826053619385)),(to_sfixed_a(3.2128631573868915e-05)),(to_sfixed_a(0.0001248792978003621)),(to_sfixed_a(9.812566713662818e-05)),(to_sfixed_a(0.007049154955893755)),(to_sfixed_a(-0.00020609052444342524)),(to_sfixed_a(-0.00041684129973873496)),(to_sfixed_a(6.679049693048e-05)),(to_sfixed_a(-0.009180126711726189)),(to_sfixed_a(0.5088933110237122)),(to_sfixed_a(-2.2918084141565487e-05)),(to_sfixed_a(-6.278615182964131e-05)),(to_sfixed_a(0.00015477077977266163)),(to_sfixed_a(-9.30573878576979e-06)),(to_sfixed_a(0.2245389074087143)),(to_sfixed_a(-0.020739654079079628)),(to_sfixed_a(-0.002891230396926403)),(to_sfixed_a(-0.3433953523635864)),(to_sfixed_a(-0.004084968939423561)),(to_sfixed_a(-0.00014610920334234834)),(to_sfixed_a(-0.0001833986898418516)),(to_sfixed_a(2.652819239301607e-05)),(to_sfixed_a(0.0007485910318791866)),(to_sfixed_a(-0.00021378116798587143)),(to_sfixed_a(-3.510285750962794e-06)),(to_sfixed_a(-0.0004300115106161684)),(to_sfixed_a(0.007644008379429579)),(to_sfixed_a(-6.693102477584034e-06)),(to_sfixed_a(0.0007618390955030918)),(to_sfixed_a(-0.0009060350130312145)),(to_sfixed_a(-0.013679110445082188)),(to_sfixed_a(-0.008351901546120644)),(to_sfixed_a(-5.374874308472499e-05)),(to_sfixed_a(-0.0015453477390110493)),(to_sfixed_a(0.28485628962516785)),(to_sfixed_a(-0.018498579040169716)),(to_sfixed_a(-0.00017788115656003356)),(to_sfixed_a(0.0025032954290509224)),(to_sfixed_a(0.41213560104370117)),(to_sfixed_a(0.19252461194992065)));

    constant weight_n2_73 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.07130806148052216)),(to_sfixed_a(-0.26704010367393494)),(to_sfixed_a(-2.3597394829266705e-06)),(to_sfixed_a(-0.00017453302280046046)),(to_sfixed_a(0.00682141724973917)),(to_sfixed_a(-6.313979247352108e-05)),(to_sfixed_a(0.008875396102666855)),(to_sfixed_a(4.2401617974974215e-05)),(to_sfixed_a(-0.0001817286538425833)),(to_sfixed_a(-0.0004124436527490616)),(to_sfixed_a(-0.0002984104212373495)),(to_sfixed_a(0.0006435967516154051)),(to_sfixed_a(-0.32106420397758484)),(to_sfixed_a(0.0029771612025797367)),(to_sfixed_a(-7.420232577715069e-06)),(to_sfixed_a(2.076192140521016e-05)),(to_sfixed_a(0.20288033783435822)),(to_sfixed_a(-0.00031215621856972575)),(to_sfixed_a(-0.0015368008753284812)),(to_sfixed_a(0.2482903152704239)),(to_sfixed_a(-6.12640506005846e-05)),(to_sfixed_a(-2.900187246268615e-05)),(to_sfixed_a(-0.00023013379541225731)),(to_sfixed_a(0.12862376868724823)),(to_sfixed_a(-0.0025175740011036396)),(to_sfixed_a(0.1003788486123085)),(to_sfixed_a(0.00015623764193151146)),(to_sfixed_a(-0.0009459140710532665)),(to_sfixed_a(0.002323969267308712)),(to_sfixed_a(6.273999315453693e-05)),(to_sfixed_a(0.20548318326473236)),(to_sfixed_a(-2.8105132514610887e-05)),(to_sfixed_a(0.001930215279571712)),(to_sfixed_a(1.7859434592537582e-05)),(to_sfixed_a(-9.799489635042846e-05)),(to_sfixed_a(0.0002221877221018076)),(to_sfixed_a(-0.024542363360524178)),(to_sfixed_a(-0.004538557957857847)),(to_sfixed_a(-0.29012900590896606)),(to_sfixed_a(6.945141649339348e-05)),(to_sfixed_a(0.00514985341578722)),(to_sfixed_a(-0.0002143307647202164)),(to_sfixed_a(-0.000175316323293373)),(to_sfixed_a(0.0003129582619294524)),(to_sfixed_a(0.003181843552738428)),(to_sfixed_a(-0.10727415978908539)),(to_sfixed_a(0.0010172968031838536)),(to_sfixed_a(0.008264485746622086)),(to_sfixed_a(9.246095578419045e-05)),(to_sfixed_a(0.005396845750510693)),(to_sfixed_a(-0.0032480645459145308)),(to_sfixed_a(-4.459930642042309e-05)),(to_sfixed_a(-5.24161514476873e-05)),(to_sfixed_a(-0.0007170190801844001)),(to_sfixed_a(0.007323772646486759)),(to_sfixed_a(7.537448254879564e-05)),(to_sfixed_a(-8.39243657537736e-05)),(to_sfixed_a(0.004168810322880745)),(to_sfixed_a(0.00024982314789667726)),(to_sfixed_a(-4.5036427763989195e-05)),(to_sfixed_a(0.001427941839210689)),(to_sfixed_a(0.0008593745296820998)),(to_sfixed_a(-0.0010556934867054224)),(to_sfixed_a(-0.08392495661973953)),(to_sfixed_a(-9.80374461505562e-05)),(to_sfixed_a(0.000902841507922858)),(to_sfixed_a(-5.49169271835126e-06)),(to_sfixed_a(0.004281917586922646)),(to_sfixed_a(-0.0002312695432920009)),(to_sfixed_a(0.0002841013192664832)),(to_sfixed_a(-0.008246603421866894)),(to_sfixed_a(-0.0006675086915493011)),(to_sfixed_a(-0.13312435150146484)),(to_sfixed_a(-0.00013025592488702387)),(to_sfixed_a(0.00022935058223083615)),(to_sfixed_a(-0.0001361090544378385)),(to_sfixed_a(-0.004346531815826893)),(to_sfixed_a(0.0039059482514858246)),(to_sfixed_a(9.241439329343848e-06)),(to_sfixed_a(0.0008664386114105582)),(to_sfixed_a(-0.00048384195542894304)),(to_sfixed_a(0.00018841135897673666)),(to_sfixed_a(0.000916977587621659)),(to_sfixed_a(-0.018208149820566177)),(to_sfixed_a(0.000119177253509406)),(to_sfixed_a(0.0005952522624284029)),(to_sfixed_a(-0.005670242942869663)),(to_sfixed_a(-8.899991371436045e-06)),(to_sfixed_a(-5.0789134547812864e-05)),(to_sfixed_a(2.110143395839259e-05)),(to_sfixed_a(0.0037640193477272987)),(to_sfixed_a(-9.425735697732307e-06)),(to_sfixed_a(-0.0007308035856112838)),(to_sfixed_a(-6.422807928174734e-05)),(to_sfixed_a(0.002449267776682973)),(to_sfixed_a(7.897950854385272e-05)),(to_sfixed_a(-0.00015361826808657497)),(to_sfixed_a(-1.5875826647970825e-05)),(to_sfixed_a(4.416420779307373e-05)),(to_sfixed_a(3.8337704609148204e-05)),(to_sfixed_a(0.22748565673828125)),(to_sfixed_a(0.001760168350301683)),(to_sfixed_a(-0.00023227071505971253)),(to_sfixed_a(0.0015826449962332845)),(to_sfixed_a(-0.4912002980709076)),(to_sfixed_a(-3.4622891689650714e-05)),(to_sfixed_a(-0.00022899534087628126)),(to_sfixed_a(-3.873818786814809e-05)),(to_sfixed_a(0.00010699018457671627)),(to_sfixed_a(0.007267562672495842)),(to_sfixed_a(0.005239322315901518)),(to_sfixed_a(0.0002383063838351518)),(to_sfixed_a(0.0009557788143865764)),(to_sfixed_a(1.6682904970366508e-05)),(to_sfixed_a(-0.0001588701270520687)),(to_sfixed_a(0.006152525078505278)),(to_sfixed_a(9.955401037586853e-05)),(to_sfixed_a(5.443789268610999e-05)),(to_sfixed_a(8.51900695124641e-05)),(to_sfixed_a(0.005020088516175747)),(to_sfixed_a(-0.00014949115575291216)),(to_sfixed_a(0.00012072952813468874)),(to_sfixed_a(-7.82954812166281e-05)),(to_sfixed_a(-0.0002557413827162236)),(to_sfixed_a(4.313907629693858e-05)),(to_sfixed_a(0.0004803033370990306)),(to_sfixed_a(0.00012745638377964497)),(to_sfixed_a(6.61585945636034e-05)),(to_sfixed_a(3.685614501591772e-05)),(to_sfixed_a(0.00021624029614031315)),(to_sfixed_a(-2.9369184630922973e-06)),(to_sfixed_a(1.892926957225427e-05)),(to_sfixed_a(-0.0004810998507309705)),(to_sfixed_a(0.25340116024017334)),(to_sfixed_a(-6.364576984196901e-05)),(to_sfixed_a(0.00011588800407480448)),(to_sfixed_a(0.007618474308401346)),(to_sfixed_a(0.00019441723998170346)),(to_sfixed_a(-1.3426142686512321e-06)),(to_sfixed_a(-0.0001519207435194403)),(to_sfixed_a(0.00023611553478986025)),(to_sfixed_a(-2.864505586330779e-05)),(to_sfixed_a(0.00017120313714258373)),(to_sfixed_a(0.0003037659334950149)),(to_sfixed_a(0.0016271035419777036)),(to_sfixed_a(0.0003128733078483492)),(to_sfixed_a(0.0002887172158807516)),(to_sfixed_a(-0.00019163276010658592)),(to_sfixed_a(0.0001297553681069985)),(to_sfixed_a(0.0002826626878231764)),(to_sfixed_a(-0.00016875640721991658)),(to_sfixed_a(-0.00015832402277737856)),(to_sfixed_a(-0.0009633708978071809)),(to_sfixed_a(2.9785282094962895e-05)),(to_sfixed_a(0.00013038062024861574)),(to_sfixed_a(-0.0004695864918176085)),(to_sfixed_a(-0.0003174608282279223)),(to_sfixed_a(-0.00030616563162766397)),(to_sfixed_a(0.00012260591029189527)),(to_sfixed_a(9.054798283614218e-06)),(to_sfixed_a(7.461186032742262e-05)),(to_sfixed_a(-7.155764615163207e-05)),(to_sfixed_a(-0.008048636838793755)),(to_sfixed_a(-0.00032825584639795125)),(to_sfixed_a(0.005019554868340492)),(to_sfixed_a(0.33421841263771057)),(to_sfixed_a(-1.6547062841709703e-05)),(to_sfixed_a(0.22900301218032837)),(to_sfixed_a(0.00020213487732689828)),(to_sfixed_a(3.0624898499809206e-05)),(to_sfixed_a(0.01338235568255186)),(to_sfixed_a(0.0010130192385986447)),(to_sfixed_a(-0.2653448283672333)),(to_sfixed_a(-4.093715688213706e-06)),(to_sfixed_a(0.2056272029876709)),(to_sfixed_a(8.617188723292202e-05)),(to_sfixed_a(0.0033470371272414923)),(to_sfixed_a(0.22881466150283813)),(to_sfixed_a(-0.2152204066514969)),(to_sfixed_a(0.3742925822734833)),(to_sfixed_a(0.0011830677976831794)),(to_sfixed_a(-0.004055663011968136)),(to_sfixed_a(5.4770312999607995e-05)),(to_sfixed_a(4.711386281996965e-06)),(to_sfixed_a(-0.000188946578418836)),(to_sfixed_a(0.0027849997859448195)),(to_sfixed_a(-0.0011514947982504964)),(to_sfixed_a(0.0005882684490643442)),(to_sfixed_a(0.00016871021944098175)),(to_sfixed_a(1.969098229892552e-05)),(to_sfixed_a(-0.000637347751762718)),(to_sfixed_a(-2.7130772650707513e-05)),(to_sfixed_a(-0.021713314577937126)),(to_sfixed_a(-0.0007401997572742403)),(to_sfixed_a(-9.287259308621287e-05)),(to_sfixed_a(0.22211405634880066)),(to_sfixed_a(-0.0002270608238177374)),(to_sfixed_a(0.0024672141298651695)),(to_sfixed_a(-0.0025088859256356955)),(to_sfixed_a(-0.00015366119623649865)),(to_sfixed_a(9.865726315183565e-05)),(to_sfixed_a(0.00013075940660201013)),(to_sfixed_a(-0.00014908172306604683)),(to_sfixed_a(-6.129402026999742e-05)),(to_sfixed_a(-0.00013044934894423932)),(to_sfixed_a(0.00040250126039609313)),(to_sfixed_a(-0.015197383239865303)),(to_sfixed_a(-2.646265784278512e-07)),(to_sfixed_a(0.002942065242677927)),(to_sfixed_a(0.00045609555672854185)),(to_sfixed_a(-0.022829586640000343)),(to_sfixed_a(-0.00021927172201685607)),(to_sfixed_a(0.0003065411583520472)),(to_sfixed_a(-0.00010247281170450151)),(to_sfixed_a(-0.00013530692376662046)),(to_sfixed_a(0.0003173867880832404)),(to_sfixed_a(-0.0016933006700128317)),(to_sfixed_a(0.19271770119667053)),(to_sfixed_a(-0.003541266079992056)),(to_sfixed_a(-2.315106030437164e-05)),(to_sfixed_a(7.459201151505113e-05)),(to_sfixed_a(0.00028667712467722595)),(to_sfixed_a(0.00029443245148286223)),(to_sfixed_a(-0.0006700289668515325)),(to_sfixed_a(-0.007707191631197929)),(to_sfixed_a(-8.315212471643463e-05)),(to_sfixed_a(-1.0761134035419673e-05)),(to_sfixed_a(-0.00023603433510288596)),(to_sfixed_a(0.01799880713224411)),(to_sfixed_a(0.008350202813744545)),(to_sfixed_a(-9.807484457269311e-05)),(to_sfixed_a(8.121787686832249e-08)),(to_sfixed_a(-6.43891398794949e-05)),(to_sfixed_a(-8.882839028956369e-05)),(to_sfixed_a(0.0007029480184428394)),(to_sfixed_a(0.25898998975753784)),(to_sfixed_a(0.0026228672359138727)),(to_sfixed_a(0.00027015211526304483)),(to_sfixed_a(-9.301802492700517e-05)),(to_sfixed_a(-2.2241132683120668e-05)),(to_sfixed_a(0.00269195344299078)),(to_sfixed_a(-6.466647027991712e-05)),(to_sfixed_a(0.003379769390448928)),(to_sfixed_a(-6.354377546813339e-06)),(to_sfixed_a(0.22092922031879425)),(to_sfixed_a(-0.0010024415096268058)),(to_sfixed_a(0.31076779961586)),(to_sfixed_a(-0.1442326456308365)),(to_sfixed_a(-9.094210690818727e-05)),(to_sfixed_a(0.0031984683591872454)),(to_sfixed_a(0.016535060480237007)),(to_sfixed_a(-1.345520286122337e-05)),(to_sfixed_a(-0.0002369120775256306)),(to_sfixed_a(-0.00014731734700035304)),(to_sfixed_a(-1.1179072316735983e-05)),(to_sfixed_a(0.0012798457173630595)),(to_sfixed_a(0.004455338232219219)),(to_sfixed_a(-2.2317391994874924e-05)),(to_sfixed_a(-0.00014657391875516623)),(to_sfixed_a(-0.00043045729398727417)),(to_sfixed_a(-0.00029142946004867554)),(to_sfixed_a(0.0025574597530066967)),(to_sfixed_a(-0.00024046497128438205)),(to_sfixed_a(-0.00011826119589386508)),(to_sfixed_a(0.00015097497089300305)),(to_sfixed_a(0.007802373263984919)),(to_sfixed_a(6.443161692004651e-05)),(to_sfixed_a(4.052784061059356e-05)),(to_sfixed_a(7.941125659272075e-07)),(to_sfixed_a(0.19939257204532623)),(to_sfixed_a(-0.010047322139143944)),(to_sfixed_a(-6.30506910965778e-05)),(to_sfixed_a(-0.00013832340482622385)),(to_sfixed_a(3.3630276448093355e-05)),(to_sfixed_a(-2.9526723665185273e-05)),(to_sfixed_a(4.299533611629158e-05)),(to_sfixed_a(0.010258854366838932)),(to_sfixed_a(0.0042177606374025345)),(to_sfixed_a(0.003952110186219215)),(to_sfixed_a(-0.002210106234997511)),(to_sfixed_a(-5.728251562686637e-05)),(to_sfixed_a(7.969517901074141e-05)),(to_sfixed_a(0.00013606503489427269)),(to_sfixed_a(-0.00012601003982126713)),(to_sfixed_a(-0.00013526080874726176)),(to_sfixed_a(0.00015559679013676941)),(to_sfixed_a(-0.31866586208343506)),(to_sfixed_a(-0.3293604254722595)),(to_sfixed_a(-0.00016597307694610208)),(to_sfixed_a(5.187372153159231e-05)),(to_sfixed_a(-0.03950994089245796)),(to_sfixed_a(0.0064814286306500435)),(to_sfixed_a(-0.00037932873237878084)),(to_sfixed_a(-0.0002870935422834009)),(to_sfixed_a(-5.438185326056555e-05)),(to_sfixed_a(0.015260054729878902)),(to_sfixed_a(0.006979756988584995)),(to_sfixed_a(-6.674964242847636e-05)),(to_sfixed_a(-0.0041160280816257)),(to_sfixed_a(-0.004910647869110107)),(to_sfixed_a(-0.12547838687896729)));

    constant weight_n2_74 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.23064076900482178)),(to_sfixed_a(0.005530684720724821)),(to_sfixed_a(0.3559834659099579)),(to_sfixed_a(0.00015378493117168546)),(to_sfixed_a(-0.0005082066054455936)),(to_sfixed_a(0.00010695469245547429)),(to_sfixed_a(0.0037707118317484856)),(to_sfixed_a(-0.00013506911636795849)),(to_sfixed_a(-4.582786641549319e-05)),(to_sfixed_a(-0.0002745077945291996)),(to_sfixed_a(-0.0004189334867987782)),(to_sfixed_a(0.013733625411987305)),(to_sfixed_a(-0.003144201124086976)),(to_sfixed_a(-0.008506955578923225)),(to_sfixed_a(-0.0001352991530438885)),(to_sfixed_a(1.920527938636951e-05)),(to_sfixed_a(0.004822126589715481)),(to_sfixed_a(0.00011283579806331545)),(to_sfixed_a(-0.011965567246079445)),(to_sfixed_a(-0.002921930281445384)),(to_sfixed_a(-0.00018313087639398873)),(to_sfixed_a(-0.00012847153993789107)),(to_sfixed_a(0.0009669377468526363)),(to_sfixed_a(-0.44657382369041443)),(to_sfixed_a(0.002006084192544222)),(to_sfixed_a(-0.004918654449284077)),(to_sfixed_a(7.938557246234268e-05)),(to_sfixed_a(0.0001404552604071796)),(to_sfixed_a(-0.006617048289626837)),(to_sfixed_a(0.0001843203790485859)),(to_sfixed_a(0.0136239780113101)),(to_sfixed_a(2.1684900275431573e-05)),(to_sfixed_a(0.002052046125754714)),(to_sfixed_a(-0.0001291548542212695)),(to_sfixed_a(0.00011453318438725546)),(to_sfixed_a(-0.0001318576978519559)),(to_sfixed_a(0.309767484664917)),(to_sfixed_a(0.17363309860229492)),(to_sfixed_a(0.0006330403848551214)),(to_sfixed_a(-0.00021317516802810133)),(to_sfixed_a(-0.12160447984933853)),(to_sfixed_a(-0.00028506090166047215)),(to_sfixed_a(-0.00012991385301575065)),(to_sfixed_a(-6.183836376294494e-06)),(to_sfixed_a(0.005311725661158562)),(to_sfixed_a(0.38597822189331055)),(to_sfixed_a(0.07687804847955704)),(to_sfixed_a(-0.00034505611984059215)),(to_sfixed_a(0.0002830014855135232)),(to_sfixed_a(-0.004873222671449184)),(to_sfixed_a(-0.0040253582410514355)),(to_sfixed_a(7.059129711706191e-05)),(to_sfixed_a(5.650726961903274e-06)),(to_sfixed_a(-0.002793853636831045)),(to_sfixed_a(0.02401728741824627)),(to_sfixed_a(-0.001379271736368537)),(to_sfixed_a(-0.0001898840127978474)),(to_sfixed_a(0.0073906672187149525)),(to_sfixed_a(-0.0001300627482123673)),(to_sfixed_a(7.523042586399242e-05)),(to_sfixed_a(0.0033152520190924406)),(to_sfixed_a(0.0004465834645088762)),(to_sfixed_a(-0.4036240577697754)),(to_sfixed_a(0.009675135836005211)),(to_sfixed_a(5.8318692026659846e-05)),(to_sfixed_a(-0.0029504098929464817)),(to_sfixed_a(0.00045824304106645286)),(to_sfixed_a(-0.005474405363202095)),(to_sfixed_a(0.0011548695620149374)),(to_sfixed_a(-1.924347088788636e-05)),(to_sfixed_a(0.0013686256716027856)),(to_sfixed_a(-0.007842881605029106)),(to_sfixed_a(0.0014240742893889546)),(to_sfixed_a(-0.00010916498285951093)),(to_sfixed_a(-6.772697088308632e-05)),(to_sfixed_a(0.00020515196956694126)),(to_sfixed_a(0.028135504573583603)),(to_sfixed_a(4.2416078940732405e-05)),(to_sfixed_a(5.7643832406029105e-05)),(to_sfixed_a(0.31811556220054626)),(to_sfixed_a(0.0024342602118849754)),(to_sfixed_a(-2.3557011445518583e-05)),(to_sfixed_a(0.31103813648223877)),(to_sfixed_a(-0.0004926291876472533)),(to_sfixed_a(-0.00012901278387289494)),(to_sfixed_a(-0.23373648524284363)),(to_sfixed_a(0.24438069760799408)),(to_sfixed_a(0.2458333522081375)),(to_sfixed_a(1.1549476766958833e-05)),(to_sfixed_a(1.5229554264806211e-05)),(to_sfixed_a(0.009149564430117607)),(to_sfixed_a(-1.0651338016032241e-05)),(to_sfixed_a(0.003649370511993766)),(to_sfixed_a(6.429114728234708e-05)),(to_sfixed_a(0.38684991002082825)),(to_sfixed_a(-9.099789167521521e-05)),(to_sfixed_a(-0.0002877347287721932)),(to_sfixed_a(-0.0004147042927797884)),(to_sfixed_a(3.836306859739125e-05)),(to_sfixed_a(3.18843376589939e-05)),(to_sfixed_a(0.004675497300922871)),(to_sfixed_a(0.008476161397993565)),(to_sfixed_a(-7.071242725942284e-05)),(to_sfixed_a(0.2688484489917755)),(to_sfixed_a(0.382743239402771)),(to_sfixed_a(-0.0005599490250460804)),(to_sfixed_a(-2.5203880795743316e-05)),(to_sfixed_a(-0.000101189871202223)),(to_sfixed_a(0.0002218517620349303)),(to_sfixed_a(-0.39921867847442627)),(to_sfixed_a(-0.4480993449687958)),(to_sfixed_a(-3.7548874388448894e-05)),(to_sfixed_a(0.09794791787862778)),(to_sfixed_a(3.904060577042401e-07)),(to_sfixed_a(-0.00030803499976173043)),(to_sfixed_a(0.0056396592408418655)),(to_sfixed_a(0.006738022901117802)),(to_sfixed_a(-0.0004050515126436949)),(to_sfixed_a(-0.00045794836478307843)),(to_sfixed_a(0.17076702415943146)),(to_sfixed_a(-3.25428118230775e-06)),(to_sfixed_a(0.00014448688307311386)),(to_sfixed_a(0.0030548064969480038)),(to_sfixed_a(-0.0002819244982674718)),(to_sfixed_a(-0.0001805057399906218)),(to_sfixed_a(-0.011539138853549957)),(to_sfixed_a(-0.007148674223572016)),(to_sfixed_a(-2.782951924018562e-06)),(to_sfixed_a(-2.2608677682001144e-05)),(to_sfixed_a(-3.903730248566717e-05)),(to_sfixed_a(-0.00013881885388400406)),(to_sfixed_a(0.0001763203472364694)),(to_sfixed_a(0.00079344492405653)),(to_sfixed_a(-0.09730114042758942)),(to_sfixed_a(7.255740638356656e-05)),(to_sfixed_a(-1.2305477866902947e-05)),(to_sfixed_a(-0.2714453339576721)),(to_sfixed_a(1.3871547707822174e-05)),(to_sfixed_a(-6.824450974818319e-05)),(to_sfixed_a(0.0001073805833584629)),(to_sfixed_a(0.002123042242601514)),(to_sfixed_a(0.00013703486183658242)),(to_sfixed_a(-3.025074693141505e-05)),(to_sfixed_a(5.77803366468288e-05)),(to_sfixed_a(0.2033350169658661)),(to_sfixed_a(3.010145155712962e-05)),(to_sfixed_a(0.0002533535589464009)),(to_sfixed_a(4.6302287955768406e-05)),(to_sfixed_a(1.7868700524559245e-05)),(to_sfixed_a(-0.005878957454115152)),(to_sfixed_a(-0.000286920927464962)),(to_sfixed_a(4.147127037867904e-05)),(to_sfixed_a(0.012032691389322281)),(to_sfixed_a(-0.0001020931958919391)),(to_sfixed_a(-6.9735266151838e-05)),(to_sfixed_a(0.3155288100242615)),(to_sfixed_a(-0.000152201610035263)),(to_sfixed_a(-0.0005739331245422363)),(to_sfixed_a(-7.36199872335419e-05)),(to_sfixed_a(2.4378325178986415e-05)),(to_sfixed_a(-2.3406377295032144e-05)),(to_sfixed_a(0.00017512243357487023)),(to_sfixed_a(-0.0006018095882609487)),(to_sfixed_a(-0.2211112678050995)),(to_sfixed_a(0.005017037969082594)),(to_sfixed_a(0.005609693005681038)),(to_sfixed_a(0.00016848790983203799)),(to_sfixed_a(0.001349292928352952)),(to_sfixed_a(-0.00017877074424177408)),(to_sfixed_a(-0.00013027331442572176)),(to_sfixed_a(0.016126668080687523)),(to_sfixed_a(0.0012126427609473467)),(to_sfixed_a(-0.007310275919735432)),(to_sfixed_a(-5.7593431847635657e-05)),(to_sfixed_a(0.002057868055999279)),(to_sfixed_a(0.0002946395834442228)),(to_sfixed_a(-0.029143113642930984)),(to_sfixed_a(-0.004116331692785025)),(to_sfixed_a(-0.006962247658520937)),(to_sfixed_a(0.003418965497985482)),(to_sfixed_a(-0.0011211868841201067)),(to_sfixed_a(0.01591426506638527)),(to_sfixed_a(-0.00023771786072757095)),(to_sfixed_a(6.560480687767267e-05)),(to_sfixed_a(3.011951775988564e-05)),(to_sfixed_a(-9.005371975945309e-05)),(to_sfixed_a(-0.17287342250347137)),(to_sfixed_a(-0.004091957118362188)),(to_sfixed_a(0.0003981199115514755)),(to_sfixed_a(-0.0015878098784014583)),(to_sfixed_a(-0.0026270970702171326)),(to_sfixed_a(0.0003195015888195485)),(to_sfixed_a(0.010606423951685429)),(to_sfixed_a(0.002454376081004739)),(to_sfixed_a(-6.791928899474442e-05)),(to_sfixed_a(-0.0029165588784962893)),(to_sfixed_a(-2.3193631932372227e-05)),(to_sfixed_a(0.0033361243549734354)),(to_sfixed_a(0.00221537658944726)),(to_sfixed_a(2.737539034569636e-05)),(to_sfixed_a(-0.00017824704991653562)),(to_sfixed_a(-3.849803761113435e-05)),(to_sfixed_a(-1.4346391253639013e-05)),(to_sfixed_a(7.061980431899428e-05)),(to_sfixed_a(8.308392716571689e-05)),(to_sfixed_a(-0.0024091152008622885)),(to_sfixed_a(0.21731555461883545)),(to_sfixed_a(-0.051004357635974884)),(to_sfixed_a(-0.042316485196352005)),(to_sfixed_a(-0.00042833026964217424)),(to_sfixed_a(0.0029950756579637527)),(to_sfixed_a(-0.00022227906447369605)),(to_sfixed_a(3.0322182283271104e-05)),(to_sfixed_a(-3.534831557772122e-05)),(to_sfixed_a(-1.6914214938879013e-05)),(to_sfixed_a(0.00018349218589719385)),(to_sfixed_a(1.6201011021621525e-05)),(to_sfixed_a(-0.0058855777606368065)),(to_sfixed_a(-0.003508979920297861)),(to_sfixed_a(0.00011365889804437757)),(to_sfixed_a(0.00013010436668992043)),(to_sfixed_a(-0.00017702396144159138)),(to_sfixed_a(-0.00015300995437428355)),(to_sfixed_a(0.00046534810098819435)),(to_sfixed_a(0.22597768902778625)),(to_sfixed_a(-0.00013060038327239454)),(to_sfixed_a(0.0001766008062986657)),(to_sfixed_a(5.158327621757053e-05)),(to_sfixed_a(0.0008982904837466776)),(to_sfixed_a(0.0025671268813312054)),(to_sfixed_a(-0.011639382690191269)),(to_sfixed_a(4.81390452478081e-05)),(to_sfixed_a(0.00018035164976026863)),(to_sfixed_a(-0.00016758398851379752)),(to_sfixed_a(0.23102135956287384)),(to_sfixed_a(0.004182429984211922)),(to_sfixed_a(0.017432963475584984)),(to_sfixed_a(-8.040491229621693e-05)),(to_sfixed_a(-6.410702917492017e-05)),(to_sfixed_a(-0.0002990980283357203)),(to_sfixed_a(-0.010163848288357258)),(to_sfixed_a(-8.393692405661568e-05)),(to_sfixed_a(0.41402173042297363)),(to_sfixed_a(-9.189943375531584e-05)),(to_sfixed_a(0.007148700300604105)),(to_sfixed_a(6.659275095444173e-05)),(to_sfixed_a(0.0032668497879058123)),(to_sfixed_a(-0.2686429023742676)),(to_sfixed_a(-0.00016604985285084695)),(to_sfixed_a(0.03124697133898735)),(to_sfixed_a(-0.0008959076949395239)),(to_sfixed_a(-6.695894990116358e-05)),(to_sfixed_a(0.4688752591609955)),(to_sfixed_a(2.4856853997334838e-05)),(to_sfixed_a(0.0003110522811766714)),(to_sfixed_a(0.006833919323980808)),(to_sfixed_a(-0.006320555228739977)),(to_sfixed_a(-0.00010185273276874796)),(to_sfixed_a(-3.845662286039442e-05)),(to_sfixed_a(-0.0015492227394133806)),(to_sfixed_a(-0.00011290617840131745)),(to_sfixed_a(-0.00021109115914441645)),(to_sfixed_a(0.0003138186875730753)),(to_sfixed_a(-0.0011396324262022972)),(to_sfixed_a(0.0002479201357346028)),(to_sfixed_a(-0.20480626821517944)),(to_sfixed_a(0.00024267687695100904)),(to_sfixed_a(3.700883826240897e-05)),(to_sfixed_a(1.7554288206156343e-05)),(to_sfixed_a(-0.0005390046280808747)),(to_sfixed_a(0.004822275601327419)),(to_sfixed_a(3.549011307768524e-05)),(to_sfixed_a(0.00030641938792541623)),(to_sfixed_a(0.00013672461500391364)),(to_sfixed_a(2.907909220084548e-06)),(to_sfixed_a(-0.0009329585009254515)),(to_sfixed_a(0.00032767068478278816)),(to_sfixed_a(-0.003731510369107127)),(to_sfixed_a(0.0020160928834229708)),(to_sfixed_a(-0.0016302444273605943)),(to_sfixed_a(-0.00010865950753213838)),(to_sfixed_a(0.00022009552048984915)),(to_sfixed_a(9.662604861659929e-05)),(to_sfixed_a(-0.003014281624928117)),(to_sfixed_a(0.00022991270816419274)),(to_sfixed_a(-0.00026536535006016493)),(to_sfixed_a(-0.0030604053754359484)),(to_sfixed_a(0.2123805731534958)),(to_sfixed_a(2.5760469725355506e-05)),(to_sfixed_a(0.3521486818790436)),(to_sfixed_a(-0.0001322641910519451)),(to_sfixed_a(-0.0005277726450003684)),(to_sfixed_a(0.001514995819889009)),(to_sfixed_a(-6.564176874235272e-05)),(to_sfixed_a(-0.0014645042829215527)),(to_sfixed_a(-0.001968357479199767)),(to_sfixed_a(0.00935695506632328)),(to_sfixed_a(0.00044492457527667284)),(to_sfixed_a(0.159155011177063)),(to_sfixed_a(-0.0044320388697087765)),(to_sfixed_a(0.010447355918586254)));

    constant weight_n2_75 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.04877933859825134)),(to_sfixed_a(0.17528852820396423)),(to_sfixed_a(0.0056683653965592384)),(to_sfixed_a(-0.00044544722186401486)),(to_sfixed_a(0.0004819793102797121)),(to_sfixed_a(-9.820362174650654e-05)),(to_sfixed_a(-0.0061363899149000645)),(to_sfixed_a(-0.000134584290208295)),(to_sfixed_a(-0.00011336844909237698)),(to_sfixed_a(-3.0113966204226017e-05)),(to_sfixed_a(-0.0001678447297308594)),(to_sfixed_a(-0.00012942112516611814)),(to_sfixed_a(0.006510118022561073)),(to_sfixed_a(0.004400618840008974)),(to_sfixed_a(0.00012127427180530503)),(to_sfixed_a(-0.00011355554306646809)),(to_sfixed_a(-0.003247942076995969)),(to_sfixed_a(0.00015213216829579324)),(to_sfixed_a(0.5759950876235962)),(to_sfixed_a(-0.0008312148274853826)),(to_sfixed_a(0.00015391557826660573)),(to_sfixed_a(-6.298239895841107e-05)),(to_sfixed_a(4.3768864998128265e-05)),(to_sfixed_a(0.0002668921952135861)),(to_sfixed_a(-0.00683684041723609)),(to_sfixed_a(-0.0004707577172666788)),(to_sfixed_a(6.602205394301564e-05)),(to_sfixed_a(0.001062476192601025)),(to_sfixed_a(0.013673897832632065)),(to_sfixed_a(-7.456492312485352e-05)),(to_sfixed_a(-0.011770679615437984)),(to_sfixed_a(-3.0185219657141715e-05)),(to_sfixed_a(0.004162647761404514)),(to_sfixed_a(0.0002021897817030549)),(to_sfixed_a(-0.00016511589637957513)),(to_sfixed_a(-0.00015351468755397946)),(to_sfixed_a(0.39312371611595154)),(to_sfixed_a(-0.3402467966079712)),(to_sfixed_a(-0.010108585469424725)),(to_sfixed_a(-1.6675738152116537e-05)),(to_sfixed_a(-0.0032992935739457607)),(to_sfixed_a(-0.00115670682862401)),(to_sfixed_a(8.99099322850816e-05)),(to_sfixed_a(0.00014719633327331394)),(to_sfixed_a(-0.00036482332507148385)),(to_sfixed_a(0.008770271204411983)),(to_sfixed_a(-0.000772498082369566)),(to_sfixed_a(0.4187409281730652)),(to_sfixed_a(-1.6254040019703098e-05)),(to_sfixed_a(0.0021564506459981203)),(to_sfixed_a(0.0030915173701941967)),(to_sfixed_a(-3.362981078680605e-05)),(to_sfixed_a(-0.00013424210192169994)),(to_sfixed_a(3.094996282015927e-05)),(to_sfixed_a(-0.0037163926754146814)),(to_sfixed_a(-0.009295446798205376)),(to_sfixed_a(-5.943191354162991e-06)),(to_sfixed_a(-0.01210982259362936)),(to_sfixed_a(9.751374454936013e-05)),(to_sfixed_a(-6.526373908855021e-05)),(to_sfixed_a(-6.135491275927052e-05)),(to_sfixed_a(-0.0005048586754128337)),(to_sfixed_a(-0.001405029557645321)),(to_sfixed_a(-0.0006930056260898709)),(to_sfixed_a(9.659372881287709e-05)),(to_sfixed_a(-0.00043735577492043376)),(to_sfixed_a(-0.00011673879635054618)),(to_sfixed_a(0.4101419746875763)),(to_sfixed_a(-0.005104747135192156)),(to_sfixed_a(0.00023842984228394926)),(to_sfixed_a(-0.007570174988359213)),(to_sfixed_a(-0.0029084498528391123)),(to_sfixed_a(0.0013837575679644942)),(to_sfixed_a(3.757626473088749e-05)),(to_sfixed_a(4.5067099563311785e-07)),(to_sfixed_a(-6.422211299650371e-05)),(to_sfixed_a(-0.0059482743963599205)),(to_sfixed_a(-0.0011072867782786489)),(to_sfixed_a(7.103079406078905e-05)),(to_sfixed_a(-0.0012695640325546265)),(to_sfixed_a(0.00014263257617130876)),(to_sfixed_a(0.00011506711598485708)),(to_sfixed_a(-0.0001381165930069983)),(to_sfixed_a(-0.0006265029078349471)),(to_sfixed_a(0.00021939282305538654)),(to_sfixed_a(-0.004387933295220137)),(to_sfixed_a(-0.00045372030581347644)),(to_sfixed_a(0.00021124296472407877)),(to_sfixed_a(-8.740271005081013e-05)),(to_sfixed_a(-0.0003048023208975792)),(to_sfixed_a(-0.013584903441369534)),(to_sfixed_a(-6.646854308201e-05)),(to_sfixed_a(-0.0027021076530218124)),(to_sfixed_a(4.82098403153941e-06)),(to_sfixed_a(0.0009104221826419234)),(to_sfixed_a(2.430094900773838e-05)),(to_sfixed_a(6.800245319027454e-05)),(to_sfixed_a(-7.321588054765016e-05)),(to_sfixed_a(0.00018991754041053355)),(to_sfixed_a(-2.4340184609172866e-05)),(to_sfixed_a(-0.0009733270271681249)),(to_sfixed_a(-0.0007782866014167666)),(to_sfixed_a(2.7172674890607595e-05)),(to_sfixed_a(-0.0028561463113874197)),(to_sfixed_a(-0.2987922430038452)),(to_sfixed_a(0.0007526531699113548)),(to_sfixed_a(-6.989216490183026e-05)),(to_sfixed_a(-1.0617550287861377e-05)),(to_sfixed_a(0.00038149007013998926)),(to_sfixed_a(-0.009264147840440273)),(to_sfixed_a(-0.004959414713084698)),(to_sfixed_a(5.5700005759717897e-05)),(to_sfixed_a(0.01330706849694252)),(to_sfixed_a(0.0001566790451761335)),(to_sfixed_a(-0.00014947204908821732)),(to_sfixed_a(-0.0018505530897527933)),(to_sfixed_a(-2.493192005204037e-05)),(to_sfixed_a(-0.0021119441371411085)),(to_sfixed_a(2.0697189029306173e-07)),(to_sfixed_a(0.013621478341519833)),(to_sfixed_a(-0.00012027121556457132)),(to_sfixed_a(-0.0002986060280818492)),(to_sfixed_a(0.0064197201281785965)),(to_sfixed_a(-0.00014889505109749734)),(to_sfixed_a(-7.46997247915715e-05)),(to_sfixed_a(0.0013934805756434798)),(to_sfixed_a(-0.0007549537112936378)),(to_sfixed_a(-0.00010638145613484085)),(to_sfixed_a(-0.00019648336456157267)),(to_sfixed_a(0.00011433311010478064)),(to_sfixed_a(-0.00010738701530499384)),(to_sfixed_a(-5.651643732562661e-06)),(to_sfixed_a(-0.001413437188602984)),(to_sfixed_a(-0.020408598706126213)),(to_sfixed_a(-0.00024745165137574077)),(to_sfixed_a(3.655689943116158e-05)),(to_sfixed_a(-0.008560610935091972)),(to_sfixed_a(-7.783350883983076e-05)),(to_sfixed_a(-4.4929314753971994e-05)),(to_sfixed_a(3.126038427581079e-05)),(to_sfixed_a(-0.0005166896735318005)),(to_sfixed_a(-5.914062057854608e-05)),(to_sfixed_a(-2.467409649398178e-05)),(to_sfixed_a(0.00018925077165476978)),(to_sfixed_a(0.00011906815780093893)),(to_sfixed_a(0.0007325666956603527)),(to_sfixed_a(3.7483187043108046e-06)),(to_sfixed_a(0.00018111641111318022)),(to_sfixed_a(1.280528522329405e-05)),(to_sfixed_a(-0.00899454951286316)),(to_sfixed_a(0.00023564860748592764)),(to_sfixed_a(0.00021251742145977914)),(to_sfixed_a(-0.001353928237222135)),(to_sfixed_a(0.00015497449203394353)),(to_sfixed_a(0.0002982483129017055)),(to_sfixed_a(-0.06293558329343796)),(to_sfixed_a(-0.00022661122784484178)),(to_sfixed_a(0.0016939020715653896)),(to_sfixed_a(-8.118974801618606e-05)),(to_sfixed_a(-4.404973878990859e-06)),(to_sfixed_a(9.45847132243216e-05)),(to_sfixed_a(8.047489973250777e-05)),(to_sfixed_a(0.001050817547366023)),(to_sfixed_a(-0.00020695161947514862)),(to_sfixed_a(-0.01102590560913086)),(to_sfixed_a(0.0005698291934095323)),(to_sfixed_a(-0.0001273356901947409)),(to_sfixed_a(0.2992860674858093)),(to_sfixed_a(0.0002389983128523454)),(to_sfixed_a(-0.00014694410492666066)),(to_sfixed_a(0.0007946465048007667)),(to_sfixed_a(-0.0036643417552113533)),(to_sfixed_a(-0.001069692661985755)),(to_sfixed_a(-0.0003050119266845286)),(to_sfixed_a(-0.00024202672648243606)),(to_sfixed_a(-0.00034640406374819577)),(to_sfixed_a(-0.0035010192077606916)),(to_sfixed_a(0.0010529417777433991)),(to_sfixed_a(-0.26817354559898376)),(to_sfixed_a(-0.007913138717412949)),(to_sfixed_a(-6.493482942460105e-05)),(to_sfixed_a(-0.010713433846831322)),(to_sfixed_a(-0.00023836438776925206)),(to_sfixed_a(0.0002907873713411391)),(to_sfixed_a(-3.859996286337264e-05)),(to_sfixed_a(-3.6459474358707666e-05)),(to_sfixed_a(0.14960148930549622)),(to_sfixed_a(0.004729305859655142)),(to_sfixed_a(-0.0006962578045204282)),(to_sfixed_a(0.00041316193528473377)),(to_sfixed_a(0.0025930586270987988)),(to_sfixed_a(0.00018236144387628883)),(to_sfixed_a(0.3330114781856537)),(to_sfixed_a(-0.25089508295059204)),(to_sfixed_a(9.823206346482038e-05)),(to_sfixed_a(0.0031557735055685043)),(to_sfixed_a(-0.00010832979751285166)),(to_sfixed_a(-0.0033610539976507425)),(to_sfixed_a(-0.0071898652240633965)),(to_sfixed_a(-2.4562479666201398e-05)),(to_sfixed_a(-0.0002184088370995596)),(to_sfixed_a(-0.00010717411350924522)),(to_sfixed_a(-0.0001621004776097834)),(to_sfixed_a(-4.394122152007185e-05)),(to_sfixed_a(2.913130447268486e-05)),(to_sfixed_a(8.5333755123429e-05)),(to_sfixed_a(-0.0004078741476405412)),(to_sfixed_a(-0.0026025203987956047)),(to_sfixed_a(-0.003555938135832548)),(to_sfixed_a(0.002815056126564741)),(to_sfixed_a(-0.0063909199088811874)),(to_sfixed_a(0.00019935952150262892)),(to_sfixed_a(-0.00022084955708123744)),(to_sfixed_a(-6.713961192872375e-05)),(to_sfixed_a(6.681743252556771e-05)),(to_sfixed_a(7.613627531100065e-05)),(to_sfixed_a(-0.001932517159730196)),(to_sfixed_a(0.001700431341305375)),(to_sfixed_a(0.0034977684263139963)),(to_sfixed_a(-9.558800957165658e-05)),(to_sfixed_a(-1.5143523341976106e-05)),(to_sfixed_a(4.458328476175666e-06)),(to_sfixed_a(-3.614499291870743e-06)),(to_sfixed_a(0.0001362880866508931)),(to_sfixed_a(0.006610007956624031)),(to_sfixed_a(-5.114779924042523e-06)),(to_sfixed_a(-8.484495629090816e-05)),(to_sfixed_a(-6.793231295887381e-05)),(to_sfixed_a(-0.18274585902690887)),(to_sfixed_a(-0.15186993777751923)),(to_sfixed_a(-0.00019657667144201696)),(to_sfixed_a(0.0002864475827664137)),(to_sfixed_a(-0.0002511770580895245)),(to_sfixed_a(-9.875649266177788e-05)),(to_sfixed_a(-0.0058913505636155605)),(to_sfixed_a(0.0037414610851556063)),(to_sfixed_a(0.1363043636083603)),(to_sfixed_a(7.163177360780537e-05)),(to_sfixed_a(0.00011677382281050086)),(to_sfixed_a(-9.920011507347226e-06)),(to_sfixed_a(-0.004309727344661951)),(to_sfixed_a(-0.00031705404398962855)),(to_sfixed_a(-0.4480675458908081)),(to_sfixed_a(0.0001539008371764794)),(to_sfixed_a(0.043899353593587875)),(to_sfixed_a(-0.012116233818233013)),(to_sfixed_a(0.0005356676992960274)),(to_sfixed_a(0.006550587248057127)),(to_sfixed_a(8.791811706032604e-05)),(to_sfixed_a(-0.007737628184258938)),(to_sfixed_a(-0.0014766284730285406)),(to_sfixed_a(-3.545460640452802e-05)),(to_sfixed_a(-0.3336794376373291)),(to_sfixed_a(0.00029124505817890167)),(to_sfixed_a(0.00022389684454537928)),(to_sfixed_a(0.007668999955058098)),(to_sfixed_a(0.0005726362578570843)),(to_sfixed_a(5.610319203697145e-05)),(to_sfixed_a(-3.1780255085323006e-05)),(to_sfixed_a(0.0032556771766394377)),(to_sfixed_a(5.753741424996406e-05)),(to_sfixed_a(-0.0028815653640776873)),(to_sfixed_a(6.507616490125656e-05)),(to_sfixed_a(-4.5806995331076905e-05)),(to_sfixed_a(0.0002295042504556477)),(to_sfixed_a(-0.005561309400945902)),(to_sfixed_a(0.00013255837257020175)),(to_sfixed_a(3.809277404798195e-05)),(to_sfixed_a(1.5653646187274717e-05)),(to_sfixed_a(-0.0008188688079826534)),(to_sfixed_a(0.38507983088493347)),(to_sfixed_a(-0.00030837111989967525)),(to_sfixed_a(0.00013574794866144657)),(to_sfixed_a(0.00010470773850101978)),(to_sfixed_a(-6.056081110727973e-05)),(to_sfixed_a(-0.0038361982442438602)),(to_sfixed_a(0.3228839039802551)),(to_sfixed_a(-0.000923818675801158)),(to_sfixed_a(0.0977601483464241)),(to_sfixed_a(0.0062822806648910046)),(to_sfixed_a(0.00012085140770068392)),(to_sfixed_a(4.68551843368914e-05)),(to_sfixed_a(-6.19676211499609e-05)),(to_sfixed_a(-0.00014523821300826967)),(to_sfixed_a(0.00016737182158976793)),(to_sfixed_a(-9.308638254879043e-05)),(to_sfixed_a(-0.002230798825621605)),(to_sfixed_a(-0.0006071706884540617)),(to_sfixed_a(0.00023975606018211693)),(to_sfixed_a(-0.00025388889480382204)),(to_sfixed_a(-0.0004241003771312535)),(to_sfixed_a(-0.007637070491909981)),(to_sfixed_a(-0.00034274079371243715)),(to_sfixed_a(-2.3628763301530853e-05)),(to_sfixed_a(-0.0005367575795389712)),(to_sfixed_a(0.019822893664240837)),(to_sfixed_a(-0.004084730986505747)),(to_sfixed_a(0.00024005463637877256)),(to_sfixed_a(-0.010298054665327072)),(to_sfixed_a(0.5839604735374451)),(to_sfixed_a(-0.012408211827278137)));

    constant weight_n2_76 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.16452278196811676)),(to_sfixed_a(0.2693217098712921)),(to_sfixed_a(0.2994874119758606)),(to_sfixed_a(-0.00010540487710386515)),(to_sfixed_a(0.3925662338733673)),(to_sfixed_a(1.1587046174099669e-05)),(to_sfixed_a(-0.00032330231624655426)),(to_sfixed_a(6.056507118046284e-06)),(to_sfixed_a(3.586531602195464e-05)),(to_sfixed_a(0.00032535596983507276)),(to_sfixed_a(0.00020166525791864842)),(to_sfixed_a(-0.0010232818312942982)),(to_sfixed_a(-0.1422458440065384)),(to_sfixed_a(0.00042721343925222754)),(to_sfixed_a(-3.131257835775614e-05)),(to_sfixed_a(-1.1417658242862672e-05)),(to_sfixed_a(0.005925765726715326)),(to_sfixed_a(3.02720618492458e-05)),(to_sfixed_a(0.24226388335227966)),(to_sfixed_a(-0.016212131828069687)),(to_sfixed_a(0.00011249048839090392)),(to_sfixed_a(6.939704326214269e-05)),(to_sfixed_a(-1.0544526958256029e-06)),(to_sfixed_a(-0.0001738598948577419)),(to_sfixed_a(0.011724048294126987)),(to_sfixed_a(0.003119697095826268)),(to_sfixed_a(2.4206285161199048e-05)),(to_sfixed_a(-0.00010195554932579398)),(to_sfixed_a(-0.0005044471472501755)),(to_sfixed_a(0.00015639681078027934)),(to_sfixed_a(0.0014353652950376272)),(to_sfixed_a(9.388149919686839e-05)),(to_sfixed_a(-0.010074689984321594)),(to_sfixed_a(6.260597729124129e-05)),(to_sfixed_a(0.00018100868328474462)),(to_sfixed_a(0.00018487172201275826)),(to_sfixed_a(0.023033490404486656)),(to_sfixed_a(-0.2959984540939331)),(to_sfixed_a(0.00128455413505435)),(to_sfixed_a(7.162717520259321e-05)),(to_sfixed_a(0.0028808547649532557)),(to_sfixed_a(0.0007527070702053607)),(to_sfixed_a(0.00011468907177913934)),(to_sfixed_a(-2.5315624952781945e-05)),(to_sfixed_a(4.088778223376721e-05)),(to_sfixed_a(0.004802437033504248)),(to_sfixed_a(0.43406081199645996)),(to_sfixed_a(2.1361738617997617e-05)),(to_sfixed_a(-0.00030675786547362804)),(to_sfixed_a(0.0006804888835176826)),(to_sfixed_a(-0.01669802889227867)),(to_sfixed_a(-0.00029450072906911373)),(to_sfixed_a(-0.00018338172230869532)),(to_sfixed_a(7.622208795510232e-05)),(to_sfixed_a(-0.17430543899536133)),(to_sfixed_a(0.09022104740142822)),(to_sfixed_a(8.264348434749991e-05)),(to_sfixed_a(-0.0005208103684708476)),(to_sfixed_a(-0.00039038664544932544)),(to_sfixed_a(-9.899747237795964e-05)),(to_sfixed_a(0.29047802090644836)),(to_sfixed_a(0.0004841781628783792)),(to_sfixed_a(0.00043183041270822287)),(to_sfixed_a(0.00637977896258235)),(to_sfixed_a(-5.781275103799999e-05)),(to_sfixed_a(0.41508835554122925)),(to_sfixed_a(-0.00013554496399592608)),(to_sfixed_a(0.15996377170085907)),(to_sfixed_a(0.00012102007167413831)),(to_sfixed_a(-7.439089677063748e-05)),(to_sfixed_a(-0.062205515801906586)),(to_sfixed_a(-0.004381400067359209)),(to_sfixed_a(0.01082267239689827)),(to_sfixed_a(0.0001159657840617001)),(to_sfixed_a(0.0004135336494073272)),(to_sfixed_a(-7.06529026501812e-05)),(to_sfixed_a(0.0009618413168936968)),(to_sfixed_a(0.0013015250442549586)),(to_sfixed_a(5.722327477997169e-05)),(to_sfixed_a(0.27069926261901855)),(to_sfixed_a(-0.0005668114172294736)),(to_sfixed_a(0.00025151786394417286)),(to_sfixed_a(0.0002504961739759892)),(to_sfixed_a(0.009639467112720013)),(to_sfixed_a(-7.1927206590771675e-06)),(to_sfixed_a(0.0017130480846390128)),(to_sfixed_a(-0.0039461879059672356)),(to_sfixed_a(-0.00020039633091073483)),(to_sfixed_a(6.489385123131797e-05)),(to_sfixed_a(-6.922610918991268e-05)),(to_sfixed_a(0.0006680248188786209)),(to_sfixed_a(0.00012961370521225035)),(to_sfixed_a(9.595750452717766e-05)),(to_sfixed_a(-1.144791895058006e-05)),(to_sfixed_a(-0.0009653489105403423)),(to_sfixed_a(5.641021562041715e-05)),(to_sfixed_a(5.2457322453847155e-05)),(to_sfixed_a(-0.000167071761097759)),(to_sfixed_a(-9.718570072436705e-05)),(to_sfixed_a(-0.00014238794392440468)),(to_sfixed_a(0.002217354718595743)),(to_sfixed_a(0.000843244546558708)),(to_sfixed_a(-6.2294457165990025e-06)),(to_sfixed_a(-0.00859521608799696)),(to_sfixed_a(0.002591185038909316)),(to_sfixed_a(0.0002890345058403909)),(to_sfixed_a(3.2149648177437484e-05)),(to_sfixed_a(-2.775632674456574e-05)),(to_sfixed_a(-0.00015727760910522193)),(to_sfixed_a(0.003119796747341752)),(to_sfixed_a(-0.21455585956573486)),(to_sfixed_a(-9.502060856902972e-05)),(to_sfixed_a(0.23762905597686768)),(to_sfixed_a(-8.574928506277502e-05)),(to_sfixed_a(3.670859587145969e-05)),(to_sfixed_a(0.0016829394735395908)),(to_sfixed_a(-0.0001025889505399391)),(to_sfixed_a(-3.7469915696419775e-05)),(to_sfixed_a(7.592231850139797e-05)),(to_sfixed_a(0.001831294153816998)),(to_sfixed_a(0.0001826146908570081)),(to_sfixed_a(0.00010360358282923698)),(to_sfixed_a(-0.00012500392040237784)),(to_sfixed_a(0.0001174011267721653)),(to_sfixed_a(-3.998559259343892e-05)),(to_sfixed_a(-0.0036529013887047768)),(to_sfixed_a(-0.0039323060773313046)),(to_sfixed_a(-0.00025132583687081933)),(to_sfixed_a(3.1451156246475875e-05)),(to_sfixed_a(0.00018034991808235645)),(to_sfixed_a(-6.705295527353883e-05)),(to_sfixed_a(-0.00015056796837598085)),(to_sfixed_a(0.0027426783926784992)),(to_sfixed_a(-0.00090707530034706)),(to_sfixed_a(-6.768238381482661e-05)),(to_sfixed_a(4.313260433264077e-06)),(to_sfixed_a(-0.002175078261643648)),(to_sfixed_a(0.0003177294274792075)),(to_sfixed_a(0.00027404187130741775)),(to_sfixed_a(-4.011832061223686e-06)),(to_sfixed_a(2.026725087489467e-05)),(to_sfixed_a(7.608570012962446e-05)),(to_sfixed_a(-1.1336647730786353e-05)),(to_sfixed_a(-0.00018017817637883127)),(to_sfixed_a(0.3282642364501953)),(to_sfixed_a(3.768836904782802e-05)),(to_sfixed_a(0.0003309951280243695)),(to_sfixed_a(0.00011746179370675236)),(to_sfixed_a(-9.306010906584561e-05)),(to_sfixed_a(0.008824440650641918)),(to_sfixed_a(-0.00011227904906263575)),(to_sfixed_a(2.03435993171297e-05)),(to_sfixed_a(-0.3542633056640625)),(to_sfixed_a(1.6399826563429087e-07)),(to_sfixed_a(0.00016818208678159863)),(to_sfixed_a(-0.18792474269866943)),(to_sfixed_a(-2.5967892725020647e-06)),(to_sfixed_a(0.00164792500436306)),(to_sfixed_a(2.0492287148954347e-05)),(to_sfixed_a(0.00012276499182917178)),(to_sfixed_a(-0.00024345410929527134)),(to_sfixed_a(0.00019126717234030366)),(to_sfixed_a(-0.2652536630630493)),(to_sfixed_a(0.0004510215949267149)),(to_sfixed_a(0.00275072711519897)),(to_sfixed_a(0.0015096795978024602)),(to_sfixed_a(0.00010200160613749176)),(to_sfixed_a(-0.0008220359450206161)),(to_sfixed_a(2.2746637114323676e-05)),(to_sfixed_a(4.781881580129266e-05)),(to_sfixed_a(-0.014573754742741585)),(to_sfixed_a(-0.13120931386947632)),(to_sfixed_a(0.00040172331500798464)),(to_sfixed_a(0.00015054222603794187)),(to_sfixed_a(-0.006459745112806559)),(to_sfixed_a(-0.0010759581346064806)),(to_sfixed_a(-0.005147216375917196)),(to_sfixed_a(0.002369967522099614)),(to_sfixed_a(0.08262284100055695)),(to_sfixed_a(-8.588054333813488e-05)),(to_sfixed_a(-0.0003365936572663486)),(to_sfixed_a(-0.013495024293661118)),(to_sfixed_a(0.0001682690781308338)),(to_sfixed_a(0.00013028195826336741)),(to_sfixed_a(-1.1420270311646163e-05)),(to_sfixed_a(0.00015868604532442987)),(to_sfixed_a(0.0026893585454672575)),(to_sfixed_a(-0.0009392115753144026)),(to_sfixed_a(0.0006147082895040512)),(to_sfixed_a(-0.002187056001275778)),(to_sfixed_a(0.0018981362227350473)),(to_sfixed_a(-0.0002194490807596594)),(to_sfixed_a(0.0029140207916498184)),(to_sfixed_a(-0.04707731679081917)),(to_sfixed_a(-2.9322800401132554e-05)),(to_sfixed_a(0.001964119030162692)),(to_sfixed_a(-1.9078135665040463e-05)),(to_sfixed_a(-0.0020740744657814503)),(to_sfixed_a(0.3686978220939636)),(to_sfixed_a(5.627977952826768e-05)),(to_sfixed_a(-4.2264218791387975e-07)),(to_sfixed_a(-0.00010272701911162585)),(to_sfixed_a(0.0001574684720253572)),(to_sfixed_a(0.0001567929284647107)),(to_sfixed_a(6.202104123076424e-05)),(to_sfixed_a(-2.0384813979035243e-05)),(to_sfixed_a(0.23176734149456024)),(to_sfixed_a(-0.0007835209253244102)),(to_sfixed_a(-0.004994560033082962)),(to_sfixed_a(-0.009316974319517612)),(to_sfixed_a(0.22671911120414734)),(to_sfixed_a(5.138383130542934e-05)),(to_sfixed_a(-0.00014801825454924256)),(to_sfixed_a(-8.573315426474437e-05)),(to_sfixed_a(-0.000162718934006989)),(to_sfixed_a(0.00027819297974929214)),(to_sfixed_a(-0.0012388259638100863)),(to_sfixed_a(-0.005690285470336676)),(to_sfixed_a(0.011916178278625011)),(to_sfixed_a(-0.00015613601135555655)),(to_sfixed_a(-0.00028732488863170147)),(to_sfixed_a(-5.544152372749522e-07)),(to_sfixed_a(0.0003070243401452899)),(to_sfixed_a(0.00030235323356464505)),(to_sfixed_a(0.0005577093688771129)),(to_sfixed_a(0.00014747760724276304)),(to_sfixed_a(-3.0728875572094694e-05)),(to_sfixed_a(4.250068741384894e-06)),(to_sfixed_a(0.000160292285727337)),(to_sfixed_a(-0.001290117739699781)),(to_sfixed_a(0.0005893795168958604)),(to_sfixed_a(-7.030636334093288e-05)),(to_sfixed_a(-9.398820111528039e-06)),(to_sfixed_a(0.00023559399414807558)),(to_sfixed_a(-0.0017827715491876006)),(to_sfixed_a(1.8840913980966434e-05)),(to_sfixed_a(-3.307060615043156e-05)),(to_sfixed_a(1.1681382602546364e-05)),(to_sfixed_a(-0.00023421653895638883)),(to_sfixed_a(-0.0003808008914347738)),(to_sfixed_a(-0.015759624540805817)),(to_sfixed_a(0.00020012045570183545)),(to_sfixed_a(0.1835630089044571)),(to_sfixed_a(6.146293162601069e-05)),(to_sfixed_a(0.19449494779109955)),(to_sfixed_a(0.4274410903453827)),(to_sfixed_a(0.000422583834733814)),(to_sfixed_a(0.5139904618263245)),(to_sfixed_a(-0.0001146181020885706)),(to_sfixed_a(-0.002231539925560355)),(to_sfixed_a(-0.00042343573295511305)),(to_sfixed_a(-1.5469631762243807e-05)),(to_sfixed_a(0.0031684560235589743)),(to_sfixed_a(6.686964479740709e-05)),(to_sfixed_a(1.760946906870231e-05)),(to_sfixed_a(0.34436723589897156)),(to_sfixed_a(-0.004140738397836685)),(to_sfixed_a(-3.754037243197672e-05)),(to_sfixed_a(6.946178473299369e-05)),(to_sfixed_a(-0.0007394255371764302)),(to_sfixed_a(0.00017481090617366135)),(to_sfixed_a(0.004155103117227554)),(to_sfixed_a(0.0001725734182400629)),(to_sfixed_a(-0.0003056743589695543)),(to_sfixed_a(0.00012957098078913987)),(to_sfixed_a(0.013474982231855392)),(to_sfixed_a(0.0001052280276780948)),(to_sfixed_a(-0.0001271830260520801)),(to_sfixed_a(-6.802837015129626e-05)),(to_sfixed_a(0.0023601220455020666)),(to_sfixed_a(0.013539686799049377)),(to_sfixed_a(6.89594162395224e-05)),(to_sfixed_a(0.0002723895595408976)),(to_sfixed_a(-1.2906129995826632e-05)),(to_sfixed_a(0.0001056739711202681)),(to_sfixed_a(0.2809591293334961)),(to_sfixed_a(-0.003058261936530471)),(to_sfixed_a(-0.0019664852879941463)),(to_sfixed_a(0.2985535264015198)),(to_sfixed_a(0.0025754068046808243)),(to_sfixed_a(6.0698657762259245e-06)),(to_sfixed_a(-0.0001016145251924172)),(to_sfixed_a(-4.1202743886969984e-05)),(to_sfixed_a(0.0006235413602553308)),(to_sfixed_a(0.00010134237527381629)),(to_sfixed_a(-0.00013782801397610456)),(to_sfixed_a(-0.0016537477495148778)),(to_sfixed_a(0.007469760254025459)),(to_sfixed_a(-4.318177525419742e-05)),(to_sfixed_a(0.19443468749523163)),(to_sfixed_a(-0.00020987897005397826)),(to_sfixed_a(0.0038315998390316963)),(to_sfixed_a(0.0015451553044840693)),(to_sfixed_a(-9.699651855044067e-07)),(to_sfixed_a(0.11231370270252228)),(to_sfixed_a(0.009474352933466434)),(to_sfixed_a(0.004513058811426163)),(to_sfixed_a(7.662994175916538e-05)),(to_sfixed_a(-0.3062015771865845)),(to_sfixed_a(-0.021941756829619408)),(to_sfixed_a(-0.0013336273841559887)));

    constant weight_n2_77 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.08949767798185349)),(to_sfixed_a(-0.004233600106090307)),(to_sfixed_a(0.003629202488809824)),(to_sfixed_a(0.0001550064916955307)),(to_sfixed_a(-0.0030292472802102566)),(to_sfixed_a(0.0002691370318643749)),(to_sfixed_a(-0.00060495879733935)),(to_sfixed_a(0.00016003244672901928)),(to_sfixed_a(4.873341822531074e-06)),(to_sfixed_a(0.00015373851056210697)),(to_sfixed_a(-0.00011570842616492882)),(to_sfixed_a(0.004427335690706968)),(to_sfixed_a(0.36115700006484985)),(to_sfixed_a(-0.5959569215774536)),(to_sfixed_a(2.335533281438984e-05)),(to_sfixed_a(1.3262528227642179e-05)),(to_sfixed_a(-0.43486759066581726)),(to_sfixed_a(-0.0001670012716203928)),(to_sfixed_a(-0.2588183879852295)),(to_sfixed_a(-0.003652665065601468)),(to_sfixed_a(-4.863213689532131e-06)),(to_sfixed_a(-1.0189731256105006e-05)),(to_sfixed_a(0.0001288544590352103)),(to_sfixed_a(0.006350739859044552)),(to_sfixed_a(0.01009416114538908)),(to_sfixed_a(-0.5398269891738892)),(to_sfixed_a(-0.00016802732716314495)),(to_sfixed_a(0.0002601461310405284)),(to_sfixed_a(-0.0017457505455240607)),(to_sfixed_a(7.017963071120903e-05)),(to_sfixed_a(-0.5006734132766724)),(to_sfixed_a(-0.00037987844552844763)),(to_sfixed_a(0.001952196704223752)),(to_sfixed_a(0.00011448063014540821)),(to_sfixed_a(-2.9595779778901488e-05)),(to_sfixed_a(0.00014083289715927094)),(to_sfixed_a(0.4463859498500824)),(to_sfixed_a(0.2171991467475891)),(to_sfixed_a(0.33567124605178833)),(to_sfixed_a(-2.156767004635185e-05)),(to_sfixed_a(-0.002059018239378929)),(to_sfixed_a(-0.16157901287078857)),(to_sfixed_a(-0.00018906423065345734)),(to_sfixed_a(0.00010389919771114364)),(to_sfixed_a(-0.010319779627025127)),(to_sfixed_a(-0.02260163240134716)),(to_sfixed_a(0.001547126448713243)),(to_sfixed_a(-0.0075711351819336414)),(to_sfixed_a(-1.6191064787562937e-05)),(to_sfixed_a(-0.001074566855095327)),(to_sfixed_a(0.012871324084699154)),(to_sfixed_a(0.004366199020296335)),(to_sfixed_a(-4.6350112825166434e-05)),(to_sfixed_a(-0.0007314853719435632)),(to_sfixed_a(-0.009628456085920334)),(to_sfixed_a(-3.2191463105846196e-05)),(to_sfixed_a(1.892432919703424e-06)),(to_sfixed_a(-0.008648591116070747)),(to_sfixed_a(3.736952203325927e-05)),(to_sfixed_a(-0.0002387634594924748)),(to_sfixed_a(-0.030818946659564972)),(to_sfixed_a(-0.0014356400351971388)),(to_sfixed_a(0.007731997407972813)),(to_sfixed_a(0.4015480875968933)),(to_sfixed_a(0.00014917843509465456)),(to_sfixed_a(-0.3107815682888031)),(to_sfixed_a(-6.93512411089614e-05)),(to_sfixed_a(-0.3305145502090454)),(to_sfixed_a(-5.565218816627748e-05)),(to_sfixed_a(0.00030772556783631444)),(to_sfixed_a(0.10755761712789536)),(to_sfixed_a(-0.015368000604212284)),(to_sfixed_a(0.2681286931037903)),(to_sfixed_a(-6.518121517729014e-05)),(to_sfixed_a(-6.900110747665167e-05)),(to_sfixed_a(-7.033672591205686e-05)),(to_sfixed_a(0.017430977895855904)),(to_sfixed_a(0.0021642560604959726)),(to_sfixed_a(-0.00021851985366083682)),(to_sfixed_a(0.2973654270172119)),(to_sfixed_a(-0.009919097647070885)),(to_sfixed_a(0.00027467746986076236)),(to_sfixed_a(0.006861306726932526)),(to_sfixed_a(0.0022425632923841476)),(to_sfixed_a(6.954435957595706e-05)),(to_sfixed_a(0.012642821297049522)),(to_sfixed_a(0.00553413201123476)),(to_sfixed_a(0.004048622213304043)),(to_sfixed_a(3.791331619140692e-05)),(to_sfixed_a(-0.00018973999249283224)),(to_sfixed_a(-0.004512502811849117)),(to_sfixed_a(-5.741013592341915e-05)),(to_sfixed_a(-0.014826709404587746)),(to_sfixed_a(-5.915186193305999e-06)),(to_sfixed_a(-0.0025847468059509993)),(to_sfixed_a(-4.827704469789751e-05)),(to_sfixed_a(0.0003092942060902715)),(to_sfixed_a(-8.311857527587563e-05)),(to_sfixed_a(-0.0001300408912356943)),(to_sfixed_a(0.00011363725934643298)),(to_sfixed_a(0.0046363468281924725)),(to_sfixed_a(-0.0007909539854153991)),(to_sfixed_a(0.00038693295209668577)),(to_sfixed_a(-0.00183375203050673)),(to_sfixed_a(0.12107542157173157)),(to_sfixed_a(-0.0014949331525713205)),(to_sfixed_a(4.386890941532329e-05)),(to_sfixed_a(3.1836207199376076e-05)),(to_sfixed_a(-5.211201641941443e-05)),(to_sfixed_a(0.0012215846218168736)),(to_sfixed_a(-0.24399025738239288)),(to_sfixed_a(0.00015003833686932921)),(to_sfixed_a(-0.001395387458615005)),(to_sfixed_a(-0.00010123633546754718)),(to_sfixed_a(5.868717562407255e-05)),(to_sfixed_a(-0.35456377267837524)),(to_sfixed_a(0.0015329369343817234)),(to_sfixed_a(-0.0013742765877395868)),(to_sfixed_a(-0.00016181661339942366)),(to_sfixed_a(-0.0034272661432623863)),(to_sfixed_a(-0.0001074797473847866)),(to_sfixed_a(0.00015722544048912823)),(to_sfixed_a(-0.0038324855268001556)),(to_sfixed_a(7.419665053021163e-05)),(to_sfixed_a(4.88331716042012e-06)),(to_sfixed_a(-0.06376084685325623)),(to_sfixed_a(-0.012884248048067093)),(to_sfixed_a(-0.00011614375398494303)),(to_sfixed_a(0.00027665821835398674)),(to_sfixed_a(3.5789307730738074e-05)),(to_sfixed_a(3.261632809881121e-05)),(to_sfixed_a(-9.506355854682624e-05)),(to_sfixed_a(-0.42790940403938293)),(to_sfixed_a(-0.009134196676313877)),(to_sfixed_a(6.310297612799332e-05)),(to_sfixed_a(6.111752009019256e-05)),(to_sfixed_a(-0.016654208302497864)),(to_sfixed_a(-0.0010752310045063496)),(to_sfixed_a(-0.00016870969557203352)),(to_sfixed_a(-0.00012964213965460658)),(to_sfixed_a(-0.0021735152695327997)),(to_sfixed_a(-7.125205593183637e-05)),(to_sfixed_a(0.00037593237357214093)),(to_sfixed_a(0.004305116832256317)),(to_sfixed_a(-0.0018268770072609186)),(to_sfixed_a(0.00021490234939847142)),(to_sfixed_a(-0.0005120012210682034)),(to_sfixed_a(7.330853259190917e-05)),(to_sfixed_a(-4.5834840420866385e-05)),(to_sfixed_a(-0.011847035028040409)),(to_sfixed_a(-2.102871803799644e-05)),(to_sfixed_a(-0.00017486052820459008)),(to_sfixed_a(0.2372484803199768)),(to_sfixed_a(1.4936493244022131e-05)),(to_sfixed_a(0.00011373143206583336)),(to_sfixed_a(0.0016411597607657313)),(to_sfixed_a(4.7825400542933494e-05)),(to_sfixed_a(0.0045721218921244144)),(to_sfixed_a(-4.5826447603758425e-05)),(to_sfixed_a(9.012910595629364e-05)),(to_sfixed_a(1.0481693607289344e-05)),(to_sfixed_a(-0.00015424411685671657)),(to_sfixed_a(0.007166841998696327)),(to_sfixed_a(0.00027434490039013326)),(to_sfixed_a(-0.003946125973016024)),(to_sfixed_a(0.006440505851060152)),(to_sfixed_a(1.3908400433138013e-05)),(to_sfixed_a(-0.2236613929271698)),(to_sfixed_a(-0.00014911065227352083)),(to_sfixed_a(6.045605186955072e-05)),(to_sfixed_a(0.004855479579418898)),(to_sfixed_a(-0.003990902099758387)),(to_sfixed_a(0.0012073490070179105)),(to_sfixed_a(7.057515904307365e-05)),(to_sfixed_a(0.03109523467719555)),(to_sfixed_a(0.0025106866378337145)),(to_sfixed_a(0.0013753476087003946)),(to_sfixed_a(-0.0018028297927230597)),(to_sfixed_a(-0.003662529867142439)),(to_sfixed_a(-0.0038223022129386663)),(to_sfixed_a(-0.0015156145673245192)),(to_sfixed_a(-0.0008373691234737635)),(to_sfixed_a(3.815411764662713e-05)),(to_sfixed_a(2.591008524177596e-05)),(to_sfixed_a(0.00011280239414190874)),(to_sfixed_a(0.0015308087458834052)),(to_sfixed_a(-0.004117737524211407)),(to_sfixed_a(-0.19577661156654358)),(to_sfixed_a(0.0010940715437754989)),(to_sfixed_a(-0.17871393263339996)),(to_sfixed_a(0.00528872013092041)),(to_sfixed_a(-0.0001783583138603717)),(to_sfixed_a(-0.002101066056638956)),(to_sfixed_a(0.16375380754470825)),(to_sfixed_a(0.0001484207750763744)),(to_sfixed_a(-0.5165566205978394)),(to_sfixed_a(-0.0003041826712433249)),(to_sfixed_a(-0.006919399369508028)),(to_sfixed_a(0.004577031824737787)),(to_sfixed_a(-1.132007673732005e-05)),(to_sfixed_a(-2.5582339731045067e-05)),(to_sfixed_a(-3.3719989005476236e-06)),(to_sfixed_a(-0.00014033036131877452)),(to_sfixed_a(-4.82905306853354e-06)),(to_sfixed_a(-0.0002424277481622994)),(to_sfixed_a(-0.0005228001391515136)),(to_sfixed_a(0.2932858169078827)),(to_sfixed_a(0.2528587281703949)),(to_sfixed_a(0.0039914632216095924)),(to_sfixed_a(0.00562703562900424)),(to_sfixed_a(0.002983552636578679)),(to_sfixed_a(0.0001715410326141864)),(to_sfixed_a(8.50578144309111e-05)),(to_sfixed_a(0.00018995969730895013)),(to_sfixed_a(-6.885335460538045e-05)),(to_sfixed_a(0.0002263198548462242)),(to_sfixed_a(0.19108472764492035)),(to_sfixed_a(0.014173830859363079)),(to_sfixed_a(0.0017476172652095556)),(to_sfixed_a(0.00018373312195762992)),(to_sfixed_a(0.00016973508172668517)),(to_sfixed_a(0.00015416393580380827)),(to_sfixed_a(1.9875878933817148e-05)),(to_sfixed_a(0.004166295286267996)),(to_sfixed_a(0.48811766505241394)),(to_sfixed_a(6.3344050431624055e-06)),(to_sfixed_a(-7.766587077639997e-05)),(to_sfixed_a(0.00016676259110681713)),(to_sfixed_a(-0.024664631113409996)),(to_sfixed_a(-0.0012157490709796548)),(to_sfixed_a(-0.011506653390824795)),(to_sfixed_a(0.00011713099956978112)),(to_sfixed_a(-0.00021348675363697112)),(to_sfixed_a(-3.873692185152322e-05)),(to_sfixed_a(0.0003112632839474827)),(to_sfixed_a(-0.0043713743798434734)),(to_sfixed_a(0.23765550553798676)),(to_sfixed_a(0.00018283385725226253)),(to_sfixed_a(-0.006596258841454983)),(to_sfixed_a(9.532051626592875e-05)),(to_sfixed_a(-0.6129531860351562)),(to_sfixed_a(0.00015966585488058627)),(to_sfixed_a(-0.018638305366039276)),(to_sfixed_a(-0.00014746030501555651)),(to_sfixed_a(-0.005227430257946253)),(to_sfixed_a(0.024176057428121567)),(to_sfixed_a(-0.43211594223976135)),(to_sfixed_a(0.2502596378326416)),(to_sfixed_a(7.058828487060964e-05)),(to_sfixed_a(-0.00791812315583229)),(to_sfixed_a(0.00039769301656633615)),(to_sfixed_a(-7.459854532498866e-05)),(to_sfixed_a(0.001257686410099268)),(to_sfixed_a(7.214499783003703e-05)),(to_sfixed_a(6.38777855783701e-05)),(to_sfixed_a(-0.0012009604834020138)),(to_sfixed_a(-8.556393731851131e-05)),(to_sfixed_a(0.0001866426318883896)),(to_sfixed_a(-5.650712409988046e-05)),(to_sfixed_a(0.0027095680125057697)),(to_sfixed_a(2.2308486222755164e-06)),(to_sfixed_a(-5.3284387831809e-05)),(to_sfixed_a(-7.079554779920727e-05)),(to_sfixed_a(-0.00011297276068944484)),(to_sfixed_a(6.555450818268582e-05)),(to_sfixed_a(0.014324069023132324)),(to_sfixed_a(0.0001291001244680956)),(to_sfixed_a(1.2046784831909463e-06)),(to_sfixed_a(8.398214413318783e-05)),(to_sfixed_a(-0.004118913784623146)),(to_sfixed_a(0.47989922761917114)),(to_sfixed_a(-0.0003786063753068447)),(to_sfixed_a(5.685573705704883e-05)),(to_sfixed_a(-0.00024132891849149019)),(to_sfixed_a(0.0002428235748084262)),(to_sfixed_a(-0.010995190590620041)),(to_sfixed_a(-0.4021638035774231)),(to_sfixed_a(-0.0017613086383789778)),(to_sfixed_a(-0.27670818567276)),(to_sfixed_a(-0.003055570414289832)),(to_sfixed_a(4.072256706422195e-05)),(to_sfixed_a(0.00022651688777841628)),(to_sfixed_a(-4.123421967960894e-05)),(to_sfixed_a(1.3893088180338964e-05)),(to_sfixed_a(0.00015224215167108923)),(to_sfixed_a(6.177219620440155e-05)),(to_sfixed_a(0.3298158645629883)),(to_sfixed_a(0.2959432005882263)),(to_sfixed_a(-4.8313850129488856e-05)),(to_sfixed_a(0.41563376784324646)),(to_sfixed_a(-0.27943849563598633)),(to_sfixed_a(-0.0059760818257927895)),(to_sfixed_a(-0.08309916406869888)),(to_sfixed_a(0.00010687710891943425)),(to_sfixed_a(0.00858012679964304)),(to_sfixed_a(0.006276977714151144)),(to_sfixed_a(-0.0058876629918813705)),(to_sfixed_a(6.224277603905648e-05)),(to_sfixed_a(-0.00535435089841485)),(to_sfixed_a(-0.008617710322141647)),(to_sfixed_a(-0.007038179785013199)));

    constant weight_n2_78 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.10383819788694382)),(to_sfixed_a(0.009521342813968658)),(to_sfixed_a(2.5331788492621854e-05)),(to_sfixed_a(0.00024111659149639308)),(to_sfixed_a(0.003810441354289651)),(to_sfixed_a(-3.0295152100734413e-05)),(to_sfixed_a(-0.0015393184730783105)),(to_sfixed_a(5.754245648859069e-06)),(to_sfixed_a(7.065772661007941e-05)),(to_sfixed_a(-0.0002439900126773864)),(to_sfixed_a(1.11880581243895e-06)),(to_sfixed_a(0.26770085096359253)),(to_sfixed_a(0.005526898428797722)),(to_sfixed_a(-0.0002381584927206859)),(to_sfixed_a(0.00024331720487680286)),(to_sfixed_a(-0.0001062646770151332)),(to_sfixed_a(-0.0022721595596522093)),(to_sfixed_a(1.3941003999207169e-05)),(to_sfixed_a(-0.01145462691783905)),(to_sfixed_a(-7.312708476092666e-05)),(to_sfixed_a(0.0002687801606953144)),(to_sfixed_a(-0.0002938128018286079)),(to_sfixed_a(0.0015938901342451572)),(to_sfixed_a(-0.0002256229054182768)),(to_sfixed_a(-0.02308550290763378)),(to_sfixed_a(-0.008505289442837238)),(to_sfixed_a(1.2579090252984315e-05)),(to_sfixed_a(-0.0034508181270211935)),(to_sfixed_a(-0.0011559100821614265)),(to_sfixed_a(0.0001694392558420077)),(to_sfixed_a(0.00433321250602603)),(to_sfixed_a(-0.0001759962469805032)),(to_sfixed_a(-0.011856774799525738)),(to_sfixed_a(-5.747332761529833e-05)),(to_sfixed_a(-0.0002750780258793384)),(to_sfixed_a(0.00021866097813472152)),(to_sfixed_a(-0.5641070604324341)),(to_sfixed_a(-0.002973885042592883)),(to_sfixed_a(-0.09904362261295319)),(to_sfixed_a(-6.961825420148671e-06)),(to_sfixed_a(0.01092721801251173)),(to_sfixed_a(0.22777453064918518)),(to_sfixed_a(-1.887016696855426e-05)),(to_sfixed_a(-0.00011100385745521635)),(to_sfixed_a(0.003452196717262268)),(to_sfixed_a(-0.3824683725833893)),(to_sfixed_a(0.009843624196946621)),(to_sfixed_a(0.009373834356665611)),(to_sfixed_a(8.746806997805834e-05)),(to_sfixed_a(0.013576092198491096)),(to_sfixed_a(0.002156279282644391)),(to_sfixed_a(-0.000480568123748526)),(to_sfixed_a(3.373806976014748e-07)),(to_sfixed_a(-0.0003098129527643323)),(to_sfixed_a(0.017077714204788208)),(to_sfixed_a(-0.007212683092802763)),(to_sfixed_a(3.790749178733677e-05)),(to_sfixed_a(0.5391330718994141)),(to_sfixed_a(-3.930521779693663e-05)),(to_sfixed_a(0.00015283437096513808)),(to_sfixed_a(0.0019761500880122185)),(to_sfixed_a(0.0029088128358125687)),(to_sfixed_a(-0.00207078387029469)),(to_sfixed_a(-0.002153246197849512)),(to_sfixed_a(0.00013530913565773517)),(to_sfixed_a(-0.0003094458079431206)),(to_sfixed_a(0.00011468239972600713)),(to_sfixed_a(0.2661505341529846)),(to_sfixed_a(-0.002950174268335104)),(to_sfixed_a(-1.2642223737202585e-05)),(to_sfixed_a(-0.742284893989563)),(to_sfixed_a(0.0007552794995717704)),(to_sfixed_a(-0.5907706618309021)),(to_sfixed_a(0.00014839284995105118)),(to_sfixed_a(-3.912078682333231e-06)),(to_sfixed_a(-0.00011641239689197391)),(to_sfixed_a(-0.000923378684092313)),(to_sfixed_a(0.0035764924250543118)),(to_sfixed_a(-0.000197227782336995)),(to_sfixed_a(-0.007974575273692608)),(to_sfixed_a(0.004818019922822714)),(to_sfixed_a(0.00012137964949943125)),(to_sfixed_a(-0.299744576215744)),(to_sfixed_a(0.005517001263797283)),(to_sfixed_a(-3.86806350434199e-05)),(to_sfixed_a(-0.004607027862221003)),(to_sfixed_a(0.0009207756374962628)),(to_sfixed_a(-0.007536135148257017)),(to_sfixed_a(0.00026442494709044695)),(to_sfixed_a(-7.143936090869829e-05)),(to_sfixed_a(0.006945946253836155)),(to_sfixed_a(0.00013075309107080102)),(to_sfixed_a(0.007294098846614361)),(to_sfixed_a(-0.00029691614327020943)),(to_sfixed_a(-0.0016210397006943822)),(to_sfixed_a(4.314748366596177e-06)),(to_sfixed_a(-3.86940773751121e-05)),(to_sfixed_a(0.00017558937543071806)),(to_sfixed_a(4.0726299630478024e-05)),(to_sfixed_a(0.00018544083286542445)),(to_sfixed_a(0.013744935393333435)),(to_sfixed_a(0.007815353572368622)),(to_sfixed_a(-0.00019951164722442627)),(to_sfixed_a(0.006791250314563513)),(to_sfixed_a(-0.5930505990982056)),(to_sfixed_a(0.1329360157251358)),(to_sfixed_a(-5.748210969613865e-05)),(to_sfixed_a(-8.65620095282793e-05)),(to_sfixed_a(-0.00028740125708281994)),(to_sfixed_a(0.0008853196050040424)),(to_sfixed_a(0.0006873732781969011)),(to_sfixed_a(1.9530438294168562e-05)),(to_sfixed_a(0.003807301400229335)),(to_sfixed_a(6.503261101897806e-05)),(to_sfixed_a(-0.00017275349819101393)),(to_sfixed_a(0.01386429462581873)),(to_sfixed_a(0.0006343546556308866)),(to_sfixed_a(0.006677001249045134)),(to_sfixed_a(-1.2573000276461244e-05)),(to_sfixed_a(0.0029378451872617006)),(to_sfixed_a(-0.00010534618922974914)),(to_sfixed_a(-6.293524347711354e-05)),(to_sfixed_a(0.007361616473644972)),(to_sfixed_a(-5.99009872530587e-05)),(to_sfixed_a(-0.00015065715706441551)),(to_sfixed_a(0.005432289559394121)),(to_sfixed_a(0.004287700168788433)),(to_sfixed_a(-0.0002862905093934387)),(to_sfixed_a(0.0003049145161639899)),(to_sfixed_a(5.765022069681436e-05)),(to_sfixed_a(0.0001666184252826497)),(to_sfixed_a(-0.00018834759248420596)),(to_sfixed_a(0.00043449990334920585)),(to_sfixed_a(0.2769472897052765)),(to_sfixed_a(-0.00011790313146775588)),(to_sfixed_a(2.3896063794381917e-06)),(to_sfixed_a(0.3247548043727875)),(to_sfixed_a(0.6198799014091492)),(to_sfixed_a(8.95458651939407e-05)),(to_sfixed_a(7.97430329839699e-05)),(to_sfixed_a(-0.007724623195827007)),(to_sfixed_a(5.105353920953348e-05)),(to_sfixed_a(-4.240755515638739e-07)),(to_sfixed_a(-0.00022347393678501248)),(to_sfixed_a(-0.00010876852320507169)),(to_sfixed_a(-0.003115789033472538)),(to_sfixed_a(-0.0013629661407321692)),(to_sfixed_a(0.00010641204426065087)),(to_sfixed_a(-0.00011570037895580754)),(to_sfixed_a(0.004168080631643534)),(to_sfixed_a(8.512244676239789e-05)),(to_sfixed_a(0.00010805096826516092)),(to_sfixed_a(-0.0025183381512761116)),(to_sfixed_a(-0.00010696740355342627)),(to_sfixed_a(1.953011451405473e-05)),(to_sfixed_a(-0.008749493397772312)),(to_sfixed_a(-0.00012312672333791852)),(to_sfixed_a(0.005376587156206369)),(to_sfixed_a(2.1118474251125008e-05)),(to_sfixed_a(-4.9955309805227444e-05)),(to_sfixed_a(-4.031922435387969e-05)),(to_sfixed_a(-0.0001064108801074326)),(to_sfixed_a(0.32881492376327515)),(to_sfixed_a(-0.0004925714456476271)),(to_sfixed_a(0.007353235501796007)),(to_sfixed_a(-0.004235394764691591)),(to_sfixed_a(4.06842736992985e-05)),(to_sfixed_a(0.258556604385376)),(to_sfixed_a(1.0421281331218779e-05)),(to_sfixed_a(0.00019023186177946627)),(to_sfixed_a(0.014215877279639244)),(to_sfixed_a(0.0022347047924995422)),(to_sfixed_a(-0.009038995951414108)),(to_sfixed_a(-0.00020527018932625651)),(to_sfixed_a(0.39091920852661133)),(to_sfixed_a(-0.0007452304707840085)),(to_sfixed_a(0.007015276234596968)),(to_sfixed_a(0.2535749673843384)),(to_sfixed_a(-0.4385201930999756)),(to_sfixed_a(-0.45725852251052856)),(to_sfixed_a(0.0003074902342632413)),(to_sfixed_a(-0.0031624173279851675)),(to_sfixed_a(-0.00022093234292697161)),(to_sfixed_a(0.00011195766273885965)),(to_sfixed_a(-2.9753136914223433e-05)),(to_sfixed_a(0.009737841784954071)),(to_sfixed_a(-0.007590349297970533)),(to_sfixed_a(-0.000755906687118113)),(to_sfixed_a(0.00014868745347484946)),(to_sfixed_a(-0.003804450621828437)),(to_sfixed_a(0.0011010951129719615)),(to_sfixed_a(4.231304046697915e-06)),(to_sfixed_a(0.009968200698494911)),(to_sfixed_a(0.000908637244720012)),(to_sfixed_a(0.00010274270607624203)),(to_sfixed_a(0.028007330372929573)),(to_sfixed_a(-3.155348531436175e-05)),(to_sfixed_a(-0.006018056534230709)),(to_sfixed_a(-0.0013532619923353195)),(to_sfixed_a(0.00019955233437940478)),(to_sfixed_a(-0.0003053369000554085)),(to_sfixed_a(-0.0001868267572717741)),(to_sfixed_a(-0.00017799930355977267)),(to_sfixed_a(-2.7470814529806376e-05)),(to_sfixed_a(-0.00024354943889193237)),(to_sfixed_a(-0.0011068300809711218)),(to_sfixed_a(0.007498641032725573)),(to_sfixed_a(0.15784120559692383)),(to_sfixed_a(0.0073079937137663364)),(to_sfixed_a(-0.002274178434163332)),(to_sfixed_a(-0.004080815240740776)),(to_sfixed_a(0.00020031261374242604)),(to_sfixed_a(-2.814449544530362e-07)),(to_sfixed_a(6.484294135589153e-05)),(to_sfixed_a(5.500978295458481e-05)),(to_sfixed_a(-0.0001554276968818158)),(to_sfixed_a(0.0003342010313645005)),(to_sfixed_a(0.08006185293197632)),(to_sfixed_a(2.4255539756268263e-05)),(to_sfixed_a(7.003858627285808e-05)),(to_sfixed_a(-0.00015124741184990853)),(to_sfixed_a(-0.00028657246730290353)),(to_sfixed_a(0.00016650558973196894)),(to_sfixed_a(-0.0029691793024539948)),(to_sfixed_a(-0.4228479862213135)),(to_sfixed_a(-3.6592973629012704e-07)),(to_sfixed_a(2.6159585104323924e-05)),(to_sfixed_a(-0.00010630321776261553)),(to_sfixed_a(0.2954760491847992)),(to_sfixed_a(-0.0017788917757570744)),(to_sfixed_a(-0.24851416051387787)),(to_sfixed_a(-0.0001682547153905034)),(to_sfixed_a(-1.0614021448418498e-06)),(to_sfixed_a(3.268098225817084e-05)),(to_sfixed_a(-0.001153472694568336)),(to_sfixed_a(0.0126345781609416)),(to_sfixed_a(0.192380890250206)),(to_sfixed_a(-3.333248969283886e-05)),(to_sfixed_a(-0.0008272123523056507)),(to_sfixed_a(0.00017640180885791779)),(to_sfixed_a(0.0067781428806483746)),(to_sfixed_a(0.00014898122753947973)),(to_sfixed_a(0.18444930016994476)),(to_sfixed_a(0.000148480583447963)),(to_sfixed_a(0.012739231809973717)),(to_sfixed_a(0.07438571006059647)),(to_sfixed_a(-0.1426268368959427)),(to_sfixed_a(0.0011357309995219111)),(to_sfixed_a(1.8400169210508466e-07)),(to_sfixed_a(0.0037364524323493242)),(to_sfixed_a(0.030229156836867332)),(to_sfixed_a(0.00012686284026131034)),(to_sfixed_a(0.0015954282134771347)),(to_sfixed_a(0.00015421077841892838)),(to_sfixed_a(0.0003710882447194308)),(to_sfixed_a(0.22704480588436127)),(to_sfixed_a(0.189675971865654)),(to_sfixed_a(3.68275614164304e-05)),(to_sfixed_a(4.8002038965933025e-06)),(to_sfixed_a(-0.021868648007512093)),(to_sfixed_a(0.00030820112442597747)),(to_sfixed_a(0.2932886779308319)),(to_sfixed_a(-9.146513184532523e-05)),(to_sfixed_a(-0.00011555009405128658)),(to_sfixed_a(0.000104550774267409)),(to_sfixed_a(0.009094123728573322)),(to_sfixed_a(0.00022500216437038034)),(to_sfixed_a(-3.666751581477001e-05)),(to_sfixed_a(-0.00014278164599090815)),(to_sfixed_a(-0.005965930409729481)),(to_sfixed_a(0.0023091849870979786)),(to_sfixed_a(2.197510184487328e-05)),(to_sfixed_a(1.5443431038875133e-05)),(to_sfixed_a(8.467325096717104e-05)),(to_sfixed_a(-5.071360646979883e-06)),(to_sfixed_a(-0.17101366817951202)),(to_sfixed_a(0.531286895275116)),(to_sfixed_a(0.48560386896133423)),(to_sfixed_a(0.006191836204379797)),(to_sfixed_a(0.002627464709803462)),(to_sfixed_a(-0.00011199861182831228)),(to_sfixed_a(-3.3851174521259964e-06)),(to_sfixed_a(-0.00015040273137856275)),(to_sfixed_a(0.00031186934211291373)),(to_sfixed_a(0.000413787376601249)),(to_sfixed_a(1.1591277143452317e-05)),(to_sfixed_a(0.0002633988915476948)),(to_sfixed_a(-0.3691607713699341)),(to_sfixed_a(-7.292822556337342e-05)),(to_sfixed_a(-0.2859739363193512)),(to_sfixed_a(-0.001488422742113471)),(to_sfixed_a(0.009971392340958118)),(to_sfixed_a(-0.003361096838489175)),(to_sfixed_a(1.3400531315710396e-06)),(to_sfixed_a(-0.0009633441222831607)),(to_sfixed_a(0.26046183705329895)),(to_sfixed_a(0.020526399835944176)),(to_sfixed_a(-5.823623723699711e-05)),(to_sfixed_a(0.1444857120513916)),(to_sfixed_a(-0.08177589625120163)),(to_sfixed_a(0.35250431299209595)));

    constant weight_n2_79 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.060581423342227936)),(to_sfixed_a(0.36663368344306946)),(to_sfixed_a(0.010465269908308983)),(to_sfixed_a(0.0002373760798946023)),(to_sfixed_a(0.002405889332294464)),(to_sfixed_a(-2.57527717621997e-05)),(to_sfixed_a(0.1936541199684143)),(to_sfixed_a(0.00021747378923464566)),(to_sfixed_a(1.157532460638322e-05)),(to_sfixed_a(-8.993006485980004e-05)),(to_sfixed_a(-2.270199911436066e-05)),(to_sfixed_a(-0.020629758015275)),(to_sfixed_a(-0.4591562747955322)),(to_sfixed_a(-0.2529982328414917)),(to_sfixed_a(9.714020416140556e-05)),(to_sfixed_a(0.00017577753169462085)),(to_sfixed_a(0.002934037707746029)),(to_sfixed_a(-0.00015183407231234014)),(to_sfixed_a(-0.010528025217354298)),(to_sfixed_a(5.970410711597651e-05)),(to_sfixed_a(0.00011476607323857024)),(to_sfixed_a(-8.646052447147667e-05)),(to_sfixed_a(-0.0001952608145074919)),(to_sfixed_a(0.3082525134086609)),(to_sfixed_a(0.2780846655368805)),(to_sfixed_a(0.017872238531708717)),(to_sfixed_a(-1.931948645506054e-08)),(to_sfixed_a(0.00034331250935792923)),(to_sfixed_a(-4.136670759180561e-05)),(to_sfixed_a(-2.328784466953948e-05)),(to_sfixed_a(-0.1521167755126953)),(to_sfixed_a(-5.912653432460502e-05)),(to_sfixed_a(-8.532636275049299e-05)),(to_sfixed_a(0.00011500081745907664)),(to_sfixed_a(5.853762559127063e-07)),(to_sfixed_a(-0.00019554329628590494)),(to_sfixed_a(-0.030328840017318726)),(to_sfixed_a(-0.016060316935181618)),(to_sfixed_a(-0.36774417757987976)),(to_sfixed_a(4.778265065397136e-05)),(to_sfixed_a(-0.0028116307221353054)),(to_sfixed_a(0.5179362297058105)),(to_sfixed_a(-2.2860134777147323e-05)),(to_sfixed_a(-0.00018388012540526688)),(to_sfixed_a(0.008783872239291668)),(to_sfixed_a(-0.43941524624824524)),(to_sfixed_a(0.29853707551956177)),(to_sfixed_a(0.0012657159240916371)),(to_sfixed_a(-0.00023072445765137672)),(to_sfixed_a(-0.0013793527614325285)),(to_sfixed_a(0.23665963113307953)),(to_sfixed_a(0.00015098685980774462)),(to_sfixed_a(-0.0001532431342639029)),(to_sfixed_a(0.0003836044343188405)),(to_sfixed_a(-0.00885696429759264)),(to_sfixed_a(6.981308979447931e-05)),(to_sfixed_a(7.124849071260542e-05)),(to_sfixed_a(-0.04082359001040459)),(to_sfixed_a(-0.00019109086133539677)),(to_sfixed_a(0.000382670114049688)),(to_sfixed_a(0.0006710940506309271)),(to_sfixed_a(0.0001668865152169019)),(to_sfixed_a(-0.00033555933623574674)),(to_sfixed_a(0.015197527594864368)),(to_sfixed_a(-6.0552203649422154e-05)),(to_sfixed_a(-0.0016138850478455424)),(to_sfixed_a(6.842192669864744e-05)),(to_sfixed_a(0.009218757040798664)),(to_sfixed_a(0.004130663815885782)),(to_sfixed_a(-0.0004240741254761815)),(to_sfixed_a(0.011203641071915627)),(to_sfixed_a(0.2774222195148468)),(to_sfixed_a(-0.00841300655156374)),(to_sfixed_a(0.00010767533240141347)),(to_sfixed_a(7.129920413717628e-05)),(to_sfixed_a(0.00020734268764499575)),(to_sfixed_a(0.3444375693798065)),(to_sfixed_a(-0.0044170706532895565)),(to_sfixed_a(-0.00010683364962460473)),(to_sfixed_a(0.1787276566028595)),(to_sfixed_a(0.0015724659897387028)),(to_sfixed_a(1.545949635328725e-05)),(to_sfixed_a(0.27519023418426514)),(to_sfixed_a(-0.037666164338588715)),(to_sfixed_a(-0.00012927020725328475)),(to_sfixed_a(0.2646133601665497)),(to_sfixed_a(-0.3045465648174286)),(to_sfixed_a(0.0005512741045095026)),(to_sfixed_a(-0.00029241980519145727)),(to_sfixed_a(-9.266455890610814e-05)),(to_sfixed_a(-0.42906466126441956)),(to_sfixed_a(-0.00011522929708007723)),(to_sfixed_a(-0.008310205303132534)),(to_sfixed_a(1.6815989511087537e-05)),(to_sfixed_a(-0.30901628732681274)),(to_sfixed_a(-9.360752301290631e-05)),(to_sfixed_a(-0.00011592552618822083)),(to_sfixed_a(-2.296437742188573e-06)),(to_sfixed_a(-1.7138991097453982e-06)),(to_sfixed_a(-9.749310265760869e-06)),(to_sfixed_a(0.387357622385025)),(to_sfixed_a(-0.014433103613555431)),(to_sfixed_a(0.0001541844685561955)),(to_sfixed_a(-0.0013743990566581488)),(to_sfixed_a(0.004991100635379553)),(to_sfixed_a(-1.1192421879968606e-05)),(to_sfixed_a(-5.163696187082678e-06)),(to_sfixed_a(1.2949458323419094e-06)),(to_sfixed_a(-2.6661335141398013e-05)),(to_sfixed_a(0.0017885632114484906)),(to_sfixed_a(-0.01750023104250431)),(to_sfixed_a(-7.030655251583084e-05)),(to_sfixed_a(0.010724418796598911)),(to_sfixed_a(-0.0002777990885078907)),(to_sfixed_a(-0.0001551563327666372)),(to_sfixed_a(-0.013563446700572968)),(to_sfixed_a(-0.01390556339174509)),(to_sfixed_a(-0.20300593972206116)),(to_sfixed_a(6.604946975130588e-05)),(to_sfixed_a(0.00027258932823315263)),(to_sfixed_a(1.1449301382526755e-05)),(to_sfixed_a(7.197332161013037e-05)),(to_sfixed_a(0.0002952358918264508)),(to_sfixed_a(-3.8980881072347984e-05)),(to_sfixed_a(-0.00029183554579503834)),(to_sfixed_a(-0.018081434071063995)),(to_sfixed_a(-0.013152186758816242)),(to_sfixed_a(0.00013306527398526669)),(to_sfixed_a(7.650574843864888e-05)),(to_sfixed_a(2.71051685558632e-05)),(to_sfixed_a(6.084957567509264e-05)),(to_sfixed_a(0.00013755033432971686)),(to_sfixed_a(-0.0011176326079294086)),(to_sfixed_a(-0.0037675744388252497)),(to_sfixed_a(-0.0001974902697838843)),(to_sfixed_a(0.00010562299576122314)),(to_sfixed_a(0.0071197315119206905)),(to_sfixed_a(0.001277604722417891)),(to_sfixed_a(7.009844557614997e-05)),(to_sfixed_a(-4.606526272254996e-05)),(to_sfixed_a(-0.07490312308073044)),(to_sfixed_a(3.2708121580071747e-06)),(to_sfixed_a(-0.0001170241812360473)),(to_sfixed_a(-0.00026351812994107604)),(to_sfixed_a(1.5480814909096807e-05)),(to_sfixed_a(-0.0006513114785775542)),(to_sfixed_a(0.0033801484387367964)),(to_sfixed_a(2.634781412780285e-05)),(to_sfixed_a(0.00016823344049043953)),(to_sfixed_a(-0.001197858597151935)),(to_sfixed_a(-0.00013022130588069558)),(to_sfixed_a(0.00023954513017088175)),(to_sfixed_a(-0.005601088982075453)),(to_sfixed_a(0.00010578506044112146)),(to_sfixed_a(0.00014408999413717538)),(to_sfixed_a(-0.14221341907978058)),(to_sfixed_a(0.0002551706857047975)),(to_sfixed_a(0.00038797594606876373)),(to_sfixed_a(5.185114059713669e-05)),(to_sfixed_a(-0.0001275136019103229)),(to_sfixed_a(-0.00021235737949609756)),(to_sfixed_a(0.00019952932780142874)),(to_sfixed_a(0.003913321997970343)),(to_sfixed_a(0.017195776104927063)),(to_sfixed_a(-0.004972459748387337)),(to_sfixed_a(0.0031446816865354776)),(to_sfixed_a(-0.0001861990604083985)),(to_sfixed_a(0.3340640962123871)),(to_sfixed_a(-0.00018106045899912715)),(to_sfixed_a(0.00010670714254956692)),(to_sfixed_a(-0.0034774430096149445)),(to_sfixed_a(0.01808025874197483)),(to_sfixed_a(0.006400062702596188)),(to_sfixed_a(-0.0002487890888005495)),(to_sfixed_a(0.5439876317977905)),(to_sfixed_a(0.011983061209321022)),(to_sfixed_a(-0.007067384198307991)),(to_sfixed_a(-0.00755904009565711)),(to_sfixed_a(0.0012418613769114017)),(to_sfixed_a(0.37268778681755066)),(to_sfixed_a(-0.0005015188944526017)),(to_sfixed_a(0.001364926341921091)),(to_sfixed_a(0.00013068267435301095)),(to_sfixed_a(-6.952141120564193e-07)),(to_sfixed_a(-7.907569670351222e-05)),(to_sfixed_a(0.0031687894370406866)),(to_sfixed_a(-0.26190418004989624)),(to_sfixed_a(-8.824731048662215e-05)),(to_sfixed_a(2.4579401724622585e-05)),(to_sfixed_a(0.001736782374791801)),(to_sfixed_a(-0.001052726642228663)),(to_sfixed_a(-0.0001725491601973772)),(to_sfixed_a(-0.011595731601119041)),(to_sfixed_a(0.18404975533485413)),(to_sfixed_a(-1.1103969882242382e-05)),(to_sfixed_a(-0.00016348378267139196)),(to_sfixed_a(2.963357837870717e-05)),(to_sfixed_a(-0.01007268950343132)),(to_sfixed_a(0.004352563060820103)),(to_sfixed_a(-0.00018235815514344722)),(to_sfixed_a(1.2613192666321993e-05)),(to_sfixed_a(-0.00019107556727249175)),(to_sfixed_a(-7.671586354263127e-05)),(to_sfixed_a(0.0003067964571528137)),(to_sfixed_a(-7.606152212247252e-05)),(to_sfixed_a(0.0012850590283051133)),(to_sfixed_a(0.2365177720785141)),(to_sfixed_a(-0.23655864596366882)),(to_sfixed_a(0.0033645331859588623)),(to_sfixed_a(0.0018219280755147338)),(to_sfixed_a(-0.3303004801273346)),(to_sfixed_a(-0.00029126345179975033)),(to_sfixed_a(-0.0001519956422271207)),(to_sfixed_a(0.0001720304717309773)),(to_sfixed_a(0.00013345539628062397)),(to_sfixed_a(2.4349370505660772e-05)),(to_sfixed_a(-0.023259466513991356)),(to_sfixed_a(-0.5236642360687256)),(to_sfixed_a(-0.004959672689437866)),(to_sfixed_a(-0.00013531309377867728)),(to_sfixed_a(0.00015340697427745908)),(to_sfixed_a(-1.9611390598583966e-05)),(to_sfixed_a(-1.8304490367881954e-05)),(to_sfixed_a(0.01162271574139595)),(to_sfixed_a(0.18740421533584595)),(to_sfixed_a(-0.00016046779637690634)),(to_sfixed_a(0.00010398670565336943)),(to_sfixed_a(-0.00011690935934893787)),(to_sfixed_a(0.0018662638030946255)),(to_sfixed_a(0.0019277505343779922)),(to_sfixed_a(-0.0012040076544508338)),(to_sfixed_a(-2.9089569579809904e-06)),(to_sfixed_a(-0.00041434826562181115)),(to_sfixed_a(6.107444642111659e-05)),(to_sfixed_a(-0.00016908897669054568)),(to_sfixed_a(0.28628814220428467)),(to_sfixed_a(-0.1753871887922287)),(to_sfixed_a(4.642012208933011e-05)),(to_sfixed_a(0.0001708328491076827)),(to_sfixed_a(3.352657950017601e-05)),(to_sfixed_a(0.1744651049375534)),(to_sfixed_a(0.00010639740503393114)),(to_sfixed_a(-0.009096463210880756)),(to_sfixed_a(4.90856655233074e-05)),(to_sfixed_a(-0.039418112486600876)),(to_sfixed_a(-0.21527931094169617)),(to_sfixed_a(0.010372444987297058)),(to_sfixed_a(-0.3416643738746643)),(to_sfixed_a(1.0984509572153911e-05)),(to_sfixed_a(0.20731666684150696)),(to_sfixed_a(-5.500995030160993e-05)),(to_sfixed_a(0.00017862292588688433)),(to_sfixed_a(-0.00017625234613660723)),(to_sfixed_a(-4.655412340071052e-06)),(to_sfixed_a(0.0005551475915126503)),(to_sfixed_a(0.4521493911743164)),(to_sfixed_a(-0.007612064480781555)),(to_sfixed_a(0.0001564616395626217)),(to_sfixed_a(-0.00023586062889080495)),(to_sfixed_a(0.0010160963283851743)),(to_sfixed_a(3.0758455977775156e-06)),(to_sfixed_a(-0.14985904097557068)),(to_sfixed_a(-0.00012848516053054482)),(to_sfixed_a(1.7525890143588185e-06)),(to_sfixed_a(-0.00010886361997108907)),(to_sfixed_a(-0.0074203647673130035)),(to_sfixed_a(-7.4548370321281254e-06)),(to_sfixed_a(9.527472138870507e-05)),(to_sfixed_a(-5.238031008047983e-06)),(to_sfixed_a(-0.24341636896133423)),(to_sfixed_a(0.0733649879693985)),(to_sfixed_a(-7.07876606611535e-05)),(to_sfixed_a(-0.00023889177828095853)),(to_sfixed_a(5.7888944866135716e-05)),(to_sfixed_a(-4.1047693230211735e-05)),(to_sfixed_a(0.4980379641056061)),(to_sfixed_a(0.009964058175683022)),(to_sfixed_a(0.00011869746231241152)),(to_sfixed_a(-0.3204112648963928)),(to_sfixed_a(0.4331158399581909)),(to_sfixed_a(0.00019335380056872964)),(to_sfixed_a(2.4736811610637233e-05)),(to_sfixed_a(-0.00011433100735303015)),(to_sfixed_a(0.0006370117771439254)),(to_sfixed_a(0.00019315133977215737)),(to_sfixed_a(0.000384340004529804)),(to_sfixed_a(0.001310691237449646)),(to_sfixed_a(-0.012814865447580814)),(to_sfixed_a(6.4582891354803e-05)),(to_sfixed_a(0.30904796719551086)),(to_sfixed_a(-0.010879483073949814)),(to_sfixed_a(-0.21004703640937805)),(to_sfixed_a(0.019085019826889038)),(to_sfixed_a(-1.5740690287202597e-05)),(to_sfixed_a(0.0233757421374321)),(to_sfixed_a(-0.008067108690738678)),(to_sfixed_a(-0.29798051714897156)),(to_sfixed_a(0.0001778046425897628)),(to_sfixed_a(0.010735894553363323)),(to_sfixed_a(0.0010624259011819959)),(to_sfixed_a(0.0014378436608240008)));

    constant weight_n2_80 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.459077388048172)),(to_sfixed_a(0.000388826010748744)),(to_sfixed_a(0.005952415056526661)),(to_sfixed_a(0.0002979316341225058)),(to_sfixed_a(0.0009549512760713696)),(to_sfixed_a(0.00016185888671316206)),(to_sfixed_a(-0.001373585662804544)),(to_sfixed_a(-5.8729165175464e-07)),(to_sfixed_a(7.3960545705631375e-06)),(to_sfixed_a(4.3081643525511026e-05)),(to_sfixed_a(-7.415347499772906e-05)),(to_sfixed_a(0.4215445816516876)),(to_sfixed_a(0.010281611233949661)),(to_sfixed_a(0.0039685796946287155)),(to_sfixed_a(-0.0003134212747681886)),(to_sfixed_a(-0.00011303540668450296)),(to_sfixed_a(-0.6882676482200623)),(to_sfixed_a(5.88414040976204e-05)),(to_sfixed_a(0.005578155629336834)),(to_sfixed_a(0.010568269528448582)),(to_sfixed_a(-0.00021391079644672573)),(to_sfixed_a(3.158519393764436e-05)),(to_sfixed_a(-0.0010736525291576982)),(to_sfixed_a(-0.3443252742290497)),(to_sfixed_a(0.0013754275860264897)),(to_sfixed_a(-0.0023839191999286413)),(to_sfixed_a(-0.00022251048358157277)),(to_sfixed_a(0.00023630031500943005)),(to_sfixed_a(-0.006857253611087799)),(to_sfixed_a(-5.7215347624151036e-05)),(to_sfixed_a(-0.3544529974460602)),(to_sfixed_a(6.536433647852391e-05)),(to_sfixed_a(-0.012992747128009796)),(to_sfixed_a(-0.0002462518750689924)),(to_sfixed_a(1.2295640772208571e-06)),(to_sfixed_a(-0.00017502460104878992)),(to_sfixed_a(0.0012613178696483374)),(to_sfixed_a(-0.17733429372310638)),(to_sfixed_a(0.040840886533260345)),(to_sfixed_a(-0.00018043041927739978)),(to_sfixed_a(0.009024766273796558)),(to_sfixed_a(0.007416196167469025)),(to_sfixed_a(-6.086849680286832e-05)),(to_sfixed_a(-7.056332106003538e-05)),(to_sfixed_a(0.00021024169109296054)),(to_sfixed_a(-0.26796892285346985)),(to_sfixed_a(-0.12974253296852112)),(to_sfixed_a(0.0005568512133322656)),(to_sfixed_a(0.00013376340211834759)),(to_sfixed_a(0.00150851730722934)),(to_sfixed_a(-0.003977901767939329)),(to_sfixed_a(2.578287967480719e-05)),(to_sfixed_a(-0.00015720214287284762)),(to_sfixed_a(0.002188229700550437)),(to_sfixed_a(-0.4614546597003937)),(to_sfixed_a(-0.003025833750143647)),(to_sfixed_a(-7.134339830372483e-05)),(to_sfixed_a(0.013853141106665134)),(to_sfixed_a(-0.00015928485663607717)),(to_sfixed_a(-0.000310627743601799)),(to_sfixed_a(-0.0004069832502864301)),(to_sfixed_a(0.0008626761846244335)),(to_sfixed_a(-0.00011372198059689254)),(to_sfixed_a(0.16063176095485687)),(to_sfixed_a(-0.00016858335584402084)),(to_sfixed_a(0.15380805730819702)),(to_sfixed_a(-0.0001368011871818453)),(to_sfixed_a(0.0020165329333394766)),(to_sfixed_a(-0.002868575043976307)),(to_sfixed_a(-2.9423332307487726e-05)),(to_sfixed_a(0.01659664511680603)),(to_sfixed_a(-0.3598019480705261)),(to_sfixed_a(-0.0025160787627100945)),(to_sfixed_a(0.00031126884277909994)),(to_sfixed_a(0.00023705651983618736)),(to_sfixed_a(-4.0727172745391726e-05)),(to_sfixed_a(0.0010538174537941813)),(to_sfixed_a(0.08583920449018478)),(to_sfixed_a(6.270612357184291e-05)),(to_sfixed_a(0.007751213852316141)),(to_sfixed_a(0.0018796056974679232)),(to_sfixed_a(-0.00010198486415902153)),(to_sfixed_a(-0.5621685981750488)),(to_sfixed_a(0.0013831217074766755)),(to_sfixed_a(3.842081787297502e-05)),(to_sfixed_a(0.000901938765309751)),(to_sfixed_a(0.01668984815478325)),(to_sfixed_a(0.0035835783928632736)),(to_sfixed_a(-4.52702515758574e-05)),(to_sfixed_a(-0.00011308798275422305)),(to_sfixed_a(-0.27325376868247986)),(to_sfixed_a(-0.000410490611102432)),(to_sfixed_a(0.005341552663594484)),(to_sfixed_a(7.788763468852267e-05)),(to_sfixed_a(0.004814197774976492)),(to_sfixed_a(-4.639998223865405e-05)),(to_sfixed_a(-0.0001355412823613733)),(to_sfixed_a(0.00013953282905276865)),(to_sfixed_a(1.6371195670217276e-06)),(to_sfixed_a(-1.2714859622064978e-05)),(to_sfixed_a(-0.014516727067530155)),(to_sfixed_a(0.005973931401968002)),(to_sfixed_a(-0.00024086817575152963)),(to_sfixed_a(0.0024930473882704973)),(to_sfixed_a(-0.0010488504776731133)),(to_sfixed_a(0.008371568284928799)),(to_sfixed_a(-2.373848474235274e-05)),(to_sfixed_a(-3.37668061547447e-05)),(to_sfixed_a(-0.0001025526289595291)),(to_sfixed_a(0.0036277000326663256)),(to_sfixed_a(-0.1554589867591858)),(to_sfixed_a(-2.4903794837882742e-05)),(to_sfixed_a(-0.011102559044957161)),(to_sfixed_a(0.00037674076156690717)),(to_sfixed_a(-0.0001372861588606611)),(to_sfixed_a(-0.0016229344764724374)),(to_sfixed_a(0.0011426092823967338)),(to_sfixed_a(0.22309720516204834)),(to_sfixed_a(6.817451503593475e-05)),(to_sfixed_a(-0.00293605774641037)),(to_sfixed_a(-0.00013952868175692856)),(to_sfixed_a(3.4717144444584846e-05)),(to_sfixed_a(-6.124304491095245e-05)),(to_sfixed_a(9.121859329752624e-05)),(to_sfixed_a(-0.0001996695646084845)),(to_sfixed_a(-0.005085028242319822)),(to_sfixed_a(0.07168912887573242)),(to_sfixed_a(1.1623204045463353e-05)),(to_sfixed_a(7.192284101620317e-05)),(to_sfixed_a(-2.9886803531553596e-05)),(to_sfixed_a(-0.00013383988698478788)),(to_sfixed_a(-0.0002981617581099272)),(to_sfixed_a(0.0007063396042212844)),(to_sfixed_a(0.0022241848055273294)),(to_sfixed_a(-0.00015772823826409876)),(to_sfixed_a(0.00018809438915923238)),(to_sfixed_a(0.33586058020591736)),(to_sfixed_a(1.499316749686841e-05)),(to_sfixed_a(0.0001060717404470779)),(to_sfixed_a(0.00020194104581605643)),(to_sfixed_a(0.0002676654257811606)),(to_sfixed_a(1.7731217667460442e-06)),(to_sfixed_a(9.829494956647977e-05)),(to_sfixed_a(-1.9242370399297215e-06)),(to_sfixed_a(-0.00011258562153670937)),(to_sfixed_a(0.00024045226746238768)),(to_sfixed_a(-0.008559064008295536)),(to_sfixed_a(-4.322909808252007e-05)),(to_sfixed_a(0.00026129884645342827)),(to_sfixed_a(0.007700543384999037)),(to_sfixed_a(0.0001273303059861064)),(to_sfixed_a(-5.830588634125888e-06)),(to_sfixed_a(-0.00045920387492515147)),(to_sfixed_a(-0.00011648941290332004)),(to_sfixed_a(-8.09258344816044e-05)),(to_sfixed_a(-0.028042610734701157)),(to_sfixed_a(0.0002982212172355503)),(to_sfixed_a(0.21809041500091553)),(to_sfixed_a(4.152339533902705e-05)),(to_sfixed_a(-4.7455319872824475e-05)),(to_sfixed_a(0.0002658574376255274)),(to_sfixed_a(-4.455967427929863e-05)),(to_sfixed_a(-0.00023725457140244544)),(to_sfixed_a(0.002995405113324523)),(to_sfixed_a(0.011722752824425697)),(to_sfixed_a(0.005439197178930044)),(to_sfixed_a(6.36764889350161e-05)),(to_sfixed_a(-0.004131961148232222)),(to_sfixed_a(6.857152038719505e-05)),(to_sfixed_a(5.660607712343335e-05)),(to_sfixed_a(0.004277522675693035)),(to_sfixed_a(-0.012699284590780735)),(to_sfixed_a(0.0012190802954137325)),(to_sfixed_a(4.5483473513741046e-05)),(to_sfixed_a(0.25167542695999146)),(to_sfixed_a(0.00012008664634777233)),(to_sfixed_a(0.00942497793585062)),(to_sfixed_a(0.0018099453300237656)),(to_sfixed_a(0.00870874710381031)),(to_sfixed_a(-0.503258466720581)),(to_sfixed_a(-8.641537715448067e-05)),(to_sfixed_a(-0.20745545625686646)),(to_sfixed_a(0.0001684415910858661)),(to_sfixed_a(-9.917770512402058e-06)),(to_sfixed_a(-0.00023086313740350306)),(to_sfixed_a(0.005265190731734037)),(to_sfixed_a(-0.0022867454681545496)),(to_sfixed_a(-0.0006819766131229699)),(to_sfixed_a(0.0023468935396522284)),(to_sfixed_a(0.00028707078308798373)),(to_sfixed_a(0.026824750006198883)),(to_sfixed_a(-0.00021517589630093426)),(to_sfixed_a(0.002182048512622714)),(to_sfixed_a(-0.0011054653441533446)),(to_sfixed_a(-0.0002709082909859717)),(to_sfixed_a(-0.4699374735355377)),(to_sfixed_a(-0.00019739892741199583)),(to_sfixed_a(-0.016602899879217148)),(to_sfixed_a(0.3621995449066162)),(to_sfixed_a(-0.00029985111905261874)),(to_sfixed_a(-3.336345616844483e-05)),(to_sfixed_a(0.00018256015027873218)),(to_sfixed_a(0.00010076382022816688)),(to_sfixed_a(-8.954836812335998e-05)),(to_sfixed_a(-0.00016728065384086221)),(to_sfixed_a(-0.0003185143868904561)),(to_sfixed_a(0.0038707812782377005)),(to_sfixed_a(0.37446945905685425)),(to_sfixed_a(-0.03758137673139572)),(to_sfixed_a(0.3613610863685608)),(to_sfixed_a(0.010959537699818611)),(to_sfixed_a(-0.00012819662515539676)),(to_sfixed_a(0.00014489583554677665)),(to_sfixed_a(-0.00016891660925466567)),(to_sfixed_a(-2.262965790578164e-05)),(to_sfixed_a(-8.181077282642946e-05)),(to_sfixed_a(-0.012236948125064373)),(to_sfixed_a(-0.005480518564581871)),(to_sfixed_a(-0.011093324050307274)),(to_sfixed_a(0.00014933929196558893)),(to_sfixed_a(-7.366437057498842e-05)),(to_sfixed_a(-5.225079075898975e-05)),(to_sfixed_a(1.738545688567683e-05)),(to_sfixed_a(0.0005539482808671892)),(to_sfixed_a(-0.018730107694864273)),(to_sfixed_a(-6.268332799663767e-05)),(to_sfixed_a(2.2239259124035016e-05)),(to_sfixed_a(3.4619049984030426e-05)),(to_sfixed_a(0.18588189780712128)),(to_sfixed_a(-0.01655307225883007)),(to_sfixed_a(0.004734036512672901)),(to_sfixed_a(-0.00010233913053525612)),(to_sfixed_a(7.659418042749166e-05)),(to_sfixed_a(0.00010287998884450644)),(to_sfixed_a(-0.004202600568532944)),(to_sfixed_a(-0.013098616153001785)),(to_sfixed_a(-0.2265346795320511)),(to_sfixed_a(-0.00016724009765312076)),(to_sfixed_a(0.00035800636396743357)),(to_sfixed_a(-0.00016127672279253602)),(to_sfixed_a(-0.013407973572611809)),(to_sfixed_a(-3.719730375451036e-05)),(to_sfixed_a(-0.431887149810791)),(to_sfixed_a(0.00018760640523396432)),(to_sfixed_a(0.19835707545280457)),(to_sfixed_a(0.3737967908382416)),(to_sfixed_a(-0.4646987020969391)),(to_sfixed_a(-0.005945142358541489)),(to_sfixed_a(0.00011334996088407934)),(to_sfixed_a(-0.007411746308207512)),(to_sfixed_a(0.017765101045370102)),(to_sfixed_a(3.703608672367409e-05)),(to_sfixed_a(0.007015959359705448)),(to_sfixed_a(-0.00020749411487486213)),(to_sfixed_a(0.0003675520420074463)),(to_sfixed_a(-0.004351034760475159)),(to_sfixed_a(0.005134006962180138)),(to_sfixed_a(-0.00018287589773535728)),(to_sfixed_a(-0.00017057059449143708)),(to_sfixed_a(-0.2431052029132843)),(to_sfixed_a(-0.0001583456469234079)),(to_sfixed_a(0.009858951903879642)),(to_sfixed_a(-7.455578452209011e-05)),(to_sfixed_a(0.0003479327424429357)),(to_sfixed_a(0.00023962119303178042)),(to_sfixed_a(0.20859284698963165)),(to_sfixed_a(-9.547144873067737e-05)),(to_sfixed_a(4.1853636503219604e-06)),(to_sfixed_a(-0.0002991396759171039)),(to_sfixed_a(0.00021778466179966927)),(to_sfixed_a(-0.006285442039370537)),(to_sfixed_a(-5.7078825193457305e-05)),(to_sfixed_a(5.697352025890723e-05)),(to_sfixed_a(0.00023909338051453233)),(to_sfixed_a(-0.0001463352527935058)),(to_sfixed_a(-0.010153360664844513)),(to_sfixed_a(-0.002864337991923094)),(to_sfixed_a(-0.13909687101840973)),(to_sfixed_a(0.0019935572054237127)),(to_sfixed_a(0.002312661614269018)),(to_sfixed_a(-0.00020008793217130005)),(to_sfixed_a(-7.091986481100321e-05)),(to_sfixed_a(-9.172537829726934e-05)),(to_sfixed_a(0.007600985001772642)),(to_sfixed_a(-6.312448385870084e-05)),(to_sfixed_a(3.071455648750998e-05)),(to_sfixed_a(0.007310671266168356)),(to_sfixed_a(0.0027130006346851587)),(to_sfixed_a(-0.00019597257778514177)),(to_sfixed_a(0.00019679567776620388)),(to_sfixed_a(-0.0006794198998250067)),(to_sfixed_a(0.007098437752574682)),(to_sfixed_a(0.32302555441856384)),(to_sfixed_a(-0.00010421633487567306)),(to_sfixed_a(-0.005897918716073036)),(to_sfixed_a(0.417621910572052)),(to_sfixed_a(0.012105755507946014)),(to_sfixed_a(-1.6208279703278095e-05)),(to_sfixed_a(0.004626519978046417)),(to_sfixed_a(0.18812699615955353)),(to_sfixed_a(0.001454163808375597)));

    constant weight_n2_81 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.19730454683303833)),(to_sfixed_a(-0.00030713988235220313)),(to_sfixed_a(-0.0024002757854759693)),(to_sfixed_a(0.00021738522627856582)),(to_sfixed_a(-0.13326925039291382)),(to_sfixed_a(0.00011473096674308181)),(to_sfixed_a(0.00609844783321023)),(to_sfixed_a(0.00016168142610695213)),(to_sfixed_a(-0.00019926762615796179)),(to_sfixed_a(0.0003142467176076025)),(to_sfixed_a(-6.73598115099594e-05)),(to_sfixed_a(0.0032087513245642185)),(to_sfixed_a(0.003141263732686639)),(to_sfixed_a(-0.00010410293907625601)),(to_sfixed_a(-0.00015793480270076543)),(to_sfixed_a(7.001435005804524e-05)),(to_sfixed_a(0.006483545992523432)),(to_sfixed_a(0.00029389167320914567)),(to_sfixed_a(-0.2551444470882416)),(to_sfixed_a(0.006039903964847326)),(to_sfixed_a(-6.354387005558237e-05)),(to_sfixed_a(7.165873103076592e-05)),(to_sfixed_a(0.005572745576500893)),(to_sfixed_a(0.46077847480773926)),(to_sfixed_a(0.012906715273857117)),(to_sfixed_a(0.19459904730319977)),(to_sfixed_a(-1.0423609637655318e-06)),(to_sfixed_a(-0.0012015787651762366)),(to_sfixed_a(-0.005594425834715366)),(to_sfixed_a(6.14546297583729e-06)),(to_sfixed_a(-0.008820770308375359)),(to_sfixed_a(-6.647518603131175e-06)),(to_sfixed_a(0.0001510905276518315)),(to_sfixed_a(-3.4271826734766364e-05)),(to_sfixed_a(-0.00011708040983648971)),(to_sfixed_a(-4.915831232210621e-05)),(to_sfixed_a(-0.5276765823364258)),(to_sfixed_a(0.2682974934577942)),(to_sfixed_a(-0.4176144301891327)),(to_sfixed_a(4.321922460803762e-05)),(to_sfixed_a(0.3422867953777313)),(to_sfixed_a(0.3275999128818512)),(to_sfixed_a(2.913904609158635e-06)),(to_sfixed_a(3.255141564295627e-05)),(to_sfixed_a(0.006474868394434452)),(to_sfixed_a(-0.6476671695709229)),(to_sfixed_a(-0.009319557808339596)),(to_sfixed_a(-0.008512207306921482)),(to_sfixed_a(-0.00011297065793769434)),(to_sfixed_a(0.011704915203154087)),(to_sfixed_a(0.00408614007756114)),(to_sfixed_a(-7.62150957598351e-05)),(to_sfixed_a(6.082050094846636e-05)),(to_sfixed_a(-0.00016946664254646748)),(to_sfixed_a(0.01208256185054779)),(to_sfixed_a(0.014995680190622807)),(to_sfixed_a(-7.141341484384611e-05)),(to_sfixed_a(-0.0035625137388706207)),(to_sfixed_a(-0.00023677220451645553)),(to_sfixed_a(-6.413149822037667e-05)),(to_sfixed_a(-0.005206454079598188)),(to_sfixed_a(-0.0004889664123766124)),(to_sfixed_a(0.003056539222598076)),(to_sfixed_a(-0.00015327722940128297)),(to_sfixed_a(5.878355295863003e-07)),(to_sfixed_a(-0.2939281463623047)),(to_sfixed_a(6.0112310166005045e-05)),(to_sfixed_a(1.6140384104801342e-06)),(to_sfixed_a(0.0300463680177927)),(to_sfixed_a(-0.0004456281312741339)),(to_sfixed_a(-0.18122559785842896)),(to_sfixed_a(-0.0010263274889439344)),(to_sfixed_a(0.006461556069552898)),(to_sfixed_a(-2.3703461920376867e-05)),(to_sfixed_a(-0.00038369448157027364)),(to_sfixed_a(-1.1061547411372885e-06)),(to_sfixed_a(0.23179861903190613)),(to_sfixed_a(0.4041981101036072)),(to_sfixed_a(2.5520952476654202e-05)),(to_sfixed_a(-0.03705504909157753)),(to_sfixed_a(-0.0006518175359815359)),(to_sfixed_a(-0.00020508554007392377)),(to_sfixed_a(0.00013201958790887147)),(to_sfixed_a(-0.2784336507320404)),(to_sfixed_a(-0.00011436177737778053)),(to_sfixed_a(0.21770377457141876)),(to_sfixed_a(-0.47475847601890564)),(to_sfixed_a(0.002839397406205535)),(to_sfixed_a(6.798170215915889e-05)),(to_sfixed_a(0.00012953311670571566)),(to_sfixed_a(-0.008502870798110962)),(to_sfixed_a(-3.924938209820539e-05)),(to_sfixed_a(-0.007593095768243074)),(to_sfixed_a(1.4251680113375187e-05)),(to_sfixed_a(-0.021426595747470856)),(to_sfixed_a(0.00011861525126732886)),(to_sfixed_a(-2.0197687263134867e-05)),(to_sfixed_a(6.2257815443445e-05)),(to_sfixed_a(0.0001912789884954691)),(to_sfixed_a(9.327734005637467e-05)),(to_sfixed_a(0.003412544960156083)),(to_sfixed_a(-0.00893645640462637)),(to_sfixed_a(-3.0352937756106257e-05)),(to_sfixed_a(-0.007458611857146025)),(to_sfixed_a(-0.31518349051475525)),(to_sfixed_a(0.008994854055345058)),(to_sfixed_a(-8.753602742217481e-06)),(to_sfixed_a(4.716347757494077e-05)),(to_sfixed_a(-6.435370596591383e-05)),(to_sfixed_a(0.003705345094203949)),(to_sfixed_a(0.0005768932169303298)),(to_sfixed_a(-0.00016875614528544247)),(to_sfixed_a(-0.6910194158554077)),(to_sfixed_a(-6.842531001893803e-05)),(to_sfixed_a(-0.0002369467547396198)),(to_sfixed_a(0.006049616727977991)),(to_sfixed_a(0.03410942479968071)),(to_sfixed_a(0.002922873944044113)),(to_sfixed_a(0.00025351191288791597)),(to_sfixed_a(0.02558782882988453)),(to_sfixed_a(-2.2714280930813402e-05)),(to_sfixed_a(-2.613465767353773e-06)),(to_sfixed_a(-0.01807466894388199)),(to_sfixed_a(-6.674219912383705e-05)),(to_sfixed_a(4.090492438990623e-06)),(to_sfixed_a(0.005822748877108097)),(to_sfixed_a(0.006230639759451151)),(to_sfixed_a(-1.1236461432417855e-06)),(to_sfixed_a(1.4919925888534635e-05)),(to_sfixed_a(-0.00022704109142068774)),(to_sfixed_a(-4.6324130380526185e-06)),(to_sfixed_a(-6.55973344692029e-05)),(to_sfixed_a(-0.0030296293552964926)),(to_sfixed_a(-0.010582247748970985)),(to_sfixed_a(0.0001066448021447286)),(to_sfixed_a(0.00022139149950817227)),(to_sfixed_a(0.47895094752311707)),(to_sfixed_a(0.23993107676506042)),(to_sfixed_a(0.00016000276082195342)),(to_sfixed_a(1.559848169563338e-05)),(to_sfixed_a(-0.010983589105308056)),(to_sfixed_a(1.9466177036520094e-05)),(to_sfixed_a(-5.460953980218619e-05)),(to_sfixed_a(9.733709885040298e-05)),(to_sfixed_a(-9.612590656615794e-05)),(to_sfixed_a(-0.0033948407508432865)),(to_sfixed_a(-0.002771661849692464)),(to_sfixed_a(-7.114923209883273e-05)),(to_sfixed_a(1.0419505997560918e-05)),(to_sfixed_a(-0.40776872634887695)),(to_sfixed_a(-7.071304571582004e-05)),(to_sfixed_a(-0.00014790697605349123)),(to_sfixed_a(0.17002195119857788)),(to_sfixed_a(-6.133102579042315e-05)),(to_sfixed_a(-0.0002807548444252461)),(to_sfixed_a(-0.011557865887880325)),(to_sfixed_a(-0.0001782740728231147)),(to_sfixed_a(0.0008811140432953835)),(to_sfixed_a(0.0006284712580963969)),(to_sfixed_a(-0.00020341029448900372)),(to_sfixed_a(-0.00010526982077863067)),(to_sfixed_a(-0.00018971173267345876)),(to_sfixed_a(0.21705031394958496)),(to_sfixed_a(0.00018361720140092075)),(to_sfixed_a(0.0007852595299482346)),(to_sfixed_a(0.2250039428472519)),(to_sfixed_a(0.00013000876060687006)),(to_sfixed_a(-0.6398687958717346)),(to_sfixed_a(4.388370143715292e-06)),(to_sfixed_a(0.00023079573293216527)),(to_sfixed_a(0.038895510137081146)),(to_sfixed_a(-0.0020744921639561653)),(to_sfixed_a(0.009044744074344635)),(to_sfixed_a(0.0004235637024976313)),(to_sfixed_a(0.015418299473822117)),(to_sfixed_a(-8.84148757904768e-05)),(to_sfixed_a(0.008021112531423569)),(to_sfixed_a(-0.0010583058465272188)),(to_sfixed_a(0.0029602604918181896)),(to_sfixed_a(0.20531871914863586)),(to_sfixed_a(-0.0025588832795619965)),(to_sfixed_a(-0.35224294662475586)),(to_sfixed_a(3.855963586829603e-05)),(to_sfixed_a(0.0003775653603952378)),(to_sfixed_a(-0.00017528471653349698)),(to_sfixed_a(0.024636641144752502)),(to_sfixed_a(-0.3472824990749359)),(to_sfixed_a(0.0013552383752539754)),(to_sfixed_a(-3.3100259315688163e-06)),(to_sfixed_a(0.0010983417741954327)),(to_sfixed_a(0.0018744160188362002)),(to_sfixed_a(0.00011238655861234292)),(to_sfixed_a(0.0005017053917981684)),(to_sfixed_a(0.265286386013031)),(to_sfixed_a(-3.8764337659813464e-05)),(to_sfixed_a(-0.30561354756355286)),(to_sfixed_a(-0.0003844864259008318)),(to_sfixed_a(-0.006628950126469135)),(to_sfixed_a(0.01228339597582817)),(to_sfixed_a(7.000208279350773e-05)),(to_sfixed_a(6.817205576226115e-05)),(to_sfixed_a(-6.698656943626702e-05)),(to_sfixed_a(0.0001749163493514061)),(to_sfixed_a(-1.1973839718848467e-05)),(to_sfixed_a(8.00727866590023e-06)),(to_sfixed_a(0.0022119979839771986)),(to_sfixed_a(0.0034165414981544018)),(to_sfixed_a(-0.0034354908857494593)),(to_sfixed_a(-0.005751828197389841)),(to_sfixed_a(-0.01040293462574482)),(to_sfixed_a(-0.5030356049537659)),(to_sfixed_a(6.29413771093823e-05)),(to_sfixed_a(-7.307274790946394e-05)),(to_sfixed_a(-0.000286368653178215)),(to_sfixed_a(0.0001714422833174467)),(to_sfixed_a(0.00010809939703904092)),(to_sfixed_a(0.5408619046211243)),(to_sfixed_a(-0.005724653601646423)),(to_sfixed_a(-0.005522406660020351)),(to_sfixed_a(-0.00014103447028901428)),(to_sfixed_a(1.3683093129657209e-05)),(to_sfixed_a(9.802822023630142e-05)),(to_sfixed_a(-4.929846545564942e-05)),(to_sfixed_a(-0.007996250875294209)),(to_sfixed_a(-0.20966501533985138)),(to_sfixed_a(0.00014174227544572204)),(to_sfixed_a(4.758150316774845e-05)),(to_sfixed_a(3.808994733844884e-05)),(to_sfixed_a(0.47140270471572876)),(to_sfixed_a(-0.012747419998049736)),(to_sfixed_a(-0.618021547794342)),(to_sfixed_a(-0.0001846526429289952)),(to_sfixed_a(-4.9877653509611264e-05)),(to_sfixed_a(-0.00021588867821265012)),(to_sfixed_a(0.0010991755407303572)),(to_sfixed_a(0.17503124475479126)),(to_sfixed_a(-0.021517740562558174)),(to_sfixed_a(-5.0830461987061426e-05)),(to_sfixed_a(-0.00233886344358325)),(to_sfixed_a(-6.606431998079643e-05)),(to_sfixed_a(0.03316815197467804)),(to_sfixed_a(0.0003057504363823682)),(to_sfixed_a(-0.01785452291369438)),(to_sfixed_a(-7.447772077284753e-06)),(to_sfixed_a(0.16197356581687927)),(to_sfixed_a(7.198925595730543e-05)),(to_sfixed_a(0.015986710786819458)),(to_sfixed_a(-0.0054267882369458675)),(to_sfixed_a(-8.567014447180554e-05)),(to_sfixed_a(-0.0013966659316793084)),(to_sfixed_a(0.015109967440366745)),(to_sfixed_a(-1.8594437278807163e-05)),(to_sfixed_a(-5.160974251339212e-05)),(to_sfixed_a(-0.00018812248890753835)),(to_sfixed_a(-0.003889220766723156)),(to_sfixed_a(0.6857001781463623)),(to_sfixed_a(0.2615126371383667)),(to_sfixed_a(5.78209146624431e-05)),(to_sfixed_a(5.645507189910859e-05)),(to_sfixed_a(-0.0013285985914990306)),(to_sfixed_a(-2.0890438463538885e-06)),(to_sfixed_a(-0.0005087212193757296)),(to_sfixed_a(7.07663712091744e-05)),(to_sfixed_a(-0.00032205969910137355)),(to_sfixed_a(-2.195847628172487e-06)),(to_sfixed_a(0.04130099341273308)),(to_sfixed_a(-3.274306436651386e-05)),(to_sfixed_a(5.8640602219384164e-05)),(to_sfixed_a(-0.0002039121463894844)),(to_sfixed_a(-0.23134078085422516)),(to_sfixed_a(-0.39565950632095337)),(to_sfixed_a(-0.00016629145829938352)),(to_sfixed_a(1.19389733299613e-05)),(to_sfixed_a(0.0001697861880529672)),(to_sfixed_a(-7.125472620828077e-05)),(to_sfixed_a(0.005021470133215189)),(to_sfixed_a(0.012387082912027836)),(to_sfixed_a(5.918621172895655e-05)),(to_sfixed_a(0.01748082973062992)),(to_sfixed_a(-0.00153604825027287)),(to_sfixed_a(-0.0001567839935887605)),(to_sfixed_a(-4.3730873585445806e-05)),(to_sfixed_a(4.6676308556925505e-05)),(to_sfixed_a(-0.002639053389430046)),(to_sfixed_a(-1.8769926100503653e-05)),(to_sfixed_a(-0.00015483421157114208)),(to_sfixed_a(-0.00028707709861919284)),(to_sfixed_a(-0.004703112877905369)),(to_sfixed_a(6.801003473810852e-05)),(to_sfixed_a(0.34202343225479126)),(to_sfixed_a(-0.008149603381752968)),(to_sfixed_a(0.01653861254453659)),(to_sfixed_a(0.010289931669831276)),(to_sfixed_a(-5.90818453929387e-05)),(to_sfixed_a(0.0026410967111587524)),(to_sfixed_a(-0.018961932510137558)),(to_sfixed_a(0.013800307177007198)),(to_sfixed_a(0.00022875687864143401)),(to_sfixed_a(-0.0027130611706525087)),(to_sfixed_a(-0.15933848917484283)),(to_sfixed_a(0.007914968766272068)));

    constant weight_n2_82 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.36742618680000305)),(to_sfixed_a(0.00011323028593324125)),(to_sfixed_a(0.00013594262418337166)),(to_sfixed_a(-8.644202898722142e-05)),(to_sfixed_a(0.0004001874476671219)),(to_sfixed_a(0.000154264344018884)),(to_sfixed_a(-0.009533138945698738)),(to_sfixed_a(-0.00024795884382911026)),(to_sfixed_a(3.071381070185453e-05)),(to_sfixed_a(0.00010094303434016183)),(to_sfixed_a(0.00026437663473188877)),(to_sfixed_a(-0.002940528793260455)),(to_sfixed_a(-0.005633702501654625)),(to_sfixed_a(0.008386441506445408)),(to_sfixed_a(6.173847214085981e-05)),(to_sfixed_a(-0.00011640239972621202)),(to_sfixed_a(-0.3150479197502136)),(to_sfixed_a(5.2401446737349033e-08)),(to_sfixed_a(0.003859525080770254)),(to_sfixed_a(-0.011413230560719967)),(to_sfixed_a(-1.7518919776193798e-05)),(to_sfixed_a(2.4506716727046296e-05)),(to_sfixed_a(-0.0023816085886210203)),(to_sfixed_a(-3.5905177355743945e-06)),(to_sfixed_a(-0.009071960113942623)),(to_sfixed_a(-0.0029660777654498816)),(to_sfixed_a(0.000172883112099953)),(to_sfixed_a(1.1071208064095117e-05)),(to_sfixed_a(0.006334078963845968)),(to_sfixed_a(-0.0001687726762611419)),(to_sfixed_a(-0.39857473969459534)),(to_sfixed_a(0.0004116878262721002)),(to_sfixed_a(-0.0005931634805165231)),(to_sfixed_a(-2.3556069209007546e-05)),(to_sfixed_a(3.857018600683659e-05)),(to_sfixed_a(-0.00010258001566398889)),(to_sfixed_a(0.18490605056285858)),(to_sfixed_a(0.009601627476513386)),(to_sfixed_a(-0.005498223472386599)),(to_sfixed_a(-4.5247979869600385e-06)),(to_sfixed_a(0.00900090578943491)),(to_sfixed_a(0.0002953497169073671)),(to_sfixed_a(3.598543116822839e-05)),(to_sfixed_a(-0.00020147293980699033)),(to_sfixed_a(-0.0016425253124907613)),(to_sfixed_a(-0.0029020574875175953)),(to_sfixed_a(-0.0011997364927083254)),(to_sfixed_a(0.005886537954211235)),(to_sfixed_a(9.998868335969746e-06)),(to_sfixed_a(0.3819068670272827)),(to_sfixed_a(-0.3018173575401306)),(to_sfixed_a(0.0007839783211238682)),(to_sfixed_a(7.135803753044456e-05)),(to_sfixed_a(0.001004534773528576)),(to_sfixed_a(-0.008228117600083351)),(to_sfixed_a(-0.008534341119229794)),(to_sfixed_a(0.00010809952800627798)),(to_sfixed_a(-0.011216294020414352)),(to_sfixed_a(0.00014246886712498963)),(to_sfixed_a(0.00016717334801796824)),(to_sfixed_a(-0.0036670530680567026)),(to_sfixed_a(-0.0015177989844232798)),(to_sfixed_a(0.0013167986180633307)),(to_sfixed_a(-0.00369746214710176)),(to_sfixed_a(0.000150089428643696)),(to_sfixed_a(0.6012421250343323)),(to_sfixed_a(-2.209267404396087e-05)),(to_sfixed_a(0.3076048493385315)),(to_sfixed_a(-0.009519458748400211)),(to_sfixed_a(8.55882462929003e-05)),(to_sfixed_a(-0.00627824617549777)),(to_sfixed_a(0.018346210941672325)),(to_sfixed_a(-0.02190636470913887)),(to_sfixed_a(-0.00014949837350286543)),(to_sfixed_a(0.00010466380626894534)),(to_sfixed_a(0.00017473756452091038)),(to_sfixed_a(-0.021330473944544792)),(to_sfixed_a(-0.003799924859777093)),(to_sfixed_a(0.00010413307609269395)),(to_sfixed_a(-0.6410173177719116)),(to_sfixed_a(-0.002850254997611046)),(to_sfixed_a(-5.2402083383640274e-05)),(to_sfixed_a(0.0031815655529499054)),(to_sfixed_a(0.00021545737399719656)),(to_sfixed_a(-1.831736881285906e-05)),(to_sfixed_a(0.0007264208979904652)),(to_sfixed_a(-0.0021990370005369186)),(to_sfixed_a(-6.735981878591701e-05)),(to_sfixed_a(0.00021790106256958097)),(to_sfixed_a(7.170946628320962e-05)),(to_sfixed_a(-0.0037841342855244875)),(to_sfixed_a(8.509978943038732e-05)),(to_sfixed_a(-0.008631259202957153)),(to_sfixed_a(7.014404400251806e-05)),(to_sfixed_a(-0.0054907421581447124)),(to_sfixed_a(3.1474210118176416e-05)),(to_sfixed_a(0.00010548772115726024)),(to_sfixed_a(-8.317107131006196e-05)),(to_sfixed_a(0.00011452993931015953)),(to_sfixed_a(0.00030647453968413174)),(to_sfixed_a(-0.00660719396546483)),(to_sfixed_a(0.00010353281686548144)),(to_sfixed_a(0.00029516126960515976)),(to_sfixed_a(-0.007210797164589167)),(to_sfixed_a(-0.007707959972321987)),(to_sfixed_a(4.8154684918699786e-05)),(to_sfixed_a(-8.449002780253068e-05)),(to_sfixed_a(-7.867746899137273e-05)),(to_sfixed_a(0.00012820113624911755)),(to_sfixed_a(-0.0046707200817763805)),(to_sfixed_a(0.1597663164138794)),(to_sfixed_a(0.00015652422735001892)),(to_sfixed_a(-0.0003394211526028812)),(to_sfixed_a(-0.00014015765918884426)),(to_sfixed_a(-0.00016551592852920294)),(to_sfixed_a(0.0036684200167655945)),(to_sfixed_a(-0.0006030616932548583)),(to_sfixed_a(-0.002904218854382634)),(to_sfixed_a(0.00016684315050952137)),(to_sfixed_a(-0.23608922958374023)),(to_sfixed_a(7.719627319602296e-05)),(to_sfixed_a(-9.788999886950478e-05)),(to_sfixed_a(-0.0005183628527447581)),(to_sfixed_a(-0.00024716914049349725)),(to_sfixed_a(0.0001302170567214489)),(to_sfixed_a(-0.00028884579660370946)),(to_sfixed_a(-0.008519412949681282)),(to_sfixed_a(-3.875956463161856e-05)),(to_sfixed_a(-1.2298303772695363e-05)),(to_sfixed_a(1.7664206097833812e-07)),(to_sfixed_a(7.095558248693123e-05)),(to_sfixed_a(-5.7244280469603837e-05)),(to_sfixed_a(0.0007443332578986883)),(to_sfixed_a(0.19570143520832062)),(to_sfixed_a(0.00016809298540465534)),(to_sfixed_a(3.084231138927862e-06)),(to_sfixed_a(-0.011393526569008827)),(to_sfixed_a(0.0002273433783557266)),(to_sfixed_a(2.038273487414699e-05)),(to_sfixed_a(6.787992606405169e-05)),(to_sfixed_a(0.10311418026685715)),(to_sfixed_a(-0.00010935959289781749)),(to_sfixed_a(0.00015522174362558872)),(to_sfixed_a(-4.804122363566421e-05)),(to_sfixed_a(-0.00016368973592761904)),(to_sfixed_a(0.00012276749475859106)),(to_sfixed_a(-0.0003022169694304466)),(to_sfixed_a(6.723732076352462e-05)),(to_sfixed_a(-6.654100434388965e-05)),(to_sfixed_a(-0.011725255288183689)),(to_sfixed_a(-2.978478732984513e-06)),(to_sfixed_a(-2.4556655262131244e-05)),(to_sfixed_a(-0.004507946316152811)),(to_sfixed_a(3.0619383323937654e-05)),(to_sfixed_a(0.00010364246554672718)),(to_sfixed_a(-0.20218540728092194)),(to_sfixed_a(0.00018733894103206694)),(to_sfixed_a(0.004326599184423685)),(to_sfixed_a(5.382819290389307e-05)),(to_sfixed_a(-0.000137026741867885)),(to_sfixed_a(0.00010683832078939304)),(to_sfixed_a(-0.00015233681187964976)),(to_sfixed_a(0.003068332327529788)),(to_sfixed_a(3.9590544474776834e-05)),(to_sfixed_a(-0.0037899294402450323)),(to_sfixed_a(-0.1918952763080597)),(to_sfixed_a(0.00038909309660084546)),(to_sfixed_a(-0.0027769843582063913)),(to_sfixed_a(-0.00010058128100354224)),(to_sfixed_a(2.6630070351529866e-05)),(to_sfixed_a(-0.16682633757591248)),(to_sfixed_a(-0.005437915213406086)),(to_sfixed_a(-0.003687492338940501)),(to_sfixed_a(7.959100184962153e-05)),(to_sfixed_a(0.002955728443339467)),(to_sfixed_a(-0.0015647426480427384)),(to_sfixed_a(-0.0023984836880117655)),(to_sfixed_a(0.000577675411477685)),(to_sfixed_a(-0.28197887539863586)),(to_sfixed_a(-0.6169329881668091)),(to_sfixed_a(0.001077391323633492)),(to_sfixed_a(0.009625455364584923)),(to_sfixed_a(7.787093636579812e-05)),(to_sfixed_a(1.8307291611563414e-05)),(to_sfixed_a(0.00015697335766162723)),(to_sfixed_a(-0.00011362937220837921)),(to_sfixed_a(-0.3640438914299011)),(to_sfixed_a(0.0004121753154322505)),(to_sfixed_a(0.0010012804996222258)),(to_sfixed_a(0.003896260168403387)),(to_sfixed_a(0.0015495273983106017)),(to_sfixed_a(0.00018680380890145898)),(to_sfixed_a(-0.30592241883277893)),(to_sfixed_a(-0.003940684720873833)),(to_sfixed_a(-0.0001562755205668509)),(to_sfixed_a(-0.38034096360206604)),(to_sfixed_a(8.100811101030558e-06)),(to_sfixed_a(-0.008702604100108147)),(to_sfixed_a(0.028648948296904564)),(to_sfixed_a(1.5247678675223142e-06)),(to_sfixed_a(-0.00027319390210323036)),(to_sfixed_a(-8.352551230927929e-05)),(to_sfixed_a(0.0002419886877760291)),(to_sfixed_a(2.339487400604412e-05)),(to_sfixed_a(2.6063280529342592e-05)),(to_sfixed_a(0.2809523940086365)),(to_sfixed_a(0.010275375097990036)),(to_sfixed_a(0.3044365346431732)),(to_sfixed_a(-0.000968850392382592)),(to_sfixed_a(0.2578470706939697)),(to_sfixed_a(-0.011744583025574684)),(to_sfixed_a(3.6370838643051684e-06)),(to_sfixed_a(-5.711299309041351e-07)),(to_sfixed_a(-9.673953172750771e-06)),(to_sfixed_a(6.466947525041178e-05)),(to_sfixed_a(0.0002001666434807703)),(to_sfixed_a(0.010767754167318344)),(to_sfixed_a(-0.00011802333756349981)),(to_sfixed_a(-0.0023784751538187265)),(to_sfixed_a(0.0001302054151892662)),(to_sfixed_a(0.00022245194122660905)),(to_sfixed_a(7.658989488845691e-05)),(to_sfixed_a(0.0002534622617531568)),(to_sfixed_a(6.672507879557088e-05)),(to_sfixed_a(0.000625012326054275)),(to_sfixed_a(0.00014920937246643007)),(to_sfixed_a(-0.00012939819134771824)),(to_sfixed_a(1.6389094525948167e-07)),(to_sfixed_a(0.0018524155020713806)),(to_sfixed_a(0.17430563271045685)),(to_sfixed_a(-0.0028138591442257166)),(to_sfixed_a(-1.1764066584873945e-05)),(to_sfixed_a(8.60091095091775e-05)),(to_sfixed_a(-3.209754140698351e-05)),(to_sfixed_a(-0.007841216400265694)),(to_sfixed_a(-0.006199117284268141)),(to_sfixed_a(0.4699595272541046)),(to_sfixed_a(1.2357377272564918e-06)),(to_sfixed_a(0.0021493996027857065)),(to_sfixed_a(0.0004462827346287668)),(to_sfixed_a(0.00021453169756568968)),(to_sfixed_a(-0.00046022055903449655)),(to_sfixed_a(-0.002754343207925558)),(to_sfixed_a(-3.6455312510952353e-05)),(to_sfixed_a(-0.08840817213058472)),(to_sfixed_a(-0.00168905989266932)),(to_sfixed_a(-0.2219811975955963)),(to_sfixed_a(0.5842064023017883)),(to_sfixed_a(-2.3945751308929175e-05)),(to_sfixed_a(-0.011457770131528378)),(to_sfixed_a(0.00018059927970170975)),(to_sfixed_a(-0.00013349879009183496)),(to_sfixed_a(0.001608927152119577)),(to_sfixed_a(-6.264685362111777e-05)),(to_sfixed_a(3.2300857128575444e-05)),(to_sfixed_a(0.0003386142780072987)),(to_sfixed_a(-0.0045958287082612514)),(to_sfixed_a(0.00023003818932920694)),(to_sfixed_a(0.00023743975907564163)),(to_sfixed_a(0.017649739980697632)),(to_sfixed_a(-2.4120850866893306e-05)),(to_sfixed_a(0.00024311717425007373)),(to_sfixed_a(3.8886635593371466e-05)),(to_sfixed_a(0.0003920658491551876)),(to_sfixed_a(0.00031938249594531953)),(to_sfixed_a(-0.01279985997825861)),(to_sfixed_a(1.9533399608917534e-05)),(to_sfixed_a(-5.379635695135221e-05)),(to_sfixed_a(-0.00018070259829983115)),(to_sfixed_a(-5.1301525672897696e-05)),(to_sfixed_a(0.22038500010967255)),(to_sfixed_a(-0.00020149863848928362)),(to_sfixed_a(0.0001281409931834787)),(to_sfixed_a(-2.919701364589855e-05)),(to_sfixed_a(2.1111578462296166e-05)),(to_sfixed_a(-0.008023764938116074)),(to_sfixed_a(-0.0001353735278826207)),(to_sfixed_a(-0.0020156074315309525)),(to_sfixed_a(-0.004948012065142393)),(to_sfixed_a(0.0009615081362426281)),(to_sfixed_a(-6.448541535064578e-05)),(to_sfixed_a(-1.8939404981210828e-05)),(to_sfixed_a(-0.00013918844342697412)),(to_sfixed_a(4.161664401181042e-05)),(to_sfixed_a(6.332444172585383e-05)),(to_sfixed_a(1.0570169251877815e-05)),(to_sfixed_a(0.0002519277622923255)),(to_sfixed_a(-0.22437074780464172)),(to_sfixed_a(3.68157125194557e-05)),(to_sfixed_a(-9.576747106621042e-05)),(to_sfixed_a(0.00030559106380678713)),(to_sfixed_a(0.3020760118961334)),(to_sfixed_a(0.15940755605697632)),(to_sfixed_a(1.851632259786129e-05)),(to_sfixed_a(0.006668898276984692)),(to_sfixed_a(0.002608007052913308)),(to_sfixed_a(-0.0013639659155160189)),(to_sfixed_a(0.00020477747602853924)),(to_sfixed_a(-0.009304987266659737)),(to_sfixed_a(-0.0035137904342263937)),(to_sfixed_a(-0.0138560114428401)));

    constant weight_n2_83 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.059866201132535934)),(to_sfixed_a(-0.00011233624536544085)),(to_sfixed_a(0.00018764007836580276)),(to_sfixed_a(0.00018779862148221582)),(to_sfixed_a(0.00018058318528346717)),(to_sfixed_a(-1.85796307050623e-06)),(to_sfixed_a(7.293615635717288e-05)),(to_sfixed_a(-0.0002451443288009614)),(to_sfixed_a(-0.00028321449644863605)),(to_sfixed_a(-0.00013626430882140994)),(to_sfixed_a(6.966409273445606e-05)),(to_sfixed_a(-7.014871516730636e-05)),(to_sfixed_a(0.0002667965891305357)),(to_sfixed_a(0.00010259730333928019)),(to_sfixed_a(-4.438572796061635e-05)),(to_sfixed_a(-4.543241811916232e-05)),(to_sfixed_a(3.8989848690107465e-05)),(to_sfixed_a(0.0001815012947190553)),(to_sfixed_a(-0.00011428205471020192)),(to_sfixed_a(7.841166370781139e-05)),(to_sfixed_a(-3.324489443912171e-05)),(to_sfixed_a(4.552252357825637e-05)),(to_sfixed_a(1.4701341569889337e-05)),(to_sfixed_a(-0.0002914436627179384)),(to_sfixed_a(-0.00024032533110585064)),(to_sfixed_a(0.00031608602148480713)),(to_sfixed_a(0.00024315033806487918)),(to_sfixed_a(-7.282272417796776e-05)),(to_sfixed_a(7.671705679968e-05)),(to_sfixed_a(-6.984776700846851e-05)),(to_sfixed_a(0.00024027161998674273)),(to_sfixed_a(-4.5185661292634904e-06)),(to_sfixed_a(0.00015524223272223026)),(to_sfixed_a(-2.4719047360122204e-05)),(to_sfixed_a(3.0138948204694316e-05)),(to_sfixed_a(0.00017401244258508086)),(to_sfixed_a(-1.8869082850869745e-05)),(to_sfixed_a(2.4246630346169695e-05)),(to_sfixed_a(9.761910769157112e-05)),(to_sfixed_a(-9.875990144792013e-06)),(to_sfixed_a(3.0110240913927555e-05)),(to_sfixed_a(0.00020037617650814354)),(to_sfixed_a(0.00015109135711099952)),(to_sfixed_a(4.3193100282223895e-05)),(to_sfixed_a(-0.00011788152187364176)),(to_sfixed_a(3.1094888981897384e-05)),(to_sfixed_a(-1.0815307177836075e-05)),(to_sfixed_a(-5.8339232055004686e-05)),(to_sfixed_a(0.00015847808390390128)),(to_sfixed_a(-0.0001466987596359104)),(to_sfixed_a(0.00012896512635052204)),(to_sfixed_a(-0.00012326615978963673)),(to_sfixed_a(4.999594239052385e-06)),(to_sfixed_a(-0.0001030758794513531)),(to_sfixed_a(-1.8162587366532534e-05)),(to_sfixed_a(-0.00023987775784917176)),(to_sfixed_a(-6.667283014394343e-05)),(to_sfixed_a(8.597358828410506e-05)),(to_sfixed_a(6.019307329552248e-05)),(to_sfixed_a(-0.00010517360351514071)),(to_sfixed_a(0.0001648096222197637)),(to_sfixed_a(0.0001357549917884171)),(to_sfixed_a(6.741298420820385e-05)),(to_sfixed_a(-9.012751979753375e-05)),(to_sfixed_a(2.08600249607116e-06)),(to_sfixed_a(2.9792801797157153e-05)),(to_sfixed_a(0.00010725504398578778)),(to_sfixed_a(-0.00017430567822884768)),(to_sfixed_a(2.4136312276823446e-05)),(to_sfixed_a(0.0002643494517542422)),(to_sfixed_a(5.6466808018740267e-05)),(to_sfixed_a(3.259629011154175e-09)),(to_sfixed_a(0.00023876060731709003)),(to_sfixed_a(0.00017281487816944718)),(to_sfixed_a(7.042459037620574e-05)),(to_sfixed_a(0.00011259419261477888)),(to_sfixed_a(9.948800652637146e-06)),(to_sfixed_a(0.00010795627167681232)),(to_sfixed_a(-3.088466473855078e-05)),(to_sfixed_a(-0.00023565496667288244)),(to_sfixed_a(-0.00011689573875628412)),(to_sfixed_a(-6.821143324486911e-05)),(to_sfixed_a(-0.000204829266294837)),(to_sfixed_a(-1.3508033589459956e-06)),(to_sfixed_a(-1.903050724649802e-05)),(to_sfixed_a(0.00011350827844580635)),(to_sfixed_a(-1.2454926036298275e-05)),(to_sfixed_a(6.844656309112906e-05)),(to_sfixed_a(0.00020444214169401675)),(to_sfixed_a(5.6864446378313005e-05)),(to_sfixed_a(-7.79697293182835e-05)),(to_sfixed_a(0.00022202415857464075)),(to_sfixed_a(-0.00010157405631616712)),(to_sfixed_a(0.00010651886987034231)),(to_sfixed_a(0.00016740764840506017)),(to_sfixed_a(-1.2194424925837666e-05)),(to_sfixed_a(-7.028922846075147e-05)),(to_sfixed_a(-3.704657137859613e-05)),(to_sfixed_a(0.00015502612222917378)),(to_sfixed_a(7.106548582669348e-05)),(to_sfixed_a(-0.00011563846055651084)),(to_sfixed_a(-0.00011313751747366041)),(to_sfixed_a(-0.0002361278748139739)),(to_sfixed_a(7.870529225328937e-05)),(to_sfixed_a(2.7652211429085582e-05)),(to_sfixed_a(-2.6241792511427775e-05)),(to_sfixed_a(4.4165150029584765e-05)),(to_sfixed_a(-0.0001559277152409777)),(to_sfixed_a(-1.1272219126112759e-05)),(to_sfixed_a(0.00015165164950303733)),(to_sfixed_a(9.403738658875227e-07)),(to_sfixed_a(0.00013406641664914787)),(to_sfixed_a(4.279873246559873e-05)),(to_sfixed_a(-0.0001532937603769824)),(to_sfixed_a(-1.5106488717719913e-06)),(to_sfixed_a(0.00018479529535397887)),(to_sfixed_a(-2.9680508305318654e-05)),(to_sfixed_a(-5.9882833738811314e-05)),(to_sfixed_a(3.829365596175194e-05)),(to_sfixed_a(-3.9132915844675153e-05)),(to_sfixed_a(1.7400940123479813e-05)),(to_sfixed_a(-0.00018868438201025128)),(to_sfixed_a(-0.00010617046791594476)),(to_sfixed_a(-7.896337046986446e-05)),(to_sfixed_a(-7.030799315543845e-05)),(to_sfixed_a(-6.80097728036344e-05)),(to_sfixed_a(-0.00011189384531462565)),(to_sfixed_a(0.00024795817444100976)),(to_sfixed_a(-0.0001271688670385629)),(to_sfixed_a(-7.011371781118214e-05)),(to_sfixed_a(-7.180833199527115e-05)),(to_sfixed_a(-0.00010579847730696201)),(to_sfixed_a(8.315519517054781e-05)),(to_sfixed_a(6.753361958544701e-07)),(to_sfixed_a(0.000129307372844778)),(to_sfixed_a(-7.002479105722159e-05)),(to_sfixed_a(-0.00016738404519855976)),(to_sfixed_a(-3.7639329093508422e-06)),(to_sfixed_a(6.514223059639335e-06)),(to_sfixed_a(0.00023701471218373626)),(to_sfixed_a(4.8973201046464965e-05)),(to_sfixed_a(0.0001907187106553465)),(to_sfixed_a(-0.0002059554390143603)),(to_sfixed_a(0.00021953796385787427)),(to_sfixed_a(9.018345735967159e-05)),(to_sfixed_a(-0.00028326865867711604)),(to_sfixed_a(-3.320059840916656e-05)),(to_sfixed_a(-0.00022756410180591047)),(to_sfixed_a(-0.00010565028060227633)),(to_sfixed_a(0.00024015840608626604)),(to_sfixed_a(-0.00021086857304908335)),(to_sfixed_a(-0.00012052751844748855)),(to_sfixed_a(-5.293343565426767e-05)),(to_sfixed_a(0.0001700255088508129)),(to_sfixed_a(-3.624544478952885e-05)),(to_sfixed_a(0.00011690022802213207)),(to_sfixed_a(1.7446691344957799e-06)),(to_sfixed_a(-0.000172157131601125)),(to_sfixed_a(0.00011655237176455557)),(to_sfixed_a(-0.00027159429737366736)),(to_sfixed_a(-4.5351043809205294e-07)),(to_sfixed_a(4.739478754345328e-06)),(to_sfixed_a(-7.643583376193419e-05)),(to_sfixed_a(-0.0001509102585259825)),(to_sfixed_a(-5.838801007485017e-05)),(to_sfixed_a(0.00014557027316186577)),(to_sfixed_a(6.692881288472563e-05)),(to_sfixed_a(-0.00017770074191503227)),(to_sfixed_a(5.793158197775483e-05)),(to_sfixed_a(0.0002950623747892678)),(to_sfixed_a(-5.8880548749584705e-05)),(to_sfixed_a(7.137260399758816e-05)),(to_sfixed_a(-0.00020020102965645492)),(to_sfixed_a(0.00012973553384654224)),(to_sfixed_a(0.0002853356418199837)),(to_sfixed_a(5.6819662859197706e-05)),(to_sfixed_a(0.00016796881391201168)),(to_sfixed_a(-5.9647500165738165e-06)),(to_sfixed_a(9.787920862436295e-05)),(to_sfixed_a(6.760485121048987e-05)),(to_sfixed_a(3.145112714264542e-05)),(to_sfixed_a(6.975750147830695e-05)),(to_sfixed_a(-0.00015124141646083444)),(to_sfixed_a(8.069226169027388e-06)),(to_sfixed_a(7.93521394371055e-05)),(to_sfixed_a(-0.00010305390605935827)),(to_sfixed_a(-7.112635648809373e-05)),(to_sfixed_a(-8.538130350643769e-05)),(to_sfixed_a(-0.0002263169299112633)),(to_sfixed_a(-0.00041676830733194947)),(to_sfixed_a(0.00019941560458391905)),(to_sfixed_a(-0.00022784204338677227)),(to_sfixed_a(-9.196769678965211e-05)),(to_sfixed_a(-0.00013731399667449296)),(to_sfixed_a(-3.9500489947386086e-05)),(to_sfixed_a(0.00011355207243468612)),(to_sfixed_a(0.00014601774455513805)),(to_sfixed_a(0.00011544092558324337)),(to_sfixed_a(-0.00016864860663190484)),(to_sfixed_a(-0.00014787045074626803)),(to_sfixed_a(-0.0001126719216699712)),(to_sfixed_a(0.00023587755276821554)),(to_sfixed_a(-4.819534660782665e-05)),(to_sfixed_a(-7.998733053682372e-05)),(to_sfixed_a(4.7726178308948874e-05)),(to_sfixed_a(-2.013843368331436e-05)),(to_sfixed_a(0.0001362746552331373)),(to_sfixed_a(-2.09314857784193e-05)),(to_sfixed_a(0.00011562589497771114)),(to_sfixed_a(0.00022241839906200767)),(to_sfixed_a(0.00015326208085753024)),(to_sfixed_a(0.00014998162805568427)),(to_sfixed_a(6.0713795392075554e-05)),(to_sfixed_a(1.5713143511675298e-05)),(to_sfixed_a(1.0469848348293453e-06)),(to_sfixed_a(-0.00011723889474524185)),(to_sfixed_a(-2.229688107036054e-06)),(to_sfixed_a(9.313298505730927e-05)),(to_sfixed_a(-0.0002468838356435299)),(to_sfixed_a(0.000247189833316952)),(to_sfixed_a(-0.00020041828975081444)),(to_sfixed_a(-0.0001426785602234304)),(to_sfixed_a(-9.016495823743753e-06)),(to_sfixed_a(0.00010824152559507638)),(to_sfixed_a(-0.0004523933748714626)),(to_sfixed_a(-8.554814849048853e-05)),(to_sfixed_a(-7.155607454478741e-05)),(to_sfixed_a(2.2630054445471615e-05)),(to_sfixed_a(-4.709208951680921e-05)),(to_sfixed_a(-9.750308527145535e-05)),(to_sfixed_a(1.1360862117726356e-05)),(to_sfixed_a(-0.00015611109847668558)),(to_sfixed_a(-1.1852538591483608e-05)),(to_sfixed_a(0.00018061662558466196)),(to_sfixed_a(0.0001289533538511023)),(to_sfixed_a(2.0198229321977124e-05)),(to_sfixed_a(0.00010128138092113659)),(to_sfixed_a(-1.655772575759329e-05)),(to_sfixed_a(0.00029991494375281036)),(to_sfixed_a(-5.1694260037038475e-06)),(to_sfixed_a(-0.00017404179379809648)),(to_sfixed_a(-0.00014821579679846764)),(to_sfixed_a(-8.181384328054264e-05)),(to_sfixed_a(1.6888821846805513e-05)),(to_sfixed_a(-2.299995321664028e-05)),(to_sfixed_a(0.0002141384029528126)),(to_sfixed_a(0.00020455448247957975)),(to_sfixed_a(0.0002982188016176224)),(to_sfixed_a(2.4457116523990408e-05)),(to_sfixed_a(4.747309139929712e-05)),(to_sfixed_a(-0.0003131665289402008)),(to_sfixed_a(0.00017807097174227238)),(to_sfixed_a(-0.00022980858921073377)),(to_sfixed_a(-0.00010237125388812274)),(to_sfixed_a(1.4830169675406069e-05)),(to_sfixed_a(0.00011195256956852973)),(to_sfixed_a(-1.7001213564071804e-05)),(to_sfixed_a(0.0001415805018041283)),(to_sfixed_a(-8.737774624023587e-05)),(to_sfixed_a(3.865941835101694e-05)),(to_sfixed_a(-0.00029470736626535654)),(to_sfixed_a(-3.714820559252985e-05)),(to_sfixed_a(-3.149130861856975e-05)),(to_sfixed_a(-0.00012927295756526291)),(to_sfixed_a(-4.281660949345678e-06)),(to_sfixed_a(-7.089781138347462e-05)),(to_sfixed_a(-0.00022341076692100614)),(to_sfixed_a(0.00012956665887031704)),(to_sfixed_a(0.00011180095316376537)),(to_sfixed_a(-0.00020572126959450543)),(to_sfixed_a(-0.00016561834490858018)),(to_sfixed_a(0.00011652577086351812)),(to_sfixed_a(6.090129318181425e-06)),(to_sfixed_a(-4.9443526222603396e-05)),(to_sfixed_a(2.4638735339976847e-05)),(to_sfixed_a(2.3640521249035373e-05)),(to_sfixed_a(-8.722557686269283e-05)),(to_sfixed_a(-4.088896093890071e-05)),(to_sfixed_a(5.795087054139003e-05)),(to_sfixed_a(0.00012746299034915864)),(to_sfixed_a(-5.731578130507842e-05)),(to_sfixed_a(9.796662197913975e-05)),(to_sfixed_a(-8.617935236543417e-07)),(to_sfixed_a(1.1891177564393729e-05)),(to_sfixed_a(-7.115615881048143e-05)),(to_sfixed_a(0.00032310461392626166)),(to_sfixed_a(0.00015681581862736493)),(to_sfixed_a(0.00014785882376600057)),(to_sfixed_a(-0.0002368787390878424)),(to_sfixed_a(2.3180411517387256e-05)),(to_sfixed_a(-0.0002966286556329578)),(to_sfixed_a(-1.1065929356846027e-05)),(to_sfixed_a(-0.0001498161582276225)),(to_sfixed_a(-7.335786358453333e-05)),(to_sfixed_a(-6.260530062718317e-05)),(to_sfixed_a(0.00012750312453135848)),(to_sfixed_a(2.0227671484462917e-06)),(to_sfixed_a(-7.73514766478911e-05)),(to_sfixed_a(3.911659223376773e-05)),(to_sfixed_a(0.00012580926704686135)),(to_sfixed_a(-0.00018356679356656969)));

    constant weight_n2_84 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.14054161310195923)),(to_sfixed_a(0.00014935355284251273)),(to_sfixed_a(-0.0005485427100211382)),(to_sfixed_a(-0.00010626696166582406)),(to_sfixed_a(0.017795182764530182)),(to_sfixed_a(-3.850090433843434e-05)),(to_sfixed_a(-0.0015869532944634557)),(to_sfixed_a(8.165562758222222e-05)),(to_sfixed_a(6.016940824338235e-05)),(to_sfixed_a(1.1320225894451141e-06)),(to_sfixed_a(0.00010974879842251539)),(to_sfixed_a(-0.0014858460053801537)),(to_sfixed_a(0.2126595824956894)),(to_sfixed_a(0.004515317268669605)),(to_sfixed_a(3.0189432436600327e-05)),(to_sfixed_a(8.539945702068508e-05)),(to_sfixed_a(0.0001053988016792573)),(to_sfixed_a(-6.899250001879409e-05)),(to_sfixed_a(0.011989698745310307)),(to_sfixed_a(0.5451145172119141)),(to_sfixed_a(-0.00016453911666758358)),(to_sfixed_a(-0.00011711417755577713)),(to_sfixed_a(-0.0007523818057961762)),(to_sfixed_a(-0.0008897182997316122)),(to_sfixed_a(-0.003694054903462529)),(to_sfixed_a(-0.0041749621741473675)),(to_sfixed_a(-0.00015118550800252706)),(to_sfixed_a(0.0008853923063725233)),(to_sfixed_a(-0.002910957206040621)),(to_sfixed_a(-0.00018655632447917014)),(to_sfixed_a(0.0026094026397913694)),(to_sfixed_a(-7.114918844308704e-05)),(to_sfixed_a(0.1888015866279602)),(to_sfixed_a(-2.835600753314793e-05)),(to_sfixed_a(0.00010455770825501531)),(to_sfixed_a(0.00017221641610376537)),(to_sfixed_a(0.0040666405111551285)),(to_sfixed_a(-0.15620163083076477)),(to_sfixed_a(-0.27146977186203003)),(to_sfixed_a(3.7332316423999146e-05)),(to_sfixed_a(-0.004568647127598524)),(to_sfixed_a(0.0016239732503890991)),(to_sfixed_a(-0.0001721050648484379)),(to_sfixed_a(0.0002342141669942066)),(to_sfixed_a(-0.1875099390745163)),(to_sfixed_a(-0.005017862655222416)),(to_sfixed_a(0.0008960051345638931)),(to_sfixed_a(-0.014546002261340618)),(to_sfixed_a(-6.391666829586029e-05)),(to_sfixed_a(-0.006758802570402622)),(to_sfixed_a(0.0005794721655547619)),(to_sfixed_a(-0.0012871884973719716)),(to_sfixed_a(0.0002688225940801203)),(to_sfixed_a(0.002446783008053899)),(to_sfixed_a(-0.005210179835557938)),(to_sfixed_a(-0.0012126057408750057)),(to_sfixed_a(-0.0001552020403323695)),(to_sfixed_a(-0.002446696860715747)),(to_sfixed_a(1.0569841833785176e-05)),(to_sfixed_a(-7.822563929948956e-05)),(to_sfixed_a(-0.0007144931005313993)),(to_sfixed_a(-0.0013530742144212127)),(to_sfixed_a(-0.0008317462634295225)),(to_sfixed_a(0.007419710513204336)),(to_sfixed_a(-0.00022730026103090495)),(to_sfixed_a(-0.00919388048350811)),(to_sfixed_a(-0.00010550308070378378)),(to_sfixed_a(0.0019614044576883316)),(to_sfixed_a(-0.00354603654704988)),(to_sfixed_a(0.00011232275574002415)),(to_sfixed_a(0.004890882410109043)),(to_sfixed_a(-0.0018267510458827019)),(to_sfixed_a(0.2110876888036728)),(to_sfixed_a(-7.071414438541979e-05)),(to_sfixed_a(-5.6925327953649685e-05)),(to_sfixed_a(6.298845983110368e-05)),(to_sfixed_a(-0.09614436328411102)),(to_sfixed_a(0.25828686356544495)),(to_sfixed_a(2.0601219148375094e-05)),(to_sfixed_a(0.022012174129486084)),(to_sfixed_a(-0.0006040803855285048)),(to_sfixed_a(-0.00011194541002623737)),(to_sfixed_a(-0.001824043458327651)),(to_sfixed_a(0.006559882778674364)),(to_sfixed_a(-0.00014779125922359526)),(to_sfixed_a(0.008965757675468922)),(to_sfixed_a(-0.01993831992149353)),(to_sfixed_a(-0.00041736342245712876)),(to_sfixed_a(7.123093382688239e-05)),(to_sfixed_a(-0.0002003332629101351)),(to_sfixed_a(0.016530655324459076)),(to_sfixed_a(-2.88133742287755e-05)),(to_sfixed_a(0.22485661506652832)),(to_sfixed_a(3.193491284037009e-05)),(to_sfixed_a(0.2721767723560333)),(to_sfixed_a(-3.0146900826366618e-05)),(to_sfixed_a(-6.968537491047755e-05)),(to_sfixed_a(2.6177367544732988e-05)),(to_sfixed_a(5.857380892848596e-05)),(to_sfixed_a(-1.727984636090696e-05)),(to_sfixed_a(-0.011624589562416077)),(to_sfixed_a(-0.00122252746950835)),(to_sfixed_a(-0.00042254605796188116)),(to_sfixed_a(0.0005286643281579018)),(to_sfixed_a(0.008535554632544518)),(to_sfixed_a(-0.16811677813529968)),(to_sfixed_a(0.00012875838729087263)),(to_sfixed_a(6.205511454027146e-05)),(to_sfixed_a(-0.0001837957534007728)),(to_sfixed_a(-0.14444129168987274)),(to_sfixed_a(0.0015550855314359069)),(to_sfixed_a(-1.6241654520854354e-05)),(to_sfixed_a(0.25339311361312866)),(to_sfixed_a(-2.9733566407230683e-05)),(to_sfixed_a(3.7299079849617556e-05)),(to_sfixed_a(0.007195711135864258)),(to_sfixed_a(0.0033204681240022182)),(to_sfixed_a(-0.004217073321342468)),(to_sfixed_a(-3.608452243497595e-05)),(to_sfixed_a(-0.0006212295265868306)),(to_sfixed_a(-3.8245212635956705e-05)),(to_sfixed_a(9.91017441265285e-06)),(to_sfixed_a(0.0025675774086266756)),(to_sfixed_a(5.1880069804610685e-05)),(to_sfixed_a(0.00015059515135362744)),(to_sfixed_a(0.23056554794311523)),(to_sfixed_a(0.006910047028213739)),(to_sfixed_a(-0.00010241138807032257)),(to_sfixed_a(-6.180698983371258e-05)),(to_sfixed_a(6.506832141894847e-05)),(to_sfixed_a(-0.0001121709865401499)),(to_sfixed_a(-4.611282201949507e-05)),(to_sfixed_a(-4.3084422941319644e-05)),(to_sfixed_a(0.013174599967896938)),(to_sfixed_a(-4.6063505578786135e-06)),(to_sfixed_a(-0.0001564708218211308)),(to_sfixed_a(-0.40718257427215576)),(to_sfixed_a(-0.00017107941675931215)),(to_sfixed_a(-4.158602678216994e-06)),(to_sfixed_a(9.174994920613244e-05)),(to_sfixed_a(-6.711269088555127e-05)),(to_sfixed_a(-0.00023249424702953547)),(to_sfixed_a(6.938633305253461e-05)),(to_sfixed_a(0.0012347609736025333)),(to_sfixed_a(-0.0016879242612048984)),(to_sfixed_a(0.003115659113973379)),(to_sfixed_a(0.0013885971857234836)),(to_sfixed_a(2.657193545019254e-05)),(to_sfixed_a(0.00011338886542944238)),(to_sfixed_a(0.003526422893628478)),(to_sfixed_a(0.00010245675366604701)),(to_sfixed_a(-2.1973828552290797e-06)),(to_sfixed_a(-0.0024232622236013412)),(to_sfixed_a(0.00025087245739996433)),(to_sfixed_a(3.754257704713382e-05)),(to_sfixed_a(-0.016926495358347893)),(to_sfixed_a(-9.581322956364602e-06)),(to_sfixed_a(-0.004808661062270403)),(to_sfixed_a(8.198575960705057e-05)),(to_sfixed_a(0.0001279084972338751)),(to_sfixed_a(-0.00024262390797957778)),(to_sfixed_a(0.00010241303243674338)),(to_sfixed_a(0.001288411789573729)),(to_sfixed_a(0.00010357380961067975)),(to_sfixed_a(-0.015290208160877228)),(to_sfixed_a(0.003746303729712963)),(to_sfixed_a(5.941909330431372e-05)),(to_sfixed_a(-0.3129376769065857)),(to_sfixed_a(4.5779888750985265e-06)),(to_sfixed_a(0.00015544501366093755)),(to_sfixed_a(-0.012517188675701618)),(to_sfixed_a(0.0013669815380126238)),(to_sfixed_a(-0.016688883304595947)),(to_sfixed_a(0.0002452404878567904)),(to_sfixed_a(-0.3317644000053406)),(to_sfixed_a(-0.004996137693524361)),(to_sfixed_a(0.18787911534309387)),(to_sfixed_a(-0.0008930756594054401)),(to_sfixed_a(-0.04358657822012901)),(to_sfixed_a(0.0031073589343577623)),(to_sfixed_a(-0.0013437489978969097)),(to_sfixed_a(0.01778835617005825)),(to_sfixed_a(-0.0002380804653512314)),(to_sfixed_a(6.734502676408738e-05)),(to_sfixed_a(2.3256732674781233e-05)),(to_sfixed_a(0.2284727394580841)),(to_sfixed_a(-0.006120759062469006)),(to_sfixed_a(0.24713213741779327)),(to_sfixed_a(0.0030018442776054144)),(to_sfixed_a(0.005407107062637806)),(to_sfixed_a(0.012088874354958534)),(to_sfixed_a(7.853604620322585e-05)),(to_sfixed_a(-0.010416229255497456)),(to_sfixed_a(0.01437093410640955)),(to_sfixed_a(-2.090570706059225e-05)),(to_sfixed_a(-0.0005789148854091763)),(to_sfixed_a(4.495041139307432e-05)),(to_sfixed_a(0.009487126022577286)),(to_sfixed_a(-0.004287916235625744)),(to_sfixed_a(5.7159995776601136e-05)),(to_sfixed_a(5.7437333452980965e-05)),(to_sfixed_a(4.483065276872367e-05)),(to_sfixed_a(-1.2070908269379288e-05)),(to_sfixed_a(-7.12581240804866e-05)),(to_sfixed_a(1.9275939848739654e-05)),(to_sfixed_a(-0.0013523069210350513)),(to_sfixed_a(-0.0023930303286761045)),(to_sfixed_a(0.025678060948848724)),(to_sfixed_a(-0.40649813413619995)),(to_sfixed_a(-0.20175467431545258)),(to_sfixed_a(0.005336340982466936)),(to_sfixed_a(-6.0044112615287304e-05)),(to_sfixed_a(2.4795222998363897e-05)),(to_sfixed_a(9.574260184308514e-05)),(to_sfixed_a(0.00021698587806895375)),(to_sfixed_a(-2.8453989216359332e-05)),(to_sfixed_a(0.002041025087237358)),(to_sfixed_a(0.00015865171735640615)),(to_sfixed_a(-0.0007464558002538979)),(to_sfixed_a(-0.00023100629914551973)),(to_sfixed_a(0.0002880091196857393)),(to_sfixed_a(0.00027334477636031806)),(to_sfixed_a(-1.2547076039481908e-05)),(to_sfixed_a(0.4337954819202423)),(to_sfixed_a(0.26706427335739136)),(to_sfixed_a(-0.00013718268019147217)),(to_sfixed_a(-2.065183434751816e-05)),(to_sfixed_a(5.980225978419185e-06)),(to_sfixed_a(-0.2482464611530304)),(to_sfixed_a(0.00021350212045945227)),(to_sfixed_a(-0.004003841895610094)),(to_sfixed_a(-8.485202852170914e-05)),(to_sfixed_a(0.00013009659596718848)),(to_sfixed_a(-2.059827238554135e-05)),(to_sfixed_a(-0.007989569567143917)),(to_sfixed_a(0.015614851377904415)),(to_sfixed_a(-0.0071547687985002995)),(to_sfixed_a(-8.478482050122693e-05)),(to_sfixed_a(0.005410567857325077)),(to_sfixed_a(-1.8759543308988214e-05)),(to_sfixed_a(0.30046898126602173)),(to_sfixed_a(8.156232070177794e-06)),(to_sfixed_a(0.31423136591911316)),(to_sfixed_a(0.00018094322877004743)),(to_sfixed_a(0.00046653312165290117)),(to_sfixed_a(-0.001537702395580709)),(to_sfixed_a(-0.06487499922513962)),(to_sfixed_a(0.39816638827323914)),(to_sfixed_a(0.00014707079390063882)),(to_sfixed_a(-0.38988396525382996)),(to_sfixed_a(-0.01867908611893654)),(to_sfixed_a(1.1628690117504448e-05)),(to_sfixed_a(-0.0004611258627846837)),(to_sfixed_a(0.0001771084644133225)),(to_sfixed_a(-4.316767444834113e-06)),(to_sfixed_a(-0.0034841857850551605)),(to_sfixed_a(-0.0017546655144542456)),(to_sfixed_a(-8.585149771533906e-06)),(to_sfixed_a(0.00016683975991327316)),(to_sfixed_a(-0.0012612289283424616)),(to_sfixed_a(-0.00031651818426325917)),(to_sfixed_a(-0.015500766225159168)),(to_sfixed_a(-0.00010608749289531261)),(to_sfixed_a(-0.00033853689092211425)),(to_sfixed_a(-6.052220851415768e-05)),(to_sfixed_a(-0.001989849144592881)),(to_sfixed_a(2.6516827347222716e-05)),(to_sfixed_a(0.00011372077278792858)),(to_sfixed_a(-6.158080941531807e-05)),(to_sfixed_a(-0.0012529336381703615)),(to_sfixed_a(0.5648377537727356)),(to_sfixed_a(0.00019662329577840865)),(to_sfixed_a(6.356067024171352e-05)),(to_sfixed_a(-0.00016707388567738235)),(to_sfixed_a(3.063331314479001e-05)),(to_sfixed_a(0.36828652024269104)),(to_sfixed_a(-0.2533215582370758)),(to_sfixed_a(-0.06806941330432892)),(to_sfixed_a(0.004333257209509611)),(to_sfixed_a(0.0021607151720672846)),(to_sfixed_a(0.00014174316311255097)),(to_sfixed_a(0.00018772164185065776)),(to_sfixed_a(0.00044995584175921977)),(to_sfixed_a(0.001409107819199562)),(to_sfixed_a(1.1515585356391966e-05)),(to_sfixed_a(0.00037707906449213624)),(to_sfixed_a(0.0005826972192153335)),(to_sfixed_a(0.4006863832473755)),(to_sfixed_a(-1.022921787807718e-05)),(to_sfixed_a(0.18757419288158417)),(to_sfixed_a(0.2918364405632019)),(to_sfixed_a(-0.012420810759067535)),(to_sfixed_a(0.003457808867096901)),(to_sfixed_a(0.00015174163854680955)),(to_sfixed_a(-0.004242993891239166)),(to_sfixed_a(-0.0008249988895840943)),(to_sfixed_a(-0.020300408825278282)),(to_sfixed_a(0.00011269650713074952)),(to_sfixed_a(-0.04062376171350479)),(to_sfixed_a(0.7634978890419006)),(to_sfixed_a(-0.011979001574218273)));

    constant weight_n2_85 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.20128607749938965)),(to_sfixed_a(0.2342565357685089)),(to_sfixed_a(0.0004053141747135669)),(to_sfixed_a(0.00011510804324643686)),(to_sfixed_a(0.0011351199354976416)),(to_sfixed_a(0.00011262287443969399)),(to_sfixed_a(-0.3487052023410797)),(to_sfixed_a(0.0001549823791719973)),(to_sfixed_a(0.00010374787962064147)),(to_sfixed_a(2.7048845367971808e-06)),(to_sfixed_a(0.000302600470604375)),(to_sfixed_a(0.01392614096403122)),(to_sfixed_a(0.006152500864118338)),(to_sfixed_a(0.024339932948350906)),(to_sfixed_a(-8.532311767339706e-05)),(to_sfixed_a(0.0002946064341813326)),(to_sfixed_a(0.008833354339003563)),(to_sfixed_a(8.417728531640023e-05)),(to_sfixed_a(0.286965012550354)),(to_sfixed_a(-0.00020995836530346423)),(to_sfixed_a(9.8936099675484e-05)),(to_sfixed_a(-2.8723879950121045e-05)),(to_sfixed_a(-0.00013074673188384622)),(to_sfixed_a(-0.0073386733420193195)),(to_sfixed_a(0.0005502818385139108)),(to_sfixed_a(-0.0021909300703555346)),(to_sfixed_a(-2.4841196136549115e-05)),(to_sfixed_a(-0.3710055649280548)),(to_sfixed_a(0.0005223563057370484)),(to_sfixed_a(6.121982005424798e-05)),(to_sfixed_a(0.0049249702133238316)),(to_sfixed_a(-5.8653335145208985e-05)),(to_sfixed_a(0.011895681731402874)),(to_sfixed_a(3.6548553907778114e-05)),(to_sfixed_a(2.370043148403056e-05)),(to_sfixed_a(-0.0002998589479830116)),(to_sfixed_a(0.4635184407234192)),(to_sfixed_a(0.0164467915892601)),(to_sfixed_a(0.24083158373832703)),(to_sfixed_a(-0.0004505031101871282)),(to_sfixed_a(0.0042246137745678425)),(to_sfixed_a(0.04348143935203552)),(to_sfixed_a(-0.00016952306032180786)),(to_sfixed_a(0.00018127736984752119)),(to_sfixed_a(0.005795920267701149)),(to_sfixed_a(0.02439606375992298)),(to_sfixed_a(-0.002687235129997134)),(to_sfixed_a(0.0005507580353878438)),(to_sfixed_a(6.764883437426761e-05)),(to_sfixed_a(-0.1599116325378418)),(to_sfixed_a(0.14346376061439514)),(to_sfixed_a(0.000864161760546267)),(to_sfixed_a(1.7883849068311974e-06)),(to_sfixed_a(0.0023481023963540792)),(to_sfixed_a(0.04591439664363861)),(to_sfixed_a(-0.009769015945494175)),(to_sfixed_a(0.00029315362917259336)),(to_sfixed_a(0.005823442712426186)),(to_sfixed_a(4.794468986801803e-05)),(to_sfixed_a(8.511403575539589e-05)),(to_sfixed_a(0.0006666409317404032)),(to_sfixed_a(0.0009612469584681094)),(to_sfixed_a(-0.0016744957538321614)),(to_sfixed_a(-0.03621261194348335)),(to_sfixed_a(-0.00023895471531432122)),(to_sfixed_a(-0.013868439942598343)),(to_sfixed_a(1.035921013681218e-05)),(to_sfixed_a(0.40478330850601196)),(to_sfixed_a(-0.0029227875638753176)),(to_sfixed_a(8.39323183754459e-06)),(to_sfixed_a(-0.06786587089300156)),(to_sfixed_a(-0.5019012093544006)),(to_sfixed_a(0.28470781445503235)),(to_sfixed_a(-4.628534225048497e-05)),(to_sfixed_a(0.00010337537969462574)),(to_sfixed_a(-0.0001366916549159214)),(to_sfixed_a(0.022664425894618034)),(to_sfixed_a(-0.0001381135662086308)),(to_sfixed_a(-6.809148180764169e-05)),(to_sfixed_a(-0.0021200350020080805)),(to_sfixed_a(-5.528676410904154e-05)),(to_sfixed_a(2.4821303668431938e-05)),(to_sfixed_a(0.024483220651745796)),(to_sfixed_a(-0.0023698078002780676)),(to_sfixed_a(-2.1996291252435185e-05)),(to_sfixed_a(-0.16848905384540558)),(to_sfixed_a(0.35869669914245605)),(to_sfixed_a(0.00834780465811491)),(to_sfixed_a(-7.1699709224049e-05)),(to_sfixed_a(3.990741970483214e-05)),(to_sfixed_a(-0.006887029390782118)),(to_sfixed_a(-6.423283775802702e-05)),(to_sfixed_a(-0.2655044198036194)),(to_sfixed_a(0.0001554932096041739)),(to_sfixed_a(0.33693358302116394)),(to_sfixed_a(0.00010707449109759182)),(to_sfixed_a(0.0001859218318713829)),(to_sfixed_a(-7.160725363064557e-05)),(to_sfixed_a(1.075044747267384e-05)),(to_sfixed_a(3.983135684393346e-06)),(to_sfixed_a(0.002918662503361702)),(to_sfixed_a(0.008341523818671703)),(to_sfixed_a(-0.00029411716968752444)),(to_sfixed_a(-0.32848843932151794)),(to_sfixed_a(-0.007618552073836327)),(to_sfixed_a(0.0008172154775820673)),(to_sfixed_a(-7.361545431194827e-05)),(to_sfixed_a(-5.2908784709870815e-05)),(to_sfixed_a(3.0735216569155455e-05)),(to_sfixed_a(-0.28540411591529846)),(to_sfixed_a(-0.0036785819102078676)),(to_sfixed_a(2.1913248929195106e-05)),(to_sfixed_a(0.2034837305545807)),(to_sfixed_a(6.301306711975485e-05)),(to_sfixed_a(-0.00022428701049648225)),(to_sfixed_a(-0.10334467887878418)),(to_sfixed_a(0.01576172187924385)),(to_sfixed_a(-0.0017336257733404636)),(to_sfixed_a(-3.986497176811099e-07)),(to_sfixed_a(-0.017915114760398865)),(to_sfixed_a(0.0001266449980903417)),(to_sfixed_a(7.15658679837361e-05)),(to_sfixed_a(0.006350470706820488)),(to_sfixed_a(-3.79121775040403e-05)),(to_sfixed_a(-5.9458201576489955e-05)),(to_sfixed_a(0.3565269410610199)),(to_sfixed_a(0.004912118893116713)),(to_sfixed_a(-0.00011568097397685051)),(to_sfixed_a(-0.0001917273475555703)),(to_sfixed_a(-6.45002000965178e-05)),(to_sfixed_a(-1.4511129847960547e-05)),(to_sfixed_a(-0.000315716490149498)),(to_sfixed_a(-0.00013601449609268457)),(to_sfixed_a(0.016498593613505363)),(to_sfixed_a(-7.220447878353298e-05)),(to_sfixed_a(4.7202076530084014e-05)),(to_sfixed_a(-0.025356391444802284)),(to_sfixed_a(0.00017070583999156952)),(to_sfixed_a(-0.00021358559024520218)),(to_sfixed_a(0.00015802509733475745)),(to_sfixed_a(0.24611525237560272)),(to_sfixed_a(3.64048573828768e-05)),(to_sfixed_a(-0.00011324630759190768)),(to_sfixed_a(0.026464004069566727)),(to_sfixed_a(-0.0045729330740869045)),(to_sfixed_a(0.005010404158383608)),(to_sfixed_a(0.0004962034290656447)),(to_sfixed_a(0.00010078713239636272)),(to_sfixed_a(0.00014003575779497623)),(to_sfixed_a(-0.014892748557031155)),(to_sfixed_a(0.0002170264779124409)),(to_sfixed_a(0.00045162817696109414)),(to_sfixed_a(0.004679224453866482)),(to_sfixed_a(0.00010365302296122536)),(to_sfixed_a(-0.00029172905487939715)),(to_sfixed_a(6.399624544428661e-05)),(to_sfixed_a(-0.00020171205687802285)),(to_sfixed_a(0.34461063146591187)),(to_sfixed_a(6.854921139165526e-06)),(to_sfixed_a(-0.00011249280214542523)),(to_sfixed_a(-2.3577522370032966e-06)),(to_sfixed_a(1.080325455404818e-05)),(to_sfixed_a(0.015744147822260857)),(to_sfixed_a(0.0017710562096908689)),(to_sfixed_a(0.0007823449559509754)),(to_sfixed_a(-0.14093875885009766)),(to_sfixed_a(-0.00041083560790866613)),(to_sfixed_a(0.39462053775787354)),(to_sfixed_a(-0.00013001347542740405)),(to_sfixed_a(0.00014187002670951188)),(to_sfixed_a(0.008679194375872612)),(to_sfixed_a(-0.004190649837255478)),(to_sfixed_a(-0.006057041697204113)),(to_sfixed_a(6.936813588254154e-05)),(to_sfixed_a(-0.005941182374954224)),(to_sfixed_a(-0.0010648377938196063)),(to_sfixed_a(-0.0025868143420666456)),(to_sfixed_a(0.0007668499602004886)),(to_sfixed_a(-0.009083010256290436)),(to_sfixed_a(-0.4871213734149933)),(to_sfixed_a(0.00039085280150175095)),(to_sfixed_a(0.46043798327445984)),(to_sfixed_a(0.00030832350603304803)),(to_sfixed_a(-4.920705396216363e-05)),(to_sfixed_a(-0.00041133392369374633)),(to_sfixed_a(-0.00015271329903043807)),(to_sfixed_a(0.3964695930480957)),(to_sfixed_a(0.00048168544890359044)),(to_sfixed_a(0.3889884054660797)),(to_sfixed_a(0.0005624178447760642)),(to_sfixed_a(0.31294283270835876)),(to_sfixed_a(-4.55184344900772e-05)),(to_sfixed_a(0.017949244007468224)),(to_sfixed_a(-0.09557370841503143)),(to_sfixed_a(-4.1444392991252244e-05)),(to_sfixed_a(-0.005734799895435572)),(to_sfixed_a(4.916222678730264e-05)),(to_sfixed_a(0.00998193584382534)),(to_sfixed_a(-0.4254993796348572)),(to_sfixed_a(2.4393375497311354e-07)),(to_sfixed_a(3.863220626953989e-06)),(to_sfixed_a(-0.0001686920877546072)),(to_sfixed_a(-3.082001057919115e-06)),(to_sfixed_a(-7.976276538101956e-05)),(to_sfixed_a(0.00011453318438725546)),(to_sfixed_a(-0.020885668694972992)),(to_sfixed_a(0.06064719706773758)),(to_sfixed_a(0.3263564109802246)),(to_sfixed_a(0.3770851194858551)),(to_sfixed_a(0.0006625856622122228)),(to_sfixed_a(-0.0006220282521098852)),(to_sfixed_a(-4.780414383276366e-05)),(to_sfixed_a(0.00023673295800108463)),(to_sfixed_a(6.542708433698863e-05)),(to_sfixed_a(-1.4840654330328107e-05)),(to_sfixed_a(0.0002836073108483106)),(to_sfixed_a(0.010095181874930859)),(to_sfixed_a(0.004614824894815683)),(to_sfixed_a(0.007460631430149078)),(to_sfixed_a(-0.00012902516755275428)),(to_sfixed_a(-0.00013657205272465944)),(to_sfixed_a(-6.94136178935878e-05)),(to_sfixed_a(3.71807036572136e-05)),(to_sfixed_a(0.0003300987009424716)),(to_sfixed_a(0.0014702974585816264)),(to_sfixed_a(2.5475492293480784e-07)),(to_sfixed_a(-2.896923979278654e-05)),(to_sfixed_a(-0.0004563575785141438)),(to_sfixed_a(-0.2922889292240143)),(to_sfixed_a(-0.20997510850429535)),(to_sfixed_a(-0.007179793436080217)),(to_sfixed_a(7.608263695146888e-05)),(to_sfixed_a(2.0532766939140856e-05)),(to_sfixed_a(0.00011211234232177958)),(to_sfixed_a(-0.13556575775146484)),(to_sfixed_a(0.019885100424289703)),(to_sfixed_a(-0.0014550811611115932)),(to_sfixed_a(-0.0002698359021451324)),(to_sfixed_a(-1.3338649296201766e-05)),(to_sfixed_a(3.509423913783394e-05)),(to_sfixed_a(-0.5781781077384949)),(to_sfixed_a(-1.8480714061297476e-05)),(to_sfixed_a(-0.12228646874427795)),(to_sfixed_a(6.830011261627078e-05)),(to_sfixed_a(0.015418345108628273)),(to_sfixed_a(0.41567495465278625)),(to_sfixed_a(-0.20977845788002014)),(to_sfixed_a(-0.2288840264081955)),(to_sfixed_a(0.00016734057862777263)),(to_sfixed_a(0.0024700849317014217)),(to_sfixed_a(-0.0006737762596458197)),(to_sfixed_a(-7.12585388100706e-05)),(to_sfixed_a(0.005962766241282225)),(to_sfixed_a(3.415047831367701e-05)),(to_sfixed_a(0.005229519680142403)),(to_sfixed_a(0.02601744420826435)),(to_sfixed_a(-0.0005590313812717795)),(to_sfixed_a(-4.806202196050435e-05)),(to_sfixed_a(-0.00014727184316143394)),(to_sfixed_a(-0.004597448278218508)),(to_sfixed_a(-0.00010609094169922173)),(to_sfixed_a(0.00013678731920663267)),(to_sfixed_a(-6.279382796492428e-05)),(to_sfixed_a(-6.691753515042365e-05)),(to_sfixed_a(0.00013098825002089143)),(to_sfixed_a(0.012364461086690426)),(to_sfixed_a(-6.627055699937046e-05)),(to_sfixed_a(-0.00010573030158411711)),(to_sfixed_a(2.3746855731587857e-05)),(to_sfixed_a(-0.2357180118560791)),(to_sfixed_a(0.01149611547589302)),(to_sfixed_a(0.0003851600631605834)),(to_sfixed_a(-4.986790008842945e-05)),(to_sfixed_a(-0.0002102509024553001)),(to_sfixed_a(-5.833753675688058e-07)),(to_sfixed_a(-0.00573402363806963)),(to_sfixed_a(0.0021540510933846235)),(to_sfixed_a(0.28446099162101746)),(to_sfixed_a(-0.002626276109367609)),(to_sfixed_a(-0.002224538242444396)),(to_sfixed_a(-6.686296546831727e-05)),(to_sfixed_a(-0.0004186522273812443)),(to_sfixed_a(0.00025198361254297197)),(to_sfixed_a(0.00039724810631014407)),(to_sfixed_a(0.00011352337605785578)),(to_sfixed_a(1.0947405826300383e-06)),(to_sfixed_a(0.35171687602996826)),(to_sfixed_a(0.024245133623480797)),(to_sfixed_a(-6.385636515915394e-05)),(to_sfixed_a(0.04625986889004707)),(to_sfixed_a(0.003789168084040284)),(to_sfixed_a(-0.010558223351836205)),(to_sfixed_a(-0.0007106172270141542)),(to_sfixed_a(0.00011274082498857751)),(to_sfixed_a(-0.0015092289540916681)),(to_sfixed_a(0.14239320158958435)),(to_sfixed_a(0.009857607074081898)),(to_sfixed_a(-5.0323385949013755e-05)),(to_sfixed_a(-0.0050416444428265095)),(to_sfixed_a(0.4290074408054352)),(to_sfixed_a(0.0024339696392416954)));

    constant weight_n2_86 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.11194605380296707)),(to_sfixed_a(-0.006075763143599033)),(to_sfixed_a(0.00019372922542970628)),(to_sfixed_a(0.00018033370724879205)),(to_sfixed_a(0.000738640665076673)),(to_sfixed_a(-0.0001394862192682922)),(to_sfixed_a(-0.004473233595490456)),(to_sfixed_a(3.5505865525919944e-05)),(to_sfixed_a(-2.6130452170036733e-05)),(to_sfixed_a(7.15803325874731e-05)),(to_sfixed_a(-1.6051788406912237e-05)),(to_sfixed_a(-0.383405476808548)),(to_sfixed_a(-0.01504733506590128)),(to_sfixed_a(-0.011031005531549454)),(to_sfixed_a(-6.32982118986547e-05)),(to_sfixed_a(-0.0002371152222622186)),(to_sfixed_a(0.10662558674812317)),(to_sfixed_a(-0.00012895003601443022)),(to_sfixed_a(-0.013499844819307327)),(to_sfixed_a(-0.006161018740385771)),(to_sfixed_a(-0.0001566489227116108)),(to_sfixed_a(-3.868692147079855e-06)),(to_sfixed_a(0.0008057450177147985)),(to_sfixed_a(-0.0009915055707097054)),(to_sfixed_a(0.004197125788778067)),(to_sfixed_a(0.012680490501224995)),(to_sfixed_a(1.8362683476880193e-05)),(to_sfixed_a(-0.2980717420578003)),(to_sfixed_a(-0.0023430988658219576)),(to_sfixed_a(6.5410858951509e-09)),(to_sfixed_a(0.3713749647140503)),(to_sfixed_a(3.41630911862012e-05)),(to_sfixed_a(-0.0011517482344061136)),(to_sfixed_a(1.3859316823072731e-06)),(to_sfixed_a(4.4502245145849884e-05)),(to_sfixed_a(-9.896996198222041e-05)),(to_sfixed_a(0.22716204822063446)),(to_sfixed_a(0.20200829207897186)),(to_sfixed_a(-0.46463313698768616)),(to_sfixed_a(-0.00044581477413885295)),(to_sfixed_a(-0.059146177023649216)),(to_sfixed_a(-0.005726139526814222)),(to_sfixed_a(-7.006134546827525e-05)),(to_sfixed_a(0.00014286238001659513)),(to_sfixed_a(-0.0015261791413649917)),(to_sfixed_a(0.3734652101993561)),(to_sfixed_a(-0.00335677620023489)),(to_sfixed_a(9.97809402178973e-05)),(to_sfixed_a(0.0001520495570730418)),(to_sfixed_a(-0.0007861083140596747)),(to_sfixed_a(0.2621566653251648)),(to_sfixed_a(-0.00018783807172439992)),(to_sfixed_a(0.0003150136035401374)),(to_sfixed_a(-0.0027070236392319202)),(to_sfixed_a(0.006219283677637577)),(to_sfixed_a(-0.1102491244673729)),(to_sfixed_a(-0.00028097385074943304)),(to_sfixed_a(-7.346221536863595e-05)),(to_sfixed_a(-2.5162473320961e-05)),(to_sfixed_a(-1.1768133845180273e-06)),(to_sfixed_a(0.002610444789752364)),(to_sfixed_a(-0.00037468134541995823)),(to_sfixed_a(0.0013335173716768622)),(to_sfixed_a(-0.0018282317323610187)),(to_sfixed_a(-7.78325556893833e-05)),(to_sfixed_a(-0.0012793963542208076)),(to_sfixed_a(-0.0002480594557709992)),(to_sfixed_a(0.009935179725289345)),(to_sfixed_a(0.006371039431542158)),(to_sfixed_a(-9.633089575800113e-06)),(to_sfixed_a(0.3514818549156189)),(to_sfixed_a(-0.003311727661639452)),(to_sfixed_a(-0.008851875551044941)),(to_sfixed_a(2.6802670618053526e-05)),(to_sfixed_a(5.859454540768638e-05)),(to_sfixed_a(2.5394219846930355e-06)),(to_sfixed_a(-0.2435666024684906)),(to_sfixed_a(0.0033748445566743612)),(to_sfixed_a(-0.00015070113295223564)),(to_sfixed_a(-0.12680411338806152)),(to_sfixed_a(-0.0003104248607996851)),(to_sfixed_a(-0.00015271673328243196)),(to_sfixed_a(0.0012326512951403856)),(to_sfixed_a(-0.005170414224267006)),(to_sfixed_a(-0.00029017377528361976)),(to_sfixed_a(-0.0032788049429655075)),(to_sfixed_a(0.5281566977500916)),(to_sfixed_a(-0.004694740753620863)),(to_sfixed_a(4.1464343667030334e-05)),(to_sfixed_a(-0.00013498785847332329)),(to_sfixed_a(-0.30601590871810913)),(to_sfixed_a(7.060663483571261e-05)),(to_sfixed_a(0.004083588719367981)),(to_sfixed_a(-6.777218368370086e-05)),(to_sfixed_a(-6.455121911130846e-05)),(to_sfixed_a(-4.888014154857956e-05)),(to_sfixed_a(0.0002473712956998497)),(to_sfixed_a(-3.18631500704214e-05)),(to_sfixed_a(-2.5901972549036145e-06)),(to_sfixed_a(0.00011242431355640292)),(to_sfixed_a(-0.0038438246119767427)),(to_sfixed_a(0.002369153080508113)),(to_sfixed_a(2.722893259488046e-05)),(to_sfixed_a(0.3021315634250641)),(to_sfixed_a(0.49319061636924744)),(to_sfixed_a(0.23334309458732605)),(to_sfixed_a(2.0312512788223103e-05)),(to_sfixed_a(2.2797494239057414e-05)),(to_sfixed_a(0.00010440080222906545)),(to_sfixed_a(-0.2872636616230011)),(to_sfixed_a(-0.08861187100410461)),(to_sfixed_a(6.732669135089964e-05)),(to_sfixed_a(0.5351644158363342)),(to_sfixed_a(2.819635847117752e-05)),(to_sfixed_a(-0.00011600545258261263)),(to_sfixed_a(-0.0025145120453089476)),(to_sfixed_a(-4.865113442065194e-05)),(to_sfixed_a(-0.0008490444160997868)),(to_sfixed_a(-3.3859469112940133e-06)),(to_sfixed_a(-0.0007093906169757247)),(to_sfixed_a(3.312921762699261e-05)),(to_sfixed_a(4.126130079384893e-05)),(to_sfixed_a(0.003012523055076599)),(to_sfixed_a(-8.531208004569635e-05)),(to_sfixed_a(4.617997183231637e-05)),(to_sfixed_a(0.1908567249774933)),(to_sfixed_a(-0.0027060036081820726)),(to_sfixed_a(6.766633305232972e-06)),(to_sfixed_a(0.0002001341781578958)),(to_sfixed_a(-8.022889232961461e-05)),(to_sfixed_a(0.0001488567650085315)),(to_sfixed_a(-0.0002003966219490394)),(to_sfixed_a(-0.002104430925101042)),(to_sfixed_a(0.0012573940912261605)),(to_sfixed_a(6.885106267873198e-05)),(to_sfixed_a(-6.429337372537702e-05)),(to_sfixed_a(-0.39885473251342773)),(to_sfixed_a(8.308676478918642e-05)),(to_sfixed_a(-1.765526394592598e-05)),(to_sfixed_a(-2.739726915024221e-05)),(to_sfixed_a(0.00046110511175356805)),(to_sfixed_a(3.8667090848321095e-05)),(to_sfixed_a(-0.00010732758528320119)),(to_sfixed_a(2.26006013690494e-05)),(to_sfixed_a(-0.0014806927647441626)),(to_sfixed_a(0.00015039366553537548)),(to_sfixed_a(0.005373399239033461)),(to_sfixed_a(-8.534688095096499e-05)),(to_sfixed_a(-5.047990271123126e-05)),(to_sfixed_a(-0.019006283953785896)),(to_sfixed_a(-1.4227851352188736e-05)),(to_sfixed_a(-1.054842141456902e-05)),(to_sfixed_a(0.003247960237786174)),(to_sfixed_a(-0.0001502867671661079)),(to_sfixed_a(-2.111131470883265e-05)),(to_sfixed_a(0.16932877898216248)),(to_sfixed_a(6.0461537941591814e-05)),(to_sfixed_a(-0.09596819430589676)),(to_sfixed_a(-4.7726651246193796e-05)),(to_sfixed_a(8.59333376865834e-05)),(to_sfixed_a(0.0001177708909381181)),(to_sfixed_a(0.00012946274364367127)),(to_sfixed_a(-0.003421621862798929)),(to_sfixed_a(-0.003197701647877693)),(to_sfixed_a(-0.0031083463691174984)),(to_sfixed_a(-0.005525683984160423)),(to_sfixed_a(0.00031087332172319293)),(to_sfixed_a(0.0045440769754350185)),(to_sfixed_a(0.0002517051761969924)),(to_sfixed_a(0.00020049842714797705)),(to_sfixed_a(-4.487654223339632e-06)),(to_sfixed_a(-0.0034969209227710962)),(to_sfixed_a(-0.005167532246559858)),(to_sfixed_a(0.0001661153946770355)),(to_sfixed_a(0.22361266613006592)),(to_sfixed_a(1.5296080164262094e-05)),(to_sfixed_a(0.3602827787399292)),(to_sfixed_a(0.24967502057552338)),(to_sfixed_a(0.14670901000499725)),(to_sfixed_a(0.24731217324733734)),(to_sfixed_a(0.0007243914296850562)),(to_sfixed_a(-0.00607592286542058)),(to_sfixed_a(0.00014611355436500162)),(to_sfixed_a(-8.2269252743572e-07)),(to_sfixed_a(-5.6360346206929535e-05)),(to_sfixed_a(-0.010582820512354374)),(to_sfixed_a(0.2215399593114853)),(to_sfixed_a(-0.0023015004117041826)),(to_sfixed_a(-0.0009053109097294509)),(to_sfixed_a(-0.00038155922084115446)),(to_sfixed_a(0.22229209542274475)),(to_sfixed_a(-0.00011576047108974308)),(to_sfixed_a(0.1553504914045334)),(to_sfixed_a(0.00014091083721723408)),(to_sfixed_a(-0.00023765102378092706)),(to_sfixed_a(-0.0016605829587206244)),(to_sfixed_a(-0.0001754346303641796)),(to_sfixed_a(-0.003871200606226921)),(to_sfixed_a(-0.30983057618141174)),(to_sfixed_a(-0.00016604826669208705)),(to_sfixed_a(-7.004426151979715e-06)),(to_sfixed_a(0.00012128661182941869)),(to_sfixed_a(0.00023486978898290545)),(to_sfixed_a(7.28682498447597e-05)),(to_sfixed_a(-3.330798426759429e-05)),(to_sfixed_a(0.0005854961345903575)),(to_sfixed_a(-0.041877277195453644)),(to_sfixed_a(-0.18622194230556488)),(to_sfixed_a(-0.003763271728530526)),(to_sfixed_a(0.0009301866521127522)),(to_sfixed_a(-0.009849360212683678)),(to_sfixed_a(-3.826537431450561e-05)),(to_sfixed_a(-0.00014928744349163026)),(to_sfixed_a(-6.0057333030272275e-05)),(to_sfixed_a(0.0001688510092208162)),(to_sfixed_a(0.00013708783080801368)),(to_sfixed_a(0.356082022190094)),(to_sfixed_a(-0.011961116455495358)),(to_sfixed_a(-0.4176783859729767)),(to_sfixed_a(-7.705901225563139e-05)),(to_sfixed_a(-1.0897445463342592e-05)),(to_sfixed_a(-5.6441815104335546e-05)),(to_sfixed_a(0.00010531915177125484)),(to_sfixed_a(2.0574170775944367e-06)),(to_sfixed_a(-0.002456313231959939)),(to_sfixed_a(0.0001487236440880224)),(to_sfixed_a(-5.6911343563115224e-05)),(to_sfixed_a(-4.204659489914775e-06)),(to_sfixed_a(-0.44794580340385437)),(to_sfixed_a(0.0029744994826614857)),(to_sfixed_a(-0.0009757229709066451)),(to_sfixed_a(6.097127334214747e-05)),(to_sfixed_a(-0.00020289275562390685)),(to_sfixed_a(-0.00010570352606009692)),(to_sfixed_a(0.0008094999939203262)),(to_sfixed_a(-0.00033027405152097344)),(to_sfixed_a(-0.5985009670257568)),(to_sfixed_a(0.00010533338354434818)),(to_sfixed_a(0.0006901281303726137)),(to_sfixed_a(0.00025149507564492524)),(to_sfixed_a(-0.005080115515738726)),(to_sfixed_a(-6.2935272580944e-05)),(to_sfixed_a(0.00016787310596555471)),(to_sfixed_a(0.0001591659674886614)),(to_sfixed_a(0.008073226548731327)),(to_sfixed_a(0.10694356262683868)),(to_sfixed_a(0.11814667284488678)),(to_sfixed_a(0.009076029062271118)),(to_sfixed_a(-0.00011391986481612548)),(to_sfixed_a(0.0029465053230524063)),(to_sfixed_a(-0.01101604476571083)),(to_sfixed_a(4.416827141540125e-05)),(to_sfixed_a(-0.008494320325553417)),(to_sfixed_a(-2.8892827685922384e-06)),(to_sfixed_a(-7.408375677186996e-05)),(to_sfixed_a(0.0187753364443779)),(to_sfixed_a(-0.006485030986368656)),(to_sfixed_a(0.00010765536717372015)),(to_sfixed_a(-0.0002648166846483946)),(to_sfixed_a(0.18859393894672394)),(to_sfixed_a(-1.5780344256199896e-05)),(to_sfixed_a(-0.005955163389444351)),(to_sfixed_a(-2.1196794477873482e-05)),(to_sfixed_a(0.0006888827192597091)),(to_sfixed_a(7.418263703584671e-05)),(to_sfixed_a(0.0007475214079022408)),(to_sfixed_a(-6.562830822076648e-05)),(to_sfixed_a(-6.385189772117883e-05)),(to_sfixed_a(2.1845666196895763e-05)),(to_sfixed_a(-0.22379259765148163)),(to_sfixed_a(0.0008055715006776154)),(to_sfixed_a(0.00018321456445846707)),(to_sfixed_a(-2.310157287865877e-05)),(to_sfixed_a(-0.00010092418233398348)),(to_sfixed_a(-1.5107194485608488e-05)),(to_sfixed_a(0.0031468523666262627)),(to_sfixed_a(0.001390855060890317)),(to_sfixed_a(0.3115714490413666)),(to_sfixed_a(-0.01083382498472929)),(to_sfixed_a(-0.014330223202705383)),(to_sfixed_a(-0.00013042772479820997)),(to_sfixed_a(1.15161674330011e-06)),(to_sfixed_a(-0.00028215927886776626)),(to_sfixed_a(-0.012812197208404541)),(to_sfixed_a(-0.0001564912381581962)),(to_sfixed_a(4.33262248407118e-05)),(to_sfixed_a(-0.008586960844695568)),(to_sfixed_a(0.0021978027652949095)),(to_sfixed_a(-0.0002124207967426628)),(to_sfixed_a(-0.1914312094449997)),(to_sfixed_a(0.0006676054326817393)),(to_sfixed_a(-0.010078205727040768)),(to_sfixed_a(0.003076596651226282)),(to_sfixed_a(6.931733514647931e-05)),(to_sfixed_a(-0.4405635893344879)),(to_sfixed_a(0.1328321397304535)),(to_sfixed_a(-0.002711439970880747)),(to_sfixed_a(0.00015125209756661206)),(to_sfixed_a(-0.014948826283216476)),(to_sfixed_a(0.29550522565841675)),(to_sfixed_a(-0.00835621077567339)));

    constant weight_n2_87 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.01753714680671692)),(to_sfixed_a(-0.0012832428328692913)),(to_sfixed_a(-0.7501499056816101)),(to_sfixed_a(1.5421537682414055e-06)),(to_sfixed_a(0.029989521950483322)),(to_sfixed_a(-0.00010525662946747616)),(to_sfixed_a(0.007882112637162209)),(to_sfixed_a(-0.00018521584570407867)),(to_sfixed_a(-0.00015353562775999308)),(to_sfixed_a(-7.147730502765626e-05)),(to_sfixed_a(0.00012740306556224823)),(to_sfixed_a(-0.0003874344693031162)),(to_sfixed_a(0.004596616141498089)),(to_sfixed_a(0.000107753679913003)),(to_sfixed_a(-0.00017486032447777689)),(to_sfixed_a(2.5878209271468222e-05)),(to_sfixed_a(0.47966113686561584)),(to_sfixed_a(-7.01696117175743e-05)),(to_sfixed_a(0.005054330453276634)),(to_sfixed_a(-0.005011211149394512)),(to_sfixed_a(-4.0679515223018825e-05)),(to_sfixed_a(1.8591985281091183e-05)),(to_sfixed_a(-0.00035154441138729453)),(to_sfixed_a(0.22398662567138672)),(to_sfixed_a(0.26491793990135193)),(to_sfixed_a(0.3352900743484497)),(to_sfixed_a(0.00010531261068535969)),(to_sfixed_a(-0.0006471279775723815)),(to_sfixed_a(0.010721644386649132)),(to_sfixed_a(-0.00021941243903711438)),(to_sfixed_a(0.37369391322135925)),(to_sfixed_a(-0.00022290171182248741)),(to_sfixed_a(0.16014093160629272)),(to_sfixed_a(-0.0001061700313584879)),(to_sfixed_a(1.9014521967619658e-05)),(to_sfixed_a(-0.00011591435031732544)),(to_sfixed_a(-0.3296383023262024)),(to_sfixed_a(0.074651800096035)),(to_sfixed_a(-0.5687326788902283)),(to_sfixed_a(0.00011382691445760429)),(to_sfixed_a(0.002506458666175604)),(to_sfixed_a(0.4263412654399872)),(to_sfixed_a(0.0002367268898524344)),(to_sfixed_a(-7.672212814213708e-05)),(to_sfixed_a(-0.0007140500238165259)),(to_sfixed_a(0.008089297451078892)),(to_sfixed_a(-0.014340457506477833)),(to_sfixed_a(0.009007963351905346)),(to_sfixed_a(-0.00010891981946770102)),(to_sfixed_a(0.013414119370281696)),(to_sfixed_a(0.4321165680885315)),(to_sfixed_a(-0.0006160663906484842)),(to_sfixed_a(-9.395483357366174e-05)),(to_sfixed_a(0.009186475537717342)),(to_sfixed_a(0.5679412484169006)),(to_sfixed_a(-0.22375960648059845)),(to_sfixed_a(-0.0001372484111925587)),(to_sfixed_a(0.006189220119267702)),(to_sfixed_a(6.292982288869098e-05)),(to_sfixed_a(-0.0002917373785749078)),(to_sfixed_a(-0.40566927194595337)),(to_sfixed_a(-0.003806505585089326)),(to_sfixed_a(-0.0002850376768037677)),(to_sfixed_a(-0.732067346572876)),(to_sfixed_a(-1.497105768066831e-05)),(to_sfixed_a(0.005424953065812588)),(to_sfixed_a(6.330995529424399e-05)),(to_sfixed_a(-0.012947160750627518)),(to_sfixed_a(0.012983664870262146)),(to_sfixed_a(0.00030179371242411435)),(to_sfixed_a(0.00879282783716917)),(to_sfixed_a(-0.0020473101176321507)),(to_sfixed_a(-0.00014669039228465408)),(to_sfixed_a(-0.00016912934370338917)),(to_sfixed_a(-0.00011067282321164384)),(to_sfixed_a(-6.052324897609651e-05)),(to_sfixed_a(0.006140605080872774)),(to_sfixed_a(0.008210200816392899)),(to_sfixed_a(7.047133840387687e-05)),(to_sfixed_a(-0.22631341218948364)),(to_sfixed_a(0.19107097387313843)),(to_sfixed_a(-6.525207572849467e-05)),(to_sfixed_a(0.318024218082428)),(to_sfixed_a(-0.3101484179496765)),(to_sfixed_a(-0.00032560178078711033)),(to_sfixed_a(0.2662920355796814)),(to_sfixed_a(-0.01252036727964878)),(to_sfixed_a(-0.005903180222958326)),(to_sfixed_a(-0.00012926390627399087)),(to_sfixed_a(0.00010814043343998492)),(to_sfixed_a(0.007285819388926029)),(to_sfixed_a(0.00014877138892188668)),(to_sfixed_a(0.4962631165981293)),(to_sfixed_a(-0.00015017094847280532)),(to_sfixed_a(0.016993243247270584)),(to_sfixed_a(8.333641017088667e-05)),(to_sfixed_a(-3.3366828574799e-05)),(to_sfixed_a(-2.8962414944544435e-05)),(to_sfixed_a(0.00016725153545849025)),(to_sfixed_a(7.876619201852009e-05)),(to_sfixed_a(-0.005666394252330065)),(to_sfixed_a(-0.00893071573227644)),(to_sfixed_a(-0.00016871263505890965)),(to_sfixed_a(-0.0011843114625662565)),(to_sfixed_a(0.011880841106176376)),(to_sfixed_a(0.0019191469764336944)),(to_sfixed_a(-2.939136902568862e-05)),(to_sfixed_a(6.84870028635487e-05)),(to_sfixed_a(0.00044994044583290815)),(to_sfixed_a(0.1551140397787094)),(to_sfixed_a(0.2066473811864853)),(to_sfixed_a(7.719360291957855e-05)),(to_sfixed_a(0.003185032634064555)),(to_sfixed_a(-2.997832780238241e-06)),(to_sfixed_a(8.906310540623963e-06)),(to_sfixed_a(0.30112171173095703)),(to_sfixed_a(-0.005149537231773138)),(to_sfixed_a(0.004346257075667381)),(to_sfixed_a(-5.696347216144204e-07)),(to_sfixed_a(0.00976615957915783)),(to_sfixed_a(-0.0002910451148636639)),(to_sfixed_a(2.752611180767417e-06)),(to_sfixed_a(0.0011348231928423047)),(to_sfixed_a(-1.785527274478227e-06)),(to_sfixed_a(-7.064913370413706e-05)),(to_sfixed_a(-0.0008392833406105638)),(to_sfixed_a(-0.004202587530016899)),(to_sfixed_a(6.995850708335638e-05)),(to_sfixed_a(5.80226733291056e-05)),(to_sfixed_a(-0.0001512592425569892)),(to_sfixed_a(0.00025090796407312155)),(to_sfixed_a(2.402414429525379e-05)),(to_sfixed_a(0.3353610336780548)),(to_sfixed_a(0.0019753912929445505)),(to_sfixed_a(-5.901165422983468e-06)),(to_sfixed_a(-0.00013346948253456503)),(to_sfixed_a(-0.002433792920783162)),(to_sfixed_a(-0.005168397910892963)),(to_sfixed_a(-2.050111652351916e-05)),(to_sfixed_a(-5.618870636681095e-05)),(to_sfixed_a(0.1866876780986786)),(to_sfixed_a(-4.572776015265845e-05)),(to_sfixed_a(-1.800665631890297e-05)),(to_sfixed_a(-1.609556784387678e-05)),(to_sfixed_a(-0.0009965873323380947)),(to_sfixed_a(0.0024815865326672792)),(to_sfixed_a(0.0015856061363592744)),(to_sfixed_a(0.00023620029969606549)),(to_sfixed_a(-4.76235436508432e-06)),(to_sfixed_a(0.0077798496931791306)),(to_sfixed_a(2.6222427550237626e-05)),(to_sfixed_a(-0.00011532891949173063)),(to_sfixed_a(0.0028246615547686815)),(to_sfixed_a(6.641687650699168e-05)),(to_sfixed_a(-2.055656659649685e-05)),(to_sfixed_a(-0.015043457970023155)),(to_sfixed_a(-0.0004194344219285995)),(to_sfixed_a(-0.011896326206624508)),(to_sfixed_a(0.00017735891742631793)),(to_sfixed_a(0.0002956193930003792)),(to_sfixed_a(-0.00010762463352875784)),(to_sfixed_a(-7.143958646338433e-05)),(to_sfixed_a(-0.004249056801199913)),(to_sfixed_a(0.3512935936450958)),(to_sfixed_a(0.2665795385837555)),(to_sfixed_a(-0.002051963470876217)),(to_sfixed_a(-2.8055677830707282e-05)),(to_sfixed_a(0.009019848890602589)),(to_sfixed_a(-2.3957174562383443e-05)),(to_sfixed_a(0.0002047852030955255)),(to_sfixed_a(0.09284961968660355)),(to_sfixed_a(0.00408389326184988)),(to_sfixed_a(-0.00046167781692929566)),(to_sfixed_a(5.696013249689713e-05)),(to_sfixed_a(0.00397430220618844)),(to_sfixed_a(0.0009007608168758452)),(to_sfixed_a(0.000855850987136364)),(to_sfixed_a(0.42158088088035583)),(to_sfixed_a(-0.26375481486320496)),(to_sfixed_a(0.2417529970407486)),(to_sfixed_a(0.00012876561959274113)),(to_sfixed_a(0.11412075906991959)),(to_sfixed_a(-0.00015136436559259892)),(to_sfixed_a(-0.00012920124572701752)),(to_sfixed_a(-0.00016859867901075631)),(to_sfixed_a(5.2099152526352555e-05)),(to_sfixed_a(-0.014267523773014545)),(to_sfixed_a(-0.0010312339290976524)),(to_sfixed_a(-0.003282288322225213)),(to_sfixed_a(0.000865457346662879)),(to_sfixed_a(-0.012021404691040516)),(to_sfixed_a(0.0003219749196432531)),(to_sfixed_a(-0.0040922751650214195)),(to_sfixed_a(0.015664519742131233)),(to_sfixed_a(-0.00020080602553207427)),(to_sfixed_a(0.6632804870605469)),(to_sfixed_a(-0.00010459705663379282)),(to_sfixed_a(-0.1913774013519287)),(to_sfixed_a(-0.012234359979629517)),(to_sfixed_a(-0.00018326427380088717)),(to_sfixed_a(-0.00020935977227054536)),(to_sfixed_a(3.0099756259005517e-05)),(to_sfixed_a(-0.0002719883341342211)),(to_sfixed_a(0.00018270855071023107)),(to_sfixed_a(1.216716191265732e-05)),(to_sfixed_a(-0.4269294738769531)),(to_sfixed_a(-0.0027574163395911455)),(to_sfixed_a(-0.41145995259284973)),(to_sfixed_a(0.002529232297092676)),(to_sfixed_a(-0.010821971110999584)),(to_sfixed_a(0.0038408380933105946)),(to_sfixed_a(7.673715299461037e-05)),(to_sfixed_a(0.00015802605776116252)),(to_sfixed_a(-6.331547047011554e-05)),(to_sfixed_a(0.00014798268966842443)),(to_sfixed_a(0.000152208172949031)),(to_sfixed_a(-0.009906169958412647)),(to_sfixed_a(0.33670735359191895)),(to_sfixed_a(-0.16549311578273773)),(to_sfixed_a(-0.00044870999408885837)),(to_sfixed_a(-5.650779348798096e-05)),(to_sfixed_a(-0.00018920065485872328)),(to_sfixed_a(1.5724785043857992e-05)),(to_sfixed_a(-0.0033423008862882853)),(to_sfixed_a(-0.01307707093656063)),(to_sfixed_a(-7.775372068863362e-05)),(to_sfixed_a(6.566732190549374e-05)),(to_sfixed_a(0.0002818201610352844)),(to_sfixed_a(-0.3043663203716278)),(to_sfixed_a(0.3183799386024475)),(to_sfixed_a(-0.0014359726337715983)),(to_sfixed_a(0.0001557761279400438)),(to_sfixed_a(0.0001416662271367386)),(to_sfixed_a(-4.811038525076583e-05)),(to_sfixed_a(0.001654339488595724)),(to_sfixed_a(0.19150684773921967)),(to_sfixed_a(-0.8233330845832825)),(to_sfixed_a(-1.4585872122552246e-05)),(to_sfixed_a(-3.8619393308181316e-05)),(to_sfixed_a(-8.306717791128904e-05)),(to_sfixed_a(-0.0003891782835125923)),(to_sfixed_a(-0.00023534164938610047)),(to_sfixed_a(0.0008103119325824082)),(to_sfixed_a(0.000113646914542187)),(to_sfixed_a(0.0030877389945089817)),(to_sfixed_a(-0.00034867069916799664)),(to_sfixed_a(0.5388301014900208)),(to_sfixed_a(0.007314910180866718)),(to_sfixed_a(-0.0001283002202399075)),(to_sfixed_a(0.002113182097673416)),(to_sfixed_a(0.006853659637272358)),(to_sfixed_a(0.0001611491315998137)),(to_sfixed_a(-0.00030093046370893717)),(to_sfixed_a(-7.874550647102296e-05)),(to_sfixed_a(0.2781100869178772)),(to_sfixed_a(0.037833571434020996)),(to_sfixed_a(0.0015543026383966208)),(to_sfixed_a(-0.00011374612950021401)),(to_sfixed_a(0.00010008273966377601)),(to_sfixed_a(0.046021319925785065)),(to_sfixed_a(6.155176379252225e-05)),(to_sfixed_a(-0.3973304331302643)),(to_sfixed_a(-0.0002133504895027727)),(to_sfixed_a(2.271361881867051e-05)),(to_sfixed_a(-0.00015826980234123766)),(to_sfixed_a(0.26233816146850586)),(to_sfixed_a(0.0001660699344938621)),(to_sfixed_a(-4.636029916582629e-05)),(to_sfixed_a(0.00024169808602891862)),(to_sfixed_a(0.001674890168942511)),(to_sfixed_a(0.010481023229658604)),(to_sfixed_a(0.0001502543454989791)),(to_sfixed_a(0.0001077835913747549)),(to_sfixed_a(-3.697481588460505e-06)),(to_sfixed_a(0.00015262103988789022)),(to_sfixed_a(0.26129934191703796)),(to_sfixed_a(-0.06848534941673279)),(to_sfixed_a(-0.008790245279669762)),(to_sfixed_a(0.000562569999601692)),(to_sfixed_a(0.001008416642434895)),(to_sfixed_a(0.00010404165368527174)),(to_sfixed_a(5.916517693549395e-06)),(to_sfixed_a(8.508504834026098e-08)),(to_sfixed_a(-0.22405731678009033)),(to_sfixed_a(3.8612641219515353e-05)),(to_sfixed_a(-8.478462405037135e-05)),(to_sfixed_a(-0.0030152862891554832)),(to_sfixed_a(0.0009600563207641244)),(to_sfixed_a(6.376780947903171e-05)),(to_sfixed_a(-0.00013555525219999254)),(to_sfixed_a(0.001853102003224194)),(to_sfixed_a(0.004711076617240906)),(to_sfixed_a(0.02260754443705082)),(to_sfixed_a(-0.0004096135962754488)),(to_sfixed_a(0.0037289063911885023)),(to_sfixed_a(0.005421699956059456)),(to_sfixed_a(0.000504323048517108)),(to_sfixed_a(0.0002876564103644341)),(to_sfixed_a(0.01927538961172104)),(to_sfixed_a(0.03840918093919754)),(to_sfixed_a(-0.07488614320755005)));

    constant weight_n2_88 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.06874671578407288)),(to_sfixed_a(0.0023667821660637856)),(to_sfixed_a(0.010207115672528744)),(to_sfixed_a(5.434839113149792e-05)),(to_sfixed_a(0.001161954365670681)),(to_sfixed_a(2.1570267563220114e-05)),(to_sfixed_a(0.002661663107573986)),(to_sfixed_a(0.00022324235760606825)),(to_sfixed_a(6.305419083219022e-05)),(to_sfixed_a(3.841618308797479e-05)),(to_sfixed_a(0.00014227414794731885)),(to_sfixed_a(-0.001491026720032096)),(to_sfixed_a(0.0005987173644825816)),(to_sfixed_a(0.10328804701566696)),(to_sfixed_a(9.2007961939089e-05)),(to_sfixed_a(-7.435706356773153e-05)),(to_sfixed_a(0.12324347347021103)),(to_sfixed_a(-0.00011671868560370058)),(to_sfixed_a(-0.005176735110580921)),(to_sfixed_a(-0.00017715948342811316)),(to_sfixed_a(-2.657072400324978e-05)),(to_sfixed_a(-1.4151723007671535e-05)),(to_sfixed_a(0.0003817327378783375)),(to_sfixed_a(0.38417747616767883)),(to_sfixed_a(0.000739111565053463)),(to_sfixed_a(0.0003653027815744281)),(to_sfixed_a(0.00020548269094433635)),(to_sfixed_a(-0.001841501914896071)),(to_sfixed_a(-5.4683401685906574e-05)),(to_sfixed_a(2.807231794577092e-06)),(to_sfixed_a(0.27219918370246887)),(to_sfixed_a(-5.0635273510124534e-05)),(to_sfixed_a(-0.014014321379363537)),(to_sfixed_a(-1.2255506590008736e-05)),(to_sfixed_a(-6.812772335251793e-05)),(to_sfixed_a(-0.0001600346149643883)),(to_sfixed_a(-0.45545724034309387)),(to_sfixed_a(-0.003440272528678179)),(to_sfixed_a(-0.0011740770423784852)),(to_sfixed_a(2.2721309505868703e-05)),(to_sfixed_a(-0.004180495627224445)),(to_sfixed_a(-0.0005116150714457035)),(to_sfixed_a(-0.0002030900795944035)),(to_sfixed_a(0.0001496560435043648)),(to_sfixed_a(0.2840852737426758)),(to_sfixed_a(-0.3546810448169708)),(to_sfixed_a(0.0005019746022298932)),(to_sfixed_a(-0.001986322458833456)),(to_sfixed_a(-0.00019103797967545688)),(to_sfixed_a(0.005542617756873369)),(to_sfixed_a(-0.006413597147911787)),(to_sfixed_a(-5.351072468329221e-05)),(to_sfixed_a(-0.0001052070947480388)),(to_sfixed_a(0.0004470670537557453)),(to_sfixed_a(0.003116349456831813)),(to_sfixed_a(-0.0012291353195905685)),(to_sfixed_a(9.407027391716838e-05)),(to_sfixed_a(0.0006877438863739371)),(to_sfixed_a(-7.118238863768056e-05)),(to_sfixed_a(6.254890467971563e-05)),(to_sfixed_a(0.2873077392578125)),(to_sfixed_a(0.0034218074288219213)),(to_sfixed_a(-0.0015301632229238749)),(to_sfixed_a(0.021924396976828575)),(to_sfixed_a(0.00017672441026661545)),(to_sfixed_a(0.20856021344661713)),(to_sfixed_a(-6.308353476924822e-05)),(to_sfixed_a(3.831181675195694e-05)),(to_sfixed_a(-7.981750241015106e-05)),(to_sfixed_a(-0.00010572317114565521)),(to_sfixed_a(-0.6670372486114502)),(to_sfixed_a(0.010899013839662075)),(to_sfixed_a(-0.38386937975883484)),(to_sfixed_a(-1.2148244422860444e-05)),(to_sfixed_a(-9.207240509567782e-05)),(to_sfixed_a(-6.604853842873126e-05)),(to_sfixed_a(0.31502875685691833)),(to_sfixed_a(0.000762264768127352)),(to_sfixed_a(-0.0002162560704164207)),(to_sfixed_a(-0.005319197662174702)),(to_sfixed_a(-6.887239578645676e-05)),(to_sfixed_a(-5.9321126173017547e-05)),(to_sfixed_a(0.0034781177528202534)),(to_sfixed_a(0.0006336129736155272)),(to_sfixed_a(-8.599908323958516e-05)),(to_sfixed_a(-0.002772229490801692)),(to_sfixed_a(-0.0002198671572841704)),(to_sfixed_a(-0.0012046379270032048)),(to_sfixed_a(4.644470027415082e-05)),(to_sfixed_a(-0.0001063846139004454)),(to_sfixed_a(0.4534641206264496)),(to_sfixed_a(-5.813136522192508e-05)),(to_sfixed_a(-0.003317194525152445)),(to_sfixed_a(6.967864464968443e-05)),(to_sfixed_a(-0.17911295592784882)),(to_sfixed_a(-0.0004918669001199305)),(to_sfixed_a(0.00017564906738698483)),(to_sfixed_a(1.45881058415398e-05)),(to_sfixed_a(-0.00026200077263638377)),(to_sfixed_a(8.420963422395289e-05)),(to_sfixed_a(-0.0032944129779934883)),(to_sfixed_a(0.0012204485246911645)),(to_sfixed_a(0.00013945400132797658)),(to_sfixed_a(0.03174504637718201)),(to_sfixed_a(-0.30226343870162964)),(to_sfixed_a(0.0003833947121165693)),(to_sfixed_a(6.375747034326196e-06)),(to_sfixed_a(-1.6536054317839444e-05)),(to_sfixed_a(-0.00019756675465032458)),(to_sfixed_a(0.000853740784805268)),(to_sfixed_a(0.0017456869827583432)),(to_sfixed_a(-6.723586557200179e-05)),(to_sfixed_a(-0.0014756462769582868)),(to_sfixed_a(0.00024497322738170624)),(to_sfixed_a(-4.0845683543011546e-05)),(to_sfixed_a(0.0013728175545111299)),(to_sfixed_a(-0.0033916952088475227)),(to_sfixed_a(0.0013410806423053145)),(to_sfixed_a(-0.00010912006837315857)),(to_sfixed_a(0.00021597396698780358)),(to_sfixed_a(-1.28697429317981e-05)),(to_sfixed_a(1.08074200397823e-05)),(to_sfixed_a(-0.0039909943006932735)),(to_sfixed_a(-0.00012602424249053001)),(to_sfixed_a(1.6963400412350893e-05)),(to_sfixed_a(0.00828083511441946)),(to_sfixed_a(0.003506104927510023)),(to_sfixed_a(3.817973265540786e-05)),(to_sfixed_a(4.980087396688759e-06)),(to_sfixed_a(-0.00015665829414501786)),(to_sfixed_a(-0.00013312484952621162)),(to_sfixed_a(0.0001865322410594672)),(to_sfixed_a(-0.002455526264384389)),(to_sfixed_a(-0.0003163152723573148)),(to_sfixed_a(-0.00015175265434663743)),(to_sfixed_a(-0.00021766213467344642)),(to_sfixed_a(0.367801696062088)),(to_sfixed_a(-0.0008188328938558698)),(to_sfixed_a(0.00017815129831433296)),(to_sfixed_a(-0.00019532660371623933)),(to_sfixed_a(-0.0011360221542418003)),(to_sfixed_a(-0.0001550941087771207)),(to_sfixed_a(0.00030654441798105836)),(to_sfixed_a(-5.03106857649982e-05)),(to_sfixed_a(0.00366249680519104)),(to_sfixed_a(0.00034584873355925083)),(to_sfixed_a(-0.00041949955630116165)),(to_sfixed_a(0.00018854642985388637)),(to_sfixed_a(-0.00014710769755765796)),(to_sfixed_a(-0.26613226532936096)),(to_sfixed_a(5.714097642339766e-05)),(to_sfixed_a(-0.000148551887832582)),(to_sfixed_a(0.00020898334332741797)),(to_sfixed_a(-0.0001468511763960123)),(to_sfixed_a(1.2885197065770626e-05)),(to_sfixed_a(0.010496732778847218)),(to_sfixed_a(-0.00015913156676106155)),(to_sfixed_a(0.002553253434598446)),(to_sfixed_a(-2.7960952138528228e-05)),(to_sfixed_a(0.00011201715824427083)),(to_sfixed_a(-0.00013080784992780536)),(to_sfixed_a(-6.916516576893628e-05)),(to_sfixed_a(-0.010664509609341621)),(to_sfixed_a(-0.00013517867773771286)),(to_sfixed_a(0.0006120299221947789)),(to_sfixed_a(-0.001976326573640108)),(to_sfixed_a(6.044624751666561e-05)),(to_sfixed_a(0.47101715207099915)),(to_sfixed_a(0.00017705745995044708)),(to_sfixed_a(-0.0001339234586339444)),(to_sfixed_a(0.0013639600947499275)),(to_sfixed_a(-0.0019070282578468323)),(to_sfixed_a(-4.605405410984531e-05)),(to_sfixed_a(-9.074864647118375e-05)),(to_sfixed_a(0.38823992013931274)),(to_sfixed_a(-9.986090299207717e-05)),(to_sfixed_a(0.020560316741466522)),(to_sfixed_a(0.33976826071739197)),(to_sfixed_a(-0.38045841455459595)),(to_sfixed_a(-0.0022123348899185658)),(to_sfixed_a(0.002464839955791831)),(to_sfixed_a(-0.015376130118966103)),(to_sfixed_a(0.00011638842261163518)),(to_sfixed_a(-5.748899275204167e-05)),(to_sfixed_a(0.0002202607283834368)),(to_sfixed_a(0.0008340962813235819)),(to_sfixed_a(0.0009473867830820382)),(to_sfixed_a(0.0013300051214173436)),(to_sfixed_a(0.0017689550295472145)),(to_sfixed_a(-0.002350522205233574)),(to_sfixed_a(3.0419229005929083e-05)),(to_sfixed_a(-5.189332296140492e-05)),(to_sfixed_a(-0.010365571826696396)),(to_sfixed_a(-0.002490777987986803)),(to_sfixed_a(-0.0001023158329189755)),(to_sfixed_a(5.771344876848161e-05)),(to_sfixed_a(0.00016659838729538023)),(to_sfixed_a(0.006644584238529205)),(to_sfixed_a(-0.00048466463340446353)),(to_sfixed_a(-1.3061187928542495e-05)),(to_sfixed_a(0.00015050293586682528)),(to_sfixed_a(0.0002968179469462484)),(to_sfixed_a(-1.6333156963810325e-05)),(to_sfixed_a(-0.0001119722073781304)),(to_sfixed_a(7.888750405982137e-05)),(to_sfixed_a(0.00028761057183146477)),(to_sfixed_a(0.0030337271746248007)),(to_sfixed_a(-0.01744861528277397)),(to_sfixed_a(0.010786166414618492)),(to_sfixed_a(0.003054010681807995)),(to_sfixed_a(-0.0013919174671173096)),(to_sfixed_a(6.25776665401645e-05)),(to_sfixed_a(-5.203117325436324e-06)),(to_sfixed_a(7.843293133191764e-06)),(to_sfixed_a(0.00031152847805060446)),(to_sfixed_a(0.0002261216868646443)),(to_sfixed_a(0.004710203967988491)),(to_sfixed_a(-0.0008131489157676697)),(to_sfixed_a(7.766287308186293e-05)),(to_sfixed_a(0.00010473205475136638)),(to_sfixed_a(0.00019511037680786103)),(to_sfixed_a(0.00020471253083087504)),(to_sfixed_a(0.00028303242288529873)),(to_sfixed_a(-0.29607558250427246)),(to_sfixed_a(-0.5058561563491821)),(to_sfixed_a(-0.00012130709365010262)),(to_sfixed_a(0.00014962763816583902)),(to_sfixed_a(-0.0002048924216069281)),(to_sfixed_a(-0.0018084964249283075)),(to_sfixed_a(0.0024831430055201054)),(to_sfixed_a(0.0005332462606020272)),(to_sfixed_a(-0.00011677867587422952)),(to_sfixed_a(-0.00010347177158109844)),(to_sfixed_a(-0.0003001876175403595)),(to_sfixed_a(0.000529309269040823)),(to_sfixed_a(0.0005965708987787366)),(to_sfixed_a(-0.006945595610886812)),(to_sfixed_a(-3.646976620075293e-05)),(to_sfixed_a(0.00031974678859114647)),(to_sfixed_a(-0.00019305438036099076)),(to_sfixed_a(-0.0005010726163163781)),(to_sfixed_a(-1.4349119737744331e-05)),(to_sfixed_a(-0.3209931552410126)),(to_sfixed_a(-6.921924068592489e-05)),(to_sfixed_a(-0.006994632072746754)),(to_sfixed_a(0.005163851659744978)),(to_sfixed_a(0.001857612980529666)),(to_sfixed_a(-0.0008875248022377491)),(to_sfixed_a(-0.000288316048681736)),(to_sfixed_a(0.38633179664611816)),(to_sfixed_a(0.0037538723554462194)),(to_sfixed_a(-0.0002263545320602134)),(to_sfixed_a(-2.5982091756304726e-05)),(to_sfixed_a(0.00024754254263825715)),(to_sfixed_a(3.778421159950085e-06)),(to_sfixed_a(0.0006948006921447814)),(to_sfixed_a(0.002485650358721614)),(to_sfixed_a(2.4044988094829023e-05)),(to_sfixed_a(-0.0001817153679439798)),(to_sfixed_a(-0.0038774514105170965)),(to_sfixed_a(0.00015006632020231336)),(to_sfixed_a(-0.0006356019875966012)),(to_sfixed_a(0.00045219974708743393)),(to_sfixed_a(-0.0001131899916799739)),(to_sfixed_a(-0.00025018653832376003)),(to_sfixed_a(-0.002678793156519532)),(to_sfixed_a(0.0002168084029108286)),(to_sfixed_a(1.6847479855641723e-05)),(to_sfixed_a(-0.00010532320447964594)),(to_sfixed_a(-0.0030999905429780483)),(to_sfixed_a(-0.010191601701080799)),(to_sfixed_a(0.00010252639185637236)),(to_sfixed_a(-0.0002734071167651564)),(to_sfixed_a(3.767314774449915e-05)),(to_sfixed_a(0.0001430611009709537)),(to_sfixed_a(0.0063584730960428715)),(to_sfixed_a(0.0029515104833990335)),(to_sfixed_a(0.19538277387619019)),(to_sfixed_a(0.002105953171849251)),(to_sfixed_a(0.002259031403809786)),(to_sfixed_a(0.000302924367133528)),(to_sfixed_a(6.805760494899005e-05)),(to_sfixed_a(-0.000201792674488388)),(to_sfixed_a(9.982217306969687e-06)),(to_sfixed_a(-4.005269147455692e-06)),(to_sfixed_a(-0.0002934451913461089)),(to_sfixed_a(-0.00011068718595197424)),(to_sfixed_a(0.004459911026060581)),(to_sfixed_a(-3.847830885206349e-05)),(to_sfixed_a(-0.2920193374156952)),(to_sfixed_a(2.41694797296077e-05)),(to_sfixed_a(0.0009322134428657591)),(to_sfixed_a(0.0007849233807064593)),(to_sfixed_a(-0.0001682589208940044)),(to_sfixed_a(0.26023441553115845)),(to_sfixed_a(0.01278930064290762)),(to_sfixed_a(0.001848897198215127)),(to_sfixed_a(0.00019430328393355012)),(to_sfixed_a(-0.0027079631108790636)),(to_sfixed_a(0.0017573584336787462)),(to_sfixed_a(0.00208604009822011)));

    constant weight_n2_89 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.03612072765827179)),(to_sfixed_a(6.889701762702316e-05)),(to_sfixed_a(-1.6135716577991843e-05)),(to_sfixed_a(0.00012984435306861997)),(to_sfixed_a(-4.082497980562039e-05)),(to_sfixed_a(0.00025064341025426984)),(to_sfixed_a(-9.378733375342563e-05)),(to_sfixed_a(-0.000322874344419688)),(to_sfixed_a(0.00010305454634362832)),(to_sfixed_a(0.000152963912114501)),(to_sfixed_a(-0.00039206710061989725)),(to_sfixed_a(0.00016465241787955165)),(to_sfixed_a(0.0001503278035670519)),(to_sfixed_a(-7.461196946678683e-05)),(to_sfixed_a(-3.223067324142903e-06)),(to_sfixed_a(-0.0001830640685511753)),(to_sfixed_a(0.00012803549179807305)),(to_sfixed_a(-8.314545266330242e-05)),(to_sfixed_a(0.00011994503438472748)),(to_sfixed_a(-1.5946978237479925e-05)),(to_sfixed_a(0.00011679398448904976)),(to_sfixed_a(-0.00011943878052989021)),(to_sfixed_a(-0.00013478941400535405)),(to_sfixed_a(4.929395799990743e-06)),(to_sfixed_a(3.223475505365059e-05)),(to_sfixed_a(-0.0002285564405610785)),(to_sfixed_a(0.0002078352845273912)),(to_sfixed_a(0.00017247811774723232)),(to_sfixed_a(5.8290497690904886e-06)),(to_sfixed_a(6.815945380367339e-05)),(to_sfixed_a(-0.00028951140120625496)),(to_sfixed_a(-3.5579578252509236e-06)),(to_sfixed_a(0.00016649148892611265)),(to_sfixed_a(-6.973020936129615e-05)),(to_sfixed_a(0.00013852117990609258)),(to_sfixed_a(3.871155786328018e-05)),(to_sfixed_a(-5.732259160140529e-05)),(to_sfixed_a(-6.724696140736341e-05)),(to_sfixed_a(-0.00029640033608302474)),(to_sfixed_a(-6.99474330758676e-05)),(to_sfixed_a(-0.0002267306699650362)),(to_sfixed_a(0.0002903435961343348)),(to_sfixed_a(6.872996891615912e-05)),(to_sfixed_a(0.00012788439926225692)),(to_sfixed_a(1.4779361663386226e-06)),(to_sfixed_a(0.0001856861199485138)),(to_sfixed_a(-7.407955854432657e-05)),(to_sfixed_a(5.05511779920198e-05)),(to_sfixed_a(-5.534305455512367e-05)),(to_sfixed_a(2.4504544853698462e-05)),(to_sfixed_a(-0.0002967653563246131)),(to_sfixed_a(8.704485662747175e-05)),(to_sfixed_a(9.101094474317506e-05)),(to_sfixed_a(-6.764993304386735e-05)),(to_sfixed_a(-6.0311565903248265e-05)),(to_sfixed_a(6.155409209895879e-05)),(to_sfixed_a(0.00031138386111706495)),(to_sfixed_a(6.962531915633008e-05)),(to_sfixed_a(-0.00024783413391560316)),(to_sfixed_a(0.00015671282017137855)),(to_sfixed_a(-0.0004103864775970578)),(to_sfixed_a(-2.0990919438190758e-05)),(to_sfixed_a(0.00010536712943576276)),(to_sfixed_a(0.0002655585412867367)),(to_sfixed_a(7.326866762014106e-05)),(to_sfixed_a(1.330390659859404e-05)),(to_sfixed_a(3.026393096661195e-05)),(to_sfixed_a(3.1096351449377835e-06)),(to_sfixed_a(1.5598561731167138e-05)),(to_sfixed_a(-1.0077950719278306e-05)),(to_sfixed_a(-9.984387361328118e-06)),(to_sfixed_a(3.796254168264568e-05)),(to_sfixed_a(0.0002111482317559421)),(to_sfixed_a(-0.00023810485436115414)),(to_sfixed_a(1.7808270058594644e-07)),(to_sfixed_a(0.0001035256136674434)),(to_sfixed_a(0.00021910945361014456)),(to_sfixed_a(-7.415001164190471e-06)),(to_sfixed_a(-0.00024031901557464153)),(to_sfixed_a(0.00012159665493527427)),(to_sfixed_a(-0.00014996808022260666)),(to_sfixed_a(-1.4132259821053594e-05)),(to_sfixed_a(-0.00010546360863372684)),(to_sfixed_a(5.693329148925841e-05)),(to_sfixed_a(6.91372188157402e-05)),(to_sfixed_a(-0.0001522829697933048)),(to_sfixed_a(3.7680365494452417e-06)),(to_sfixed_a(0.0003196320903953165)),(to_sfixed_a(8.404436084674671e-05)),(to_sfixed_a(-0.00010531961015658453)),(to_sfixed_a(0.0002266780356876552)),(to_sfixed_a(-0.0001963756512850523)),(to_sfixed_a(-0.0001829505490604788)),(to_sfixed_a(0.00011565486784093082)),(to_sfixed_a(-2.4324384867213666e-05)),(to_sfixed_a(0.00029880882357247174)),(to_sfixed_a(0.00016725307796150446)),(to_sfixed_a(3.892874883604236e-05)),(to_sfixed_a(-0.00022153167810756713)),(to_sfixed_a(-0.000106118168332614)),(to_sfixed_a(-0.00024350198509637266)),(to_sfixed_a(-0.00023709087690804154)),(to_sfixed_a(-9.632878209231421e-05)),(to_sfixed_a(0.00037760817212983966)),(to_sfixed_a(4.3013333197450265e-05)),(to_sfixed_a(-9.891096851788461e-06)),(to_sfixed_a(5.8596095186658204e-05)),(to_sfixed_a(-7.43611017242074e-05)),(to_sfixed_a(4.673511648434214e-05)),(to_sfixed_a(0.00017509181634522974)),(to_sfixed_a(-0.00017089555331040174)),(to_sfixed_a(4.428432657732628e-05)),(to_sfixed_a(-0.00014657192514277995)),(to_sfixed_a(-0.00022215649369172752)),(to_sfixed_a(-0.00018737699429038912)),(to_sfixed_a(4.396223448566161e-05)),(to_sfixed_a(-0.00020855374168604612)),(to_sfixed_a(-3.776869925786741e-05)),(to_sfixed_a(6.611809658352286e-05)),(to_sfixed_a(-0.00011769535194616765)),(to_sfixed_a(-0.0002208515943493694)),(to_sfixed_a(0.0003071035898756236)),(to_sfixed_a(7.63856660341844e-05)),(to_sfixed_a(-0.00030822743428871036)),(to_sfixed_a(0.00010254255175823346)),(to_sfixed_a(-6.73414979246445e-06)),(to_sfixed_a(2.230617610621266e-06)),(to_sfixed_a(2.7746791602112353e-06)),(to_sfixed_a(7.257387915160507e-05)),(to_sfixed_a(-8.567585609853268e-07)),(to_sfixed_a(1.6860685718711466e-06)),(to_sfixed_a(6.572713027708232e-05)),(to_sfixed_a(8.497658564010635e-05)),(to_sfixed_a(-0.0001128126896219328)),(to_sfixed_a(-4.822197661269456e-05)),(to_sfixed_a(-0.0001289883366553113)),(to_sfixed_a(9.012120426632464e-05)),(to_sfixed_a(0.0001500649523222819)),(to_sfixed_a(-0.00018398815882392228)),(to_sfixed_a(8.250462997239083e-07)),(to_sfixed_a(-0.0002452070184517652)),(to_sfixed_a(0.00011748790711862966)),(to_sfixed_a(0.0003886207123287022)),(to_sfixed_a(-6.738062074873596e-05)),(to_sfixed_a(-7.037619798211381e-05)),(to_sfixed_a(0.00013702866272069514)),(to_sfixed_a(-0.0001176066798507236)),(to_sfixed_a(-1.9087536202277988e-05)),(to_sfixed_a(0.00015827383322175592)),(to_sfixed_a(-4.883653309661895e-05)),(to_sfixed_a(3.218881829525344e-05)),(to_sfixed_a(0.00017329634283669293)),(to_sfixed_a(0.00017535149527247995)),(to_sfixed_a(-7.00742966728285e-05)),(to_sfixed_a(-0.00016419001622125506)),(to_sfixed_a(6.145394581835717e-05)),(to_sfixed_a(4.588825686369091e-05)),(to_sfixed_a(-1.1108408216387033e-05)),(to_sfixed_a(6.844867311883718e-05)),(to_sfixed_a(-0.000272571574896574)),(to_sfixed_a(-0.00013500118802767247)),(to_sfixed_a(-0.00041629280894994736)),(to_sfixed_a(-0.00022565768449567258)),(to_sfixed_a(8.02217036834918e-05)),(to_sfixed_a(-9.10947856027633e-05)),(to_sfixed_a(0.00015523380716331303)),(to_sfixed_a(-0.00012858310947194695)),(to_sfixed_a(0.00010727354674600065)),(to_sfixed_a(-4.692616857937537e-05)),(to_sfixed_a(-5.768506525782868e-05)),(to_sfixed_a(-0.00012080872693331912)),(to_sfixed_a(-0.0002768073754850775)),(to_sfixed_a(-5.855961353518069e-05)),(to_sfixed_a(-2.0842890080530196e-07)),(to_sfixed_a(-6.275861233007163e-05)),(to_sfixed_a(0.0002963231527246535)),(to_sfixed_a(6.737536750733852e-06)),(to_sfixed_a(2.8731825295835733e-05)),(to_sfixed_a(7.002049096627161e-05)),(to_sfixed_a(2.667814987944439e-05)),(to_sfixed_a(-0.0002482210984453559)),(to_sfixed_a(2.3997039534151554e-05)),(to_sfixed_a(5.176199192646891e-05)),(to_sfixed_a(1.5227105905069038e-05)),(to_sfixed_a(-0.00024013451184146106)),(to_sfixed_a(1.7762213246896863e-05)),(to_sfixed_a(-4.8957903345581144e-05)),(to_sfixed_a(0.0001478803314967081)),(to_sfixed_a(-0.00018207557150162756)),(to_sfixed_a(6.294957711361349e-05)),(to_sfixed_a(-5.7935743825510144e-05)),(to_sfixed_a(-0.0001515306648798287)),(to_sfixed_a(-0.00023553062055725604)),(to_sfixed_a(2.3471875465475023e-05)),(to_sfixed_a(4.4764557969756424e-05)),(to_sfixed_a(-7.876966265030205e-05)),(to_sfixed_a(-1.672350481385365e-05)),(to_sfixed_a(1.5382771380245686e-05)),(to_sfixed_a(0.00021930961520411074)),(to_sfixed_a(-2.96569342026487e-05)),(to_sfixed_a(1.4053111954126507e-06)),(to_sfixed_a(0.00029424933018162847)),(to_sfixed_a(-7.298671698663384e-05)),(to_sfixed_a(1.0135408956557512e-06)),(to_sfixed_a(0.00015006955072749406)),(to_sfixed_a(-0.00011457000073278323)),(to_sfixed_a(3.753071359824389e-05)),(to_sfixed_a(3.099906462011859e-05)),(to_sfixed_a(-0.00010598258813843131)),(to_sfixed_a(-1.1491629265947267e-05)),(to_sfixed_a(0.0001334378612227738)),(to_sfixed_a(1.9297891412861645e-05)),(to_sfixed_a(-0.0001507624110672623)),(to_sfixed_a(-1.2216805771458894e-05)),(to_sfixed_a(0.00013018102617934346)),(to_sfixed_a(0.00013516141916625202)),(to_sfixed_a(-6.005787872709334e-05)),(to_sfixed_a(-0.0001064277530531399)),(to_sfixed_a(-0.00021392152120824903)),(to_sfixed_a(-0.00022611864551436156)),(to_sfixed_a(-0.0003013969399034977)),(to_sfixed_a(6.785481673432514e-06)),(to_sfixed_a(-1.5383033314719796e-05)),(to_sfixed_a(5.240253813099116e-06)),(to_sfixed_a(-5.261419573798776e-06)),(to_sfixed_a(-0.00011348578846082091)),(to_sfixed_a(0.00011737868044292554)),(to_sfixed_a(6.024881440680474e-05)),(to_sfixed_a(0.00030574382981285453)),(to_sfixed_a(-9.9582157417899e-06)),(to_sfixed_a(7.446940435329452e-05)),(to_sfixed_a(-0.0002869179006665945)),(to_sfixed_a(0.0002864756970666349)),(to_sfixed_a(6.946177745703608e-05)),(to_sfixed_a(-7.229782931972295e-05)),(to_sfixed_a(0.0002518881228752434)),(to_sfixed_a(-3.331076368340291e-05)),(to_sfixed_a(9.138270252151415e-05)),(to_sfixed_a(-5.777664773631841e-05)),(to_sfixed_a(0.0001388436503475532)),(to_sfixed_a(-7.010975241428241e-05)),(to_sfixed_a(-3.0535207770299166e-05)),(to_sfixed_a(-0.00011540757259353995)),(to_sfixed_a(-0.00011650552187347785)),(to_sfixed_a(0.00010588264558464289)),(to_sfixed_a(-0.00010490330896573141)),(to_sfixed_a(-1.7897880752570927e-05)),(to_sfixed_a(-2.9307091608643532e-05)),(to_sfixed_a(-0.00014955594087950885)),(to_sfixed_a(-0.00015700147196184844)),(to_sfixed_a(8.494868234265596e-05)),(to_sfixed_a(-6.497862341348082e-05)),(to_sfixed_a(4.7757450374774635e-05)),(to_sfixed_a(-4.3210187868680805e-05)),(to_sfixed_a(0.00016454467549920082)),(to_sfixed_a(-0.0002611349045764655)),(to_sfixed_a(5.782834705314599e-05)),(to_sfixed_a(0.00013075079186819494)),(to_sfixed_a(0.00015634894953109324)),(to_sfixed_a(-0.0001358662557322532)),(to_sfixed_a(-0.00016631597827654332)),(to_sfixed_a(6.544629286509007e-05)),(to_sfixed_a(-0.0002000277891056612)),(to_sfixed_a(5.0591730541782454e-05)),(to_sfixed_a(0.00017357405158691108)),(to_sfixed_a(-0.00011320693010929972)),(to_sfixed_a(-8.635938866063952e-05)),(to_sfixed_a(0.00013093264715280384)),(to_sfixed_a(-1.2432472431100905e-05)),(to_sfixed_a(-0.0001281589939026162)),(to_sfixed_a(-7.466891111107543e-05)),(to_sfixed_a(-1.902158692246303e-05)),(to_sfixed_a(6.887942436151206e-05)),(to_sfixed_a(0.00010186730651184916)),(to_sfixed_a(7.239389378810301e-05)),(to_sfixed_a(1.4798948541283607e-05)),(to_sfixed_a(0.0001709410862531513)),(to_sfixed_a(6.022339221090078e-06)),(to_sfixed_a(-0.000303450069623068)),(to_sfixed_a(0.00011696561705321074)),(to_sfixed_a(0.0001677248510532081)),(to_sfixed_a(-6.2697072280570865e-06)),(to_sfixed_a(-2.5584267859812826e-07)),(to_sfixed_a(0.0001681880239630118)),(to_sfixed_a(0.00018193310825154185)),(to_sfixed_a(-0.00042607064824551344)),(to_sfixed_a(5.954180596745573e-05)),(to_sfixed_a(0.00013672221393790096)),(to_sfixed_a(-6.952373223612085e-05)),(to_sfixed_a(0.00011207604984520003)),(to_sfixed_a(1.7904158085002564e-05)),(to_sfixed_a(-0.00014674250269308686)),(to_sfixed_a(3.534779534675181e-05)),(to_sfixed_a(-2.39826476899907e-07)),(to_sfixed_a(-1.127687210100703e-05)),(to_sfixed_a(2.6836307370103896e-05)),(to_sfixed_a(-6.824910087743774e-05)),(to_sfixed_a(-4.8599031288176775e-06)),(to_sfixed_a(2.0165316527709365e-07)),(to_sfixed_a(-0.00010296780965290964)),(to_sfixed_a(7.137241482269019e-05)));

    constant weight_n2_90 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.34999996423721313)),(to_sfixed_a(0.008995883166790009)),(to_sfixed_a(-0.0007983936229720712)),(to_sfixed_a(-6.952474359422922e-05)),(to_sfixed_a(0.007241773884743452)),(to_sfixed_a(-0.0001562577235745266)),(to_sfixed_a(0.347756564617157)),(to_sfixed_a(-0.0001466814283048734)),(to_sfixed_a(-2.679813769645989e-05)),(to_sfixed_a(-0.00016463131760247052)),(to_sfixed_a(0.0004474472953006625)),(to_sfixed_a(0.000831994169857353)),(to_sfixed_a(-0.3832781910896301)),(to_sfixed_a(-0.0022356275003403425)),(to_sfixed_a(-5.5782627896405756e-05)),(to_sfixed_a(-3.270343586336821e-05)),(to_sfixed_a(0.5102249979972839)),(to_sfixed_a(8.344269735971466e-05)),(to_sfixed_a(0.4725106358528137)),(to_sfixed_a(-0.04848243296146393)),(to_sfixed_a(-0.00027897642576135695)),(to_sfixed_a(-0.00014854760956950486)),(to_sfixed_a(-0.0022388685029000044)),(to_sfixed_a(-5.842333484906703e-05)),(to_sfixed_a(0.4245030879974365)),(to_sfixed_a(0.0032773197162896395)),(to_sfixed_a(1.2401887943269685e-05)),(to_sfixed_a(3.690143785206601e-05)),(to_sfixed_a(0.009018431417644024)),(to_sfixed_a(-0.00011321240162942559)),(to_sfixed_a(-0.0040106442756950855)),(to_sfixed_a(-9.264171967515722e-05)),(to_sfixed_a(0.00048151781084015965)),(to_sfixed_a(-3.001609366037883e-05)),(to_sfixed_a(-3.854118403978646e-05)),(to_sfixed_a(-0.0001896177273010835)),(to_sfixed_a(0.0026615001261234283)),(to_sfixed_a(0.0073342109099030495)),(to_sfixed_a(0.02336963079869747)),(to_sfixed_a(-0.00011624252510955557)),(to_sfixed_a(0.0050676846876740456)),(to_sfixed_a(-0.0008996768738143146)),(to_sfixed_a(-6.751857290510088e-05)),(to_sfixed_a(-0.00023314358259085566)),(to_sfixed_a(-0.005732954945415258)),(to_sfixed_a(-0.0009815531084313989)),(to_sfixed_a(0.008060017600655556)),(to_sfixed_a(0.004024626687169075)),(to_sfixed_a(0.00017505305004306138)),(to_sfixed_a(-0.2747490406036377)),(to_sfixed_a(-0.00035291409585624933)),(to_sfixed_a(-0.0002005214337259531)),(to_sfixed_a(2.4146531359292567e-05)),(to_sfixed_a(0.01142912358045578)),(to_sfixed_a(-0.003622286021709442)),(to_sfixed_a(-0.10630075633525848)),(to_sfixed_a(2.406923158559948e-06)),(to_sfixed_a(-0.0003250125446356833)),(to_sfixed_a(-0.00024671980645507574)),(to_sfixed_a(0.00011719533358700573)),(to_sfixed_a(-0.0028784458991140127)),(to_sfixed_a(-0.004924634471535683)),(to_sfixed_a(-0.29878753423690796)),(to_sfixed_a(0.04484409838914871)),(to_sfixed_a(2.9341827030293643e-06)),(to_sfixed_a(-0.001161443768069148)),(to_sfixed_a(-7.163757982198149e-05)),(to_sfixed_a(0.001811790163628757)),(to_sfixed_a(0.002954090479761362)),(to_sfixed_a(0.0003036519919987768)),(to_sfixed_a(0.25502994656562805)),(to_sfixed_a(-0.009575916454195976)),(to_sfixed_a(-0.00019212599727325141)),(to_sfixed_a(0.00011757558968383819)),(to_sfixed_a(-2.7469686756376177e-06)),(to_sfixed_a(-0.00022547133266925812)),(to_sfixed_a(-0.015227880328893661)),(to_sfixed_a(0.003363613272085786)),(to_sfixed_a(-6.977158773224801e-05)),(to_sfixed_a(0.005782911088317633)),(to_sfixed_a(-0.0032299570739269257)),(to_sfixed_a(-8.671850082464516e-07)),(to_sfixed_a(-0.0011191965313628316)),(to_sfixed_a(0.0025391618255525827)),(to_sfixed_a(3.109486715402454e-05)),(to_sfixed_a(0.25821903347969055)),(to_sfixed_a(0.40151190757751465)),(to_sfixed_a(0.1607377827167511)),(to_sfixed_a(1.1810101568698883e-05)),(to_sfixed_a(-0.00024726902483962476)),(to_sfixed_a(-0.00126751943025738)),(to_sfixed_a(-4.8330875870306045e-06)),(to_sfixed_a(-0.003241753438487649)),(to_sfixed_a(-6.664905959041789e-05)),(to_sfixed_a(0.002699659438803792)),(to_sfixed_a(0.00014365582319442183)),(to_sfixed_a(-6.497011781902984e-05)),(to_sfixed_a(-0.00011266475485172123)),(to_sfixed_a(1.0006260708905756e-07)),(to_sfixed_a(5.8844721934292465e-05)),(to_sfixed_a(-0.0005880914977751672)),(to_sfixed_a(-0.000991301261819899)),(to_sfixed_a(6.971174298087135e-05)),(to_sfixed_a(-0.3924270570278168)),(to_sfixed_a(0.03534400835633278)),(to_sfixed_a(5.156177212484181e-05)),(to_sfixed_a(0.00013542422675527632)),(to_sfixed_a(-7.960552466101944e-05)),(to_sfixed_a(-0.00019185716519132257)),(to_sfixed_a(0.27098748087882996)),(to_sfixed_a(-0.009968003258109093)),(to_sfixed_a(4.877911123912781e-07)),(to_sfixed_a(0.34119197726249695)),(to_sfixed_a(-0.00026553956558927894)),(to_sfixed_a(-1.0961011867038906e-06)),(to_sfixed_a(0.006403392180800438)),(to_sfixed_a(0.000549978984054178)),(to_sfixed_a(-0.0001452674769097939)),(to_sfixed_a(6.197825132403523e-05)),(to_sfixed_a(0.007433594204485416)),(to_sfixed_a(0.0003019087598659098)),(to_sfixed_a(-6.000122084515169e-05)),(to_sfixed_a(0.0031006301287561655)),(to_sfixed_a(0.00015610389527864754)),(to_sfixed_a(-0.000166448880918324)),(to_sfixed_a(-0.0010306155309081078)),(to_sfixed_a(0.00386973493732512)),(to_sfixed_a(7.066567923175171e-05)),(to_sfixed_a(0.00013806969218421727)),(to_sfixed_a(2.6046291168313473e-06)),(to_sfixed_a(-0.00010597251093713567)),(to_sfixed_a(-0.00014719023602083325)),(to_sfixed_a(0.0016653880011290312)),(to_sfixed_a(0.28915926814079285)),(to_sfixed_a(6.153830327093601e-06)),(to_sfixed_a(1.0136489436263219e-05)),(to_sfixed_a(-0.0015166293596848845)),(to_sfixed_a(-0.0005651055835187435)),(to_sfixed_a(-2.736778696998954e-07)),(to_sfixed_a(-6.265618139877915e-05)),(to_sfixed_a(-0.0005259586614556611)),(to_sfixed_a(5.477659942698665e-05)),(to_sfixed_a(-1.1430976883275434e-05)),(to_sfixed_a(-7.278061093529686e-05)),(to_sfixed_a(-0.0016995702171698213)),(to_sfixed_a(0.003588475054129958)),(to_sfixed_a(0.0017842589877545834)),(to_sfixed_a(7.2953407652676105e-06)),(to_sfixed_a(-0.00018325414566788822)),(to_sfixed_a(0.0013226348673924804)),(to_sfixed_a(-6.180554919410497e-06)),(to_sfixed_a(0.00010744674364104867)),(to_sfixed_a(0.0022599671501666307)),(to_sfixed_a(-0.0002976249670609832)),(to_sfixed_a(3.725876013049856e-05)),(to_sfixed_a(0.13626451790332794)),(to_sfixed_a(-0.00016909702389966697)),(to_sfixed_a(0.0011235473211854696)),(to_sfixed_a(-5.734166734328028e-06)),(to_sfixed_a(5.5284308473346755e-05)),(to_sfixed_a(-0.00014994523371569812)),(to_sfixed_a(-0.00015079707372933626)),(to_sfixed_a(0.0032767511438578367)),(to_sfixed_a(0.000347750261425972)),(to_sfixed_a(0.000527341035194695)),(to_sfixed_a(0.0006895042024552822)),(to_sfixed_a(-0.00010438114986754954)),(to_sfixed_a(0.00576564809307456)),(to_sfixed_a(-0.0002480066323187202)),(to_sfixed_a(-1.1555806850083172e-05)),(to_sfixed_a(-0.5829349160194397)),(to_sfixed_a(0.0006014800746925175)),(to_sfixed_a(0.0018530349479988217)),(to_sfixed_a(0.00010725209722295403)),(to_sfixed_a(0.002526924479752779)),(to_sfixed_a(-0.0022670335602015257)),(to_sfixed_a(-0.010659760795533657)),(to_sfixed_a(-0.0004991978057660162)),(to_sfixed_a(-0.5485532879829407)),(to_sfixed_a(0.3422817587852478)),(to_sfixed_a(0.0001100789086194709)),(to_sfixed_a(0.005501497071236372)),(to_sfixed_a(0.00021666844259016216)),(to_sfixed_a(-0.00028825041954405606)),(to_sfixed_a(8.155271643772721e-06)),(to_sfixed_a(6.516746361739933e-05)),(to_sfixed_a(0.18760491907596588)),(to_sfixed_a(0.003726822789758444)),(to_sfixed_a(-1.27000967040658e-05)),(to_sfixed_a(0.0051720039919018745)),(to_sfixed_a(0.0004960647784173489)),(to_sfixed_a(8.227187936427072e-05)),(to_sfixed_a(0.04376501590013504)),(to_sfixed_a(-0.0017307654488831758)),(to_sfixed_a(0.00010583629773464054)),(to_sfixed_a(0.002376002725213766)),(to_sfixed_a(3.660787479020655e-05)),(to_sfixed_a(-0.00028126631514169276)),(to_sfixed_a(-0.010560265742242336)),(to_sfixed_a(-0.00018059922149404883)),(to_sfixed_a(-2.8011956601403654e-05)),(to_sfixed_a(-6.663560634478927e-05)),(to_sfixed_a(0.00030654409783892334)),(to_sfixed_a(0.00010316280531696975)),(to_sfixed_a(0.0001079783178283833)),(to_sfixed_a(0.00148022233042866)),(to_sfixed_a(-0.014189316891133785)),(to_sfixed_a(-0.030884642153978348)),(to_sfixed_a(-0.051702480763196945)),(to_sfixed_a(0.015217484906315804)),(to_sfixed_a(-0.00011965323938056827)),(to_sfixed_a(-8.468705345876515e-07)),(to_sfixed_a(-3.44500585924834e-06)),(to_sfixed_a(-0.00010898172331508249)),(to_sfixed_a(3.815839590970427e-07)),(to_sfixed_a(-0.0004517444467637688)),(to_sfixed_a(-7.77783861849457e-05)),(to_sfixed_a(0.21151615679264069)),(to_sfixed_a(0.012157067656517029)),(to_sfixed_a(-6.958529411349446e-06)),(to_sfixed_a(0.00013676095113623887)),(to_sfixed_a(7.731383084319532e-05)),(to_sfixed_a(0.0001294564426643774)),(to_sfixed_a(0.00045316381147131324)),(to_sfixed_a(-0.14706233143806458)),(to_sfixed_a(0.00023622237495146692)),(to_sfixed_a(-0.0003844235616270453)),(to_sfixed_a(0.00011375146277714521)),(to_sfixed_a(-0.00444530975073576)),(to_sfixed_a(-0.25593289732933044)),(to_sfixed_a(0.006716730538755655)),(to_sfixed_a(4.996145435143262e-06)),(to_sfixed_a(9.9067525297869e-05)),(to_sfixed_a(-0.000159441027790308)),(to_sfixed_a(-0.003266579005867243)),(to_sfixed_a(0.00028057958115823567)),(to_sfixed_a(0.041879553347826004)),(to_sfixed_a(-2.0703781046904624e-05)),(to_sfixed_a(0.0013972477754577994)),(to_sfixed_a(-1.6106932889670134e-06)),(to_sfixed_a(0.004746321123093367)),(to_sfixed_a(0.00011355915921740234)),(to_sfixed_a(-0.4915298819541931)),(to_sfixed_a(0.00014682364417240024)),(to_sfixed_a(0.22717882692813873)),(to_sfixed_a(0.001692021731287241)),(to_sfixed_a(0.6638005375862122)),(to_sfixed_a(0.002894619945436716)),(to_sfixed_a(-0.00013681285781785846)),(to_sfixed_a(0.2115190178155899)),(to_sfixed_a(-0.002958361292257905)),(to_sfixed_a(0.00012933177640661597)),(to_sfixed_a(-0.00016685274022165686)),(to_sfixed_a(-0.0001086939373635687)),(to_sfixed_a(-0.00032439519418403506)),(to_sfixed_a(-0.2692335844039917)),(to_sfixed_a(-0.3293164372444153)),(to_sfixed_a(-0.00010231410851702094)),(to_sfixed_a(0.0001260123390238732)),(to_sfixed_a(-0.00041350460378453135)),(to_sfixed_a(-4.490854553296231e-05)),(to_sfixed_a(-0.2627393901348114)),(to_sfixed_a(0.00013122570817358792)),(to_sfixed_a(0.00010078912600874901)),(to_sfixed_a(-0.00017567683244124055)),(to_sfixed_a(-0.00021599885076284409)),(to_sfixed_a(2.2767817426938564e-05)),(to_sfixed_a(-2.3540997062809765e-07)),(to_sfixed_a(-5.794248136226088e-05)),(to_sfixed_a(0.041782669723033905)),(to_sfixed_a(0.006351520773023367)),(to_sfixed_a(-0.00017060263780876994)),(to_sfixed_a(-7.329306390602142e-05)),(to_sfixed_a(0.00010236575326416641)),(to_sfixed_a(0.00011019327212125063)),(to_sfixed_a(0.004978662822395563)),(to_sfixed_a(0.003532635048031807)),(to_sfixed_a(-0.00539100356400013)),(to_sfixed_a(0.006380733102560043)),(to_sfixed_a(0.0018480572616681457)),(to_sfixed_a(-0.0002964842424262315)),(to_sfixed_a(0.00023754512949381024)),(to_sfixed_a(-2.7729300200007856e-05)),(to_sfixed_a(0.0003245555271860212)),(to_sfixed_a(2.2607946448260918e-05)),(to_sfixed_a(-1.7293787095695734e-06)),(to_sfixed_a(9.183413567370735e-06)),(to_sfixed_a(-0.011569026857614517)),(to_sfixed_a(-0.00044220403651706874)),(to_sfixed_a(0.00255887140519917)),(to_sfixed_a(0.003106840653344989)),(to_sfixed_a(0.1919817477464676)),(to_sfixed_a(0.007509094197303057)),(to_sfixed_a(0.00015592521231155843)),(to_sfixed_a(0.0031525520607829094)),(to_sfixed_a(0.0025349589996039867)),(to_sfixed_a(-0.0035032855812460184)),(to_sfixed_a(-8.76322083058767e-05)),(to_sfixed_a(-0.0017007880378514528)),(to_sfixed_a(0.15509535372257233)),(to_sfixed_a(-0.006495609413832426)));

    constant weight_n2_91 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.011748701333999634)),(to_sfixed_a(0.0009626122191548347)),(to_sfixed_a(0.0008973328513093293)),(to_sfixed_a(1.422295463271439e-05)),(to_sfixed_a(0.000808662036433816)),(to_sfixed_a(-0.00013509424752555788)),(to_sfixed_a(-0.000123189965961501)),(to_sfixed_a(8.310785779030994e-05)),(to_sfixed_a(-0.00023896837956272066)),(to_sfixed_a(-0.0001470165589125827)),(to_sfixed_a(2.547039184719324e-05)),(to_sfixed_a(0.0010255291126668453)),(to_sfixed_a(-0.013020014390349388)),(to_sfixed_a(-0.004160420037806034)),(to_sfixed_a(-6.007774572935887e-05)),(to_sfixed_a(-0.00028905842918902636)),(to_sfixed_a(0.18395964801311493)),(to_sfixed_a(9.370419138576835e-05)),(to_sfixed_a(0.14916887879371643)),(to_sfixed_a(-0.005016193725168705)),(to_sfixed_a(4.500073555391282e-05)),(to_sfixed_a(-9.194274753099307e-05)),(to_sfixed_a(0.00016521917132195085)),(to_sfixed_a(-0.006057885475456715)),(to_sfixed_a(0.0015005867462605238)),(to_sfixed_a(-0.0003113849088549614)),(to_sfixed_a(0.00020602569566108286)),(to_sfixed_a(0.0008329435950145125)),(to_sfixed_a(0.0003702231333591044)),(to_sfixed_a(0.00011650154192466289)),(to_sfixed_a(0.00012115256686229259)),(to_sfixed_a(-4.706930121756159e-05)),(to_sfixed_a(-0.005706273019313812)),(to_sfixed_a(-0.00021164440840948373)),(to_sfixed_a(5.589208740275353e-06)),(to_sfixed_a(0.00013881945051252842)),(to_sfixed_a(0.017148621380329132)),(to_sfixed_a(-0.16131319105625153)),(to_sfixed_a(-0.00022230867762118578)),(to_sfixed_a(0.0001398917374899611)),(to_sfixed_a(-0.33016353845596313)),(to_sfixed_a(-0.0018431926146149635)),(to_sfixed_a(-7.517149788327515e-05)),(to_sfixed_a(-7.025616650935262e-05)),(to_sfixed_a(9.320032404502854e-06)),(to_sfixed_a(0.001842379686422646)),(to_sfixed_a(-0.00014152421499602497)),(to_sfixed_a(0.0023956596851348877)),(to_sfixed_a(0.00011426446144469082)),(to_sfixed_a(-0.0029825158417224884)),(to_sfixed_a(0.0008581032161600888)),(to_sfixed_a(0.0005994071252644062)),(to_sfixed_a(-3.9167149225249887e-05)),(to_sfixed_a(0.0002551862271502614)),(to_sfixed_a(-0.008253967389464378)),(to_sfixed_a(-0.0018093858379870653)),(to_sfixed_a(-0.00018014886882156134)),(to_sfixed_a(0.0004486257676035166)),(to_sfixed_a(-6.0290614783298224e-05)),(to_sfixed_a(-0.00015437034016940743)),(to_sfixed_a(0.0020608403719961643)),(to_sfixed_a(-0.00016135723853949457)),(to_sfixed_a(0.00046251670573838055)),(to_sfixed_a(0.0010724249295890331)),(to_sfixed_a(0.00017332323477603495)),(to_sfixed_a(0.20173802971839905)),(to_sfixed_a(1.0059682608698495e-05)),(to_sfixed_a(-0.0028396728448569775)),(to_sfixed_a(8.593194070272148e-05)),(to_sfixed_a(-5.849435183336027e-05)),(to_sfixed_a(0.0013742432929575443)),(to_sfixed_a(0.0008526094607077539)),(to_sfixed_a(0.10034853219985962)),(to_sfixed_a(-1.129370866692625e-05)),(to_sfixed_a(0.00011912740592379123)),(to_sfixed_a(-4.436542803887278e-05)),(to_sfixed_a(-0.0009232918964698911)),(to_sfixed_a(0.0005970866186544299)),(to_sfixed_a(-5.416892236098647e-05)),(to_sfixed_a(-0.0001092588936444372)),(to_sfixed_a(0.0001681245194049552)),(to_sfixed_a(-0.00012892414815723896)),(to_sfixed_a(0.0005158072453923523)),(to_sfixed_a(0.0011109558399766684)),(to_sfixed_a(0.00030811221222393215)),(to_sfixed_a(0.001214119023643434)),(to_sfixed_a(-0.007141763810068369)),(to_sfixed_a(0.0008594001410529017)),(to_sfixed_a(-5.123187293065712e-05)),(to_sfixed_a(-0.00011309038382023573)),(to_sfixed_a(0.001440596068277955)),(to_sfixed_a(7.695555541431531e-05)),(to_sfixed_a(0.0017795967869460583)),(to_sfixed_a(-0.00012916269770357758)),(to_sfixed_a(0.36249983310699463)),(to_sfixed_a(-0.00010521471267566085)),(to_sfixed_a(2.989698259625584e-05)),(to_sfixed_a(-0.00025126885157078505)),(to_sfixed_a(0.00028197941719554365)),(to_sfixed_a(-2.4322671379195526e-06)),(to_sfixed_a(0.0003347611636854708)),(to_sfixed_a(0.0009111920953728259)),(to_sfixed_a(-1.9839644664898515e-06)),(to_sfixed_a(-0.00016018559108488262)),(to_sfixed_a(0.002703750506043434)),(to_sfixed_a(0.0005269546527415514)),(to_sfixed_a(0.00030096093541942537)),(to_sfixed_a(-0.00011312344577163458)),(to_sfixed_a(-0.0003867574851028621)),(to_sfixed_a(0.0009802093263715506)),(to_sfixed_a(-0.40403395891189575)),(to_sfixed_a(-0.00011205117334611714)),(to_sfixed_a(-0.00015166669618338346)),(to_sfixed_a(-0.00017457656213082373)),(to_sfixed_a(-0.00010691281931940466)),(to_sfixed_a(0.0023584768641740084)),(to_sfixed_a(-0.0006999021279625595)),(to_sfixed_a(-3.491837560432032e-05)),(to_sfixed_a(0.000173346750671044)),(to_sfixed_a(-0.006280485074967146)),(to_sfixed_a(-0.00011344396625645459)),(to_sfixed_a(-1.219565820065327e-05)),(to_sfixed_a(0.00044923374662175775)),(to_sfixed_a(0.00011357428593328223)),(to_sfixed_a(0.00016947995754890144)),(to_sfixed_a(-0.00015638260811101645)),(to_sfixed_a(0.0019149752333760262)),(to_sfixed_a(0.0001707777555566281)),(to_sfixed_a(-1.3173281331546605e-05)),(to_sfixed_a(-4.081884981133044e-07)),(to_sfixed_a(0.00015034162788651884)),(to_sfixed_a(4.0907616494223475e-07)),(to_sfixed_a(0.0003286387072876096)),(to_sfixed_a(0.0024906727485358715)),(to_sfixed_a(1.4913384802639484e-06)),(to_sfixed_a(0.00010359013685956597)),(to_sfixed_a(0.003396501298993826)),(to_sfixed_a(-9.843150473898277e-05)),(to_sfixed_a(-1.1429554433561862e-05)),(to_sfixed_a(0.0001508756831753999)),(to_sfixed_a(-2.1074170945212245e-05)),(to_sfixed_a(0.0004470851563382894)),(to_sfixed_a(-0.0001295888505410403)),(to_sfixed_a(9.49637615121901e-05)),(to_sfixed_a(-2.8082395147066563e-06)),(to_sfixed_a(-2.234756902907975e-05)),(to_sfixed_a(-2.468455204507336e-05)),(to_sfixed_a(0.0001899988710647449)),(to_sfixed_a(0.000113509529910516)),(to_sfixed_a(-4.0373670344706625e-05)),(to_sfixed_a(0.00027135221171192825)),(to_sfixed_a(0.00017682448378764093)),(to_sfixed_a(8.658620208734646e-05)),(to_sfixed_a(-1.1845582776004449e-05)),(to_sfixed_a(0.00023797358153387904)),(to_sfixed_a(-0.001168587477877736)),(to_sfixed_a(-0.00016721428255550563)),(to_sfixed_a(-0.0006755740032531321)),(to_sfixed_a(-5.562771184486337e-05)),(to_sfixed_a(-0.00017543967987876385)),(to_sfixed_a(0.00012749414599966258)),(to_sfixed_a(3.267763531766832e-06)),(to_sfixed_a(0.0019991733133792877)),(to_sfixed_a(0.0002081787388306111)),(to_sfixed_a(-0.0010682932334020734)),(to_sfixed_a(0.0005807943525724113)),(to_sfixed_a(6.804466102039441e-05)),(to_sfixed_a(0.0010873153805732727)),(to_sfixed_a(3.89264605473727e-05)),(to_sfixed_a(-0.00020048805163241923)),(to_sfixed_a(0.0006981816259212792)),(to_sfixed_a(-2.662494807736948e-05)),(to_sfixed_a(-0.00020125934679526836)),(to_sfixed_a(-0.00013561599189415574)),(to_sfixed_a(-0.024209540337324142)),(to_sfixed_a(1.8483729945728555e-05)),(to_sfixed_a(-0.0020095109939575195)),(to_sfixed_a(0.0016391262179240584)),(to_sfixed_a(-0.010870442725718021)),(to_sfixed_a(0.0013940819771960378)),(to_sfixed_a(0.0009587852982804179)),(to_sfixed_a(0.0006632445147261024)),(to_sfixed_a(-6.607925752177835e-05)),(to_sfixed_a(-8.978608821053058e-05)),(to_sfixed_a(-0.00013213575584813952)),(to_sfixed_a(0.00023874620092101395)),(to_sfixed_a(0.0013101856457069516)),(to_sfixed_a(0.0006175680900923908)),(to_sfixed_a(-0.00013069499982520938)),(to_sfixed_a(-4.228411489748396e-05)),(to_sfixed_a(-0.016349175944924355)),(to_sfixed_a(0.00018642710347194225)),(to_sfixed_a(0.0013537092600017786)),(to_sfixed_a(0.0022106515243649483)),(to_sfixed_a(-0.0002451069885864854)),(to_sfixed_a(0.00022177401115186512)),(to_sfixed_a(7.238877878990024e-05)),(to_sfixed_a(2.9385555535554886e-05)),(to_sfixed_a(0.00033949140924960375)),(to_sfixed_a(0.00010172116162721068)),(to_sfixed_a(0.00023224408505484462)),(to_sfixed_a(0.0002823626564349979)),(to_sfixed_a(-8.308541146107018e-05)),(to_sfixed_a(0.0002922256535384804)),(to_sfixed_a(9.247040725313127e-05)),(to_sfixed_a(6.813713844167069e-05)),(to_sfixed_a(-0.0007567162392660975)),(to_sfixed_a(-0.002382952719926834)),(to_sfixed_a(0.0008918905514292419)),(to_sfixed_a(2.027592927333899e-06)),(to_sfixed_a(-0.0064404490403831005)),(to_sfixed_a(-9.987672819988802e-05)),(to_sfixed_a(6.0609232605202124e-05)),(to_sfixed_a(8.304696530103683e-05)),(to_sfixed_a(1.9857398001477122e-06)),(to_sfixed_a(7.606358849443495e-05)),(to_sfixed_a(-6.380701051966753e-06)),(to_sfixed_a(0.0012337386142462492)),(to_sfixed_a(-0.003439187305048108)),(to_sfixed_a(0.00018719627405516803)),(to_sfixed_a(-7.14271591277793e-05)),(to_sfixed_a(7.062160148052499e-05)),(to_sfixed_a(-7.150015153456479e-05)),(to_sfixed_a(-2.838146610883996e-05)),(to_sfixed_a(0.27342936396598816)),(to_sfixed_a(-1.8369100871495903e-06)),(to_sfixed_a(-5.708840035367757e-05)),(to_sfixed_a(1.0950156138278544e-05)),(to_sfixed_a(-0.08233920484781265)),(to_sfixed_a(-0.0009188373223878443)),(to_sfixed_a(0.003172691445797682)),(to_sfixed_a(-0.0001059536516549997)),(to_sfixed_a(0.0003153387806378305)),(to_sfixed_a(-4.47034472017549e-06)),(to_sfixed_a(5.391923332354054e-05)),(to_sfixed_a(-0.0001462075742892921)),(to_sfixed_a(0.0019729435443878174)),(to_sfixed_a(0.00015642453217878938)),(to_sfixed_a(-0.00018954166444018483)),(to_sfixed_a(-6.750845204805955e-05)),(to_sfixed_a(-9.34308918658644e-05)),(to_sfixed_a(0.00012753508053719997)),(to_sfixed_a(0.0003581643686629832)),(to_sfixed_a(-0.0002928363101091236)),(to_sfixed_a(0.0008804980898275971)),(to_sfixed_a(-3.701010064105503e-05)),(to_sfixed_a(0.0016907905228435993)),(to_sfixed_a(0.0018890111241489649)),(to_sfixed_a(2.3204429453471676e-05)),(to_sfixed_a(-9.691900049801916e-05)),(to_sfixed_a(0.0003343548742122948)),(to_sfixed_a(-0.00013501665671356022)),(to_sfixed_a(0.0003972767444793135)),(to_sfixed_a(-0.00011655157140921801)),(to_sfixed_a(0.00019814661936834455)),(to_sfixed_a(-7.914623711258173e-05)),(to_sfixed_a(-0.00725628761574626)),(to_sfixed_a(-1.9156492271577008e-05)),(to_sfixed_a(-5.530164344236255e-06)),(to_sfixed_a(0.1790526658296585)),(to_sfixed_a(0.0001717672566883266)),(to_sfixed_a(0.0005440001259557903)),(to_sfixed_a(-0.0002309454430360347)),(to_sfixed_a(0.00033249345142394304)),(to_sfixed_a(6.271267193369567e-05)),(to_sfixed_a(-3.932173422072083e-05)),(to_sfixed_a(7.161525718402117e-05)),(to_sfixed_a(-0.00016332042287103832)),(to_sfixed_a(0.00013638101518154144)),(to_sfixed_a(0.00033105252077803016)),(to_sfixed_a(0.0048246076330542564)),(to_sfixed_a(-2.049418253591284e-05)),(to_sfixed_a(-0.00030771922320127487)),(to_sfixed_a(4.068117414135486e-05)),(to_sfixed_a(9.346805018140003e-05)),(to_sfixed_a(-0.0006903134053573012)),(to_sfixed_a(0.0021161455661058426)),(to_sfixed_a(-5.8284844271838665e-05)),(to_sfixed_a(0.0013638150412589312)),(to_sfixed_a(0.0012954875128343701)),(to_sfixed_a(0.00014630270015913993)),(to_sfixed_a(0.00029194989474490285)),(to_sfixed_a(-8.886454452294856e-06)),(to_sfixed_a(-0.008924315683543682)),(to_sfixed_a(6.321343971649185e-05)),(to_sfixed_a(7.8826371463947e-05)),(to_sfixed_a(-0.0016882981872186065)),(to_sfixed_a(0.00022262676793616265)),(to_sfixed_a(-9.779963875189424e-06)),(to_sfixed_a(0.0019677337259054184)),(to_sfixed_a(0.0007814886048436165)),(to_sfixed_a(-8.347077528014779e-05)),(to_sfixed_a(0.0005294120637699962)),(to_sfixed_a(0.00011662447650451213)),(to_sfixed_a(0.000854849407915026)),(to_sfixed_a(-0.005133009050041437)),(to_sfixed_a(0.0007486058166250587)),(to_sfixed_a(3.971209662267938e-05)),(to_sfixed_a(-0.002750437706708908)),(to_sfixed_a(-0.007664048578590155)),(to_sfixed_a(0.0011941551929339767)));

    constant weight_n2_92 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.41708341240882874)),(to_sfixed_a(-0.045987412333488464)),(to_sfixed_a(-0.0032608909532427788)),(to_sfixed_a(6.320769898593426e-07)),(to_sfixed_a(-0.008265466429293156)),(to_sfixed_a(-0.00011233532859478146)),(to_sfixed_a(-0.009152733720839024)),(to_sfixed_a(0.00013402814511209726)),(to_sfixed_a(-0.00010669781477190554)),(to_sfixed_a(-0.00014926522271707654)),(to_sfixed_a(-0.00010783308243844658)),(to_sfixed_a(-0.031058045104146004)),(to_sfixed_a(-0.006877577397972345)),(to_sfixed_a(0.001591916079632938)),(to_sfixed_a(0.0001808523666113615)),(to_sfixed_a(6.079044396756217e-07)),(to_sfixed_a(-0.014679986983537674)),(to_sfixed_a(0.00010156893404200673)),(to_sfixed_a(0.002927914960309863)),(to_sfixed_a(0.004676260519772768)),(to_sfixed_a(4.348301445133984e-05)),(to_sfixed_a(0.00019573629833757877)),(to_sfixed_a(-1.3480632333084941e-05)),(to_sfixed_a(0.0017810333520174026)),(to_sfixed_a(-0.0096860621124506)),(to_sfixed_a(-0.0005039084353484213)),(to_sfixed_a(3.6151817766949534e-05)),(to_sfixed_a(-0.00023435463663190603)),(to_sfixed_a(-0.0013032385613769293)),(to_sfixed_a(-2.797688648570329e-05)),(to_sfixed_a(-0.006086953449994326)),(to_sfixed_a(-1.9819377484964207e-05)),(to_sfixed_a(-0.003066104371100664)),(to_sfixed_a(5.835351112182252e-05)),(to_sfixed_a(-0.00011555308446986601)),(to_sfixed_a(0.0003123974602203816)),(to_sfixed_a(-0.012097816914319992)),(to_sfixed_a(-0.08025165647268295)),(to_sfixed_a(-0.006922573316842318)),(to_sfixed_a(-2.9766197258140892e-05)),(to_sfixed_a(-0.010851524770259857)),(to_sfixed_a(0.006239766720682383)),(to_sfixed_a(-0.00014585521421395242)),(to_sfixed_a(-8.749469998292625e-06)),(to_sfixed_a(-0.09209395200014114)),(to_sfixed_a(-0.01979142054915428)),(to_sfixed_a(-0.0034664447885006666)),(to_sfixed_a(-0.003912223502993584)),(to_sfixed_a(-0.00019220897229388356)),(to_sfixed_a(-0.00696773873642087)),(to_sfixed_a(-0.6040251851081848)),(to_sfixed_a(-3.7065110518597066e-05)),(to_sfixed_a(5.6696750107221305e-05)),(to_sfixed_a(-0.001908021979033947)),(to_sfixed_a(-0.013859191909432411)),(to_sfixed_a(-0.005177756305783987)),(to_sfixed_a(-0.00011214325786568224)),(to_sfixed_a(-0.009031391702592373)),(to_sfixed_a(-0.00011566847388166934)),(to_sfixed_a(1.8316088244318962e-05)),(to_sfixed_a(-0.009728462435305119)),(to_sfixed_a(0.170720636844635)),(to_sfixed_a(-0.001248981337994337)),(to_sfixed_a(-0.013733187690377235)),(to_sfixed_a(0.00017884024418890476)),(to_sfixed_a(0.0025648181326687336)),(to_sfixed_a(6.951912655495107e-05)),(to_sfixed_a(-0.0004735890543088317)),(to_sfixed_a(-0.004197688773274422)),(to_sfixed_a(-0.00011361097858753055)),(to_sfixed_a(-0.04973527044057846)),(to_sfixed_a(-0.0007744646281935275)),(to_sfixed_a(-0.010378253646194935)),(to_sfixed_a(-5.618316208710894e-05)),(to_sfixed_a(-0.00010654432117007673)),(to_sfixed_a(-0.0001516568154329434)),(to_sfixed_a(-0.001424035057425499)),(to_sfixed_a(-0.007931876927614212)),(to_sfixed_a(7.940069190226495e-05)),(to_sfixed_a(-0.3557591438293457)),(to_sfixed_a(-0.011991111561655998)),(to_sfixed_a(-1.1718315363395959e-05)),(to_sfixed_a(-0.0014156410470604897)),(to_sfixed_a(-0.0022768559865653515)),(to_sfixed_a(2.884346031351015e-05)),(to_sfixed_a(-0.004559300374239683)),(to_sfixed_a(0.003919479437172413)),(to_sfixed_a(-0.2611096203327179)),(to_sfixed_a(-3.071545506827533e-05)),(to_sfixed_a(-2.3265602067112923e-05)),(to_sfixed_a(-0.0029453278984874487)),(to_sfixed_a(1.0306081094313413e-05)),(to_sfixed_a(-0.008472444489598274)),(to_sfixed_a(7.367753278231248e-05)),(to_sfixed_a(-0.0025238923262804747)),(to_sfixed_a(-1.2784556020051241e-05)),(to_sfixed_a(-7.12647961336188e-05)),(to_sfixed_a(-1.2118456652387977e-05)),(to_sfixed_a(0.0001552049070596695)),(to_sfixed_a(-7.953217573231086e-05)),(to_sfixed_a(-0.0017234513070434332)),(to_sfixed_a(-0.0022297799587249756)),(to_sfixed_a(0.0001541859091958031)),(to_sfixed_a(-0.005971906706690788)),(to_sfixed_a(-0.021120639517903328)),(to_sfixed_a(-0.3312487304210663)),(to_sfixed_a(3.974189894506708e-06)),(to_sfixed_a(-0.00014064252900425345)),(to_sfixed_a(-0.00012847979087382555)),(to_sfixed_a(0.20710483193397522)),(to_sfixed_a(0.5158164501190186)),(to_sfixed_a(-3.0075618269620463e-05)),(to_sfixed_a(-0.0023272731341421604)),(to_sfixed_a(-6.281315290834755e-05)),(to_sfixed_a(-0.00014833835302852094)),(to_sfixed_a(-0.027620146051049232)),(to_sfixed_a(0.0060166665352880955)),(to_sfixed_a(0.144237220287323)),(to_sfixed_a(-3.058828951907344e-06)),(to_sfixed_a(-0.00021832509082742035)),(to_sfixed_a(0.00024216082238126546)),(to_sfixed_a(2.4307420972036198e-05)),(to_sfixed_a(-0.006745899561792612)),(to_sfixed_a(-8.991867071017623e-05)),(to_sfixed_a(3.8945065170992166e-05)),(to_sfixed_a(0.0034236754290759563)),(to_sfixed_a(0.5197188258171082)),(to_sfixed_a(-0.00023559674446005374)),(to_sfixed_a(-0.00029255080153234303)),(to_sfixed_a(-1.6548310668440536e-06)),(to_sfixed_a(-0.0002043947170022875)),(to_sfixed_a(7.2010065196082e-05)),(to_sfixed_a(-0.0005956231616437435)),(to_sfixed_a(-0.028635812923312187)),(to_sfixed_a(-0.00019973293819930404)),(to_sfixed_a(0.00016864435747265816)),(to_sfixed_a(-0.011252916418015957)),(to_sfixed_a(-9.345672151539475e-05)),(to_sfixed_a(3.0704468372277915e-05)),(to_sfixed_a(3.6875324440188706e-05)),(to_sfixed_a(-0.0004311562515795231)),(to_sfixed_a(5.7903169363271445e-05)),(to_sfixed_a(-0.0002108710614265874)),(to_sfixed_a(4.387208173284307e-05)),(to_sfixed_a(0.21151156723499298)),(to_sfixed_a(-0.0004296520201023668)),(to_sfixed_a(-8.541136048734188e-05)),(to_sfixed_a(0.0001510394795332104)),(to_sfixed_a(0.0002509369805920869)),(to_sfixed_a(-0.0025934195145964622)),(to_sfixed_a(5.0032649596687406e-05)),(to_sfixed_a(-4.761459422297776e-07)),(to_sfixed_a(0.0008200600859709084)),(to_sfixed_a(-3.9986101910471916e-05)),(to_sfixed_a(-0.00018048704077955335)),(to_sfixed_a(-0.0067601497285068035)),(to_sfixed_a(3.777834353968501e-05)),(to_sfixed_a(8.653031545691192e-05)),(to_sfixed_a(7.418366294587031e-06)),(to_sfixed_a(2.282497371197678e-05)),(to_sfixed_a(4.576535866362974e-05)),(to_sfixed_a(9.853829396888614e-08)),(to_sfixed_a(0.0008091232739388943)),(to_sfixed_a(0.0002989159256685525)),(to_sfixed_a(-0.0004074445751029998)),(to_sfixed_a(-0.0004943466046825051)),(to_sfixed_a(-0.0001309469371335581)),(to_sfixed_a(-0.6635953783988953)),(to_sfixed_a(-4.595619975589216e-05)),(to_sfixed_a(-0.00042175970156677067)),(to_sfixed_a(-0.007599617820233107)),(to_sfixed_a(-0.00020404842507559806)),(to_sfixed_a(0.16571711003780365)),(to_sfixed_a(-4.021429049316794e-05)),(to_sfixed_a(-0.519849956035614)),(to_sfixed_a(-0.0025665410794317722)),(to_sfixed_a(-0.0001867062965175137)),(to_sfixed_a(-0.22693586349487305)),(to_sfixed_a(-0.21014109253883362)),(to_sfixed_a(-0.0071174632757902145)),(to_sfixed_a(9.412199142389e-05)),(to_sfixed_a(-0.01843724399805069)),(to_sfixed_a(6.400077836588025e-07)),(to_sfixed_a(0.00015779249952174723)),(to_sfixed_a(0.00016724148008506745)),(to_sfixed_a(-0.008418052457273006)),(to_sfixed_a(-0.011591056361794472)),(to_sfixed_a(0.002794816391542554)),(to_sfixed_a(0.00633217254653573)),(to_sfixed_a(0.004730953834950924)),(to_sfixed_a(0.013663452118635178)),(to_sfixed_a(0.00015399206313304603)),(to_sfixed_a(-0.008154502138495445)),(to_sfixed_a(-0.007467071060091257)),(to_sfixed_a(0.00016655099170748144)),(to_sfixed_a(3.8131278415676206e-05)),(to_sfixed_a(-0.00010068002302432433)),(to_sfixed_a(-0.002310203853994608)),(to_sfixed_a(-0.007847066037356853)),(to_sfixed_a(0.00019565486581996083)),(to_sfixed_a(0.0001013561268337071)),(to_sfixed_a(-8.968608744908124e-05)),(to_sfixed_a(-0.000449889077572152)),(to_sfixed_a(-0.00018664698291104287)),(to_sfixed_a(0.00013635987124871463)),(to_sfixed_a(0.0008515706285834312)),(to_sfixed_a(-0.0009165071533061564)),(to_sfixed_a(0.032019734382629395)),(to_sfixed_a(-5.5050451919669285e-05)),(to_sfixed_a(0.00014721808838658035)),(to_sfixed_a(0.001277248258702457)),(to_sfixed_a(0.00013210708857513964)),(to_sfixed_a(-0.00023687387874815613)),(to_sfixed_a(0.0001252333604497835)),(to_sfixed_a(-6.852387741673738e-05)),(to_sfixed_a(-3.194367673131637e-05)),(to_sfixed_a(0.002686743624508381)),(to_sfixed_a(-0.32928913831710815)),(to_sfixed_a(0.0019248173339292407)),(to_sfixed_a(-3.0071088986005634e-05)),(to_sfixed_a(-6.756297807442024e-05)),(to_sfixed_a(3.2816351449582726e-05)),(to_sfixed_a(2.402157406322658e-06)),(to_sfixed_a(-0.00023955953656695783)),(to_sfixed_a(-0.012166537344455719)),(to_sfixed_a(7.741311128484085e-05)),(to_sfixed_a(-0.00019721627177204937)),(to_sfixed_a(0.0002932208590209484)),(to_sfixed_a(0.0001055652683135122)),(to_sfixed_a(-0.0066890413872897625)),(to_sfixed_a(-0.006558158900588751)),(to_sfixed_a(0.00027876629610545933)),(to_sfixed_a(-0.00019641799735836685)),(to_sfixed_a(-0.00013048594701103866)),(to_sfixed_a(-0.004720093682408333)),(to_sfixed_a(0.0005466067814268172)),(to_sfixed_a(0.37218403816223145)),(to_sfixed_a(1.808422530302778e-05)),(to_sfixed_a(0.002027107635512948)),(to_sfixed_a(-4.143294063396752e-06)),(to_sfixed_a(-0.004993612878024578)),(to_sfixed_a(9.892569505609572e-05)),(to_sfixed_a(-0.0031429638620465994)),(to_sfixed_a(-0.00010766007471829653)),(to_sfixed_a(-0.005277839954942465)),(to_sfixed_a(-0.00094894680660218)),(to_sfixed_a(-0.1818760484457016)),(to_sfixed_a(0.5075873732566833)),(to_sfixed_a(-0.00016801941092126071)),(to_sfixed_a(-0.01508881151676178)),(to_sfixed_a(-0.019194692373275757)),(to_sfixed_a(-0.000175066918018274)),(to_sfixed_a(0.001468475442379713)),(to_sfixed_a(2.3366170353256166e-05)),(to_sfixed_a(-9.717619104776531e-05)),(to_sfixed_a(-0.010794584639370441)),(to_sfixed_a(0.002537994645535946)),(to_sfixed_a(-3.417313564568758e-06)),(to_sfixed_a(-0.00020331956329755485)),(to_sfixed_a(-0.0020575341768562794)),(to_sfixed_a(7.021590135991573e-05)),(to_sfixed_a(-0.00030565151246264577)),(to_sfixed_a(3.9081438444554806e-05)),(to_sfixed_a(5.77784376218915e-05)),(to_sfixed_a(0.00032101868418976665)),(to_sfixed_a(-0.012485206127166748)),(to_sfixed_a(3.398003173060715e-06)),(to_sfixed_a(4.0852464735507965e-06)),(to_sfixed_a(-0.00011664150952128693)),(to_sfixed_a(0.003313204739242792)),(to_sfixed_a(-0.022194597870111465)),(to_sfixed_a(0.0001126510469475761)),(to_sfixed_a(-7.610101602040231e-05)),(to_sfixed_a(-0.00019940134370699525)),(to_sfixed_a(0.00020488408335950226)),(to_sfixed_a(-0.010112732648849487)),(to_sfixed_a(-0.00885837059468031)),(to_sfixed_a(-0.375163733959198)),(to_sfixed_a(0.025199219584465027)),(to_sfixed_a(-0.21136406064033508)),(to_sfixed_a(-0.00029723928309977055)),(to_sfixed_a(4.822482151212171e-05)),(to_sfixed_a(-0.00014739451580680907)),(to_sfixed_a(0.006074142176657915)),(to_sfixed_a(5.3856128943152726e-06)),(to_sfixed_a(-0.0003001305740326643)),(to_sfixed_a(0.001955756451934576)),(to_sfixed_a(0.44483044743537903)),(to_sfixed_a(-0.0002939679252449423)),(to_sfixed_a(-0.00011161647125845775)),(to_sfixed_a(-0.0009833276271820068)),(to_sfixed_a(0.29182106256484985)),(to_sfixed_a(-0.010684012435376644)),(to_sfixed_a(-0.00010821767500601709)),(to_sfixed_a(-0.0054971883073449135)),(to_sfixed_a(-0.02058170922100544)),(to_sfixed_a(0.2598566710948944)),(to_sfixed_a(0.00013660802505910397)),(to_sfixed_a(-0.019657853990793228)),(to_sfixed_a(0.2298518717288971)),(to_sfixed_a(-0.02096925675868988)));

    constant weight_n2_93 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.5257804989814758)),(to_sfixed_a(-0.3866516947746277)),(to_sfixed_a(-0.2897908091545105)),(to_sfixed_a(2.7213405701331794e-05)),(to_sfixed_a(0.004795533139258623)),(to_sfixed_a(0.00013300568389240652)),(to_sfixed_a(-0.00017290376126766205)),(to_sfixed_a(-0.00010251091589452699)),(to_sfixed_a(0.00017925605061464012)),(to_sfixed_a(-1.1249620001763105e-05)),(to_sfixed_a(-0.0001563607802381739)),(to_sfixed_a(-0.36253196001052856)),(to_sfixed_a(-0.005008125212043524)),(to_sfixed_a(-0.0008517430978827178)),(to_sfixed_a(-0.0001712620141915977)),(to_sfixed_a(-7.339069270528853e-05)),(to_sfixed_a(0.47232165932655334)),(to_sfixed_a(-9.391034836880863e-06)),(to_sfixed_a(0.27843037247657776)),(to_sfixed_a(-0.004773790016770363)),(to_sfixed_a(-0.0001573379267938435)),(to_sfixed_a(-0.00042127567576244473)),(to_sfixed_a(-0.0033692484721541405)),(to_sfixed_a(-0.0035351000260561705)),(to_sfixed_a(0.35235217213630676)),(to_sfixed_a(0.012460661120712757)),(to_sfixed_a(-0.0002045372675638646)),(to_sfixed_a(0.18727652728557587)),(to_sfixed_a(0.10187462717294693)),(to_sfixed_a(0.00014744323561899364)),(to_sfixed_a(-0.006101015955209732)),(to_sfixed_a(7.753227691864595e-05)),(to_sfixed_a(0.0013888663379475474)),(to_sfixed_a(-0.0001459817576687783)),(to_sfixed_a(-2.9407263355096802e-05)),(to_sfixed_a(0.00028690171893686056)),(to_sfixed_a(0.22488199174404144)),(to_sfixed_a(0.00047932181041687727)),(to_sfixed_a(0.00421031704172492)),(to_sfixed_a(-7.11856409907341e-06)),(to_sfixed_a(-0.005471029784530401)),(to_sfixed_a(-0.3799852430820465)),(to_sfixed_a(-0.00013889928231947124)),(to_sfixed_a(-0.0001144074703915976)),(to_sfixed_a(-0.007731557358056307)),(to_sfixed_a(-0.0032337915617972612)),(to_sfixed_a(0.005610638298094273)),(to_sfixed_a(0.0004144478007219732)),(to_sfixed_a(0.0003017557319253683)),(to_sfixed_a(0.004573362413793802)),(to_sfixed_a(0.00571855902671814)),(to_sfixed_a(0.004097575321793556)),(to_sfixed_a(-1.0559815564192832e-05)),(to_sfixed_a(0.005105608608573675)),(to_sfixed_a(-0.3910626173019409)),(to_sfixed_a(0.0007942271186038852)),(to_sfixed_a(0.00012017827248200774)),(to_sfixed_a(-0.006369822658598423)),(to_sfixed_a(-1.2094969861209393e-06)),(to_sfixed_a(-0.00020932278130203485)),(to_sfixed_a(-0.008424262516200542)),(to_sfixed_a(-0.006493284832686186)),(to_sfixed_a(-0.0010911053977906704)),(to_sfixed_a(-0.0007263884181156754)),(to_sfixed_a(0.00017892284085974097)),(to_sfixed_a(0.18999066948890686)),(to_sfixed_a(-0.00012184598745079711)),(to_sfixed_a(-0.0004615956568159163)),(to_sfixed_a(0.00265420856885612)),(to_sfixed_a(-1.3497265172190964e-05)),(to_sfixed_a(0.009308628737926483)),(to_sfixed_a(0.0017489709425717592)),(to_sfixed_a(-0.0009529422386549413)),(to_sfixed_a(0.0002978098636958748)),(to_sfixed_a(-1.6593243344686925e-05)),(to_sfixed_a(-6.777464295737445e-05)),(to_sfixed_a(-0.007034063804894686)),(to_sfixed_a(0.13561595976352692)),(to_sfixed_a(0.00031261343974620104)),(to_sfixed_a(-0.7874126434326172)),(to_sfixed_a(-0.008170543238520622)),(to_sfixed_a(-4.648354661185294e-06)),(to_sfixed_a(-0.5343663096427917)),(to_sfixed_a(0.19111645221710205)),(to_sfixed_a(0.00028729200130328536)),(to_sfixed_a(0.25837910175323486)),(to_sfixed_a(-0.01600983552634716)),(to_sfixed_a(-0.00013627453881781548)),(to_sfixed_a(8.915230864658952e-07)),(to_sfixed_a(-0.00010604305134620517)),(to_sfixed_a(-0.0013769996585324407)),(to_sfixed_a(3.046539131901227e-05)),(to_sfixed_a(-0.009826076216995716)),(to_sfixed_a(-8.777817129157484e-06)),(to_sfixed_a(-0.007412903942167759)),(to_sfixed_a(0.00011324984370730817)),(to_sfixed_a(-3.8040452636778355e-05)),(to_sfixed_a(-1.931687438627705e-05)),(to_sfixed_a(0.00022104292293079197)),(to_sfixed_a(6.665242835879326e-05)),(to_sfixed_a(0.00031023117480799556)),(to_sfixed_a(-0.004502346273511648)),(to_sfixed_a(0.000102154393971432)),(to_sfixed_a(-0.25614219903945923)),(to_sfixed_a(0.001535361516289413)),(to_sfixed_a(-0.00017855153419077396)),(to_sfixed_a(-0.00019501637143548578)),(to_sfixed_a(4.45814584963955e-05)),(to_sfixed_a(6.702256359858438e-05)),(to_sfixed_a(0.29153406620025635)),(to_sfixed_a(0.2421385794878006)),(to_sfixed_a(-0.00011575400276342407)),(to_sfixed_a(0.010628716088831425)),(to_sfixed_a(-0.00024751314776949584)),(to_sfixed_a(-4.39267823821865e-05)),(to_sfixed_a(0.003433349309489131)),(to_sfixed_a(-0.41252657771110535)),(to_sfixed_a(-0.0015676890034228563)),(to_sfixed_a(0.00031014042906463146)),(to_sfixed_a(-0.3105895221233368)),(to_sfixed_a(-7.866046507842839e-05)),(to_sfixed_a(6.741679680999368e-05)),(to_sfixed_a(-0.0011580759892240167)),(to_sfixed_a(-0.0001052758889272809)),(to_sfixed_a(-1.3736178516410291e-05)),(to_sfixed_a(0.026163378730416298)),(to_sfixed_a(0.34880828857421875)),(to_sfixed_a(0.00016236874216701835)),(to_sfixed_a(-8.264726056950167e-05)),(to_sfixed_a(-5.4340489441528916e-08)),(to_sfixed_a(-0.0002369149588048458)),(to_sfixed_a(0.00025176815688610077)),(to_sfixed_a(0.005340604577213526)),(to_sfixed_a(0.4118819832801819)),(to_sfixed_a(6.16317629464902e-05)),(to_sfixed_a(0.00016892848361749202)),(to_sfixed_a(-0.007732004392892122)),(to_sfixed_a(-0.00013244316505733877)),(to_sfixed_a(9.610014967620373e-05)),(to_sfixed_a(7.091526640579104e-05)),(to_sfixed_a(0.2922380268573761)),(to_sfixed_a(2.7075679099652916e-05)),(to_sfixed_a(-7.898746116552502e-05)),(to_sfixed_a(1.9703691577888094e-05)),(to_sfixed_a(0.003511507762596011)),(to_sfixed_a(-0.34692490100860596)),(to_sfixed_a(0.0030347334686666727)),(to_sfixed_a(-0.0001823311613406986)),(to_sfixed_a(6.991930422373116e-05)),(to_sfixed_a(-0.11729542165994644)),(to_sfixed_a(0.00017471426690462977)),(to_sfixed_a(0.00012800472904928029)),(to_sfixed_a(-0.0006316156941466033)),(to_sfixed_a(0.0004096670018043369)),(to_sfixed_a(6.417484837584198e-05)),(to_sfixed_a(-0.1754780113697052)),(to_sfixed_a(5.7279394241049886e-06)),(to_sfixed_a(-0.00519245071336627)),(to_sfixed_a(0.0014630926307290792)),(to_sfixed_a(-6.278492219280452e-05)),(to_sfixed_a(-6.610204582102597e-05)),(to_sfixed_a(-0.0002468108432367444)),(to_sfixed_a(-0.2983544170856476)),(to_sfixed_a(0.30135026574134827)),(to_sfixed_a(0.1510189026594162)),(to_sfixed_a(-0.00033852600608952343)),(to_sfixed_a(0.0001529590372228995)),(to_sfixed_a(-0.0003249679575674236)),(to_sfixed_a(2.4974844563985243e-05)),(to_sfixed_a(-2.5549677957314998e-05)),(to_sfixed_a(-0.520470917224884)),(to_sfixed_a(0.006213049404323101)),(to_sfixed_a(0.003174131503328681)),(to_sfixed_a(0.00022190442541614175)),(to_sfixed_a(0.00024700158974155784)),(to_sfixed_a(0.0009559144964441657)),(to_sfixed_a(-0.19571691751480103)),(to_sfixed_a(0.0015804092399775982)),(to_sfixed_a(-0.006029761396348476)),(to_sfixed_a(0.012863462790846825)),(to_sfixed_a(7.444585935445502e-05)),(to_sfixed_a(0.24697059392929077)),(to_sfixed_a(1.983225956792012e-05)),(to_sfixed_a(-3.1286952435038984e-05)),(to_sfixed_a(-0.0002478883252479136)),(to_sfixed_a(-0.00014700759493280202)),(to_sfixed_a(0.3695927560329437)),(to_sfixed_a(0.0027862703427672386)),(to_sfixed_a(0.00159578793682158)),(to_sfixed_a(-0.30704471468925476)),(to_sfixed_a(-0.010789964348077774)),(to_sfixed_a(-0.0003007999330293387)),(to_sfixed_a(0.0017153708031401038)),(to_sfixed_a(-0.008314279839396477)),(to_sfixed_a(-0.00011782596993725747)),(to_sfixed_a(0.00028542557265609503)),(to_sfixed_a(-8.121738210320473e-05)),(to_sfixed_a(0.004610100761055946)),(to_sfixed_a(0.0017998357070609927)),(to_sfixed_a(-0.00012931278615724295)),(to_sfixed_a(-0.00011607789201661944)),(to_sfixed_a(0.00010579406807664782)),(to_sfixed_a(-5.9320904256310314e-05)),(to_sfixed_a(1.2503362086135894e-05)),(to_sfixed_a(6.499716255348176e-05)),(to_sfixed_a(0.008069758303463459)),(to_sfixed_a(-0.000742643722333014)),(to_sfixed_a(0.009916694834828377)),(to_sfixed_a(0.004500677343457937)),(to_sfixed_a(0.00525107653811574)),(to_sfixed_a(-0.008685065433382988)),(to_sfixed_a(4.5698841859120876e-05)),(to_sfixed_a(-0.0001494984026066959)),(to_sfixed_a(-2.1633679352817126e-05)),(to_sfixed_a(-3.5039367503486574e-05)),(to_sfixed_a(-7.647038728464395e-06)),(to_sfixed_a(0.0022600325755774975)),(to_sfixed_a(0.23697082698345184)),(to_sfixed_a(0.45507049560546875)),(to_sfixed_a(0.00019965405226685107)),(to_sfixed_a(-0.00017161763389594853)),(to_sfixed_a(0.00017804827075451612)),(to_sfixed_a(3.705567360157147e-05)),(to_sfixed_a(-0.2534858286380768)),(to_sfixed_a(-0.00960569642484188)),(to_sfixed_a(0.0001068713390850462)),(to_sfixed_a(-8.83068423718214e-06)),(to_sfixed_a(0.00010118785576196387)),(to_sfixed_a(-0.0015725737903267145)),(to_sfixed_a(0.0039015349466353655)),(to_sfixed_a(0.007193674799054861)),(to_sfixed_a(2.0152292563579977e-06)),(to_sfixed_a(0.00042465643491595984)),(to_sfixed_a(2.5217705115210265e-05)),(to_sfixed_a(-0.004672070033848286)),(to_sfixed_a(-0.0028126174584031105)),(to_sfixed_a(-0.0036763837561011314)),(to_sfixed_a(0.00016646756557747722)),(to_sfixed_a(0.0024211006239056587)),(to_sfixed_a(0.00012049678480252624)),(to_sfixed_a(-0.26777583360671997)),(to_sfixed_a(-0.00028847946668975055)),(to_sfixed_a(-0.7529109120368958)),(to_sfixed_a(-0.0002175217668991536)),(to_sfixed_a(0.007576559670269489)),(to_sfixed_a(0.0018040018621832132)),(to_sfixed_a(0.6849409341812134)),(to_sfixed_a(0.0037038768641650677)),(to_sfixed_a(-8.366005204152316e-05)),(to_sfixed_a(-0.006336574908345938)),(to_sfixed_a(-0.006646694149821997)),(to_sfixed_a(0.00018077983986586332)),(to_sfixed_a(-0.5514408946037292)),(to_sfixed_a(-2.3742217308608815e-05)),(to_sfixed_a(0.00013338035205379128)),(to_sfixed_a(-0.20481568574905396)),(to_sfixed_a(-0.2409057766199112)),(to_sfixed_a(0.0001524482504464686)),(to_sfixed_a(0.0002426475693937391)),(to_sfixed_a(0.007357540540397167)),(to_sfixed_a(-1.1889431334566325e-05)),(to_sfixed_a(0.0010588821023702621)),(to_sfixed_a(-5.86573441978544e-05)),(to_sfixed_a(-3.610846761148423e-05)),(to_sfixed_a(7.319540600292385e-05)),(to_sfixed_a(0.3184258043766022)),(to_sfixed_a(-0.00015664324746467173)),(to_sfixed_a(0.00010665251465979964)),(to_sfixed_a(0.00016911982675082982)),(to_sfixed_a(0.010006970725953579)),(to_sfixed_a(0.00044377348967827857)),(to_sfixed_a(-2.849660813808441e-05)),(to_sfixed_a(8.946049638325348e-05)),(to_sfixed_a(-7.038265175651759e-05)),(to_sfixed_a(-2.8917718736920506e-05)),(to_sfixed_a(0.00903488788753748)),(to_sfixed_a(0.007509937044233084)),(to_sfixed_a(-0.24780285358428955)),(to_sfixed_a(0.008198144845664501)),(to_sfixed_a(-0.00013691867934539914)),(to_sfixed_a(-2.2122791051515378e-05)),(to_sfixed_a(-0.00016760558355599642)),(to_sfixed_a(-9.158485772786662e-05)),(to_sfixed_a(0.010727379471063614)),(to_sfixed_a(6.33113959338516e-05)),(to_sfixed_a(0.00019901814812328666)),(to_sfixed_a(-0.00461970642209053)),(to_sfixed_a(0.007837696932256222)),(to_sfixed_a(-0.00011632200767053291)),(to_sfixed_a(-0.004026112612336874)),(to_sfixed_a(0.0014064216520637274)),(to_sfixed_a(0.0025025689974427223)),(to_sfixed_a(0.3409927487373352)),(to_sfixed_a(-0.00028754674713127315)),(to_sfixed_a(0.028280463069677353)),(to_sfixed_a(-0.01553255133330822)),(to_sfixed_a(-0.010718378238379955)),(to_sfixed_a(0.00015288864960893989)),(to_sfixed_a(-0.00233598449267447)),(to_sfixed_a(0.3881088197231293)),(to_sfixed_a(-0.009553481824696064)));

    constant weight_n2_94 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.020030740648508072)),(to_sfixed_a(-0.00014703237684443593)),(to_sfixed_a(-6.368580216076225e-05)),(to_sfixed_a(-0.00016640857211314142)),(to_sfixed_a(-4.6975463192211464e-05)),(to_sfixed_a(1.751716627040878e-05)),(to_sfixed_a(3.9880600525066257e-05)),(to_sfixed_a(-0.0004173459892626852)),(to_sfixed_a(-0.0002502068236935884)),(to_sfixed_a(-8.411530870944262e-06)),(to_sfixed_a(-6.481961463578045e-05)),(to_sfixed_a(-6.726910942234099e-05)),(to_sfixed_a(-0.00013418136222753674)),(to_sfixed_a(9.455416147829965e-05)),(to_sfixed_a(1.1488940799608827e-05)),(to_sfixed_a(-0.00017676420975476503)),(to_sfixed_a(4.852085476159118e-05)),(to_sfixed_a(-0.00029014065512456)),(to_sfixed_a(-0.00013967763516120613)),(to_sfixed_a(0.00015686475671827793)),(to_sfixed_a(0.00012133143900427967)),(to_sfixed_a(-0.00011451276805019006)),(to_sfixed_a(-0.00030033604707568884)),(to_sfixed_a(-0.0001918063499033451)),(to_sfixed_a(2.517008761060424e-05)),(to_sfixed_a(5.69043550058268e-05)),(to_sfixed_a(8.551230712328106e-05)),(to_sfixed_a(-0.0001057506597135216)),(to_sfixed_a(-4.006919334642589e-05)),(to_sfixed_a(-0.00015767847071401775)),(to_sfixed_a(-3.792272036662325e-05)),(to_sfixed_a(-0.00011230187374167144)),(to_sfixed_a(0.00015516339044552296)),(to_sfixed_a(0.00015716953203082085)),(to_sfixed_a(0.00024339236551895738)),(to_sfixed_a(0.0001697381230769679)),(to_sfixed_a(-0.00016516968025825918)),(to_sfixed_a(-0.00024545955238863826)),(to_sfixed_a(-0.00025093590375036)),(to_sfixed_a(6.512930849567056e-05)),(to_sfixed_a(-0.00012980260362382978)),(to_sfixed_a(0.0001174634016933851)),(to_sfixed_a(-0.0002371145092183724)),(to_sfixed_a(0.00018568808445706964)),(to_sfixed_a(-0.00011389357678126544)),(to_sfixed_a(-1.964484908967279e-06)),(to_sfixed_a(6.0464524722192436e-05)),(to_sfixed_a(-0.0004249626072123647)),(to_sfixed_a(-0.00010672252392396331)),(to_sfixed_a(0.00015217791951727122)),(to_sfixed_a(-0.00024030826170928776)),(to_sfixed_a(6.828444020356983e-05)),(to_sfixed_a(0.00013984543329570442)),(to_sfixed_a(-3.145740265608765e-05)),(to_sfixed_a(0.0002910229086410254)),(to_sfixed_a(6.19732090854086e-05)),(to_sfixed_a(-0.00020535514340735972)),(to_sfixed_a(9.165596566163003e-07)),(to_sfixed_a(-3.792455390794203e-05)),(to_sfixed_a(-9.757188672665507e-05)),(to_sfixed_a(-5.976077591185458e-05)),(to_sfixed_a(-1.1980846466030926e-06)),(to_sfixed_a(-5.966343087493442e-05)),(to_sfixed_a(-0.00012972600234206766)),(to_sfixed_a(0.00016952719306573272)),(to_sfixed_a(7.324983016587794e-06)),(to_sfixed_a(1.1612428352236748e-05)),(to_sfixed_a(3.004894097102806e-05)),(to_sfixed_a(9.948023216566071e-05)),(to_sfixed_a(0.00011513286881381646)),(to_sfixed_a(0.00010300169378751889)),(to_sfixed_a(-0.00029407895635813475)),(to_sfixed_a(-0.000206269440241158)),(to_sfixed_a(-0.00023589315242134035)),(to_sfixed_a(-4.494664608500898e-06)),(to_sfixed_a(0.00019007349328603595)),(to_sfixed_a(-6.465284241130576e-05)),(to_sfixed_a(-5.235347634879872e-05)),(to_sfixed_a(-0.00019514450104907155)),(to_sfixed_a(-4.363941843621433e-05)),(to_sfixed_a(9.079311712412164e-05)),(to_sfixed_a(0.00015124156197998673)),(to_sfixed_a(-0.00010099664359586313)),(to_sfixed_a(-0.0003752534685190767)),(to_sfixed_a(0.00010756415576906875)),(to_sfixed_a(6.53169845463708e-05)),(to_sfixed_a(9.388574835611507e-05)),(to_sfixed_a(6.0447466239565983e-05)),(to_sfixed_a(-6.14030723227188e-05)),(to_sfixed_a(-0.00042094034142792225)),(to_sfixed_a(0.00015219561464618891)),(to_sfixed_a(-4.802001058124006e-06)),(to_sfixed_a(0.00030502540175803006)),(to_sfixed_a(-5.65852751606144e-05)),(to_sfixed_a(0.00011718568566720933)),(to_sfixed_a(-7.02358884154819e-05)),(to_sfixed_a(-0.00011602778977248818)),(to_sfixed_a(-0.00020012867753393948)),(to_sfixed_a(0.00016771614900790155)),(to_sfixed_a(-8.827796409605071e-05)),(to_sfixed_a(-3.998626925749704e-05)),(to_sfixed_a(0.0001957825879799202)),(to_sfixed_a(-6.508191290777177e-05)),(to_sfixed_a(-3.6540346627589315e-05)),(to_sfixed_a(-0.00029224948957562447)),(to_sfixed_a(-3.869165084324777e-06)),(to_sfixed_a(2.311680873390287e-05)),(to_sfixed_a(2.2925953089725226e-05)),(to_sfixed_a(-0.00010815741552505642)),(to_sfixed_a(-5.6435950682498515e-05)),(to_sfixed_a(5.528364272322506e-05)),(to_sfixed_a(-0.00018928031204268336)),(to_sfixed_a(-0.00011439424270065501)),(to_sfixed_a(7.470595301128924e-05)),(to_sfixed_a(0.00010110855509992689)),(to_sfixed_a(0.0001165184221463278)),(to_sfixed_a(1.4769975678063929e-05)),(to_sfixed_a(-1.360877649858594e-05)),(to_sfixed_a(-0.00010279950947733596)),(to_sfixed_a(-0.00013536016922444105)),(to_sfixed_a(-3.577665484044701e-05)),(to_sfixed_a(-2.926353772636503e-06)),(to_sfixed_a(3.351743725943379e-05)),(to_sfixed_a(-6.100136670283973e-05)),(to_sfixed_a(-0.0001054998574545607)),(to_sfixed_a(4.33490531577263e-05)),(to_sfixed_a(7.073736196616665e-05)),(to_sfixed_a(1.5715864719823003e-05)),(to_sfixed_a(0.00025126844411715865)),(to_sfixed_a(-9.83606805675663e-05)),(to_sfixed_a(0.000128680287161842)),(to_sfixed_a(-0.000235742365475744)),(to_sfixed_a(0.00025163416285067797)),(to_sfixed_a(-0.00016210752073675394)),(to_sfixed_a(6.060003215679899e-05)),(to_sfixed_a(-6.345389556372538e-05)),(to_sfixed_a(-0.00011346806422807276)),(to_sfixed_a(-0.0001333302352577448)),(to_sfixed_a(6.144179496914148e-05)),(to_sfixed_a(-0.00015391779015772045)),(to_sfixed_a(-3.2547170121688396e-05)),(to_sfixed_a(0.00020045760902576149)),(to_sfixed_a(0.00011387287668185309)),(to_sfixed_a(-0.00013714977831114084)),(to_sfixed_a(-1.169349707197398e-05)),(to_sfixed_a(0.00010511759319342673)),(to_sfixed_a(0.00011325864761602134)),(to_sfixed_a(-0.00019868288654834032)),(to_sfixed_a(-8.170028013410047e-05)),(to_sfixed_a(-3.0411654734052718e-05)),(to_sfixed_a(-5.13727827637922e-05)),(to_sfixed_a(0.0002980113495141268)),(to_sfixed_a(0.0001660371635807678)),(to_sfixed_a(-0.00011570002243388444)),(to_sfixed_a(-2.3650576622458175e-05)),(to_sfixed_a(6.556962034665048e-05)),(to_sfixed_a(1.5666038962081075e-05)),(to_sfixed_a(0.00024753439356572926)),(to_sfixed_a(4.667323082685471e-06)),(to_sfixed_a(-0.0001056630426319316)),(to_sfixed_a(1.2108284863643348e-06)),(to_sfixed_a(7.109773287083954e-05)),(to_sfixed_a(-0.00014971132623031735)),(to_sfixed_a(4.517743946053088e-06)),(to_sfixed_a(7.61107075959444e-05)),(to_sfixed_a(-2.397316347924061e-05)),(to_sfixed_a(7.162563997553661e-05)),(to_sfixed_a(6.651750300079584e-05)),(to_sfixed_a(0.0001128963558585383)),(to_sfixed_a(9.152262646239251e-05)),(to_sfixed_a(2.4451532226521522e-05)),(to_sfixed_a(1.4796154573559761e-05)),(to_sfixed_a(7.106387056410313e-05)),(to_sfixed_a(5.7266159274149686e-05)),(to_sfixed_a(-7.754882972221822e-05)),(to_sfixed_a(0.00024692912120372057)),(to_sfixed_a(-0.00017685539205558598)),(to_sfixed_a(2.626013883855194e-05)),(to_sfixed_a(0.00024028075858950615)),(to_sfixed_a(7.755181286484003e-06)),(to_sfixed_a(5.070287443231791e-07)),(to_sfixed_a(-0.00023066213179845363)),(to_sfixed_a(4.508815982262604e-05)),(to_sfixed_a(2.6827248802874237e-05)),(to_sfixed_a(0.0002956184034701437)),(to_sfixed_a(-1.7713347915560007e-05)),(to_sfixed_a(0.00010028912947745994)),(to_sfixed_a(0.00030460464768111706)),(to_sfixed_a(-3.1379629945149645e-05)),(to_sfixed_a(2.4590892280684784e-05)),(to_sfixed_a(1.1751435522455722e-05)),(to_sfixed_a(-6.413160008378327e-05)),(to_sfixed_a(-6.041665983502753e-05)),(to_sfixed_a(5.684815550921485e-05)),(to_sfixed_a(0.00012986885849386454)),(to_sfixed_a(0.00029337703017517924)),(to_sfixed_a(-1.9824667106149718e-05)),(to_sfixed_a(-6.116293661762029e-06)),(to_sfixed_a(-4.1468272684141994e-05)),(to_sfixed_a(7.040506170596927e-05)),(to_sfixed_a(0.00021102810569573194)),(to_sfixed_a(-0.0001851091510616243)),(to_sfixed_a(4.810336395166814e-05)),(to_sfixed_a(-7.860842015361413e-05)),(to_sfixed_a(8.198731666198e-05)),(to_sfixed_a(-2.2861797333462164e-05)),(to_sfixed_a(-0.00027985236374661326)),(to_sfixed_a(7.097044726833701e-05)),(to_sfixed_a(-2.809134457493201e-05)),(to_sfixed_a(-0.000181529248948209)),(to_sfixed_a(3.038993600057438e-05)),(to_sfixed_a(-9.348544699605554e-05)),(to_sfixed_a(-0.0003175794845446944)),(to_sfixed_a(0.00015414085646625608)),(to_sfixed_a(6.367434980347753e-05)),(to_sfixed_a(-0.00021830963669344783)),(to_sfixed_a(-0.00040985405212268233)),(to_sfixed_a(-0.00020634123939089477)),(to_sfixed_a(0.000182771313120611)),(to_sfixed_a(-0.0002058512473013252)),(to_sfixed_a(-0.0003101033216807991)),(to_sfixed_a(-6.92307876306586e-05)),(to_sfixed_a(-7.080016075633466e-05)),(to_sfixed_a(-7.18779192538932e-05)),(to_sfixed_a(-2.438969022477977e-05)),(to_sfixed_a(-0.0002861459506675601)),(to_sfixed_a(-0.0001169554961961694)),(to_sfixed_a(-2.6766509108711034e-05)),(to_sfixed_a(-0.00016602297546342015)),(to_sfixed_a(-6.601722998311743e-05)),(to_sfixed_a(2.048273745458573e-05)),(to_sfixed_a(0.00022491900017485023)),(to_sfixed_a(0.00023710561799816787)),(to_sfixed_a(-0.00013936249888502061)),(to_sfixed_a(-0.000154849563841708)),(to_sfixed_a(0.0002830150770023465)),(to_sfixed_a(-2.3736465664114803e-06)),(to_sfixed_a(-0.0004597283841576427)),(to_sfixed_a(8.609956421423703e-05)),(to_sfixed_a(2.203903568442911e-05)),(to_sfixed_a(4.089944195584394e-05)),(to_sfixed_a(0.00017353170551359653)),(to_sfixed_a(0.00021381370606832206)),(to_sfixed_a(-0.00012845141463913023)),(to_sfixed_a(-4.4748481741407886e-05)),(to_sfixed_a(3.680880035972223e-05)),(to_sfixed_a(-0.0001564351696288213)),(to_sfixed_a(-0.00016672458150424063)),(to_sfixed_a(-4.2324463720433414e-05)),(to_sfixed_a(-8.63818422658369e-06)),(to_sfixed_a(6.184927769936621e-07)),(to_sfixed_a(-0.00011243623885093257)),(to_sfixed_a(0.0001502603990957141)),(to_sfixed_a(-0.00016716946265660226)),(to_sfixed_a(-3.067013676627539e-05)),(to_sfixed_a(3.716530045494437e-05)),(to_sfixed_a(-1.0609001037664711e-05)),(to_sfixed_a(-0.00014303573698271066)),(to_sfixed_a(-0.00015762312978040427)),(to_sfixed_a(-4.717170668300241e-05)),(to_sfixed_a(0.00011366192484274507)),(to_sfixed_a(1.3313139788806438e-05)),(to_sfixed_a(1.605191209819168e-05)),(to_sfixed_a(8.588706259615719e-05)),(to_sfixed_a(-8.85532790562138e-06)),(to_sfixed_a(-7.08811276126653e-05)),(to_sfixed_a(4.523291136138141e-05)),(to_sfixed_a(-0.00011696379806380719)),(to_sfixed_a(6.9086738221813e-05)),(to_sfixed_a(0.00010137547360500321)),(to_sfixed_a(-1.567357685416937e-05)),(to_sfixed_a(-0.00013776813284493983)),(to_sfixed_a(-0.00018272419401910156)),(to_sfixed_a(0.0003147335664834827)),(to_sfixed_a(-8.04442897788249e-05)),(to_sfixed_a(8.494086068822071e-05)),(to_sfixed_a(-1.994924241444096e-05)),(to_sfixed_a(3.4747619793051854e-05)),(to_sfixed_a(-0.00011600787547649816)),(to_sfixed_a(0.00045222806511446834)),(to_sfixed_a(-2.9416813049465418e-05)),(to_sfixed_a(-4.988090950064361e-06)),(to_sfixed_a(-0.00018155438010580838)),(to_sfixed_a(-0.00019895390141755342)),(to_sfixed_a(-6.208203558344394e-06)),(to_sfixed_a(4.390785761643201e-07)),(to_sfixed_a(-0.00012890752987004817)),(to_sfixed_a(0.00021199806360527873)),(to_sfixed_a(0.00015152685227803886)),(to_sfixed_a(-4.982008249498904e-06)),(to_sfixed_a(2.1903157175984234e-05)),(to_sfixed_a(9.258438512915745e-05)),(to_sfixed_a(-2.709958062041551e-05)),(to_sfixed_a(0.00010766653576865792)),(to_sfixed_a(0.00019646289001684636)),(to_sfixed_a(9.587978638592176e-06)),(to_sfixed_a(0.00011950186308240518)),(to_sfixed_a(0.00010216756345471367)),(to_sfixed_a(4.301800800021738e-07)),(to_sfixed_a(1.4499164535664022e-08)),(to_sfixed_a(5.505557055585086e-06)));

    constant weight_n2_95 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.04632433503866196)),(to_sfixed_a(0.0006353548378683627)),(to_sfixed_a(0.3880881369113922)),(to_sfixed_a(-0.00030203373171389103)),(to_sfixed_a(-0.01019266340881586)),(to_sfixed_a(-4.820066169486381e-05)),(to_sfixed_a(0.004613249562680721)),(to_sfixed_a(-0.00021931160881649703)),(to_sfixed_a(6.060211671865545e-05)),(to_sfixed_a(-2.4501874577254057e-05)),(to_sfixed_a(0.00010644969734130427)),(to_sfixed_a(0.0017318606842309237)),(to_sfixed_a(0.003927523735910654)),(to_sfixed_a(7.33745691832155e-05)),(to_sfixed_a(-6.512526306323707e-05)),(to_sfixed_a(3.796961027546786e-05)),(to_sfixed_a(0.03184691444039345)),(to_sfixed_a(0.00010176482464885339)),(to_sfixed_a(-0.003811583621427417)),(to_sfixed_a(-0.001797133474610746)),(to_sfixed_a(0.00017862836830317974)),(to_sfixed_a(-2.5016910512931645e-05)),(to_sfixed_a(-1.738269565976225e-05)),(to_sfixed_a(0.0010364447953179479)),(to_sfixed_a(0.002871548291295767)),(to_sfixed_a(0.0036296546459198)),(to_sfixed_a(-6.837381079094484e-07)),(to_sfixed_a(-0.00042310310527682304)),(to_sfixed_a(-0.00735895149409771)),(to_sfixed_a(5.0783804908860475e-05)),(to_sfixed_a(0.006036385428160429)),(to_sfixed_a(3.636713881860487e-05)),(to_sfixed_a(-0.0030394101049751043)),(to_sfixed_a(-3.8107638829387724e-05)),(to_sfixed_a(-0.00010257362009724602)),(to_sfixed_a(-0.00022861828620079905)),(to_sfixed_a(0.008018900640308857)),(to_sfixed_a(0.29327043890953064)),(to_sfixed_a(0.005157288163900375)),(to_sfixed_a(-6.572566780960187e-05)),(to_sfixed_a(0.03190529718995094)),(to_sfixed_a(0.001323952223174274)),(to_sfixed_a(5.886147846467793e-06)),(to_sfixed_a(6.740017852280289e-05)),(to_sfixed_a(0.0009125579963438213)),(to_sfixed_a(-0.0073093813844025135)),(to_sfixed_a(0.0011472089681774378)),(to_sfixed_a(-0.005115285981446505)),(to_sfixed_a(0.0002197780559072271)),(to_sfixed_a(0.0005819867947138846)),(to_sfixed_a(0.0033519468270242214)),(to_sfixed_a(-0.0002948118490166962)),(to_sfixed_a(1.996922947000712e-06)),(to_sfixed_a(0.0003388980112504214)),(to_sfixed_a(0.28727203607559204)),(to_sfixed_a(-0.002144369063898921)),(to_sfixed_a(0.00011317322787363082)),(to_sfixed_a(0.0017329882830381393)),(to_sfixed_a(0.0001538298383820802)),(to_sfixed_a(-0.00013839606253895909)),(to_sfixed_a(-0.0011493598576635122)),(to_sfixed_a(-0.00040264983545057476)),(to_sfixed_a(-0.002162666991353035)),(to_sfixed_a(0.011469938792288303)),(to_sfixed_a(-0.00021790768369100988)),(to_sfixed_a(0.0011763276997953653)),(to_sfixed_a(-0.000453800312243402)),(to_sfixed_a(-0.49199527502059937)),(to_sfixed_a(-0.002838714048266411)),(to_sfixed_a(-0.00010637619561748579)),(to_sfixed_a(-0.0029906234703958035)),(to_sfixed_a(-0.5380804538726807)),(to_sfixed_a(0.012501358985900879)),(to_sfixed_a(1.1053045454900712e-05)),(to_sfixed_a(3.0217706807889044e-06)),(to_sfixed_a(0.00021039272542111576)),(to_sfixed_a(0.0019746345933526754)),(to_sfixed_a(0.001921534538269043)),(to_sfixed_a(2.3552376660518348e-05)),(to_sfixed_a(0.40482035279273987)),(to_sfixed_a(-0.1859021633863449)),(to_sfixed_a(-0.000151242216816172)),(to_sfixed_a(-0.001701264176517725)),(to_sfixed_a(0.001812923583202064)),(to_sfixed_a(-1.9331127987243235e-07)),(to_sfixed_a(0.0032722260802984238)),(to_sfixed_a(0.0021332930773496628)),(to_sfixed_a(9.529110684525222e-05)),(to_sfixed_a(0.00016085982497315854)),(to_sfixed_a(6.787209713365883e-05)),(to_sfixed_a(-0.48418116569519043)),(to_sfixed_a(-7.135961641324684e-05)),(to_sfixed_a(0.0009784927824512124)),(to_sfixed_a(9.800789848668501e-05)),(to_sfixed_a(-0.0026105036959052086)),(to_sfixed_a(1.0569141522864811e-05)),(to_sfixed_a(-0.00011748667748179287)),(to_sfixed_a(-6.397283868864179e-06)),(to_sfixed_a(0.0001272518711630255)),(to_sfixed_a(-1.6480538761243224e-05)),(to_sfixed_a(0.0031627642456442118)),(to_sfixed_a(0.0004566196585074067)),(to_sfixed_a(-2.3428066924680024e-05)),(to_sfixed_a(0.30094361305236816)),(to_sfixed_a(0.004012723453342915)),(to_sfixed_a(0.0015025349566712976)),(to_sfixed_a(-1.1221709428355098e-06)),(to_sfixed_a(2.5221197574865073e-06)),(to_sfixed_a(-3.5354478313820437e-05)),(to_sfixed_a(0.002308688359335065)),(to_sfixed_a(-0.0005707534728571773)),(to_sfixed_a(9.511118696536869e-05)),(to_sfixed_a(-0.004322139546275139)),(to_sfixed_a(0.00016811152454465628)),(to_sfixed_a(2.6684370823204517e-05)),(to_sfixed_a(0.00014189540524967015)),(to_sfixed_a(0.3244370222091675)),(to_sfixed_a(-0.00018209079280495644)),(to_sfixed_a(3.653497697087005e-05)),(to_sfixed_a(0.3011033535003662)),(to_sfixed_a(4.733301466330886e-06)),(to_sfixed_a(-1.3484292139764875e-05)),(to_sfixed_a(-0.006910794880241156)),(to_sfixed_a(0.00011197808635188267)),(to_sfixed_a(6.222003139555454e-05)),(to_sfixed_a(0.3380853831768036)),(to_sfixed_a(-0.001533702714368701)),(to_sfixed_a(4.5100961870048195e-05)),(to_sfixed_a(-0.00023119806428439915)),(to_sfixed_a(3.30436960211955e-05)),(to_sfixed_a(-7.445917435688898e-05)),(to_sfixed_a(0.00013099139323458076)),(to_sfixed_a(0.00014075872604735196)),(to_sfixed_a(0.005150269716978073)),(to_sfixed_a(0.00017654418479651213)),(to_sfixed_a(9.356135706184432e-05)),(to_sfixed_a(0.21010355651378632)),(to_sfixed_a(-0.00013611276517622173)),(to_sfixed_a(0.00011326602543704212)),(to_sfixed_a(-0.00011922864359803498)),(to_sfixed_a(-0.240640789270401)),(to_sfixed_a(-0.00013582114479504526)),(to_sfixed_a(-0.00011179152352269739)),(to_sfixed_a(0.00012179023906355724)),(to_sfixed_a(0.0001785849017323926)),(to_sfixed_a(-0.0049444399774074554)),(to_sfixed_a(-0.002474412089213729)),(to_sfixed_a(6.751900218660012e-05)),(to_sfixed_a(0.0002512522623874247)),(to_sfixed_a(0.003806786611676216)),(to_sfixed_a(3.041571835638024e-05)),(to_sfixed_a(-3.6365458072395995e-05)),(to_sfixed_a(-0.0021268874406814575)),(to_sfixed_a(6.0052982007618994e-05)),(to_sfixed_a(0.00016782332386355847)),(to_sfixed_a(0.019383404403924942)),(to_sfixed_a(-4.412533598951995e-06)),(to_sfixed_a(-0.0031338229309767485)),(to_sfixed_a(-0.0001879239862319082)),(to_sfixed_a(-0.00015678089403081685)),(to_sfixed_a(2.7204347134102136e-05)),(to_sfixed_a(-0.00010612082405714318)),(to_sfixed_a(0.0013496222672984004)),(to_sfixed_a(-0.0005772352451458573)),(to_sfixed_a(0.004261308815330267)),(to_sfixed_a(0.0060316091403365135)),(to_sfixed_a(6.480466981884092e-05)),(to_sfixed_a(-0.005848037078976631)),(to_sfixed_a(-9.368237806484103e-05)),(to_sfixed_a(-0.00010337789717596024)),(to_sfixed_a(0.2564460039138794)),(to_sfixed_a(0.00030200337641872466)),(to_sfixed_a(0.006798254791647196)),(to_sfixed_a(-5.7465302234049886e-05)),(to_sfixed_a(0.4098411500453949)),(to_sfixed_a(0.002094342140480876)),(to_sfixed_a(0.00045418483205139637)),(to_sfixed_a(-0.008918684907257557)),(to_sfixed_a(0.15770591795444489)),(to_sfixed_a(-0.40232041478157043)),(to_sfixed_a(-0.001080062473192811)),(to_sfixed_a(0.00348276156000793)),(to_sfixed_a(2.3664877517148852e-05)),(to_sfixed_a(2.9786897357553244e-06)),(to_sfixed_a(-0.00024169062089640647)),(to_sfixed_a(0.007368938066065311)),(to_sfixed_a(-0.002320545958355069)),(to_sfixed_a(-0.0008600849541835487)),(to_sfixed_a(3.26475128531456e-06)),(to_sfixed_a(0.0005997074767947197)),(to_sfixed_a(0.1849922090768814)),(to_sfixed_a(-4.6772176574449986e-05)),(to_sfixed_a(0.5233888030052185)),(to_sfixed_a(-0.00593539047986269)),(to_sfixed_a(7.451781129930168e-06)),(to_sfixed_a(-0.000533487182110548)),(to_sfixed_a(-0.00011383432138245553)),(to_sfixed_a(0.002588193165138364)),(to_sfixed_a(0.00835387036204338)),(to_sfixed_a(-0.00031270916224457324)),(to_sfixed_a(1.4931814803276211e-05)),(to_sfixed_a(-0.00014869323058519512)),(to_sfixed_a(-0.00017736965673975646)),(to_sfixed_a(-0.000221622409299016)),(to_sfixed_a(0.00018418159743305296)),(to_sfixed_a(0.00018725424888543785)),(to_sfixed_a(0.004557267762720585)),(to_sfixed_a(-0.0923897922039032)),(to_sfixed_a(-0.0009352302295155823)),(to_sfixed_a(-0.00790572538971901)),(to_sfixed_a(-0.3651418387889862)),(to_sfixed_a(6.719466182403266e-05)),(to_sfixed_a(0.00016832599067129195)),(to_sfixed_a(-5.168270581634715e-05)),(to_sfixed_a(-1.280612195841968e-06)),(to_sfixed_a(-0.0001687262556515634)),(to_sfixed_a(-0.011506851762533188)),(to_sfixed_a(0.0013725265162065625)),(to_sfixed_a(-0.01691386103630066)),(to_sfixed_a(0.0004518437199294567)),(to_sfixed_a(-0.0003826524189207703)),(to_sfixed_a(-6.890633812872693e-05)),(to_sfixed_a(-2.734655572567135e-05)),(to_sfixed_a(1.0370898962719366e-05)),(to_sfixed_a(0.00018746723071672022)),(to_sfixed_a(-0.00011412690219003707)),(to_sfixed_a(5.3212716011330485e-06)),(to_sfixed_a(7.001826452324167e-05)),(to_sfixed_a(0.00593594228848815)),(to_sfixed_a(0.0005369822029024363)),(to_sfixed_a(-0.21839295327663422)),(to_sfixed_a(-0.00018260163778904825)),(to_sfixed_a(-0.0004152712062932551)),(to_sfixed_a(-5.77215978410095e-05)),(to_sfixed_a(0.001423488138243556)),(to_sfixed_a(-0.007733053993433714)),(to_sfixed_a(0.005906557664275169)),(to_sfixed_a(4.489615821512416e-05)),(to_sfixed_a(0.00017936389485839754)),(to_sfixed_a(-0.00020011948072351515)),(to_sfixed_a(0.0008926004520617425)),(to_sfixed_a(0.0002799434296321124)),(to_sfixed_a(-0.005067511927336454)),(to_sfixed_a(5.870847962796688e-05)),(to_sfixed_a(0.4397049844264984)),(to_sfixed_a(-0.0018559558084234595)),(to_sfixed_a(-0.4380561411380768)),(to_sfixed_a(-0.011193177662789822)),(to_sfixed_a(3.855426621157676e-05)),(to_sfixed_a(0.003999421838670969)),(to_sfixed_a(0.01384802907705307)),(to_sfixed_a(6.158334144856781e-05)),(to_sfixed_a(0.3923236131668091)),(to_sfixed_a(-0.00013887640670873225)),(to_sfixed_a(-0.015420207753777504)),(to_sfixed_a(-0.014421642757952213)),(to_sfixed_a(0.0003807164030149579)),(to_sfixed_a(-0.00018029191414825618)),(to_sfixed_a(0.00017578070401214063)),(to_sfixed_a(-0.006532966159284115)),(to_sfixed_a(6.508415390271693e-05)),(to_sfixed_a(0.00039522111183032393)),(to_sfixed_a(-0.00031366702751256526)),(to_sfixed_a(1.7903003026731312e-06)),(to_sfixed_a(7.610696775373071e-05)),(to_sfixed_a(0.33254292607307434)),(to_sfixed_a(-6.90935121383518e-05)),(to_sfixed_a(0.00020546818268485367)),(to_sfixed_a(0.00023790134582668543)),(to_sfixed_a(0.001153241260908544)),(to_sfixed_a(0.006672809366136789)),(to_sfixed_a(0.00016715309175197035)),(to_sfixed_a(-7.043643563520163e-06)),(to_sfixed_a(-0.0001011730419122614)),(to_sfixed_a(0.00011459951929282397)),(to_sfixed_a(-0.002699541626498103)),(to_sfixed_a(-0.0007959427312016487)),(to_sfixed_a(0.004000375978648663)),(to_sfixed_a(-0.5321429967880249)),(to_sfixed_a(0.002773334039375186)),(to_sfixed_a(-7.348656072281301e-05)),(to_sfixed_a(0.00020473661425057799)),(to_sfixed_a(0.0002032347401836887)),(to_sfixed_a(0.0005471167387440801)),(to_sfixed_a(-5.822141974931583e-05)),(to_sfixed_a(0.00028688344173133373)),(to_sfixed_a(0.00010062273941002786)),(to_sfixed_a(-0.0036994097754359245)),(to_sfixed_a(-6.016221232130192e-05)),(to_sfixed_a(-0.5294000506401062)),(to_sfixed_a(-0.0012164554791525006)),(to_sfixed_a(0.00785957183688879)),(to_sfixed_a(-0.34181293845176697)),(to_sfixed_a(-0.00024582818150520325)),(to_sfixed_a(-0.003328859806060791)),(to_sfixed_a(0.40912482142448425)),(to_sfixed_a(0.008162355981767178)),(to_sfixed_a(0.0002157991984859109)),(to_sfixed_a(0.0013820405583828688)),(to_sfixed_a(-0.0025060568004846573)),(to_sfixed_a(0.007513978984206915)));

    constant weight_n2_96 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.1269640028476715)),(to_sfixed_a(-0.0008691004477441311)),(to_sfixed_a(0.2095245122909546)),(to_sfixed_a(-2.3429369321092963e-05)),(to_sfixed_a(-0.19574543833732605)),(to_sfixed_a(-4.118899232707918e-05)),(to_sfixed_a(0.01294793002307415)),(to_sfixed_a(-0.0003005112521350384)),(to_sfixed_a(7.647647726116702e-05)),(to_sfixed_a(0.00014005295815877616)),(to_sfixed_a(-6.430079520214349e-05)),(to_sfixed_a(0.06105672940611839)),(to_sfixed_a(0.009795697405934334)),(to_sfixed_a(-0.00017780790221877396)),(to_sfixed_a(0.00010882067726925015)),(to_sfixed_a(1.0291238140780479e-05)),(to_sfixed_a(-0.0009211471187882125)),(to_sfixed_a(-0.00044726365013048053)),(to_sfixed_a(-0.4555032551288605)),(to_sfixed_a(-8.159592834999785e-05)),(to_sfixed_a(0.00010589725570753217)),(to_sfixed_a(8.203278412111104e-06)),(to_sfixed_a(8.640492160338908e-05)),(to_sfixed_a(0.0744323581457138)),(to_sfixed_a(-0.0025852653197944164)),(to_sfixed_a(0.0019164530094712973)),(to_sfixed_a(0.0003214685129933059)),(to_sfixed_a(0.1023188903927803)),(to_sfixed_a(0.0005332690780051053)),(to_sfixed_a(-0.00016872171545401216)),(to_sfixed_a(-0.010995850898325443)),(to_sfixed_a(6.458334610215388e-06)),(to_sfixed_a(-0.006233438849449158)),(to_sfixed_a(-0.00011403219832573086)),(to_sfixed_a(-7.185875438153744e-05)),(to_sfixed_a(0.0003925918717868626)),(to_sfixed_a(-1.0572218894958496)),(to_sfixed_a(0.08647645264863968)),(to_sfixed_a(-0.4932961165904999)),(to_sfixed_a(-3.0609411624027416e-05)),(to_sfixed_a(-0.002913586562499404)),(to_sfixed_a(0.0011411102022975683)),(to_sfixed_a(-4.279008862795308e-06)),(to_sfixed_a(-9.588722605258226e-06)),(to_sfixed_a(0.004769360180944204)),(to_sfixed_a(-0.004113327711820602)),(to_sfixed_a(0.029139328747987747)),(to_sfixed_a(0.005938924849033356)),(to_sfixed_a(-4.348775837570429e-05)),(to_sfixed_a(0.0023572572972625494)),(to_sfixed_a(0.008003546856343746)),(to_sfixed_a(-0.0004741643206216395)),(to_sfixed_a(-3.804672451224178e-05)),(to_sfixed_a(-0.001808962901122868)),(to_sfixed_a(-0.002646662527695298)),(to_sfixed_a(-0.3763596713542938)),(to_sfixed_a(-0.0001598045346327126)),(to_sfixed_a(-0.008147209882736206)),(to_sfixed_a(-0.00015001953579485416)),(to_sfixed_a(6.983135244809091e-05)),(to_sfixed_a(0.010700583457946777)),(to_sfixed_a(-0.0011103819124400616)),(to_sfixed_a(-0.06511241942644119)),(to_sfixed_a(-0.001468468690291047)),(to_sfixed_a(2.973462687805295e-05)),(to_sfixed_a(-0.06068139895796776)),(to_sfixed_a(0.0002487747115083039)),(to_sfixed_a(-0.3563235402107239)),(to_sfixed_a(-0.000705558923073113)),(to_sfixed_a(-2.639374724822119e-05)),(to_sfixed_a(-0.01783393695950508)),(to_sfixed_a(0.5754032135009766)),(to_sfixed_a(0.0018188898684456944)),(to_sfixed_a(-5.261710612103343e-06)),(to_sfixed_a(-1.1613778042374179e-05)),(to_sfixed_a(-6.03022999712266e-05)),(to_sfixed_a(0.18971893191337585)),(to_sfixed_a(-0.007204144261777401)),(to_sfixed_a(-3.244755498599261e-05)),(to_sfixed_a(-0.002805443713441491)),(to_sfixed_a(0.010330883786082268)),(to_sfixed_a(-0.00014621097943745553)),(to_sfixed_a(-0.006279889494180679)),(to_sfixed_a(-0.3792998790740967)),(to_sfixed_a(-0.0003107674128841609)),(to_sfixed_a(0.18415427207946777)),(to_sfixed_a(-0.0014041434042155743)),(to_sfixed_a(-0.0038977533113211393)),(to_sfixed_a(0.0002231755934190005)),(to_sfixed_a(-1.9727303879335523e-06)),(to_sfixed_a(-0.35189393162727356)),(to_sfixed_a(5.667285586241633e-05)),(to_sfixed_a(-0.002414656337350607)),(to_sfixed_a(-9.776801016414538e-05)),(to_sfixed_a(-0.3726077377796173)),(to_sfixed_a(-4.442358113010414e-05)),(to_sfixed_a(2.5150318833766505e-05)),(to_sfixed_a(-1.6482626961078495e-06)),(to_sfixed_a(-0.00010837958689080551)),(to_sfixed_a(-0.0002810733567457646)),(to_sfixed_a(-0.00380337075330317)),(to_sfixed_a(0.15094716846942902)),(to_sfixed_a(-0.00021456333342939615)),(to_sfixed_a(-0.0013718587579205632)),(to_sfixed_a(-0.593654215335846)),(to_sfixed_a(0.002035564510151744)),(to_sfixed_a(0.00011541548883542418)),(to_sfixed_a(7.00065866112709e-05)),(to_sfixed_a(-1.806571162887849e-05)),(to_sfixed_a(0.19040986895561218)),(to_sfixed_a(0.1997632533311844)),(to_sfixed_a(-1.6357240383513272e-05)),(to_sfixed_a(-0.003715686034411192)),(to_sfixed_a(0.00024674879387021065)),(to_sfixed_a(-0.000380326877348125)),(to_sfixed_a(-0.24120433628559113)),(to_sfixed_a(-0.014555469155311584)),(to_sfixed_a(-0.06395798176527023)),(to_sfixed_a(0.00012068379146512598)),(to_sfixed_a(0.00034444211632944643)),(to_sfixed_a(-0.00025139315403066576)),(to_sfixed_a(2.216904249507934e-06)),(to_sfixed_a(0.0024037440307438374)),(to_sfixed_a(1.4604360330849886e-05)),(to_sfixed_a(4.7678695409558713e-05)),(to_sfixed_a(0.0005188114591874182)),(to_sfixed_a(-0.013566287234425545)),(to_sfixed_a(-0.0002919763792306185)),(to_sfixed_a(-0.00028907356318086386)),(to_sfixed_a(-1.6700134437996894e-05)),(to_sfixed_a(7.251478382386267e-05)),(to_sfixed_a(0.0002320755593245849)),(to_sfixed_a(-0.004202817101031542)),(to_sfixed_a(0.3507038354873657)),(to_sfixed_a(0.00010758775897556916)),(to_sfixed_a(-7.865873340051621e-05)),(to_sfixed_a(0.30823859572410583)),(to_sfixed_a(0.4104311466217041)),(to_sfixed_a(-4.258429544279352e-05)),(to_sfixed_a(0.00020438572391867638)),(to_sfixed_a(-0.008918507024645805)),(to_sfixed_a(0.00015679288480896503)),(to_sfixed_a(-0.00011717986490111798)),(to_sfixed_a(-0.00033377506770193577)),(to_sfixed_a(-0.00013092928566038609)),(to_sfixed_a(0.2883898913860321)),(to_sfixed_a(-0.0003791067865677178)),(to_sfixed_a(0.00026289306697435677)),(to_sfixed_a(-0.00015431178326252848)),(to_sfixed_a(-0.13538412749767303)),(to_sfixed_a(7.544289837824181e-05)),(to_sfixed_a(1.7926955479197204e-05)),(to_sfixed_a(-0.013437798246741295)),(to_sfixed_a(5.274283466860652e-06)),(to_sfixed_a(3.8917845813557506e-05)),(to_sfixed_a(-0.0030563261825591326)),(to_sfixed_a(-5.872057954547927e-05)),(to_sfixed_a(-0.0031894503626972437)),(to_sfixed_a(-9.057395800482482e-06)),(to_sfixed_a(2.4105665943352506e-05)),(to_sfixed_a(-6.063360342523083e-05)),(to_sfixed_a(-8.685209468239918e-05)),(to_sfixed_a(0.07201363891363144)),(to_sfixed_a(-0.002969966270029545)),(to_sfixed_a(-0.010248418897390366)),(to_sfixed_a(-0.0024859467521309853)),(to_sfixed_a(-0.0001759752631187439)),(to_sfixed_a(0.022680852562189102)),(to_sfixed_a(0.00018154791905544698)),(to_sfixed_a(0.00011544025619514287)),(to_sfixed_a(0.11796707659959793)),(to_sfixed_a(-0.001987300580367446)),(to_sfixed_a(-0.00424979766830802)),(to_sfixed_a(5.434994818642735e-07)),(to_sfixed_a(0.35648491978645325)),(to_sfixed_a(-0.0037438683211803436)),(to_sfixed_a(0.008944250643253326)),(to_sfixed_a(0.017645521089434624)),(to_sfixed_a(0.21271061897277832)),(to_sfixed_a(0.4040180742740631)),(to_sfixed_a(-0.008630623109638691)),(to_sfixed_a(-0.27399304509162903)),(to_sfixed_a(0.00018252336303703487)),(to_sfixed_a(-4.299741704016924e-06)),(to_sfixed_a(9.03769068827387e-06)),(to_sfixed_a(-0.4777281880378723)),(to_sfixed_a(-0.0004893475561402738)),(to_sfixed_a(-0.42518535256385803)),(to_sfixed_a(6.429164932342246e-05)),(to_sfixed_a(0.0025207537692040205)),(to_sfixed_a(0.3943055272102356)),(to_sfixed_a(6.697175558656454e-05)),(to_sfixed_a(-0.025192683562636375)),(to_sfixed_a(0.33799201250076294)),(to_sfixed_a(-2.5802815798670053e-05)),(to_sfixed_a(0.00698309950530529)),(to_sfixed_a(6.823881267337129e-05)),(to_sfixed_a(-0.009549528360366821)),(to_sfixed_a(0.01592940092086792)),(to_sfixed_a(8.462867845082656e-05)),(to_sfixed_a(-7.066330726956949e-05)),(to_sfixed_a(2.930601840489544e-05)),(to_sfixed_a(-0.00018552366236690432)),(to_sfixed_a(0.00013332493836060166)),(to_sfixed_a(0.00016664368740748614)),(to_sfixed_a(0.0017090887995436788)),(to_sfixed_a(0.0046833232045173645)),(to_sfixed_a(0.13123756647109985)),(to_sfixed_a(0.32468003034591675)),(to_sfixed_a(-0.0029588735196739435)),(to_sfixed_a(-0.31287527084350586)),(to_sfixed_a(-0.0002251764526590705)),(to_sfixed_a(0.00021791565814055502)),(to_sfixed_a(-6.292561010923237e-05)),(to_sfixed_a(8.371614967472851e-05)),(to_sfixed_a(1.0732037480920553e-08)),(to_sfixed_a(-0.017980726435780525)),(to_sfixed_a(0.004593249410390854)),(to_sfixed_a(-3.228618879802525e-05)),(to_sfixed_a(0.00013851301628164947)),(to_sfixed_a(-0.0002358277270104736)),(to_sfixed_a(-0.0001369862729916349)),(to_sfixed_a(0.00020504550775513053)),(to_sfixed_a(0.0004441722412593663)),(to_sfixed_a(0.28936949372291565)),(to_sfixed_a(6.235175533220172e-05)),(to_sfixed_a(3.1276431400328875e-05)),(to_sfixed_a(-6.865625618956983e-05)),(to_sfixed_a(0.19184543192386627)),(to_sfixed_a(0.4065763056278229)),(to_sfixed_a(-0.0004929401911795139)),(to_sfixed_a(-0.00013389963714871556)),(to_sfixed_a(-0.0001262175792362541)),(to_sfixed_a(-3.9584701880812645e-06)),(to_sfixed_a(-0.011854632757604122)),(to_sfixed_a(-0.019722292199730873)),(to_sfixed_a(0.005423021502792835)),(to_sfixed_a(-0.00012668329873122275)),(to_sfixed_a(0.004940680228173733)),(to_sfixed_a(8.967149187810719e-05)),(to_sfixed_a(-0.007224951405078173)),(to_sfixed_a(-1.5690835425630212e-05)),(to_sfixed_a(-0.01255420409142971)),(to_sfixed_a(-0.00011341279605403543)),(to_sfixed_a(0.13124725222587585)),(to_sfixed_a(-0.008950300514698029)),(to_sfixed_a(0.31506839394569397)),(to_sfixed_a(0.00450383685529232)),(to_sfixed_a(6.946859502932057e-05)),(to_sfixed_a(-0.06514324992895126)),(to_sfixed_a(0.003360247705131769)),(to_sfixed_a(3.934848791686818e-05)),(to_sfixed_a(-0.0014376959297806025)),(to_sfixed_a(-0.00022836732387077063)),(to_sfixed_a(-0.006278630346059799)),(to_sfixed_a(0.26472434401512146)),(to_sfixed_a(0.30296558141708374)),(to_sfixed_a(0.00013689493061974645)),(to_sfixed_a(2.9212591471150517e-05)),(to_sfixed_a(-0.1916414052248001)),(to_sfixed_a(0.00015288364375010133)),(to_sfixed_a(-0.012800437398254871)),(to_sfixed_a(6.534568819915876e-05)),(to_sfixed_a(-0.0009456605766899884)),(to_sfixed_a(7.555981574114412e-05)),(to_sfixed_a(-0.010560081340372562)),(to_sfixed_a(7.576542702736333e-05)),(to_sfixed_a(-0.0003111058322247118)),(to_sfixed_a(-1.038773189065978e-05)),(to_sfixed_a(-0.008210064843297005)),(to_sfixed_a(0.0061768763698637486)),(to_sfixed_a(5.9775818954221904e-05)),(to_sfixed_a(-8.030520984902978e-05)),(to_sfixed_a(0.0002943958679679781)),(to_sfixed_a(3.164755253237672e-05)),(to_sfixed_a(-0.31183314323425293)),(to_sfixed_a(0.011471612378954887)),(to_sfixed_a(0.018640680238604546)),(to_sfixed_a(0.01279165968298912)),(to_sfixed_a(0.0009610026609152555)),(to_sfixed_a(-2.885008871089667e-05)),(to_sfixed_a(0.00015073304530233145)),(to_sfixed_a(-1.34103320306167e-05)),(to_sfixed_a(-0.004400391131639481)),(to_sfixed_a(-2.209806552855298e-05)),(to_sfixed_a(7.474242011085153e-06)),(to_sfixed_a(-8.21111025288701e-05)),(to_sfixed_a(-0.20015288889408112)),(to_sfixed_a(-6.776781810913235e-05)),(to_sfixed_a(0.0021090770605951548)),(to_sfixed_a(-0.004675749689340591)),(to_sfixed_a(0.0020261977333575487)),(to_sfixed_a(0.0059884474612772465)),(to_sfixed_a(0.00012793263886123896)),(to_sfixed_a(0.004920169245451689)),(to_sfixed_a(-0.008698733523488045)),(to_sfixed_a(-0.17787925899028778)),(to_sfixed_a(0.00023118220269680023)),(to_sfixed_a(0.00786169059574604)),(to_sfixed_a(-0.7095603346824646)),(to_sfixed_a(0.01162412017583847)));

    constant weight_n2_97 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(-0.23141902685165405)),(to_sfixed_a(0.11885395646095276)),(to_sfixed_a(0.00013483337534125894)),(to_sfixed_a(-0.00020516464428510517)),(to_sfixed_a(-0.001013271976262331)),(to_sfixed_a(-1.899037670227699e-06)),(to_sfixed_a(0.3770414888858795)),(to_sfixed_a(-5.553643859457225e-06)),(to_sfixed_a(1.1197844287380576e-05)),(to_sfixed_a(0.00010107877460541204)),(to_sfixed_a(-0.00021664443193003535)),(to_sfixed_a(-0.012279397808015347)),(to_sfixed_a(-0.2596679925918579)),(to_sfixed_a(-0.005929878912866116)),(to_sfixed_a(1.4588396879844368e-05)),(to_sfixed_a(0.00024273377493955195)),(to_sfixed_a(-0.003456281963735819)),(to_sfixed_a(-4.990797606296837e-07)),(to_sfixed_a(-0.06624829769134521)),(to_sfixed_a(-0.006772737484425306)),(to_sfixed_a(0.0001780730381142348)),(to_sfixed_a(2.974956078105606e-05)),(to_sfixed_a(-0.00014069114695303142)),(to_sfixed_a(0.26378118991851807)),(to_sfixed_a(0.37520831823349)),(to_sfixed_a(-0.013962933793663979)),(to_sfixed_a(-6.215705070644617e-06)),(to_sfixed_a(0.0005498624523170292)),(to_sfixed_a(3.045744961127639e-06)),(to_sfixed_a(-3.0256680474849418e-05)),(to_sfixed_a(0.29815253615379333)),(to_sfixed_a(-4.8042144044302404e-05)),(to_sfixed_a(0.007859391160309315)),(to_sfixed_a(0.0001361908216495067)),(to_sfixed_a(-0.0003112399426754564)),(to_sfixed_a(-0.00020519270037766546)),(to_sfixed_a(-0.01220778189599514)),(to_sfixed_a(-0.2951447367668152)),(to_sfixed_a(-0.03470547869801521)),(to_sfixed_a(0.00015077779244165868)),(to_sfixed_a(0.0036926553584635258)),(to_sfixed_a(-0.019886570051312447)),(to_sfixed_a(-0.0001350856473436579)),(to_sfixed_a(-1.5781115507707e-05)),(to_sfixed_a(0.0142295490950346)),(to_sfixed_a(0.01750330999493599)),(to_sfixed_a(0.6489782929420471)),(to_sfixed_a(0.0005052564083598554)),(to_sfixed_a(6.665766704827547e-05)),(to_sfixed_a(0.4397922456264496)),(to_sfixed_a(0.2633000910282135)),(to_sfixed_a(-0.005454410798847675)),(to_sfixed_a(-0.00011980303679592907)),(to_sfixed_a(-0.009167936630547047)),(to_sfixed_a(0.006524510681629181)),(to_sfixed_a(-0.007084162440150976)),(to_sfixed_a(0.0001896530156955123)),(to_sfixed_a(0.007116908673197031)),(to_sfixed_a(0.0002958661352749914)),(to_sfixed_a(0.00024403989664278924)),(to_sfixed_a(0.01351907942444086)),(to_sfixed_a(-0.00010515256872167811)),(to_sfixed_a(0.000296772486763075)),(to_sfixed_a(0.00024689172278158367)),(to_sfixed_a(6.948832742637023e-05)),(to_sfixed_a(-0.20760829746723175)),(to_sfixed_a(0.00038943259278312325)),(to_sfixed_a(-0.0037335322704166174)),(to_sfixed_a(0.3418678045272827)),(to_sfixed_a(0.00021953225950710475)),(to_sfixed_a(-0.17005282640457153)),(to_sfixed_a(-0.0024584459606558084)),(to_sfixed_a(-0.0032582345884293318)),(to_sfixed_a(3.6364319385029376e-05)),(to_sfixed_a(8.393546158913523e-05)),(to_sfixed_a(-5.9986381529597566e-05)),(to_sfixed_a(0.00306294159963727)),(to_sfixed_a(-0.3139446973800659)),(to_sfixed_a(-0.00011275921860942617)),(to_sfixed_a(-0.012019741348922253)),(to_sfixed_a(0.01030071172863245)),(to_sfixed_a(2.779663191176951e-05)),(to_sfixed_a(0.2995597720146179)),(to_sfixed_a(-0.01201251894235611)),(to_sfixed_a(1.1032927432097495e-05)),(to_sfixed_a(0.003913315013051033)),(to_sfixed_a(-0.3989294171333313)),(to_sfixed_a(-0.0018135304562747478)),(to_sfixed_a(6.057324571884237e-05)),(to_sfixed_a(9.113558189710602e-05)),(to_sfixed_a(0.2723468840122223)),(to_sfixed_a(-5.996967956889421e-06)),(to_sfixed_a(0.00874802190810442)),(to_sfixed_a(-0.00011342061043251306)),(to_sfixed_a(0.0003105882497038692)),(to_sfixed_a(-3.350422775838524e-05)),(to_sfixed_a(-0.00020757369929924607)),(to_sfixed_a(-3.95057286368683e-05)),(to_sfixed_a(6.025817128829658e-06)),(to_sfixed_a(-0.0001036203175317496)),(to_sfixed_a(-0.00317291053943336)),(to_sfixed_a(0.0057176873087882996)),(to_sfixed_a(-0.00021341160754673183)),(to_sfixed_a(0.01063053123652935)),(to_sfixed_a(0.19414280354976654)),(to_sfixed_a(0.37253260612487793)),(to_sfixed_a(2.5216744688805193e-05)),(to_sfixed_a(-3.880549411405809e-05)),(to_sfixed_a(-2.2046242520445958e-05)),(to_sfixed_a(0.009584366343915462)),(to_sfixed_a(0.0028045405633747578)),(to_sfixed_a(0.00011564187298063189)),(to_sfixed_a(3.306294820504263e-05)),(to_sfixed_a(0.00011206141789443791)),(to_sfixed_a(-1.2657674233196303e-06)),(to_sfixed_a(-0.7170672416687012)),(to_sfixed_a(-0.00012901335139758885)),(to_sfixed_a(0.002569204196333885)),(to_sfixed_a(-3.6689030821435153e-05)),(to_sfixed_a(9.300222154706717e-05)),(to_sfixed_a(6.972685514483601e-05)),(to_sfixed_a(0.00024431338533759117)),(to_sfixed_a(0.007739727851003408)),(to_sfixed_a(-0.00014120832202024758)),(to_sfixed_a(0.00011307247041258961)),(to_sfixed_a(-0.554070234298706)),(to_sfixed_a(0.061004888266325)),(to_sfixed_a(-0.00016777135897427797)),(to_sfixed_a(-0.0004169110907241702)),(to_sfixed_a(-0.00012077923747710884)),(to_sfixed_a(0.00015508485375903547)),(to_sfixed_a(0.00017803366063162684)),(to_sfixed_a(-0.00995729025453329)),(to_sfixed_a(0.00690151983872056)),(to_sfixed_a(0.00010134656622540206)),(to_sfixed_a(0.00020009014406241477)),(to_sfixed_a(0.019984019920229912)),(to_sfixed_a(-6.113741255830973e-05)),(to_sfixed_a(1.1651580280158669e-05)),(to_sfixed_a(4.2633473640307784e-07)),(to_sfixed_a(0.0048105851747095585)),(to_sfixed_a(0.00022275513038039207)),(to_sfixed_a(0.00021819151879753917)),(to_sfixed_a(0.00016932730795815587)),(to_sfixed_a(-0.000418465759139508)),(to_sfixed_a(1.2976673133380245e-05)),(to_sfixed_a(0.026308316737413406)),(to_sfixed_a(-4.5995169784873724e-05)),(to_sfixed_a(-6.019996362738311e-06)),(to_sfixed_a(-0.009001616388559341)),(to_sfixed_a(4.4096064812038094e-05)),(to_sfixed_a(4.3526739318622276e-05)),(to_sfixed_a(0.0005296862800605595)),(to_sfixed_a(-0.00010588634177111089)),(to_sfixed_a(-0.00015536131104454398)),(to_sfixed_a(-0.30577221512794495)),(to_sfixed_a(9.986302757170051e-06)),(to_sfixed_a(0.05384393408894539)),(to_sfixed_a(-9.846459579421207e-05)),(to_sfixed_a(3.733061384991743e-05)),(to_sfixed_a(0.00011628773791017011)),(to_sfixed_a(0.00023116184456739575)),(to_sfixed_a(-0.00033554001129232347)),(to_sfixed_a(-0.001835643663071096)),(to_sfixed_a(-0.007776721380650997)),(to_sfixed_a(-0.0021083110477775335)),(to_sfixed_a(0.0001349036901956424)),(to_sfixed_a(0.004398969002068043)),(to_sfixed_a(-0.00018171951523981988)),(to_sfixed_a(3.675564585137181e-05)),(to_sfixed_a(-0.005272765178233385)),(to_sfixed_a(0.27578845620155334)),(to_sfixed_a(0.2423713505268097)),(to_sfixed_a(-3.1836410926189274e-05)),(to_sfixed_a(0.22512036561965942)),(to_sfixed_a(-0.00029561572591774166)),(to_sfixed_a(3.844790262519382e-05)),(to_sfixed_a(0.00047723978059366345)),(to_sfixed_a(-0.014197560027241707)),(to_sfixed_a(-0.26923489570617676)),(to_sfixed_a(-6.382470746757463e-05)),(to_sfixed_a(-0.00448789494112134)),(to_sfixed_a(0.00023285803035832942)),(to_sfixed_a(4.3483858462423086e-05)),(to_sfixed_a(0.00023729739768896252)),(to_sfixed_a(0.0001142672190326266)),(to_sfixed_a(-0.6550447344779968)),(to_sfixed_a(-0.0072255926206707954)),(to_sfixed_a(-0.006170038133859634)),(to_sfixed_a(0.5596655607223511)),(to_sfixed_a(-0.0010075995232909918)),(to_sfixed_a(-0.0001465700479457155)),(to_sfixed_a(-0.4528810679912567)),(to_sfixed_a(0.014962038956582546)),(to_sfixed_a(-0.00018292796448804438)),(to_sfixed_a(-0.3927047550678253)),(to_sfixed_a(-0.00016884587239474058)),(to_sfixed_a(0.0015872330404818058)),(to_sfixed_a(-0.00809481181204319)),(to_sfixed_a(-6.472550012404099e-05)),(to_sfixed_a(-6.595902959816158e-05)),(to_sfixed_a(-0.00022972984879743308)),(to_sfixed_a(-0.00019226089352741838)),(to_sfixed_a(0.00020176109683234245)),(to_sfixed_a(-0.00010545945406192914)),(to_sfixed_a(0.39639490842819214)),(to_sfixed_a(-0.00490706879645586)),(to_sfixed_a(-0.11690068989992142)),(to_sfixed_a(-0.0004844556387979537)),(to_sfixed_a(-2.6709691155701876e-05)),(to_sfixed_a(-0.034743182361125946)),(to_sfixed_a(0.00020115691586397588)),(to_sfixed_a(-0.0001961579837370664)),(to_sfixed_a(-6.329706957330927e-05)),(to_sfixed_a(-8.13203223515302e-06)),(to_sfixed_a(-0.0001371429389109835)),(to_sfixed_a(-0.0008903901325538754)),(to_sfixed_a(-0.21017882227897644)),(to_sfixed_a(-0.006530470680445433)),(to_sfixed_a(-0.00018900074064731598)),(to_sfixed_a(-3.183024819009006e-05)),(to_sfixed_a(0.00017532295896671712)),(to_sfixed_a(4.74863190902397e-06)),(to_sfixed_a(3.812667273450643e-06)),(to_sfixed_a(-0.10805176943540573)),(to_sfixed_a(-6.261280213948339e-05)),(to_sfixed_a(5.7137192925438285e-05)),(to_sfixed_a(0.0002938990364782512)),(to_sfixed_a(0.49923861026763916)),(to_sfixed_a(0.13296175003051758)),(to_sfixed_a(0.29209595918655396)),(to_sfixed_a(-7.739437569398433e-05)),(to_sfixed_a(-1.7635647964198142e-05)),(to_sfixed_a(0.00017389291315339506)),(to_sfixed_a(0.46152570843696594)),(to_sfixed_a(0.0035082008689641953)),(to_sfixed_a(0.0012994850985705853)),(to_sfixed_a(0.00011691037798300385)),(to_sfixed_a(-0.00210391147993505)),(to_sfixed_a(3.915953857358545e-05)),(to_sfixed_a(-0.015688985586166382)),(to_sfixed_a(0.00025578943314030766)),(to_sfixed_a(0.50534588098526)),(to_sfixed_a(-4.535129482974298e-05)),(to_sfixed_a(-0.4170364737510681)),(to_sfixed_a(0.31863072514533997)),(to_sfixed_a(-0.011429200880229473)),(to_sfixed_a(0.44473662972450256)),(to_sfixed_a(-0.00010544608085183427)),(to_sfixed_a(0.012773939408361912)),(to_sfixed_a(0.001296140137128532)),(to_sfixed_a(-0.00013649935135617852)),(to_sfixed_a(9.325033897766843e-05)),(to_sfixed_a(-0.00012170102854724973)),(to_sfixed_a(4.957935743732378e-05)),(to_sfixed_a(0.0014114173827692866)),(to_sfixed_a(-0.005647640209645033)),(to_sfixed_a(0.0001021335119730793)),(to_sfixed_a(-4.304018511902541e-05)),(to_sfixed_a(0.0028527406975626945)),(to_sfixed_a(1.8387734598945826e-05)),(to_sfixed_a(-0.0019898144528269768)),(to_sfixed_a(-0.00023263772891368717)),(to_sfixed_a(3.427783667575568e-06)),(to_sfixed_a(-6.75684423185885e-05)),(to_sfixed_a(-0.001450550858862698)),(to_sfixed_a(0.00010594353079795837)),(to_sfixed_a(2.9769824323011562e-05)),(to_sfixed_a(-7.444024959113449e-05)),(to_sfixed_a(-0.001688036834821105)),(to_sfixed_a(-0.0024998141452670097)),(to_sfixed_a(-0.00019859211170114577)),(to_sfixed_a(-6.311987817753106e-06)),(to_sfixed_a(0.00012724933912977576)),(to_sfixed_a(6.449000647990033e-05)),(to_sfixed_a(-0.005189951043576002)),(to_sfixed_a(0.2708762288093567)),(to_sfixed_a(0.23300272226333618)),(to_sfixed_a(0.0024294659961014986)),(to_sfixed_a(-0.0031358569394797087)),(to_sfixed_a(-3.2468640711158514e-05)),(to_sfixed_a(-0.00015531069948337972)),(to_sfixed_a(0.00019086833344772458)),(to_sfixed_a(5.221751780482009e-05)),(to_sfixed_a(-6.742196273989975e-05)),(to_sfixed_a(-0.00013047367974650115)),(to_sfixed_a(0.0012533603003248572)),(to_sfixed_a(0.0026220891159027815)),(to_sfixed_a(0.00011419306974858046)),(to_sfixed_a(-0.0006971515249460936)),(to_sfixed_a(-0.29996126890182495)),(to_sfixed_a(0.22598987817764282)),(to_sfixed_a(-0.018502408638596535)),(to_sfixed_a(-2.8067617677152157e-05)),(to_sfixed_a(-0.0012723295949399471)),(to_sfixed_a(4.883421934209764e-05)),(to_sfixed_a(0.11493009328842163)),(to_sfixed_a(0.00016703920846339315)),(to_sfixed_a(-0.0013525437097996473)),(to_sfixed_a(0.0024063533637672663)),(to_sfixed_a(0.1391083151102066)));

    constant weight_n2_98 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.4892161786556244)),(to_sfixed_a(-0.36527755856513977)),(to_sfixed_a(-0.6017817854881287)),(to_sfixed_a(-0.000251480785664171)),(to_sfixed_a(0.00033176096621900797)),(to_sfixed_a(0.0001296409172937274)),(to_sfixed_a(0.0003674043982755393)),(to_sfixed_a(1.1462470865808427e-05)),(to_sfixed_a(-5.094441803521477e-05)),(to_sfixed_a(-0.00015528142102994025)),(to_sfixed_a(0.00026248363428749144)),(to_sfixed_a(-0.31993088126182556)),(to_sfixed_a(-0.0006826769094914198)),(to_sfixed_a(0.01115801464766264)),(to_sfixed_a(9.310356836067513e-05)),(to_sfixed_a(6.8210756580811e-05)),(to_sfixed_a(-0.027163783088326454)),(to_sfixed_a(-7.246815948747098e-05)),(to_sfixed_a(0.0037689879536628723)),(to_sfixed_a(-0.0002447644073981792)),(to_sfixed_a(-0.00016789302753750235)),(to_sfixed_a(0.00010956081678159535)),(to_sfixed_a(-0.0002506173332221806)),(to_sfixed_a(0.0004050518327858299)),(to_sfixed_a(0.0008233898552134633)),(to_sfixed_a(4.7470366553170606e-05)),(to_sfixed_a(0.00010426988592371345)),(to_sfixed_a(3.429908974794671e-05)),(to_sfixed_a(0.27435022592544556)),(to_sfixed_a(-2.608183422125876e-06)),(to_sfixed_a(-0.27626675367355347)),(to_sfixed_a(-0.00018651687423698604)),(to_sfixed_a(-0.001516216667369008)),(to_sfixed_a(5.1123060984537005e-06)),(to_sfixed_a(-3.652734085335396e-05)),(to_sfixed_a(-1.3769997167401016e-05)),(to_sfixed_a(0.16694572567939758)),(to_sfixed_a(-0.001979326130822301)),(to_sfixed_a(0.006428475491702557)),(to_sfixed_a(0.0001283736783079803)),(to_sfixed_a(0.24206964671611786)),(to_sfixed_a(0.004939838778227568)),(to_sfixed_a(0.00023893913021311164)),(to_sfixed_a(-0.00017705137724988163)),(to_sfixed_a(-0.008296534419059753)),(to_sfixed_a(-0.017275745049118996)),(to_sfixed_a(-0.49875491857528687)),(to_sfixed_a(-0.0029216923285275698)),(to_sfixed_a(8.53941819514148e-05)),(to_sfixed_a(0.0012538135051727295)),(to_sfixed_a(0.011220172978937626)),(to_sfixed_a(-0.00036618250305764377)),(to_sfixed_a(-2.1889660274609923e-05)),(to_sfixed_a(0.0014288723468780518)),(to_sfixed_a(-0.1279737949371338)),(to_sfixed_a(0.005832526367157698)),(to_sfixed_a(5.832680471939966e-07)),(to_sfixed_a(-0.002207996789366007)),(to_sfixed_a(-1.1245199857512489e-05)),(to_sfixed_a(2.4454995582345873e-05)),(to_sfixed_a(-0.005306886043399572)),(to_sfixed_a(0.00011419501970522106)),(to_sfixed_a(-0.00027441655402071774)),(to_sfixed_a(-0.020807411521673203)),(to_sfixed_a(0.00010307988850399852)),(to_sfixed_a(0.22336852550506592)),(to_sfixed_a(6.529468373628333e-05)),(to_sfixed_a(0.0015960672171786427)),(to_sfixed_a(0.0003291968605481088)),(to_sfixed_a(-0.00017431596643291414)),(to_sfixed_a(0.014709370210766792)),(to_sfixed_a(0.012707805261015892)),(to_sfixed_a(-3.371161801624112e-05)),(to_sfixed_a(0.0004584754060488194)),(to_sfixed_a(-0.00016250723274424672)),(to_sfixed_a(0.00015432883810717613)),(to_sfixed_a(-0.34384623169898987)),(to_sfixed_a(0.1572183072566986)),(to_sfixed_a(3.229353387723677e-05)),(to_sfixed_a(-0.43202999234199524)),(to_sfixed_a(-0.00486797234043479)),(to_sfixed_a(3.0304421670734882e-05)),(to_sfixed_a(-0.398379385471344)),(to_sfixed_a(0.0008546859608031809)),(to_sfixed_a(-3.858418494928628e-05)),(to_sfixed_a(-4.500809154706076e-05)),(to_sfixed_a(0.5856648683547974)),(to_sfixed_a(0.00011671489482978359)),(to_sfixed_a(5.716155283153057e-05)),(to_sfixed_a(-7.228853064589202e-05)),(to_sfixed_a(0.015420523472130299)),(to_sfixed_a(-0.00041264755418524146)),(to_sfixed_a(-0.01182658039033413)),(to_sfixed_a(-0.00022970998543314636)),(to_sfixed_a(-0.010670553892850876)),(to_sfixed_a(1.7693833797238767e-05)),(to_sfixed_a(0.00010109358845511451)),(to_sfixed_a(-7.787689537508413e-05)),(to_sfixed_a(0.00015459457063116133)),(to_sfixed_a(-0.00017405538528691977)),(to_sfixed_a(7.078994531184435e-05)),(to_sfixed_a(-0.001610330305993557)),(to_sfixed_a(0.0003005467588081956)),(to_sfixed_a(-0.004561553243547678)),(to_sfixed_a(0.0024039142299443483)),(to_sfixed_a(-0.0007120780064724386)),(to_sfixed_a(-9.848400804912671e-05)),(to_sfixed_a(7.145700510591269e-05)),(to_sfixed_a(-1.3561118976213038e-05)),(to_sfixed_a(-0.003139782464131713)),(to_sfixed_a(-0.002535028848797083)),(to_sfixed_a(0.0002167350467061624)),(to_sfixed_a(0.00012951971439179033)),(to_sfixed_a(0.00023929028247948736)),(to_sfixed_a(0.00017114450747612864)),(to_sfixed_a(0.18016740679740906)),(to_sfixed_a(0.00011907612497452646)),(to_sfixed_a(8.556002285331488e-05)),(to_sfixed_a(0.00020455649064388126)),(to_sfixed_a(0.0008621212327852845)),(to_sfixed_a(0.0001659585104789585)),(to_sfixed_a(7.038261537672952e-05)),(to_sfixed_a(-0.006170019973069429)),(to_sfixed_a(8.554449595976621e-05)),(to_sfixed_a(3.0770243029110134e-05)),(to_sfixed_a(0.003276463830843568)),(to_sfixed_a(0.0033985183108597994)),(to_sfixed_a(0.0002499200636520982)),(to_sfixed_a(-5.011702160118148e-05)),(to_sfixed_a(0.00025071221170946956)),(to_sfixed_a(7.021697820164263e-05)),(to_sfixed_a(-0.00017213365936186165)),(to_sfixed_a(0.00024374431814067066)),(to_sfixed_a(-0.027573667466640472)),(to_sfixed_a(0.00016537836927454919)),(to_sfixed_a(1.1903339327545837e-06)),(to_sfixed_a(-0.011781474575400352)),(to_sfixed_a(-0.00018342991825193167)),(to_sfixed_a(0.00019736554531846195)),(to_sfixed_a(-0.00011372414155630395)),(to_sfixed_a(-0.002560774562880397)),(to_sfixed_a(-6.696397031191736e-05)),(to_sfixed_a(-6.46730768494308e-07)),(to_sfixed_a(2.5328730771434493e-05)),(to_sfixed_a(9.416689863428473e-06)),(to_sfixed_a(-9.81779012363404e-05)),(to_sfixed_a(0.0022194753400981426)),(to_sfixed_a(0.00017313846910838038)),(to_sfixed_a(4.403812999953516e-05)),(to_sfixed_a(0.00342165632173419)),(to_sfixed_a(-0.00023993068316485733)),(to_sfixed_a(0.00011253480624873191)),(to_sfixed_a(-0.0003951377875637263)),(to_sfixed_a(0.000116905321192462)),(to_sfixed_a(-7.7517019235529e-05)),(to_sfixed_a(0.0018333616899326444)),(to_sfixed_a(-0.0001562488469062373)),(to_sfixed_a(0.002978062490001321)),(to_sfixed_a(-4.467442340683192e-05)),(to_sfixed_a(-7.786028436385095e-05)),(to_sfixed_a(-4.44909674115479e-05)),(to_sfixed_a(-8.269526006188244e-07)),(to_sfixed_a(0.004455029033124447)),(to_sfixed_a(0.0007826965884305537)),(to_sfixed_a(0.0026426357217133045)),(to_sfixed_a(-0.0003933734551537782)),(to_sfixed_a(0.00015824197907932103)),(to_sfixed_a(0.2505352795124054)),(to_sfixed_a(0.00015310361050069332)),(to_sfixed_a(-3.6843914131168276e-05)),(to_sfixed_a(-0.00048679340397939086)),(to_sfixed_a(0.0003346044395584613)),(to_sfixed_a(0.00027110864175483584)),(to_sfixed_a(-3.0431845516432077e-05)),(to_sfixed_a(0.00030555337434634566)),(to_sfixed_a(0.00035381896304897964)),(to_sfixed_a(-0.34267255663871765)),(to_sfixed_a(-0.0002562030276749283)),(to_sfixed_a(0.0014002067036926746)),(to_sfixed_a(0.004089618567377329)),(to_sfixed_a(-4.232288119965233e-05)),(to_sfixed_a(0.010167159140110016)),(to_sfixed_a(-0.00017748872051015496)),(to_sfixed_a(0.00019208328740205616)),(to_sfixed_a(-6.434386159526184e-05)),(to_sfixed_a(-4.223869109409861e-05)),(to_sfixed_a(0.009688030928373337)),(to_sfixed_a(0.004975954536348581)),(to_sfixed_a(0.007990123704075813)),(to_sfixed_a(-0.16899380087852478)),(to_sfixed_a(0.0014097903622314334)),(to_sfixed_a(2.5628178264014423e-05)),(to_sfixed_a(-0.003963016904890537)),(to_sfixed_a(-0.007045583333820105)),(to_sfixed_a(-8.268941746791825e-05)),(to_sfixed_a(0.0003111725964117795)),(to_sfixed_a(-2.814919571392238e-05)),(to_sfixed_a(0.0009333681082352996)),(to_sfixed_a(0.010214493609964848)),(to_sfixed_a(-8.003026596270502e-05)),(to_sfixed_a(-1.2785902072209865e-05)),(to_sfixed_a(4.2130210204049945e-05)),(to_sfixed_a(-4.637894016923383e-05)),(to_sfixed_a(-8.153700764523819e-05)),(to_sfixed_a(3.358863978064619e-05)),(to_sfixed_a(0.003926421049982309)),(to_sfixed_a(-0.2013278752565384)),(to_sfixed_a(-0.0038663160521537066)),(to_sfixed_a(0.25147655606269836)),(to_sfixed_a(0.0024740842636674643)),(to_sfixed_a(0.003459411906078458)),(to_sfixed_a(0.00030947968480177224)),(to_sfixed_a(7.249755435623229e-05)),(to_sfixed_a(9.6401825430803e-05)),(to_sfixed_a(0.00016582751413807273)),(to_sfixed_a(0.00016592608881182969)),(to_sfixed_a(0.003913550172001123)),(to_sfixed_a(0.36957848072052)),(to_sfixed_a(0.015561604872345924)),(to_sfixed_a(-8.143833838403225e-07)),(to_sfixed_a(5.6829383538570255e-05)),(to_sfixed_a(-4.685512976720929e-06)),(to_sfixed_a(3.704741902765818e-05)),(to_sfixed_a(3.147327515762299e-05)),(to_sfixed_a(0.013343996368348598)),(to_sfixed_a(3.7771169445477426e-05)),(to_sfixed_a(2.4230579583672807e-05)),(to_sfixed_a(0.0001086747579392977)),(to_sfixed_a(-0.1411631554365158)),(to_sfixed_a(-0.00013814278645440936)),(to_sfixed_a(0.004128903150558472)),(to_sfixed_a(-0.00014391867443919182)),(to_sfixed_a(4.765672201756388e-05)),(to_sfixed_a(0.00021397579985205084)),(to_sfixed_a(-0.004582524299621582)),(to_sfixed_a(-0.004736663773655891)),(to_sfixed_a(-0.004387305583804846)),(to_sfixed_a(-0.0001555388153064996)),(to_sfixed_a(0.004108214285224676)),(to_sfixed_a(-1.6131889424286783e-07)),(to_sfixed_a(-0.27793052792549133)),(to_sfixed_a(5.1447856094455346e-05)),(to_sfixed_a(-0.4282519817352295)),(to_sfixed_a(0.0001569160958752036)),(to_sfixed_a(0.008536523208022118)),(to_sfixed_a(0.0016485049854964018)),(to_sfixed_a(-0.0037658517248928547)),(to_sfixed_a(-0.0027196297887712717)),(to_sfixed_a(-6.767624290660024e-05)),(to_sfixed_a(-0.012870069593191147)),(to_sfixed_a(-0.006085430271923542)),(to_sfixed_a(0.0001344291231362149)),(to_sfixed_a(0.00031811301596462727)),(to_sfixed_a(8.144073945004493e-06)),(to_sfixed_a(-0.24526429176330566)),(to_sfixed_a(-0.2895813584327698)),(to_sfixed_a(0.005013967864215374)),(to_sfixed_a(5.325615711626597e-05)),(to_sfixed_a(2.4712313461350277e-05)),(to_sfixed_a(0.00034882526961155236)),(to_sfixed_a(0.00024849671171978116)),(to_sfixed_a(0.00010718576959334314)),(to_sfixed_a(-9.216833859682083e-06)),(to_sfixed_a(-1.865820013335906e-05)),(to_sfixed_a(-0.00016710386262275279)),(to_sfixed_a(-0.0009054768015630543)),(to_sfixed_a(-0.00030904693994671106)),(to_sfixed_a(-9.402262367075309e-05)),(to_sfixed_a(3.640351496869698e-05)),(to_sfixed_a(0.00039160437881946564)),(to_sfixed_a(-0.00750504108145833)),(to_sfixed_a(2.7906326067750342e-05)),(to_sfixed_a(0.00013678264804184437)),(to_sfixed_a(-9.120747563429177e-05)),(to_sfixed_a(-2.9665170586667955e-06)),(to_sfixed_a(8.569309284212068e-05)),(to_sfixed_a(0.000537739833816886)),(to_sfixed_a(0.0004572496982291341)),(to_sfixed_a(0.0041574896313250065)),(to_sfixed_a(-0.30383726954460144)),(to_sfixed_a(-0.0001281610457226634)),(to_sfixed_a(1.651295315241441e-05)),(to_sfixed_a(0.00019701075507327914)),(to_sfixed_a(0.0005587504711002111)),(to_sfixed_a(0.0001286293991142884)),(to_sfixed_a(-0.0004136851930525154)),(to_sfixed_a(0.000563751847948879)),(to_sfixed_a(5.951007187832147e-05)),(to_sfixed_a(-2.852770921890624e-05)),(to_sfixed_a(-0.002027926268056035)),(to_sfixed_a(0.0005419125081971288)),(to_sfixed_a(-0.0019599893130362034)),(to_sfixed_a(-0.0022668878082185984)),(to_sfixed_a(-2.3900291125755757e-05)),(to_sfixed_a(0.1314830482006073)),(to_sfixed_a(0.0002727079263422638)),(to_sfixed_a(-0.007173359859734774)),(to_sfixed_a(7.066489342832938e-05)),(to_sfixed_a(0.004462711047381163)),(to_sfixed_a(0.3712695240974426)),(to_sfixed_a(-0.014903665520250797)));

    constant weight_n2_99 : sfixed_bus_array(300 downto 0) := ((to_sfixed_a(0.30035343766212463)),(to_sfixed_a(0.000461979623651132)),(to_sfixed_a(-0.0006685827393084764)),(to_sfixed_a(-0.000377038202714175)),(to_sfixed_a(0.008156852796673775)),(to_sfixed_a(-0.0001272608496947214)),(to_sfixed_a(-7.70512706367299e-05)),(to_sfixed_a(-9.873371163848788e-05)),(to_sfixed_a(2.9369006369961426e-05)),(to_sfixed_a(2.294443766004406e-05)),(to_sfixed_a(5.867919389856979e-05)),(to_sfixed_a(-0.025575270876288414)),(to_sfixed_a(-0.38180410861968994)),(to_sfixed_a(-0.001915331813506782)),(to_sfixed_a(0.00030782242538407445)),(to_sfixed_a(-0.00011052915942855179)),(to_sfixed_a(0.2524738311767578)),(to_sfixed_a(0.00022223444830160588)),(to_sfixed_a(-0.009313133545219898)),(to_sfixed_a(-0.009608536027371883)),(to_sfixed_a(-4.331304808147252e-06)),(to_sfixed_a(9.66036895988509e-06)),(to_sfixed_a(-0.0001051759027177468)),(to_sfixed_a(0.22261755168437958)),(to_sfixed_a(-0.00020518248493317515)),(to_sfixed_a(0.0009838936384767294)),(to_sfixed_a(-7.637156522832811e-05)),(to_sfixed_a(4.5894557842984796e-05)),(to_sfixed_a(0.0005880353855900466)),(to_sfixed_a(0.00016699093976058066)),(to_sfixed_a(0.0014550628839060664)),(to_sfixed_a(-1.0044812370324507e-05)),(to_sfixed_a(-0.001307008438743651)),(to_sfixed_a(0.00037932483246549964)),(to_sfixed_a(7.404306234093383e-05)),(to_sfixed_a(0.0002915484947152436)),(to_sfixed_a(0.0017987480387091637)),(to_sfixed_a(-0.00015310243179555982)),(to_sfixed_a(-0.0028737338725477457)),(to_sfixed_a(0.00010595013736747205)),(to_sfixed_a(0.03285670652985573)),(to_sfixed_a(-0.003265788545832038)),(to_sfixed_a(-3.2709813240217045e-05)),(to_sfixed_a(-0.00014804273087065667)),(to_sfixed_a(0.322843074798584)),(to_sfixed_a(-0.005921349860727787)),(to_sfixed_a(0.0003447030612733215)),(to_sfixed_a(-0.0003762636915780604)),(to_sfixed_a(-1.5991186955943704e-05)),(to_sfixed_a(-0.0008273949497379363)),(to_sfixed_a(0.0034899262245744467)),(to_sfixed_a(3.7655161577276886e-05)),(to_sfixed_a(-2.5739354896359146e-05)),(to_sfixed_a(0.0007661270210519433)),(to_sfixed_a(0.011916776187717915)),(to_sfixed_a(-0.0008748272666707635)),(to_sfixed_a(-3.221263250452466e-05)),(to_sfixed_a(-0.0006988599780015647)),(to_sfixed_a(-8.504414290655404e-05)),(to_sfixed_a(-6.846552423667163e-05)),(to_sfixed_a(0.0002066373999696225)),(to_sfixed_a(0.00032902491511777043)),(to_sfixed_a(-0.0013064203085377812)),(to_sfixed_a(-0.292063444852829)),(to_sfixed_a(2.524632145650685e-05)),(to_sfixed_a(0.2654470205307007)),(to_sfixed_a(0.0002483030839357525)),(to_sfixed_a(-0.0021982956677675247)),(to_sfixed_a(0.0002989376662299037)),(to_sfixed_a(-0.00010053481673821807)),(to_sfixed_a(0.00694514624774456)),(to_sfixed_a(0.46763256192207336)),(to_sfixed_a(0.002014008816331625)),(to_sfixed_a(-0.00023720780154690146)),(to_sfixed_a(9.718910587253049e-05)),(to_sfixed_a(-0.00011745209485525265)),(to_sfixed_a(0.40931037068367004)),(to_sfixed_a(-0.00422251271083951)),(to_sfixed_a(8.012240868993104e-05)),(to_sfixed_a(0.0010460972553119063)),(to_sfixed_a(0.0006059210281819105)),(to_sfixed_a(6.791068881284446e-05)),(to_sfixed_a(-0.0015777521766722202)),(to_sfixed_a(0.002057971665635705)),(to_sfixed_a(0.0001495414471719414)),(to_sfixed_a(0.15820841491222382)),(to_sfixed_a(-0.00903230719268322)),(to_sfixed_a(-7.036203896859661e-06)),(to_sfixed_a(-0.00021087288041599095)),(to_sfixed_a(-0.00011412370076868683)),(to_sfixed_a(-0.0008292656275443733)),(to_sfixed_a(7.600418757647276e-05)),(to_sfixed_a(-0.0015401460696011782)),(to_sfixed_a(9.357402450405061e-05)),(to_sfixed_a(0.00040811015060171485)),(to_sfixed_a(-2.051324918284081e-05)),(to_sfixed_a(-2.4860637495294213e-06)),(to_sfixed_a(1.0788036888698116e-05)),(to_sfixed_a(0.00016496612806804478)),(to_sfixed_a(1.0182106052525342e-05)),(to_sfixed_a(-1.701368273643311e-05)),(to_sfixed_a(-9.710265294415876e-05)),(to_sfixed_a(-0.00013384060002863407)),(to_sfixed_a(-0.008634747937321663)),(to_sfixed_a(0.31748566031455994)),(to_sfixed_a(-8.662394247949123e-05)),(to_sfixed_a(5.935771332588047e-05)),(to_sfixed_a(5.585404869634658e-05)),(to_sfixed_a(-7.134798215702176e-05)),(to_sfixed_a(-0.0019502906361594796)),(to_sfixed_a(0.0021795041393488646)),(to_sfixed_a(-7.882146746851504e-05)),(to_sfixed_a(-0.00043594243470579386)),(to_sfixed_a(0.00030205296934582293)),(to_sfixed_a(4.451143104233779e-05)),(to_sfixed_a(0.002418826799839735)),(to_sfixed_a(-0.0010952276643365622)),(to_sfixed_a(0.18010331690311432)),(to_sfixed_a(-2.9739036108367145e-05)),(to_sfixed_a(-0.38714364171028137)),(to_sfixed_a(-0.00015512722893618047)),(to_sfixed_a(9.670630242908373e-05)),(to_sfixed_a(-0.0002844286209437996)),(to_sfixed_a(6.395934906322509e-05)),(to_sfixed_a(-0.00015450581850018352)),(to_sfixed_a(-0.00029249119688756764)),(to_sfixed_a(0.0026100222021341324)),(to_sfixed_a(-4.850400728173554e-06)),(to_sfixed_a(-4.4897326006321236e-05)),(to_sfixed_a(-4.5855995267629623e-07)),(to_sfixed_a(3.714812555699609e-05)),(to_sfixed_a(0.00014930943143554032)),(to_sfixed_a(0.0006736959330737591)),(to_sfixed_a(0.003364736447110772)),(to_sfixed_a(0.0002499204420018941)),(to_sfixed_a(-6.036547711119056e-05)),(to_sfixed_a(0.05161191523075104)),(to_sfixed_a(-3.8633465010207146e-05)),(to_sfixed_a(-0.0001960594963748008)),(to_sfixed_a(2.9072522011119872e-05)),(to_sfixed_a(-0.0004897105973213911)),(to_sfixed_a(-0.00011706026998581365)),(to_sfixed_a(-4.273862577974796e-05)),(to_sfixed_a(2.1904055756749585e-05)),(to_sfixed_a(-0.00010775164264487103)),(to_sfixed_a(1.2825308658648282e-05)),(to_sfixed_a(-0.0001767008361639455)),(to_sfixed_a(8.641881868243217e-05)),(to_sfixed_a(-7.490170537494123e-05)),(to_sfixed_a(-0.004094335250556469)),(to_sfixed_a(-1.7083773855119944e-05)),(to_sfixed_a(6.783152639400214e-05)),(to_sfixed_a(-0.00010599872621241957)),(to_sfixed_a(-0.00010848298552446067)),(to_sfixed_a(0.00017129532352555543)),(to_sfixed_a(0.15446507930755615)),(to_sfixed_a(-3.2588512112852186e-05)),(to_sfixed_a(-0.00354961515404284)),(to_sfixed_a(4.634581273421645e-05)),(to_sfixed_a(0.00010012292477767915)),(to_sfixed_a(-0.0002892670745495707)),(to_sfixed_a(-6.839314301032573e-05)),(to_sfixed_a(0.000757515721488744)),(to_sfixed_a(0.0001884621597127989)),(to_sfixed_a(0.35160866379737854)),(to_sfixed_a(-0.0004453505971468985)),(to_sfixed_a(0.00045060255797579885)),(to_sfixed_a(0.00012104538473067805)),(to_sfixed_a(-0.00017780651978682727)),(to_sfixed_a(0.00016900910122785717)),(to_sfixed_a(-0.5506992340087891)),(to_sfixed_a(-0.00012636787141673267)),(to_sfixed_a(1.770536255207844e-05)),(to_sfixed_a(1.886237077997066e-05)),(to_sfixed_a(-0.007631960324943066)),(to_sfixed_a(-4.4710657675750554e-05)),(to_sfixed_a(-0.27365007996559143)),(to_sfixed_a(0.25608721375465393)),(to_sfixed_a(-0.00802198238670826)),(to_sfixed_a(0.5154061913490295)),(to_sfixed_a(0.0006759206880815327)),(to_sfixed_a(-0.003126956755295396)),(to_sfixed_a(-4.094902396900579e-05)),(to_sfixed_a(-3.303551784483716e-05)),(to_sfixed_a(-2.9078000807203352e-05)),(to_sfixed_a(-6.632617441937327e-05)),(to_sfixed_a(0.010491080582141876)),(to_sfixed_a(0.0020590878557413816)),(to_sfixed_a(-8.643321052659303e-05)),(to_sfixed_a(-3.793568248511292e-05)),(to_sfixed_a(-0.013600409030914307)),(to_sfixed_a(4.291661025490612e-05)),(to_sfixed_a(-0.29623812437057495)),(to_sfixed_a(0.22353392839431763)),(to_sfixed_a(-0.00017419160576537251)),(to_sfixed_a(0.0003719716041814536)),(to_sfixed_a(2.4120276066241786e-05)),(to_sfixed_a(0.002584129571914673)),(to_sfixed_a(-0.0004908589762635529)),(to_sfixed_a(-0.00020026932179462165)),(to_sfixed_a(0.00011345373786753044)),(to_sfixed_a(1.6626801880192943e-05)),(to_sfixed_a(0.00015859481936786324)),(to_sfixed_a(-6.831968494225293e-05)),(to_sfixed_a(0.00014644392649643123)),(to_sfixed_a(0.002615497447550297)),(to_sfixed_a(7.281760917976499e-05)),(to_sfixed_a(0.11492214351892471)),(to_sfixed_a(0.1755593866109848)),(to_sfixed_a(0.17858029901981354)),(to_sfixed_a(-0.00952945463359356)),(to_sfixed_a(-0.0004450474225450307)),(to_sfixed_a(-0.00019166438141837716)),(to_sfixed_a(1.0321135050617158e-05)),(to_sfixed_a(-0.0001766662171576172)),(to_sfixed_a(-7.018634642008692e-05)),(to_sfixed_a(0.0003140583576168865)),(to_sfixed_a(0.002772929146885872)),(to_sfixed_a(0.004931629169732332)),(to_sfixed_a(0.00015747180441394448)),(to_sfixed_a(-7.831687980797142e-06)),(to_sfixed_a(6.942032632650807e-05)),(to_sfixed_a(0.00015405676094815135)),(to_sfixed_a(-1.9169880033587106e-05)),(to_sfixed_a(0.44230329990386963)),(to_sfixed_a(-0.0001374419080093503)),(to_sfixed_a(-0.00011692442058119923)),(to_sfixed_a(3.345048753544688e-05)),(to_sfixed_a(0.10223506391048431)),(to_sfixed_a(-0.0009027792839333415)),(to_sfixed_a(0.42010411620140076)),(to_sfixed_a(0.00020118615066166967)),(to_sfixed_a(-0.0002864630369003862)),(to_sfixed_a(-0.00024438570835627615)),(to_sfixed_a(-0.0003571399429347366)),(to_sfixed_a(0.0003321791300550103)),(to_sfixed_a(-0.0025601775851100683)),(to_sfixed_a(-6.73479080433026e-05)),(to_sfixed_a(5.217327270656824e-05)),(to_sfixed_a(0.000163281278219074)),(to_sfixed_a(0.001141039072535932)),(to_sfixed_a(6.92751127644442e-05)),(to_sfixed_a(-0.1746227741241455)),(to_sfixed_a(-4.460227501112968e-06)),(to_sfixed_a(-0.0702044814825058)),(to_sfixed_a(-0.0013428095262497663)),(to_sfixed_a(0.4422045052051544)),(to_sfixed_a(0.01857718452811241)),(to_sfixed_a(1.9558952772058547e-05)),(to_sfixed_a(-0.009159300476312637)),(to_sfixed_a(0.0007784998160786927)),(to_sfixed_a(-5.909695755690336e-05)),(to_sfixed_a(0.0007120900554582477)),(to_sfixed_a(-2.2989352146396413e-05)),(to_sfixed_a(5.780028004664928e-06)),(to_sfixed_a(-0.25969821214675903)),(to_sfixed_a(-0.004737451206892729)),(to_sfixed_a(0.0001743861212162301)),(to_sfixed_a(-2.9126385925337672e-06)),(to_sfixed_a(-0.0003695389023050666)),(to_sfixed_a(9.80929471552372e-05)),(to_sfixed_a(-0.21065795421600342)),(to_sfixed_a(-0.000246467039687559)),(to_sfixed_a(0.00045088506885804236)),(to_sfixed_a(0.00024306614068336785)),(to_sfixed_a(0.002015241188928485)),(to_sfixed_a(-0.00022845632338430732)),(to_sfixed_a(-4.5556589611805975e-06)),(to_sfixed_a(6.797620153520256e-05)),(to_sfixed_a(0.3711185157299042)),(to_sfixed_a(0.011126893572509289)),(to_sfixed_a(-0.00024835619842633605)),(to_sfixed_a(2.2781889128964394e-05)),(to_sfixed_a(-6.776375812478364e-05)),(to_sfixed_a(-5.488065653480589e-06)),(to_sfixed_a(-0.3606738746166229)),(to_sfixed_a(0.00019360646547283977)),(to_sfixed_a(0.002134669106453657)),(to_sfixed_a(0.4340098798274994)),(to_sfixed_a(0.44263342022895813)),(to_sfixed_a(0.00028918759198859334)),(to_sfixed_a(-0.00025439480668865144)),(to_sfixed_a(7.102893141563982e-05)),(to_sfixed_a(-0.01134900376200676)),(to_sfixed_a(-5.243462510406971e-05)),(to_sfixed_a(-7.498296326957643e-05)),(to_sfixed_a(-0.0044653648510575294)),(to_sfixed_a(0.003580136224627495)),(to_sfixed_a(1.0979783837683499e-05)),(to_sfixed_a(-0.001292300526984036)),(to_sfixed_a(-0.0006156474119052291)),(to_sfixed_a(-0.00010471649875398725)),(to_sfixed_a(0.004794255364686251)),(to_sfixed_a(-2.150671207346022e-06)),(to_sfixed_a(0.0016152022872120142)),(to_sfixed_a(-0.00027389515889808536)),(to_sfixed_a(6.7056120315101e-05)),(to_sfixed_a(0.000168528436915949)),(to_sfixed_a(-0.007147282361984253)),(to_sfixed_a(-0.0024599775206297636)),(to_sfixed_a(-0.0016054688021540642)));


    constant weight_n3_0 : sfixed_bus_array(100 downto 0) := ((to_sfixed_a(-0.04710623621940613)),(to_sfixed_a(0.3763449490070343)),(to_sfixed_a(-0.7617764472961426)),(to_sfixed_a(0.4409821629524231)),(to_sfixed_a(0.0001300221192650497)),(to_sfixed_a(0.00015652738511562347)),(to_sfixed_a(0.40391218662261963)),(to_sfixed_a(-0.2840213179588318)),(to_sfixed_a(-0.10695584118366241)),(to_sfixed_a(4.31457010563463e-06)),(to_sfixed_a(-0.13787254691123962)),(to_sfixed_a(0.04132073000073433)),(to_sfixed_a(0.556298553943634)),(to_sfixed_a(0.030569227412343025)),(to_sfixed_a(-0.4266444444656372)),(to_sfixed_a(0.0019841166213154793)),(to_sfixed_a(-0.7434200644493103)),(to_sfixed_a(-0.7760781645774841)),(to_sfixed_a(-0.009446082636713982)),(to_sfixed_a(-0.8929973840713501)),(to_sfixed_a(1.422857167199254e-05)),(to_sfixed_a(-0.25395315885543823)),(to_sfixed_a(-0.4154244661331177)),(to_sfixed_a(-0.8685311675071716)),(to_sfixed_a(1.733101817080751e-05)),(to_sfixed_a(-0.329542338848114)),(to_sfixed_a(0.32824504375457764)),(to_sfixed_a(0.23624159395694733)),(to_sfixed_a(-0.43029969930648804)),(to_sfixed_a(-0.2693560719490051)),(to_sfixed_a(0.3176901340484619)),(to_sfixed_a(-1.0483064651489258)),(to_sfixed_a(-0.9791849255561829)),(to_sfixed_a(0.7979064583778381)),(to_sfixed_a(0.15571264922618866)),(to_sfixed_a(8.7624357547611e-07)),(to_sfixed_a(0.00022130478464532644)),(to_sfixed_a(0.4782354533672333)),(to_sfixed_a(-0.8895567655563354)),(to_sfixed_a(-0.5480548143386841)),(to_sfixed_a(-0.6267082691192627)),(to_sfixed_a(0.077970951795578)),(to_sfixed_a(6.754342757631093e-05)),(to_sfixed_a(0.03548820689320564)),(to_sfixed_a(-0.1397372931241989)),(to_sfixed_a(0.42480310797691345)),(to_sfixed_a(0.4264323115348816)),(to_sfixed_a(-0.37304842472076416)),(to_sfixed_a(-0.20360834896564484)),(to_sfixed_a(0.3267320990562439)),(to_sfixed_a(0.31235942244529724)),(to_sfixed_a(0.18552708625793457)),(to_sfixed_a(0.45368799567222595)),(to_sfixed_a(0.1901344656944275)),(to_sfixed_a(0.3460409641265869)),(to_sfixed_a(-0.026460113003849983)),(to_sfixed_a(0.19638189673423767)),(to_sfixed_a(-0.24961169064044952)),(to_sfixed_a(0.3460686504840851)),(to_sfixed_a(0.23853875696659088)),(to_sfixed_a(0.33994024991989136)),(to_sfixed_a(-0.00042916671372950077)),(to_sfixed_a(0.1708698868751526)),(to_sfixed_a(-0.10271141678094864)),(to_sfixed_a(0.0797453224658966)),(to_sfixed_a(0.015079135075211525)),(to_sfixed_a(-0.13844531774520874)),(to_sfixed_a(-0.0001132836114265956)),(to_sfixed_a(-0.0034344512969255447)),(to_sfixed_a(-0.25852131843566895)),(to_sfixed_a(0.31689056754112244)),(to_sfixed_a(0.14611753821372986)),(to_sfixed_a(0.3796303868293762)),(to_sfixed_a(0.12109557539224625)),(to_sfixed_a(-0.40405258536338806)),(to_sfixed_a(0.26492342352867126)),(to_sfixed_a(-0.6543368697166443)),(to_sfixed_a(0.13724003732204437)),(to_sfixed_a(0.3397751450538635)),(to_sfixed_a(0.04532172903418541)),(to_sfixed_a(-0.5592487454414368)),(to_sfixed_a(0.3962065577507019)),(to_sfixed_a(0.4146696925163269)),(to_sfixed_a(-0.4014270007610321)),(to_sfixed_a(0.00014716581790708005)),(to_sfixed_a(0.3174712657928467)),(to_sfixed_a(0.19808393716812134)),(to_sfixed_a(0.36742103099823)),(to_sfixed_a(-0.8598566651344299)),(to_sfixed_a(-0.1838712990283966)),(to_sfixed_a(0.00011374332098057494)),(to_sfixed_a(-0.433421790599823)),(to_sfixed_a(0.15760689973831177)),(to_sfixed_a(-0.07914464175701141)),(to_sfixed_a(-0.6302826404571533)),(to_sfixed_a(-6.378423131536692e-05)),(to_sfixed_a(0.17099612951278687)),(to_sfixed_a(0.35187825560569763)),(to_sfixed_a(-0.752302885055542)),(to_sfixed_a(0.26524534821510315)),(to_sfixed_a(-0.5792188048362732)));

    constant weight_n3_1 : sfixed_bus_array(100 downto 0) := ((to_sfixed_a(-0.29839757084846497)),(to_sfixed_a(-0.2937825620174408)),(to_sfixed_a(0.21300749480724335)),(to_sfixed_a(-0.012257945723831654)),(to_sfixed_a(0.0001470471324864775)),(to_sfixed_a(-0.00015719102520961314)),(to_sfixed_a(-1.0493649244308472)),(to_sfixed_a(-0.37903815507888794)),(to_sfixed_a(-0.00028018414741382003)),(to_sfixed_a(-0.00019548214913811535)),(to_sfixed_a(0.22879904508590698)),(to_sfixed_a(-0.6502016186714172)),(to_sfixed_a(-0.04232430085539818)),(to_sfixed_a(0.5192570090293884)),(to_sfixed_a(-0.24087314307689667)),(to_sfixed_a(0.38930773735046387)),(to_sfixed_a(0.3631878197193146)),(to_sfixed_a(-0.0375785231590271)),(to_sfixed_a(0.16721607744693756)),(to_sfixed_a(-0.05633193999528885)),(to_sfixed_a(2.075776683341246e-05)),(to_sfixed_a(-1.043148398399353)),(to_sfixed_a(0.18889528512954712)),(to_sfixed_a(0.18394704163074493)),(to_sfixed_a(7.224678847705945e-05)),(to_sfixed_a(-1.105270504951477)),(to_sfixed_a(-0.918992817401886)),(to_sfixed_a(-0.2999286949634552)),(to_sfixed_a(-0.3988117575645447)),(to_sfixed_a(0.2387736290693283)),(to_sfixed_a(-0.22427108883857727)),(to_sfixed_a(-0.3403360843658447)),(to_sfixed_a(0.10330092161893845)),(to_sfixed_a(0.5482797026634216)),(to_sfixed_a(0.9388211369514465)),(to_sfixed_a(-9.995291475206614e-05)),(to_sfixed_a(0.38210541009902954)),(to_sfixed_a(-0.1012345403432846)),(to_sfixed_a(0.2356419861316681)),(to_sfixed_a(-0.01824277453124523)),(to_sfixed_a(-0.09510163217782974)),(to_sfixed_a(-0.06820076704025269)),(to_sfixed_a(-2.107038744725287e-05)),(to_sfixed_a(-0.0012398118851706386)),(to_sfixed_a(0.10025772452354431)),(to_sfixed_a(0.06502222269773483)),(to_sfixed_a(-0.013082110323011875)),(to_sfixed_a(0.47002795338630676)),(to_sfixed_a(-0.09687507152557373)),(to_sfixed_a(-0.36304163932800293)),(to_sfixed_a(-0.29217061400413513)),(to_sfixed_a(-0.6964177489280701)),(to_sfixed_a(-0.14498241245746613)),(to_sfixed_a(0.21057555079460144)),(to_sfixed_a(0.20220492780208588)),(to_sfixed_a(0.038760218769311905)),(to_sfixed_a(-0.3219139873981476)),(to_sfixed_a(-0.0035186957102268934)),(to_sfixed_a(-0.1780935525894165)),(to_sfixed_a(0.12902845442295074)),(to_sfixed_a(0.0061125424690544605)),(to_sfixed_a(0.3048047423362732)),(to_sfixed_a(-0.44689255952835083)),(to_sfixed_a(0.311125248670578)),(to_sfixed_a(0.10502580553293228)),(to_sfixed_a(-0.6004634499549866)),(to_sfixed_a(0.42719316482543945)),(to_sfixed_a(-1.122952380683273e-05)),(to_sfixed_a(-0.12068583816289902)),(to_sfixed_a(0.14971554279327393)),(to_sfixed_a(0.0023129405453801155)),(to_sfixed_a(0.15481090545654297)),(to_sfixed_a(-0.0062409755773842335)),(to_sfixed_a(-0.8479071855545044)),(to_sfixed_a(0.17209124565124512)),(to_sfixed_a(0.013452956452965736)),(to_sfixed_a(0.11286912858486176)),(to_sfixed_a(0.10247360169887543)),(to_sfixed_a(-1.052510380744934)),(to_sfixed_a(0.3732805848121643)),(to_sfixed_a(0.13111914694309235)),(to_sfixed_a(0.12257011234760284)),(to_sfixed_a(-0.19690684974193573)),(to_sfixed_a(-0.16809998452663422)),(to_sfixed_a(-0.00013544327521231025)),(to_sfixed_a(-0.6833446621894836)),(to_sfixed_a(0.24959403276443481)),(to_sfixed_a(-0.6028320789337158)),(to_sfixed_a(-0.6662129759788513)),(to_sfixed_a(0.2255038022994995)),(to_sfixed_a(0.00011389065184630454)),(to_sfixed_a(-0.20575018227100372)),(to_sfixed_a(0.08582509309053421)),(to_sfixed_a(-0.6326587796211243)),(to_sfixed_a(-0.6519720554351807)),(to_sfixed_a(-2.9507153158192523e-05)),(to_sfixed_a(1.894012348202523e-05)),(to_sfixed_a(0.5721070766448975)),(to_sfixed_a(0.588867723941803)),(to_sfixed_a(-0.33286115527153015)),(to_sfixed_a(0.22069187462329865)));

    constant weight_n3_2 : sfixed_bus_array(100 downto 0) := ((to_sfixed_a(-0.04567766934633255)),(to_sfixed_a(-0.3719732165336609)),(to_sfixed_a(0.2164086103439331)),(to_sfixed_a(-0.28230464458465576)),(to_sfixed_a(-0.00017337511235382408)),(to_sfixed_a(-7.776396523695439e-05)),(to_sfixed_a(0.11960052698850632)),(to_sfixed_a(0.06724271923303604)),(to_sfixed_a(0.5639423131942749)),(to_sfixed_a(0.00022457893646787852)),(to_sfixed_a(0.36213839054107666)),(to_sfixed_a(-0.0034812455996870995)),(to_sfixed_a(-0.1074049323797226)),(to_sfixed_a(-0.5462525486946106)),(to_sfixed_a(0.08418375998735428)),(to_sfixed_a(-0.6354975700378418)),(to_sfixed_a(0.1206170916557312)),(to_sfixed_a(0.21121004223823547)),(to_sfixed_a(-0.24122704565525055)),(to_sfixed_a(-0.4089210033416748)),(to_sfixed_a(-0.0001048082485795021)),(to_sfixed_a(-0.29202035069465637)),(to_sfixed_a(-0.749655544757843)),(to_sfixed_a(0.21333745121955872)),(to_sfixed_a(-0.00013928221596870571)),(to_sfixed_a(0.23479339480400085)),(to_sfixed_a(0.04653739556670189)),(to_sfixed_a(-0.445159375667572)),(to_sfixed_a(-0.06635205447673798)),(to_sfixed_a(0.33333200216293335)),(to_sfixed_a(-0.2852790057659149)),(to_sfixed_a(0.01703648827970028)),(to_sfixed_a(0.5013839602470398)),(to_sfixed_a(-0.4865361452102661)),(to_sfixed_a(-0.8789671063423157)),(to_sfixed_a(-0.0001166290749097243)),(to_sfixed_a(-0.8689758777618408)),(to_sfixed_a(-0.028454752638936043)),(to_sfixed_a(0.31131383776664734)),(to_sfixed_a(-0.3092220425605774)),(to_sfixed_a(0.31546640396118164)),(to_sfixed_a(0.2706781029701233)),(to_sfixed_a(-0.05471564084291458)),(to_sfixed_a(0.12430910766124725)),(to_sfixed_a(-0.7832139730453491)),(to_sfixed_a(0.1474241465330124)),(to_sfixed_a(0.4077550768852234)),(to_sfixed_a(-0.2527550756931305)),(to_sfixed_a(0.00516738323494792)),(to_sfixed_a(0.21164624392986298)),(to_sfixed_a(0.2214745730161667)),(to_sfixed_a(-0.6073875427246094)),(to_sfixed_a(0.07476125657558441)),(to_sfixed_a(0.267482191324234)),(to_sfixed_a(0.31157568097114563)),(to_sfixed_a(-0.5578645467758179)),(to_sfixed_a(-0.011529149487614632)),(to_sfixed_a(-0.6457159519195557)),(to_sfixed_a(0.33731892704963684)),(to_sfixed_a(0.21108131110668182)),(to_sfixed_a(-0.3144342601299286)),(to_sfixed_a(-0.06782159954309464)),(to_sfixed_a(0.034287869930267334)),(to_sfixed_a(-0.11157676577568054)),(to_sfixed_a(-0.3241826891899109)),(to_sfixed_a(0.3343013525009155)),(to_sfixed_a(0.5410431623458862)),(to_sfixed_a(-1.1533764336491004e-05)),(to_sfixed_a(-0.22227700054645538)),(to_sfixed_a(0.18768669664859772)),(to_sfixed_a(0.16782540082931519)),(to_sfixed_a(-0.06181421875953674)),(to_sfixed_a(0.20904263854026794)),(to_sfixed_a(0.16927187144756317)),(to_sfixed_a(-0.3299201428890228)),(to_sfixed_a(0.1643693894147873)),(to_sfixed_a(-0.254702091217041)),(to_sfixed_a(0.1479976773262024)),(to_sfixed_a(0.2326970398426056)),(to_sfixed_a(-0.3517605662345886)),(to_sfixed_a(-0.16307292878627777)),(to_sfixed_a(-0.053437668830156326)),(to_sfixed_a(0.006415600888431072)),(to_sfixed_a(0.3040844202041626)),(to_sfixed_a(-3.724861016962677e-05)),(to_sfixed_a(0.2608039379119873)),(to_sfixed_a(-0.1636972576379776)),(to_sfixed_a(-0.3277636468410492)),(to_sfixed_a(0.501321017742157)),(to_sfixed_a(0.006549194920808077)),(to_sfixed_a(6.058723738533445e-05)),(to_sfixed_a(-0.8060452342033386)),(to_sfixed_a(0.02126026153564453)),(to_sfixed_a(0.27664750814437866)),(to_sfixed_a(-0.5126999616622925)),(to_sfixed_a(-0.0001466807589167729)),(to_sfixed_a(-0.6499677896499634)),(to_sfixed_a(0.16541148722171783)),(to_sfixed_a(0.611630380153656)),(to_sfixed_a(-0.09904738515615463)),(to_sfixed_a(0.10077879577875137)));

    constant weight_n3_3 : sfixed_bus_array(100 downto 0) := ((to_sfixed_a(-0.00612062681466341)),(to_sfixed_a(-0.6480770707130432)),(to_sfixed_a(0.10939638316631317)),(to_sfixed_a(0.6351779103279114)),(to_sfixed_a(0.0003889766230713576)),(to_sfixed_a(-9.609411063138396e-05)),(to_sfixed_a(-0.23910614848136902)),(to_sfixed_a(0.24895694851875305)),(to_sfixed_a(0.005492630880326033)),(to_sfixed_a(0.000109576947579626)),(to_sfixed_a(0.3855794072151184)),(to_sfixed_a(0.060337234288454056)),(to_sfixed_a(0.1461547166109085)),(to_sfixed_a(0.6108322143554688)),(to_sfixed_a(0.34351879358291626)),(to_sfixed_a(-0.7334631681442261)),(to_sfixed_a(-0.6085143089294434)),(to_sfixed_a(0.28997182846069336)),(to_sfixed_a(0.16736584901809692)),(to_sfixed_a(-0.15224239230155945)),(to_sfixed_a(9.754298662301153e-05)),(to_sfixed_a(0.7517185211181641)),(to_sfixed_a(0.12215588986873627)),(to_sfixed_a(-0.35362377762794495)),(to_sfixed_a(0.00015212985454127192)),(to_sfixed_a(0.0007045947713777423)),(to_sfixed_a(0.2967103123664856)),(to_sfixed_a(0.20046940445899963)),(to_sfixed_a(0.20176219940185547)),(to_sfixed_a(-0.49042025208473206)),(to_sfixed_a(-0.2840542495250702)),(to_sfixed_a(0.8959931135177612)),(to_sfixed_a(0.31113964319229126)),(to_sfixed_a(0.08561151474714279)),(to_sfixed_a(0.24842800199985504)),(to_sfixed_a(8.504706784151495e-06)),(to_sfixed_a(0.016794569790363312)),(to_sfixed_a(-0.16484951972961426)),(to_sfixed_a(-0.38046684861183167)),(to_sfixed_a(-0.43778762221336365)),(to_sfixed_a(-0.3304799497127533)),(to_sfixed_a(0.25321224331855774)),(to_sfixed_a(1.4721041225129738e-05)),(to_sfixed_a(0.12885160744190216)),(to_sfixed_a(-0.006006479728966951)),(to_sfixed_a(-0.6888360381126404)),(to_sfixed_a(-0.27255305647850037)),(to_sfixed_a(0.0131282489746809)),(to_sfixed_a(0.2506294846534729)),(to_sfixed_a(0.2693009078502655)),(to_sfixed_a(-0.12858368456363678)),(to_sfixed_a(0.32727670669555664)),(to_sfixed_a(-0.3351289927959442)),(to_sfixed_a(0.06104421615600586)),(to_sfixed_a(-0.19972197711467743)),(to_sfixed_a(-0.162917822599411)),(to_sfixed_a(-0.5561903715133667)),(to_sfixed_a(-0.9192735552787781)),(to_sfixed_a(-0.2353581339120865)),(to_sfixed_a(0.12886226177215576)),(to_sfixed_a(0.14225523173809052)),(to_sfixed_a(-0.9693158864974976)),(to_sfixed_a(-0.1455555260181427)),(to_sfixed_a(0.1883147805929184)),(to_sfixed_a(-0.3469448387622833)),(to_sfixed_a(-0.4642559885978699)),(to_sfixed_a(-0.74592125415802)),(to_sfixed_a(-0.00025131157599389553)),(to_sfixed_a(0.35679370164871216)),(to_sfixed_a(0.022164950147271156)),(to_sfixed_a(-0.2816550135612488)),(to_sfixed_a(-0.18428850173950195)),(to_sfixed_a(0.1228313222527504)),(to_sfixed_a(-0.0005628320504911244)),(to_sfixed_a(0.14787395298480988)),(to_sfixed_a(-0.033234309405088425)),(to_sfixed_a(0.14841608703136444)),(to_sfixed_a(0.2644636034965515)),(to_sfixed_a(-0.31242018938064575)),(to_sfixed_a(-0.9911337494850159)),(to_sfixed_a(0.3223003149032593)),(to_sfixed_a(-0.4550703465938568)),(to_sfixed_a(0.646187961101532)),(to_sfixed_a(-0.24184666574001312)),(to_sfixed_a(6.958243466215208e-05)),(to_sfixed_a(0.2789382338523865)),(to_sfixed_a(-0.30756911635398865)),(to_sfixed_a(-0.15178510546684265)),(to_sfixed_a(0.2678009569644928)),(to_sfixed_a(-0.5025453567504883)),(to_sfixed_a(7.153309707064182e-05)),(to_sfixed_a(0.3227294385433197)),(to_sfixed_a(0.09724339097738266)),(to_sfixed_a(0.45321735739707947)),(to_sfixed_a(0.2794533371925354)),(to_sfixed_a(-0.00020387909899000078)),(to_sfixed_a(-0.27010858058929443)),(to_sfixed_a(-0.4821440577507019)),(to_sfixed_a(-0.59548419713974)),(to_sfixed_a(-0.5401647090911865)),(to_sfixed_a(0.2364727407693863)));

    constant weight_n3_4 : sfixed_bus_array(100 downto 0) := ((to_sfixed_a(0.05248969793319702)),(to_sfixed_a(0.0915345847606659)),(to_sfixed_a(0.2916190028190613)),(to_sfixed_a(0.33772721886634827)),(to_sfixed_a(2.6486821298021823e-05)),(to_sfixed_a(6.425958417821676e-05)),(to_sfixed_a(-0.0025257328525185585)),(to_sfixed_a(-0.46359777450561523)),(to_sfixed_a(-0.4825516939163208)),(to_sfixed_a(0.00014830072177574039)),(to_sfixed_a(-0.2759740650653839)),(to_sfixed_a(0.3086990714073181)),(to_sfixed_a(-0.2042360156774521)),(to_sfixed_a(-0.12074330449104309)),(to_sfixed_a(-0.2717209458351135)),(to_sfixed_a(0.16558773815631866)),(to_sfixed_a(-0.28848734498023987)),(to_sfixed_a(-0.26215559244155884)),(to_sfixed_a(-0.08258985728025436)),(to_sfixed_a(0.2629663050174713)),(to_sfixed_a(-0.00019692037312779576)),(to_sfixed_a(-0.02990632876753807)),(to_sfixed_a(0.03329626843333244)),(to_sfixed_a(0.12287761270999908)),(to_sfixed_a(-5.460002284962684e-06)),(to_sfixed_a(0.12163049727678299)),(to_sfixed_a(-0.4509333372116089)),(to_sfixed_a(-0.2749398648738861)),(to_sfixed_a(0.021733593195676804)),(to_sfixed_a(-0.21040409803390503)),(to_sfixed_a(0.3486599326133728)),(to_sfixed_a(-0.6478060483932495)),(to_sfixed_a(0.10598240047693253)),(to_sfixed_a(-0.5556161999702454)),(to_sfixed_a(-0.9547532796859741)),(to_sfixed_a(6.457621930167079e-05)),(to_sfixed_a(0.25997021794319153)),(to_sfixed_a(0.15241797268390656)),(to_sfixed_a(-0.07910297065973282)),(to_sfixed_a(0.02714228630065918)),(to_sfixed_a(-0.25541725754737854)),(to_sfixed_a(0.15588398277759552)),(to_sfixed_a(-0.002540708752349019)),(to_sfixed_a(-0.18216350674629211)),(to_sfixed_a(-0.09539999067783356)),(to_sfixed_a(0.385105699300766)),(to_sfixed_a(0.07795794308185577)),(to_sfixed_a(0.18089048564434052)),(to_sfixed_a(0.18061600625514984)),(to_sfixed_a(-0.9778957366943359)),(to_sfixed_a(0.3276362121105194)),(to_sfixed_a(-0.15530027449131012)),(to_sfixed_a(-0.2629523277282715)),(to_sfixed_a(0.3396676778793335)),(to_sfixed_a(-0.5788315534591675)),(to_sfixed_a(-0.3935467600822449)),(to_sfixed_a(0.23374144732952118)),(to_sfixed_a(0.46429702639579773)),(to_sfixed_a(0.44421273469924927)),(to_sfixed_a(-0.04402035102248192)),(to_sfixed_a(0.2587847411632538)),(to_sfixed_a(0.06265582889318466)),(to_sfixed_a(0.14803391695022583)),(to_sfixed_a(-0.3387676179409027)),(to_sfixed_a(0.24620331823825836)),(to_sfixed_a(0.2281365543603897)),(to_sfixed_a(0.2525556981563568)),(to_sfixed_a(6.958001176826656e-05)),(to_sfixed_a(-0.16644319891929626)),(to_sfixed_a(0.013551031239330769)),(to_sfixed_a(-0.046899717301130295)),(to_sfixed_a(-0.8177963495254517)),(to_sfixed_a(-0.22364066541194916)),(to_sfixed_a(-0.47321367263793945)),(to_sfixed_a(0.30501970648765564)),(to_sfixed_a(-0.7205824255943298)),(to_sfixed_a(-0.24807138741016388)),(to_sfixed_a(-0.4121374189853668)),(to_sfixed_a(-0.27612608671188354)),(to_sfixed_a(0.3604657053947449)),(to_sfixed_a(0.4128926396369934)),(to_sfixed_a(0.006296674255281687)),(to_sfixed_a(0.6281859278678894)),(to_sfixed_a(-0.42006057500839233)),(to_sfixed_a(0.0001163178458227776)),(to_sfixed_a(-0.7507311105728149)),(to_sfixed_a(-1.0762388706207275)),(to_sfixed_a(-0.1773327887058258)),(to_sfixed_a(0.370973140001297)),(to_sfixed_a(0.25042128562927246)),(to_sfixed_a(-0.0002457096124999225)),(to_sfixed_a(0.09743745625019073)),(to_sfixed_a(-0.30849528312683105)),(to_sfixed_a(-0.24610871076583862)),(to_sfixed_a(0.11763749271631241)),(to_sfixed_a(-1.0446208762004972e-05)),(to_sfixed_a(0.3324810564517975)),(to_sfixed_a(0.5371590256690979)),(to_sfixed_a(-0.2658017873764038)),(to_sfixed_a(-0.1047181636095047)),(to_sfixed_a(0.19366022944450378)));

    constant weight_n3_5 : sfixed_bus_array(100 downto 0) := ((to_sfixed_a(-0.24494393169879913)),(to_sfixed_a(0.14721466600894928)),(to_sfixed_a(0.00734536349773407)),(to_sfixed_a(-0.3840744197368622)),(to_sfixed_a(-2.728057006606832e-05)),(to_sfixed_a(6.16060133324936e-05)),(to_sfixed_a(-0.07649382203817368)),(to_sfixed_a(0.014320873655378819)),(to_sfixed_a(-0.03622042387723923)),(to_sfixed_a(0.00011229767551412806)),(to_sfixed_a(-0.595202624797821)),(to_sfixed_a(0.27501192688941956)),(to_sfixed_a(0.026873312890529633)),(to_sfixed_a(-0.4984382092952728)),(to_sfixed_a(-0.2328297644853592)),(to_sfixed_a(-0.0008734696311876178)),(to_sfixed_a(0.4641610085964203)),(to_sfixed_a(0.019160035997629166)),(to_sfixed_a(-0.7108851671218872)),(to_sfixed_a(-0.5213403701782227)),(to_sfixed_a(1.521624653832987e-06)),(to_sfixed_a(0.06347030401229858)),(to_sfixed_a(0.39885690808296204)),(to_sfixed_a(0.3820946216583252)),(to_sfixed_a(7.708804332651198e-07)),(to_sfixed_a(0.17051757872104645)),(to_sfixed_a(0.1393313854932785)),(to_sfixed_a(0.2623165249824524)),(to_sfixed_a(0.003976140171289444)),(to_sfixed_a(-0.016391010954976082)),(to_sfixed_a(-0.3719802498817444)),(to_sfixed_a(-0.31657013297080994)),(to_sfixed_a(-0.2329099178314209)),(to_sfixed_a(0.018302643671631813)),(to_sfixed_a(0.5150874853134155)),(to_sfixed_a(0.00044294889084994793)),(to_sfixed_a(-0.3044734299182892)),(to_sfixed_a(-0.03400295600295067)),(to_sfixed_a(0.5426263213157654)),(to_sfixed_a(0.501980185508728)),(to_sfixed_a(0.0745469480752945)),(to_sfixed_a(0.3559316396713257)),(to_sfixed_a(-0.11426171660423279)),(to_sfixed_a(-0.2922905683517456)),(to_sfixed_a(0.41940823197364807)),(to_sfixed_a(-0.2416885793209076)),(to_sfixed_a(0.187583789229393)),(to_sfixed_a(-0.5527265667915344)),(to_sfixed_a(-1.0702999830245972)),(to_sfixed_a(0.17523641884326935)),(to_sfixed_a(0.3886815905570984)),(to_sfixed_a(0.3771229088306427)),(to_sfixed_a(0.4537293314933777)),(to_sfixed_a(-0.7813844680786133)),(to_sfixed_a(-0.5304717421531677)),(to_sfixed_a(0.1346733272075653)),(to_sfixed_a(0.006847635842859745)),(to_sfixed_a(-0.16929173469543457)),(to_sfixed_a(-0.9254948496818542)),(to_sfixed_a(-0.2475799024105072)),(to_sfixed_a(-0.4278689920902252)),(to_sfixed_a(-0.1107986718416214)),(to_sfixed_a(0.06748627871274948)),(to_sfixed_a(0.4323270916938782)),(to_sfixed_a(0.055334046483039856)),(to_sfixed_a(-0.0683533325791359)),(to_sfixed_a(-0.38989436626434326)),(to_sfixed_a(-4.3840027501573786e-05)),(to_sfixed_a(-0.6730365753173828)),(to_sfixed_a(-0.0030950915534049273)),(to_sfixed_a(-0.5787881016731262)),(to_sfixed_a(0.01953776367008686)),(to_sfixed_a(-0.4403042197227478)),(to_sfixed_a(0.12239938229322433)),(to_sfixed_a(0.11202526837587357)),(to_sfixed_a(-0.25240007042884827)),(to_sfixed_a(0.18485617637634277)),(to_sfixed_a(0.22447086870670319)),(to_sfixed_a(-0.2968589961528778)),(to_sfixed_a(-0.22458641231060028)),(to_sfixed_a(0.21375620365142822)),(to_sfixed_a(-0.4261672794818878)),(to_sfixed_a(-0.5585716962814331)),(to_sfixed_a(0.29642730951309204)),(to_sfixed_a(0.00025500921765342355)),(to_sfixed_a(0.04367583617568016)),(to_sfixed_a(0.26387014985084534)),(to_sfixed_a(0.35392066836357117)),(to_sfixed_a(0.49298742413520813)),(to_sfixed_a(0.1165127381682396)),(to_sfixed_a(-6.414762901840732e-05)),(to_sfixed_a(0.24620625376701355)),(to_sfixed_a(0.20493052899837494)),(to_sfixed_a(-0.18867413699626923)),(to_sfixed_a(0.35200372338294983)),(to_sfixed_a(0.00012882670853286982)),(to_sfixed_a(-0.7504703402519226)),(to_sfixed_a(0.07796712964773178)),(to_sfixed_a(-0.43867260217666626)),(to_sfixed_a(0.12420059740543365)),(to_sfixed_a(0.1756058633327484)));

    constant weight_n3_6 : sfixed_bus_array(100 downto 0) := ((to_sfixed_a(0.03408895805478096)),(to_sfixed_a(-0.00952710397541523)),(to_sfixed_a(-0.6830865144729614)),(to_sfixed_a(-0.5927482843399048)),(to_sfixed_a(3.407953045098111e-05)),(to_sfixed_a(0.0001317444402957335)),(to_sfixed_a(0.36434754729270935)),(to_sfixed_a(-0.32223939895629883)),(to_sfixed_a(-0.4257223904132843)),(to_sfixed_a(0.00021595902217086405)),(to_sfixed_a(-0.07782499492168427)),(to_sfixed_a(0.11613515764474869)),(to_sfixed_a(0.023617273196578026)),(to_sfixed_a(1.8393080608802848e-05)),(to_sfixed_a(-0.04401237890124321)),(to_sfixed_a(-0.35573700070381165)),(to_sfixed_a(-0.19760455191135406)),(to_sfixed_a(-0.9594861268997192)),(to_sfixed_a(-0.8114367127418518)),(to_sfixed_a(-0.25539663434028625)),(to_sfixed_a(-5.7213386753574014e-05)),(to_sfixed_a(-0.19715313613414764)),(to_sfixed_a(0.1974637806415558)),(to_sfixed_a(-0.1164369136095047)),(to_sfixed_a(-0.00029082331457175314)),(to_sfixed_a(-1.1138505935668945)),(to_sfixed_a(-0.09090390056371689)),(to_sfixed_a(-0.38808223605155945)),(to_sfixed_a(0.2140834927558899)),(to_sfixed_a(0.2524182200431824)),(to_sfixed_a(0.5355889201164246)),(to_sfixed_a(-0.22521501779556274)),(to_sfixed_a(0.15419092774391174)),(to_sfixed_a(0.2693191170692444)),(to_sfixed_a(0.28480276465415955)),(to_sfixed_a(0.00017919926904141903)),(to_sfixed_a(-0.017594249919056892)),(to_sfixed_a(0.014638882130384445)),(to_sfixed_a(0.15776585042476654)),(to_sfixed_a(-0.3775596618652344)),(to_sfixed_a(-0.018925737589597702)),(to_sfixed_a(0.20183825492858887)),(to_sfixed_a(-1.4746898159501143e-05)),(to_sfixed_a(0.21576376259326935)),(to_sfixed_a(0.39930105209350586)),(to_sfixed_a(-0.7555854916572571)),(to_sfixed_a(-0.27038466930389404)),(to_sfixed_a(0.2454451471567154)),(to_sfixed_a(-0.38118377327919006)),(to_sfixed_a(-0.04280134662985802)),(to_sfixed_a(0.19717897474765778)),(to_sfixed_a(0.3862743079662323)),(to_sfixed_a(-0.15444038808345795)),(to_sfixed_a(-0.99162757396698)),(to_sfixed_a(0.3088991641998291)),(to_sfixed_a(0.2369721680879593)),(to_sfixed_a(0.20182016491889954)),(to_sfixed_a(0.48561355471611023)),(to_sfixed_a(-0.5401318669319153)),(to_sfixed_a(0.06158645451068878)),(to_sfixed_a(0.4007931649684906)),(to_sfixed_a(-0.05398125201463699)),(to_sfixed_a(0.36335489153862)),(to_sfixed_a(-0.2719925343990326)),(to_sfixed_a(0.25011855363845825)),(to_sfixed_a(-0.30000725388526917)),(to_sfixed_a(0.3284212350845337)),(to_sfixed_a(-3.9972044760361314e-05)),(to_sfixed_a(-0.19173240661621094)),(to_sfixed_a(-0.017773183062672615)),(to_sfixed_a(-0.3297441005706787)),(to_sfixed_a(0.10729890316724777)),(to_sfixed_a(-0.49014759063720703)),(to_sfixed_a(0.3269561529159546)),(to_sfixed_a(0.002884868299588561)),(to_sfixed_a(-0.6571505069732666)),(to_sfixed_a(0.20266802608966827)),(to_sfixed_a(0.2871066927909851)),(to_sfixed_a(-0.1732713282108307)),(to_sfixed_a(0.48339781165122986)),(to_sfixed_a(-0.4797428250312805)),(to_sfixed_a(0.4140034317970276)),(to_sfixed_a(-0.1770997941493988)),(to_sfixed_a(0.3572477698326111)),(to_sfixed_a(0.00016514002345502377)),(to_sfixed_a(0.3510878384113312)),(to_sfixed_a(0.16838419437408447)),(to_sfixed_a(-0.9166480302810669)),(to_sfixed_a(-0.4803932011127472)),(to_sfixed_a(0.040730200707912445)),(to_sfixed_a(-0.00011364171223249286)),(to_sfixed_a(-0.2602718472480774)),(to_sfixed_a(-0.1155131533741951)),(to_sfixed_a(0.32994014024734497)),(to_sfixed_a(-0.43216201663017273)),(to_sfixed_a(-1.6797399439383298e-05)),(to_sfixed_a(-0.06987618654966354)),(to_sfixed_a(-0.21835310757160187)),(to_sfixed_a(0.17840056121349335)),(to_sfixed_a(0.0029421327635645866)),(to_sfixed_a(-0.8953529596328735)));

    constant weight_n3_7 : sfixed_bus_array(100 downto 0) := ((to_sfixed_a(-0.3414101004600525)),(to_sfixed_a(0.28119945526123047)),(to_sfixed_a(0.2067217081785202)),(to_sfixed_a(-0.2177887260913849)),(to_sfixed_a(0.00016770962974987924)),(to_sfixed_a(-9.070852684089914e-05)),(to_sfixed_a(-0.20015883445739746)),(to_sfixed_a(0.06850757449865341)),(to_sfixed_a(-0.7282559275627136)),(to_sfixed_a(-0.000161607182235457)),(to_sfixed_a(0.437915563583374)),(to_sfixed_a(-0.4691062271595001)),(to_sfixed_a(-1.1563191413879395)),(to_sfixed_a(0.7187780737876892)),(to_sfixed_a(-0.34266817569732666)),(to_sfixed_a(0.14933770895004272)),(to_sfixed_a(-0.20464731752872467)),(to_sfixed_a(-0.22180813550949097)),(to_sfixed_a(-0.0069189234636723995)),(to_sfixed_a(0.34597837924957275)),(to_sfixed_a(-6.826667231507599e-07)),(to_sfixed_a(0.07217399030923843)),(to_sfixed_a(-0.33571934700012207)),(to_sfixed_a(0.14620772004127502)),(to_sfixed_a(-0.00010359084990341216)),(to_sfixed_a(0.35833024978637695)),(to_sfixed_a(0.14358912408351898)),(to_sfixed_a(0.1181216612458229)),(to_sfixed_a(0.00025058252504095435)),(to_sfixed_a(0.07321150600910187)),(to_sfixed_a(-0.5117992758750916)),(to_sfixed_a(-0.34880736470222473)),(to_sfixed_a(0.33425748348236084)),(to_sfixed_a(-0.35027381777763367)),(to_sfixed_a(-0.542334258556366)),(to_sfixed_a(3.716207720572129e-05)),(to_sfixed_a(0.2882145345211029)),(to_sfixed_a(0.0008713702554814517)),(to_sfixed_a(0.19732359051704407)),(to_sfixed_a(0.4369317889213562)),(to_sfixed_a(0.3770480751991272)),(to_sfixed_a(-0.37310782074928284)),(to_sfixed_a(5.4984866437735036e-05)),(to_sfixed_a(0.031887177377939224)),(to_sfixed_a(0.4237240254878998)),(to_sfixed_a(-0.6794252395629883)),(to_sfixed_a(-0.856515645980835)),(to_sfixed_a(0.28310060501098633)),(to_sfixed_a(0.2734401822090149)),(to_sfixed_a(-0.5926557779312134)),(to_sfixed_a(-1.0748432874679565)),(to_sfixed_a(0.29376304149627686)),(to_sfixed_a(0.02322430908679962)),(to_sfixed_a(0.2778467833995819)),(to_sfixed_a(0.1130412369966507)),(to_sfixed_a(0.20826850831508636)),(to_sfixed_a(0.0051545328460633755)),(to_sfixed_a(-0.490401953458786)),(to_sfixed_a(-0.20815199613571167)),(to_sfixed_a(-0.21031306684017181)),(to_sfixed_a(-1.13694429397583)),(to_sfixed_a(0.09881105273962021)),(to_sfixed_a(0.4377237856388092)),(to_sfixed_a(-0.7901729941368103)),(to_sfixed_a(-0.22944553196430206)),(to_sfixed_a(0.34418484568595886)),(to_sfixed_a(-0.308906614780426)),(to_sfixed_a(-5.536498065339401e-06)),(to_sfixed_a(0.02599085122346878)),(to_sfixed_a(-0.262637734413147)),(to_sfixed_a(0.10064568370580673)),(to_sfixed_a(0.2496112734079361)),(to_sfixed_a(-0.020405398681759834)),(to_sfixed_a(0.16745436191558838)),(to_sfixed_a(-0.3331564664840698)),(to_sfixed_a(0.23516377806663513)),(to_sfixed_a(0.2250065952539444)),(to_sfixed_a(-0.1007133349776268)),(to_sfixed_a(0.377093642950058)),(to_sfixed_a(-0.32263079285621643)),(to_sfixed_a(0.49280813336372375)),(to_sfixed_a(0.15369336307048798)),(to_sfixed_a(-0.029999645426869392)),(to_sfixed_a(-0.24622566998004913)),(to_sfixed_a(4.4094638724345714e-05)),(to_sfixed_a(0.026212241500616074)),(to_sfixed_a(0.3221421539783478)),(to_sfixed_a(0.2574298083782196)),(to_sfixed_a(-0.4809767007827759)),(to_sfixed_a(-1.0462443828582764)),(to_sfixed_a(6.472489621955901e-05)),(to_sfixed_a(0.2141096293926239)),(to_sfixed_a(0.043769557029008865)),(to_sfixed_a(-0.18326495587825775)),(to_sfixed_a(-0.40406283736228943)),(to_sfixed_a(-6.366703019011766e-05)),(to_sfixed_a(0.4005279242992401)),(to_sfixed_a(0.3955240845680237)),(to_sfixed_a(0.26174160838127136)),(to_sfixed_a(-0.41347768902778625)),(to_sfixed_a(0.14889536798000336)));

    constant weight_n3_8 : sfixed_bus_array(100 downto 0) := ((to_sfixed_a(0.6426519155502319)),(to_sfixed_a(-0.8405122756958008)),(to_sfixed_a(0.01940959319472313)),(to_sfixed_a(-0.44530731439590454)),(to_sfixed_a(-4.247848119121045e-05)),(to_sfixed_a(0.00021916523110121489)),(to_sfixed_a(0.3019644021987915)),(to_sfixed_a(0.30512282252311707)),(to_sfixed_a(0.46171170473098755)),(to_sfixed_a(0.0003114459686912596)),(to_sfixed_a(-0.16895395517349243)),(to_sfixed_a(-0.27391284704208374)),(to_sfixed_a(0.02029799483716488)),(to_sfixed_a(-0.9821906089782715)),(to_sfixed_a(0.2857450842857361)),(to_sfixed_a(-0.0695529505610466)),(to_sfixed_a(0.3304980397224426)),(to_sfixed_a(-0.027420923113822937)),(to_sfixed_a(0.22261051833629608)),(to_sfixed_a(0.37585899233818054)),(to_sfixed_a(3.080338137806393e-05)),(to_sfixed_a(0.08669039607048035)),(to_sfixed_a(0.37382417917251587)),(to_sfixed_a(-0.43126749992370605)),(to_sfixed_a(-1.2853633961640298e-05)),(to_sfixed_a(-0.07006387412548065)),(to_sfixed_a(0.18412216007709503)),(to_sfixed_a(0.001248365850187838)),(to_sfixed_a(0.216574564576149)),(to_sfixed_a(0.18046694993972778)),(to_sfixed_a(-0.7076109647750854)),(to_sfixed_a(-0.047408200800418854)),(to_sfixed_a(-0.6070911884307861)),(to_sfixed_a(0.027549346908926964)),(to_sfixed_a(-0.32167261838912964)),(to_sfixed_a(-2.2527514374814928e-05)),(to_sfixed_a(-0.2334016114473343)),(to_sfixed_a(-0.5927971005439758)),(to_sfixed_a(-0.4435617923736572)),(to_sfixed_a(-0.05552647262811661)),(to_sfixed_a(-0.43915677070617676)),(to_sfixed_a(-0.08156965672969818)),(to_sfixed_a(6.912188837304711e-05)),(to_sfixed_a(0.18611660599708557)),(to_sfixed_a(-0.07514756172895432)),(to_sfixed_a(0.4014458954334259)),(to_sfixed_a(-0.2695533037185669)),(to_sfixed_a(-0.992247998714447)),(to_sfixed_a(0.3249672055244446)),(to_sfixed_a(0.15989115834236145)),(to_sfixed_a(0.008378442376852036)),(to_sfixed_a(-0.26200857758522034)),(to_sfixed_a(-1.0758588314056396)),(to_sfixed_a(-0.12515823543071747)),(to_sfixed_a(0.26756206154823303)),(to_sfixed_a(0.37329092621803284)),(to_sfixed_a(0.38196679949760437)),(to_sfixed_a(0.3756644129753113)),(to_sfixed_a(0.2092021107673645)),(to_sfixed_a(0.1987428069114685)),(to_sfixed_a(0.2595367431640625)),(to_sfixed_a(-0.4876076281070709)),(to_sfixed_a(-0.4810134768486023)),(to_sfixed_a(-0.7269073724746704)),(to_sfixed_a(-0.30437830090522766)),(to_sfixed_a(-0.2972984313964844)),(to_sfixed_a(-0.23549513518810272)),(to_sfixed_a(-9.095383575186133e-07)),(to_sfixed_a(-0.25565049052238464)),(to_sfixed_a(-0.3651729226112366)),(to_sfixed_a(-0.47237348556518555)),(to_sfixed_a(-0.10354266315698624)),(to_sfixed_a(0.0656202957034111)),(to_sfixed_a(-0.08846694231033325)),(to_sfixed_a(-0.08334402740001678)),(to_sfixed_a(-0.28231891989707947)),(to_sfixed_a(0.2244614213705063)),(to_sfixed_a(0.03076845034956932)),(to_sfixed_a(0.32831379771232605)),(to_sfixed_a(-0.047479767352342606)),(to_sfixed_a(-0.42202526330947876)),(to_sfixed_a(0.3184395432472229)),(to_sfixed_a(0.5072726607322693)),(to_sfixed_a(0.3646731972694397)),(to_sfixed_a(0.0001474782038712874)),(to_sfixed_a(0.06357524544000626)),(to_sfixed_a(0.3399309813976288)),(to_sfixed_a(-0.08719035238027573)),(to_sfixed_a(-0.700587272644043)),(to_sfixed_a(0.04022608697414398)),(to_sfixed_a(6.111963011790067e-05)),(to_sfixed_a(0.2855077385902405)),(to_sfixed_a(0.1893940567970276)),(to_sfixed_a(0.21168562769889832)),(to_sfixed_a(0.49429643154144287)),(to_sfixed_a(-0.0004119219374842942)),(to_sfixed_a(-0.41652923822402954)),(to_sfixed_a(-0.4837641716003418)),(to_sfixed_a(-0.8213343620300293)),(to_sfixed_a(0.3793204724788666)),(to_sfixed_a(0.35834261775016785)));

    constant weight_n3_9 : sfixed_bus_array(100 downto 0) := ((to_sfixed_a(0.08569824695587158)),(to_sfixed_a(0.3506328761577606)),(to_sfixed_a(-0.11578129976987839)),(to_sfixed_a(0.23575517535209656)),(to_sfixed_a(0.00015071041707415134)),(to_sfixed_a(-0.00010133082105312496)),(to_sfixed_a(0.3998717963695526)),(to_sfixed_a(0.22007504105567932)),(to_sfixed_a(-0.6375741958618164)),(to_sfixed_a(6.225862307474017e-05)),(to_sfixed_a(-1.1131325960159302)),(to_sfixed_a(0.35999006032943726)),(to_sfixed_a(0.31174883246421814)),(to_sfixed_a(-0.40139317512512207)),(to_sfixed_a(-0.4858134090900421)),(to_sfixed_a(0.03995184227824211)),(to_sfixed_a(0.11807803064584732)),(to_sfixed_a(0.3383883237838745)),(to_sfixed_a(0.3151725232601166)),(to_sfixed_a(0.3039608299732208)),(to_sfixed_a(2.7636997401714325e-06)),(to_sfixed_a(-0.6699275970458984)),(to_sfixed_a(-0.43309593200683594)),(to_sfixed_a(0.1648501455783844)),(to_sfixed_a(-7.382650801446289e-05)),(to_sfixed_a(0.35187846422195435)),(to_sfixed_a(0.06682047247886658)),(to_sfixed_a(0.037500523030757904)),(to_sfixed_a(0.001487975474447012)),(to_sfixed_a(0.49931785464286804)),(to_sfixed_a(0.38299375772476196)),(to_sfixed_a(0.07180514186620712)),(to_sfixed_a(-0.07713834196329117)),(to_sfixed_a(-0.5745607018470764)),(to_sfixed_a(-0.049347881227731705)),(to_sfixed_a(-0.0001655307860346511)),(to_sfixed_a(0.2819756269454956)),(to_sfixed_a(0.2544442117214203)),(to_sfixed_a(-0.5417556762695312)),(to_sfixed_a(0.08936959505081177)),(to_sfixed_a(0.4612025022506714)),(to_sfixed_a(-1.1338969469070435)),(to_sfixed_a(0.0536949560046196)),(to_sfixed_a(-0.015646716579794884)),(to_sfixed_a(-0.4831271469593048)),(to_sfixed_a(0.33968836069107056)),(to_sfixed_a(0.21940365433692932)),(to_sfixed_a(0.3366902470588684)),(to_sfixed_a(0.16800245642662048)),(to_sfixed_a(0.0542965866625309)),(to_sfixed_a(-0.5240541100502014)),(to_sfixed_a(-0.3843759298324585)),(to_sfixed_a(0.20069536566734314)),(to_sfixed_a(0.04169082269072533)),(to_sfixed_a(-0.007219257764518261)),(to_sfixed_a(0.23004558682441711)),(to_sfixed_a(0.058047596365213394)),(to_sfixed_a(0.33906909823417664)),(to_sfixed_a(0.22176560759544373)),(to_sfixed_a(-0.8153958320617676)),(to_sfixed_a(-0.030045580118894577)),(to_sfixed_a(0.7424807548522949)),(to_sfixed_a(0.22817817330360413)),(to_sfixed_a(0.2230636179447174)),(to_sfixed_a(0.15959182381629944)),(to_sfixed_a(0.3090600371360779)),(to_sfixed_a(-0.5989579558372498)),(to_sfixed_a(-0.00037717242958024144)),(to_sfixed_a(0.33674532175064087)),(to_sfixed_a(-0.004859771579504013)),(to_sfixed_a(0.3260008692741394)),(to_sfixed_a(-0.11325535923242569)),(to_sfixed_a(-0.14174386858940125)),(to_sfixed_a(-0.03705822303891182)),(to_sfixed_a(0.1057250127196312)),(to_sfixed_a(-0.13635662198066711)),(to_sfixed_a(-0.07893925160169601)),(to_sfixed_a(-0.6314873695373535)),(to_sfixed_a(-0.05060531198978424)),(to_sfixed_a(-0.5609336495399475)),(to_sfixed_a(-0.6941792964935303)),(to_sfixed_a(-0.8229686617851257)),(to_sfixed_a(-0.7862907648086548)),(to_sfixed_a(-0.5048548579216003)),(to_sfixed_a(7.021768396953121e-05)),(to_sfixed_a(0.18110206723213196)),(to_sfixed_a(-0.38241344690322876)),(to_sfixed_a(0.2872520983219147)),(to_sfixed_a(0.28659647703170776)),(to_sfixed_a(0.011108818463981152)),(to_sfixed_a(3.318168455734849e-05)),(to_sfixed_a(0.23555833101272583)),(to_sfixed_a(-0.04785829782485962)),(to_sfixed_a(0.08290141075849533)),(to_sfixed_a(0.19211067259311676)),(to_sfixed_a(-0.00018402133719064295)),(to_sfixed_a(-0.013119801878929138)),(to_sfixed_a(-0.7500252723693848)),(to_sfixed_a(-0.47694161534309387)),(to_sfixed_a(-0.05029291659593582)),(to_sfixed_a(0.1416090428829193)));




end package weights_constants;
