

package model_weights;


logic signed [31:0] VT_0 [37][37] ='{
{32'h80000000 , 32'h00000070 , 32'hFFFFFFB3 , 32'h0000004A , 32'h00000006 , 32'hFFFFFFFA , 32'h00000019 , 32'hFFFFFFF4 , 32'h00000017 , 32'h00000007 , 32'hFFFFFFFF , 32'hFFFFFFFB , 32'h00000005 , 32'h00000000 , 32'hFFFFFFFD , 32'h00000004 , 32'hFFFFFFFF , 32'h00000002 , 32'h00000005 , 32'hFFFFFFF4 , 32'h00000000 , 32'hFFFFFFFB , 32'hFFFFFFFE , 32'h00000000 , 32'hFFFFFFFD , 32'h0000000A , 32'h00000003 , 32'hFFFFFFF3 , 32'h00000001 , 32'hFFFFFFF9 , 32'h00000005 , 32'h00000000 , 32'h00000005 , 32'h00000000 , 32'hFFFFFFFC , 32'h00000002 , 32'h00000000} , 
{32'h00000070 , 32'h80000000 , 32'hFFFFFFF0 , 32'h0000000A , 32'h00000047 , 32'h00000029 , 32'h0000001B , 32'h00000005 , 32'hFFFFFFF0 , 32'h00000000 , 32'hFFFFFFFB , 32'hFFFFFFEC , 32'h00000000 , 32'h00000007 , 32'h00000009 , 32'h0000000A , 32'hFFFFFFFE , 32'h00000003 , 32'h00000009 , 32'h00000009 , 32'hFFFFFFFB , 32'h00000001 , 32'hFFFFFFFA , 32'hFFFFFFFE , 32'hFFFFFFFF , 32'hFFFFFFF6 , 32'hFFFFFFFC , 32'h00000000 , 32'h00000000 , 32'hFFFFFFFF , 32'h00000000 , 32'h00000005 , 32'hFFFFFFF9 , 32'hFFFFFFF3 , 32'hFFFFFFF8 , 32'h00000007 , 32'hFFFFFFFD} , 
{32'hFFFFFFB3 , 32'h0000000E , 32'h80000000 , 32'h00000085 , 32'hFFFFFF88 , 32'h0000004F , 32'hFFFFFFF6 , 32'h0000000C , 32'hFFFFFFF9 , 32'h0000000A , 32'hFFFFFFEC , 32'h0000000B , 32'hFFFFFFF8 , 32'hFFFFFFFB , 32'h00000009 , 32'h00000012 , 32'h00000010 , 32'hFFFFFFEB , 32'hFFFFFFF0 , 32'hFFFFFFFD , 32'hFFFFFFF9 , 32'h00000003 , 32'h00000000 , 32'h00000000 , 32'h00000005 , 32'hFFFFFFF4 , 32'hFFFFFFF3 , 32'hFFFFFFFE , 32'h00000002 , 32'hFFFFFFF7 , 32'hFFFFFFFF , 32'h00000004 , 32'h00000008 , 32'hFFFFFFFD , 32'hFFFFFFFE , 32'hFFFFFFFC , 32'hFFFFFFFD} , 
{32'h0000004A , 32'hFFFFFFF4 , 32'hFFFFFF79 , 32'h80000000 , 32'h000000B7 , 32'hFFFFFF76 , 32'hFFFFFFA3 , 32'hFFFFFFFF , 32'hFFFFFFF1 , 32'h0000001E , 32'h00000009 , 32'hFFFFFFEF , 32'h0000000A , 32'h00000005 , 32'hFFFFFFFB , 32'hFFFFFFE4 , 32'hFFFFFFFC , 32'hFFFFFFF4 , 32'hFFFFFFFD , 32'hFFFFFFFF , 32'h00000013 , 32'h00000003 , 32'h00000005 , 32'hFFFFFFF5 , 32'hFFFFFFF6 , 32'h00000004 , 32'h0000000A , 32'h00000004 , 32'h00000008 , 32'hFFFFFFFB , 32'h0000000B , 32'hFFFFFFFE , 32'h00000000 , 32'hFFFFFFFC , 32'hFFFFFFFB , 32'h00000000 , 32'hFFFFFFFC} , 
{32'hFFFFFFF8 , 32'h00000047 , 32'hFFFFFF88 , 32'h000000B7 , 32'h80000000 , 32'hFFFFFDDE , 32'hFFFFFFF7 , 32'hFFFFFFF9 , 32'h0000000A , 32'hFFFFFFE0 , 32'hFFFFFFE5 , 32'hFFFFFFE1 , 32'h00000000 , 32'h00000001 , 32'h00000001 , 32'hFFFFFFF0 , 32'h0000000C , 32'hFFFFFFFF , 32'hFFFFFFF7 , 32'hFFFFFFFD , 32'h00000002 , 32'hFFFFFFFA , 32'hFFFFFFFB , 32'hFFFFFFFD , 32'hFFFFFFF7 , 32'hFFFFFFFD , 32'h00000000 , 32'hFFFFFFFB , 32'hFFFFFFF9 , 32'h00000004 , 32'h00000000 , 32'hFFFFFFFE , 32'hFFFFFFFB , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'hFFFFFFF7} , 
{32'h00000004 , 32'h00000029 , 32'h0000004F , 32'hFFFFFF76 , 32'h00000220 , 32'h80000000 , 32'h0000000F , 32'hFFFFFFEC , 32'hFFFFFFF7 , 32'h00000006 , 32'hFFFFFFC8 , 32'hFFFFFFF1 , 32'hFFFFFFFD , 32'hFFFFFFF0 , 32'h00000009 , 32'h0000001F , 32'h0000000E , 32'hFFFFFFFE , 32'h00000006 , 32'h00000000 , 32'hFFFFFFFE , 32'hFFFFFFFB , 32'hFFFFFFFE , 32'h00000002 , 32'hFFFFFFFE , 32'hFFFFFFFA , 32'hFFFFFFFF , 32'h00000004 , 32'h00000001 , 32'hFFFFFFFB , 32'hFFFFFFFA , 32'hFFFFFFFF , 32'h00000000 , 32'h00000008 , 32'h00000003 , 32'h00000000 , 32'h00000001} , 
{32'hFFFFFFE5 , 32'h0000001B , 32'hFFFFFFF6 , 32'hFFFFFFA3 , 32'h00000007 , 32'hFFFFFFEF , 32'h80000000 , 32'h00000024 , 32'hFFFFFFEE , 32'h00000003 , 32'h00000000 , 32'h00000004 , 32'h00000000 , 32'hFFFFFFDD , 32'hFFFFFFE3 , 32'h00000003 , 32'hFFFFFFF1 , 32'h00000018 , 32'hFFFFFFFC , 32'hFFFFFFFB , 32'h00000006 , 32'hFFFFFFF8 , 32'hFFFFFFFD , 32'h00000006 , 32'h00000007 , 32'hFFFFFFFB , 32'hFFFFFFF7 , 32'h00000004 , 32'h0000000F , 32'h00000004 , 32'hFFFFFFF7 , 32'h00000000 , 32'hFFFFFFFE , 32'h00000002 , 32'hFFFFFFF3 , 32'h00000001 , 32'hFFFFFFFA} , 
{32'h0000000A , 32'h00000005 , 32'h0000000C , 32'hFFFFFFFF , 32'h00000005 , 32'h00000012 , 32'hFFFFFFDA , 32'h80000000 , 32'h00000015 , 32'h00000025 , 32'hFFFFFFC3 , 32'hFFFFFFF5 , 32'h00000014 , 32'hFFFFFFEF , 32'hFFFFFFD9 , 32'hFFFFFFF8 , 32'hFFFFFFEB , 32'h0000000D , 32'h00000004 , 32'hFFFFFFE6 , 32'hFFFFFFF1 , 32'hFFFFFFEE , 32'hFFFFFFF7 , 32'hFFFFFFEF , 32'h00000002 , 32'h00000016 , 32'hFFFFFFE7 , 32'h00000002 , 32'h00000008 , 32'h00000000 , 32'hFFFFFFFA , 32'hFFFFFFFB , 32'h00000004 , 32'h00000001 , 32'hFFFFFFF5 , 32'h0000000A , 32'h00000004} , 
{32'hFFFFFFE7 , 32'hFFFFFFF0 , 32'hFFFFFFF9 , 32'hFFFFFFF1 , 32'hFFFFFFF4 , 32'h00000007 , 32'h00000010 , 32'hFFFFFFE9 , 32'h80000000 , 32'h0000009A , 32'h00000090 , 32'h0000001E , 32'hFFFFFFF1 , 32'hFFFFFFEE , 32'h00000008 , 32'hFFFFFFE7 , 32'h00000014 , 32'hFFFFFFF7 , 32'h00000019 , 32'h0000000F , 32'h0000000A , 32'hFFFFFFFD , 32'hFFFFFFFB , 32'h00000015 , 32'h0000000B , 32'hFFFFFFFF , 32'h00000016 , 32'h0000000F , 32'h0000000C , 32'hFFFFFFF7 , 32'hFFFFFFFE , 32'h0000000A , 32'h00000000 , 32'hFFFFFFFC , 32'h00000000 , 32'hFFFFFFFC , 32'hFFFFFFFB} , 
{32'h00000007 , 32'hFFFFFFFF , 32'hFFFFFFF4 , 32'hFFFFFFE0 , 32'hFFFFFFE0 , 32'h00000006 , 32'h00000003 , 32'h00000025 , 32'h0000009A , 32'h80000000 , 32'hFFFFFF12 , 32'hFFFFFFB2 , 32'h00000027 , 32'h00000053 , 32'hFFFFFFFD , 32'h00000001 , 32'hFFFFFFFE , 32'hFFFFFFFA , 32'hFFFFFFE9 , 32'hFFFFFFDE , 32'h00000014 , 32'hFFFFFFF8 , 32'h00000005 , 32'hFFFFFFD6 , 32'h00000000 , 32'hFFFFFFF6 , 32'hFFFFFFF5 , 32'h00000004 , 32'hFFFFFFFD , 32'hFFFFFFF4 , 32'h00000002 , 32'h00000008 , 32'hFFFFFFF3 , 32'hFFFFFFFC , 32'hFFFFFFF3 , 32'h00000000 , 32'h00000007} , 
{32'h00000000 , 32'hFFFFFFFB , 32'hFFFFFFEC , 32'h00000009 , 32'h00000019 , 32'h00000036 , 32'hFFFFFFFE , 32'h0000003B , 32'hFFFFFF6E , 32'hFFFFFF12 , 32'h80000000 , 32'hFFFFFFD7 , 32'hFFFFFFDB , 32'h00000028 , 32'h0000000E , 32'h00000001 , 32'h0000001E , 32'hFFFFFFFA , 32'hFFFFFFF2 , 32'hFFFFFFF7 , 32'h0000000C , 32'h00000015 , 32'h00000002 , 32'hFFFFFFF5 , 32'h00000008 , 32'hFFFFFFFE , 32'h00000012 , 32'h00000001 , 32'h00000002 , 32'hFFFFFFF8 , 32'hFFFFFFFE , 32'h00000000 , 32'hFFFFFFFE , 32'hFFFFFFEF , 32'hFFFFFFF9 , 32'hFFFFFFFD , 32'h00000004} , 
{32'hFFFFFFFB , 32'h00000012 , 32'hFFFFFFF3 , 32'h0000000F , 32'hFFFFFFE1 , 32'hFFFFFFF1 , 32'h00000004 , 32'hFFFFFFF5 , 32'h0000001E , 32'h0000004C , 32'hFFFFFFD7 , 32'h80000000 , 32'hFFFFFFAE , 32'h00000000 , 32'h0000000E , 32'h0000002D , 32'h0000000C , 32'hFFFFFFE0 , 32'h00000020 , 32'hFFFFFFC2 , 32'h00000009 , 32'hFFFFFFEE , 32'h00000016 , 32'hFFFFFFF1 , 32'hFFFFFFFE , 32'hFFFFFFFD , 32'hFFFFFFFA , 32'hFFFFFFF1 , 32'h00000017 , 32'h00000004 , 32'h00000005 , 32'h00000004 , 32'hFFFFFFEB , 32'hFFFFFFFA , 32'hFFFFFFFE , 32'h00000006 , 32'hFFFFFFFF} , 
{32'hFFFFFFF9 , 32'h00000000 , 32'hFFFFFFF8 , 32'h0000000A , 32'hFFFFFFFF , 32'h00000001 , 32'hFFFFFFFE , 32'hFFFFFFEA , 32'h0000000D , 32'h00000027 , 32'h00000023 , 32'hFFFFFFAE , 32'h80000000 , 32'h00000114 , 32'h0000006C , 32'hFFFFFF8C , 32'h00000032 , 32'hFFFFFFF9 , 32'h00000001 , 32'h00000032 , 32'hFFFFFFEC , 32'h0000000A , 32'h00000000 , 32'hFFFFFFFB , 32'h00000000 , 32'h00000017 , 32'hFFFFFFE6 , 32'h0000000A , 32'hFFFFFFFA , 32'h00000004 , 32'hFFFFFFF7 , 32'hFFFFFFF2 , 32'h00000017 , 32'h00000006 , 32'h00000001 , 32'h0000000D , 32'hFFFFFFFC} , 
{32'hFFFFFFFE , 32'h00000007 , 32'hFFFFFFFB , 32'h00000005 , 32'hFFFFFFFD , 32'h0000000E , 32'h00000021 , 32'h0000000F , 32'h00000010 , 32'h00000053 , 32'hFFFFFFD6 , 32'h00000000 , 32'hFFFFFEEA , 32'h80000000 , 32'hFFFFFE80 , 32'h00000032 , 32'h00000049 , 32'h0000001D , 32'hFFFFFFF0 , 32'hFFFFFFBC , 32'h00000023 , 32'h0000001D , 32'h00000000 , 32'hFFFFFFF8 , 32'hFFFFFFFF , 32'h0000000E , 32'h00000007 , 32'hFFFFFFEB , 32'h00000014 , 32'h0000000A , 32'hFFFFFFED , 32'h00000018 , 32'h00000008 , 32'h00000001 , 32'h0000000A , 32'h0000000E , 32'hFFFFFFF6} , 
{32'h00000001 , 32'h00000009 , 32'h00000009 , 32'hFFFFFFFB , 32'hFFFFFFFD , 32'hFFFFFFF5 , 32'h0000001B , 32'h00000025 , 32'hFFFFFFF6 , 32'hFFFFFFFD , 32'hFFFFFFF0 , 32'h0000000E , 32'hFFFFFF92 , 32'h0000017E , 32'h80000000 , 32'hFFFFFFC8 , 32'h0000003A , 32'hFFFFFFE9 , 32'hFFFFFFE7 , 32'hFFFFFFF8 , 32'h0000000C , 32'hFFFFFFE6 , 32'hFFFFFFF3 , 32'hFFFFFFEF , 32'hFFFFFFE1 , 32'h00000006 , 32'hFFFFFFF9 , 32'h00000022 , 32'h00000019 , 32'h0000000C , 32'hFFFFFFFA , 32'hFFFFFFFB , 32'hFFFFFFF9 , 32'h00000000 , 32'hFFFFFFFD , 32'hFFFFFFFB , 32'hFFFFFFF1} , 
{32'h00000004 , 32'hFFFFFFF4 , 32'hFFFFFFEC , 32'h0000001A , 32'hFFFFFFF0 , 32'h0000001F , 32'h00000003 , 32'hFFFFFFF8 , 32'hFFFFFFE7 , 32'hFFFFFFFD , 32'h00000001 , 32'hFFFFFFD1 , 32'hFFFFFF8C , 32'h00000032 , 32'hFFFFFFC8 , 32'h80000000 , 32'hFFFFFF88 , 32'hFFFFFFF8 , 32'hFFFFFFFA , 32'hFFFFFFB7 , 32'h0000001A , 32'hFFFFFFED , 32'hFFFFFFF4 , 32'h0000000B , 32'h00000014 , 32'h00000013 , 32'h00000011 , 32'h00000001 , 32'h00000000 , 32'h00000001 , 32'h00000007 , 32'h00000000 , 32'hFFFFFFF7 , 32'h0000000D , 32'hFFFFFFF5 , 32'hFFFFFFFB , 32'h00000000} , 
{32'h00000000 , 32'hFFFFFFFE , 32'h00000010 , 32'hFFFFFFFC , 32'hFFFFFFF2 , 32'hFFFFFFF0 , 32'h0000000D , 32'h00000013 , 32'hFFFFFFEA , 32'hFFFFFFFE , 32'hFFFFFFE0 , 32'h0000000C , 32'hFFFFFFCC , 32'hFFFFFFB5 , 32'hFFFFFFC4 , 32'hFFFFFF88 , 32'h80000000 , 32'h0000003B , 32'h00000023 , 32'hFFFFFFDD , 32'h0000003B , 32'hFFFFFFC8 , 32'hFFFFFFE1 , 32'h00000007 , 32'hFFFFFFE4 , 32'hFFFFFFED , 32'h0000001B , 32'hFFFFFFF8 , 32'h0000000A , 32'h00000000 , 32'h00000009 , 32'hFFFFFFED , 32'h00000001 , 32'h00000003 , 32'h00000008 , 32'hFFFFFFE9 , 32'h00000018} , 
{32'h00000002 , 32'hFFFFFFFB , 32'h00000013 , 32'h0000000A , 32'hFFFFFFFF , 32'hFFFFFFFE , 32'h00000018 , 32'h0000000D , 32'hFFFFFFF7 , 32'h00000004 , 32'hFFFFFFFA , 32'h0000001E , 32'hFFFFFFF9 , 32'h0000001D , 32'hFFFFFFE9 , 32'h00000006 , 32'h0000003B , 32'h80000000 , 32'h0000007F , 32'hFFFFFFEF , 32'h00000011 , 32'h0000002F , 32'hFFFFFFF6 , 32'hFFFFFFE7 , 32'hFFFFFFF6 , 32'h00000004 , 32'hFFFFFFEB , 32'h00000000 , 32'hFFFFFFF3 , 32'h00000010 , 32'h00000009 , 32'hFFFFFFF9 , 32'h00000007 , 32'h00000000 , 32'hFFFFFFFF , 32'hFFFFFFFD , 32'h00000000} , 
{32'hFFFFFFF9 , 32'h00000009 , 32'hFFFFFFF0 , 32'hFFFFFFFD , 32'h00000007 , 32'hFFFFFFF8 , 32'h00000002 , 32'hFFFFFFFA , 32'hFFFFFFE5 , 32'hFFFFFFE9 , 32'h0000000C , 32'h00000020 , 32'hFFFFFFFD , 32'h0000000E , 32'h00000017 , 32'hFFFFFFFA , 32'hFFFFFFDB , 32'h0000007F , 32'h80000000 , 32'h00000136 , 32'hFFFFFF81 , 32'hFFFFFFE0 , 32'hFFFFFFD3 , 32'hFFFFFFEF , 32'h0000001B , 32'hFFFFFFF8 , 32'h00000007 , 32'h00000001 , 32'h00000009 , 32'h00000003 , 32'h00000002 , 32'hFFFFFFEE , 32'hFFFFFFF6 , 32'h0000001B , 32'hFFFFFFFD , 32'hFFFFFFFD , 32'h00000004} , 
{32'hFFFFFFF4 , 32'hFFFFFFF5 , 32'h00000001 , 32'h00000000 , 32'hFFFFFFFD , 32'h00000000 , 32'hFFFFFFFB , 32'hFFFFFFE6 , 32'h0000000F , 32'h00000020 , 32'hFFFFFFF7 , 32'h0000003C , 32'h00000032 , 32'hFFFFFFBC , 32'hFFFFFFF8 , 32'h00000047 , 32'hFFFFFFDD , 32'h0000000F , 32'h00000136 , 32'h80000000 , 32'h00000121 , 32'hFFFFFFE2 , 32'hFFFFFFC4 , 32'h00000009 , 32'h0000000D , 32'h00000017 , 32'hFFFFFFFD , 32'h00000008 , 32'hFFFFFFDD , 32'h00000007 , 32'h00000007 , 32'h00000001 , 32'hFFFFFFF1 , 32'h00000013 , 32'h00000000 , 32'hFFFFFFF9 , 32'hFFFFFFF7} , 
{32'h00000000 , 32'h00000003 , 32'h00000005 , 32'hFFFFFFEB , 32'h00000002 , 32'hFFFFFFFE , 32'h00000006 , 32'hFFFFFFF1 , 32'h0000000A , 32'hFFFFFFEA , 32'h0000000C , 32'hFFFFFFF5 , 32'hFFFFFFEC , 32'h00000023 , 32'h0000000C , 32'hFFFFFFE4 , 32'h0000003B , 32'hFFFFFFED , 32'hFFFFFF81 , 32'hFFFFFEDD , 32'h80000000 , 32'hFFFFFF78 , 32'h00000011 , 32'h00000027 , 32'hFFFFFFF1 , 32'h00000018 , 32'h00000008 , 32'h00000004 , 32'h00000007 , 32'h00000014 , 32'h00000012 , 32'hFFFFFFF2 , 32'h00000001 , 32'h00000000 , 32'h00000016 , 32'hFFFFFFFD , 32'h00000008} , 
{32'h00000003 , 32'h00000001 , 32'h00000003 , 32'h00000003 , 32'h00000004 , 32'h00000003 , 32'h00000006 , 32'h00000010 , 32'h00000001 , 32'hFFFFFFF8 , 32'hFFFFFFE9 , 32'hFFFFFFEE , 32'hFFFFFFF4 , 32'hFFFFFFE1 , 32'h00000018 , 32'hFFFFFFED , 32'h00000036 , 32'h0000002F , 32'h0000001E , 32'hFFFFFFE2 , 32'hFFFFFF78 , 32'h80000000 , 32'hFFFFFF1B , 32'h00000044 , 32'h0000000F , 32'hFFFFFFBB , 32'hFFFFFFE6 , 32'h00000006 , 32'h00000017 , 32'hFFFFFFFF , 32'h00000003 , 32'hFFFFFFF1 , 32'h00000006 , 32'hFFFFFFF9 , 32'hFFFFFFEB , 32'hFFFFFFF8 , 32'hFFFFFFF4} , 
{32'h00000000 , 32'hFFFFFFFA , 32'h00000000 , 32'h00000005 , 32'h00000003 , 32'h00000000 , 32'h00000001 , 32'h00000007 , 32'h00000003 , 32'h00000005 , 32'hFFFFFFFC , 32'h00000016 , 32'hFFFFFFFE , 32'hFFFFFFFE , 32'h0000000B , 32'hFFFFFFF4 , 32'h0000001D , 32'hFFFFFFF6 , 32'h0000002B , 32'hFFFFFFC4 , 32'h00000011 , 32'h000000E3 , 32'h80000000 , 32'hFFFFFE59 , 32'hFFFFFF83 , 32'hFFFFFFCA , 32'hFFFFFFBE , 32'hFFFFFFB3 , 32'hFFFFFFC9 , 32'h00000011 , 32'h0000000C , 32'h00000003 , 32'h00000014 , 32'hFFFFFFE1 , 32'h00000027 , 32'hFFFFFFD1 , 32'h00000010} , 
{32'h00000000 , 32'h00000000 , 32'hFFFFFFFF , 32'h00000009 , 32'hFFFFFFFD , 32'h00000002 , 32'h00000006 , 32'hFFFFFFEF , 32'h00000015 , 32'h00000028 , 32'hFFFFFFF5 , 32'h0000000D , 32'hFFFFFFFB , 32'hFFFFFFF8 , 32'hFFFFFFEF , 32'hFFFFFFF3 , 32'h00000007 , 32'h00000017 , 32'hFFFFFFEF , 32'hFFFFFFF5 , 32'hFFFFFFD7 , 32'h00000044 , 32'hFFFFFE59 , 32'h80000000 , 32'h00000017 , 32'hFFFFFFAC , 32'h00000039 , 32'hFFFFFFDD , 32'hFFFFFFCB , 32'h00000000 , 32'h0000001E , 32'hFFFFFFFB , 32'hFFFFFFEE , 32'hFFFFFFBE , 32'hFFFFFFF6 , 32'h0000000D , 32'h00000007} , 
{32'h00000001 , 32'hFFFFFFFF , 32'h00000005 , 32'hFFFFFFF6 , 32'h00000007 , 32'h00000000 , 32'hFFFFFFF7 , 32'hFFFFFFFC , 32'hFFFFFFF3 , 32'h00000000 , 32'hFFFFFFF6 , 32'hFFFFFFFE , 32'hFFFFFFFE , 32'h00000000 , 32'h0000001D , 32'h00000014 , 32'h0000001A , 32'hFFFFFFF6 , 32'hFFFFFFE3 , 32'h0000000D , 32'hFFFFFFF1 , 32'hFFFFFFEF , 32'h0000007B , 32'h00000017 , 32'h80000000 , 32'hFFFFFF73 , 32'h0000009A , 32'hFFFFFF2A , 32'h00000059 , 32'h00000014 , 32'hFFFFFFED , 32'h0000002D , 32'hFFFFFFFF , 32'hFFFFFFF5 , 32'hFFFFFFD2 , 32'hFFFFFFDA , 32'hFFFFFFFF} , 
{32'hFFFFFFF4 , 32'hFFFFFFF6 , 32'hFFFFFFF4 , 32'h00000004 , 32'h00000001 , 32'h00000004 , 32'h00000003 , 32'hFFFFFFE8 , 32'h00000000 , 32'hFFFFFFF6 , 32'h00000000 , 32'hFFFFFFFD , 32'hFFFFFFE7 , 32'hFFFFFFF0 , 32'hFFFFFFF8 , 32'h00000013 , 32'h00000011 , 32'h00000004 , 32'h00000006 , 32'h00000017 , 32'h00000018 , 32'h00000043 , 32'h00000034 , 32'hFFFFFFAC , 32'h0000008B , 32'h80000000 , 32'hFFFFFF32 , 32'h00000182 , 32'hFFFFFFE1 , 32'hFFFFFFD6 , 32'hFFFFFFB9 , 32'hFFFFFFD8 , 32'h00000013 , 32'h00000024 , 32'hFFFFFFF1 , 32'h00000017 , 32'hFFFFFFFC} , 
{32'hFFFFFFFB , 32'hFFFFFFFC , 32'hFFFFFFF3 , 32'h0000000A , 32'hFFFFFFFF , 32'h00000000 , 32'h00000007 , 32'h00000017 , 32'hFFFFFFE8 , 32'hFFFFFFF5 , 32'hFFFFFFEC , 32'hFFFFFFFA , 32'h00000018 , 32'hFFFFFFF7 , 32'h00000005 , 32'h00000011 , 32'hFFFFFFE3 , 32'hFFFFFFEB , 32'hFFFFFFF7 , 32'hFFFFFFFD , 32'h00000008 , 32'h00000018 , 32'h00000040 , 32'h00000039 , 32'hFFFFFF64 , 32'h000000CC , 32'h80000000 , 32'h00000194 , 32'h00000014 , 32'h00000029 , 32'hFFFFFFAE , 32'h00000064 , 32'h00000021 , 32'h00000021 , 32'hFFFFFFF4 , 32'h00000007 , 32'hFFFFFFE8} , 
{32'h0000000B , 32'h00000000 , 32'hFFFFFFFE , 32'h00000004 , 32'h00000003 , 32'hFFFFFFFA , 32'hFFFFFFFA , 32'hFFFFFFFC , 32'hFFFFFFEF , 32'h00000004 , 32'hFFFFFFFD , 32'hFFFFFFF1 , 32'hFFFFFFF4 , 32'h00000013 , 32'hFFFFFFDC , 32'h00000001 , 32'h00000006 , 32'h00000000 , 32'hFFFFFFFD , 32'h00000008 , 32'h00000004 , 32'hFFFFFFF8 , 32'h0000004B , 32'hFFFFFFDD , 32'h000000D4 , 32'hFFFFFE7C , 32'hFFFFFE6A , 32'h80000000 , 32'h000000FB , 32'hFFFFFFA4 , 32'hFFFFFFAA , 32'hFFFFFFFC , 32'hFFFFFFDC , 32'h00000012 , 32'h0000000B , 32'hFFFFFFEF , 32'hFFFFFFD8} , 
{32'h00000001 , 32'hFFFFFFFF , 32'hFFFFFFFC , 32'hFFFFFFF6 , 32'hFFFFFFF9 , 32'h00000001 , 32'h0000000F , 32'h00000008 , 32'h0000000C , 32'h00000001 , 32'h00000002 , 32'hFFFFFFE7 , 32'hFFFFFFFA , 32'h00000014 , 32'h00000019 , 32'hFFFFFFFF , 32'h0000000A , 32'h0000000B , 32'h00000009 , 32'h00000021 , 32'hFFFFFFF7 , 32'h00000017 , 32'hFFFFFFC9 , 32'h00000033 , 32'h00000059 , 32'hFFFFFFE1 , 32'h00000014 , 32'h000000FB , 32'h80000000 , 32'h000000B8 , 32'h00000041 , 32'hFFFFFF95 , 32'hFFFFFFED , 32'h0000000F , 32'h0000002E , 32'hFFFFFFEE , 32'h00000000} , 
{32'h00000005 , 32'hFFFFFFFF , 32'hFFFFFFF7 , 32'hFFFFFFFB , 32'hFFFFFFFA , 32'h00000003 , 32'hFFFFFFFA , 32'hFFFFFFFE , 32'h00000007 , 32'hFFFFFFF4 , 32'h00000006 , 32'h00000004 , 32'hFFFFFFFA , 32'hFFFFFFF4 , 32'hFFFFFFF2 , 32'h00000001 , 32'hFFFFFFFE , 32'h00000010 , 32'hFFFFFFFB , 32'h00000007 , 32'h00000014 , 32'h00000000 , 32'hFFFFFFED , 32'h00000000 , 32'hFFFFFFEA , 32'h00000028 , 32'hFFFFFFD5 , 32'h0000005A , 32'h000000B8 , 32'h80000000 , 32'h0000024A , 32'h00000000 , 32'hFFFFFF90 , 32'h0000007B , 32'hFFFFFFC0 , 32'hFFFFFFBD , 32'h00000021} , 
{32'hFFFFFFF9 , 32'h00000000 , 32'hFFFFFFFF , 32'h0000000B , 32'hFFFFFFFE , 32'h00000004 , 32'h00000007 , 32'h00000004 , 32'h00000000 , 32'h00000002 , 32'h00000000 , 32'h00000005 , 32'h00000007 , 32'h00000011 , 32'h00000004 , 32'h00000007 , 32'hFFFFFFF5 , 32'h00000009 , 32'hFFFFFFFC , 32'h00000007 , 32'h00000012 , 32'hFFFFFFFB , 32'hFFFFFFF2 , 32'h0000001E , 32'h00000011 , 32'h00000045 , 32'h00000050 , 32'h00000054 , 32'h00000041 , 32'hFFFFFDB4 , 32'h80000000 , 32'hFFFFFECB , 32'h000000A3 , 32'hFFFFFFCE , 32'h00000064 , 32'hFFFFFFB5 , 32'hFFFFFFF8} , 
{32'hFFFFFFFE , 32'h00000005 , 32'h00000004 , 32'hFFFFFFFE , 32'h00000000 , 32'h00000000 , 32'hFFFFFFFF , 32'h00000003 , 32'hFFFFFFF4 , 32'h00000008 , 32'hFFFFFFFF , 32'h00000004 , 32'h0000000C , 32'hFFFFFFE6 , 32'h00000003 , 32'h00000000 , 32'h00000011 , 32'hFFFFFFF9 , 32'h00000010 , 32'h00000001 , 32'hFFFFFFF2 , 32'h0000000D , 32'hFFFFFFFB , 32'hFFFFFFFB , 32'hFFFFFFD1 , 32'h00000026 , 32'hFFFFFF9A , 32'h00000002 , 32'hFFFFFF95 , 32'hFFFFFFFE , 32'h00000133 , 32'h80000000 , 32'hFFFFFFFA , 32'hFFFFFFB0 , 32'hFFFFFFAD , 32'hFFFFFFA3 , 32'hFFFFFFDB} , 
{32'hFFFFFFF9 , 32'hFFFFFFF9 , 32'h00000008 , 32'h00000000 , 32'h00000003 , 32'hFFFFFFFE , 32'h00000000 , 32'hFFFFFFFA , 32'hFFFFFFFF , 32'hFFFFFFF3 , 32'h00000000 , 32'hFFFFFFEB , 32'hFFFFFFE7 , 32'hFFFFFFF6 , 32'h00000005 , 32'hFFFFFFF7 , 32'hFFFFFFFD , 32'h00000007 , 32'h00000008 , 32'hFFFFFFF1 , 32'h00000001 , 32'hFFFFFFF8 , 32'hFFFFFFEA , 32'hFFFFFFEE , 32'h00000000 , 32'hFFFFFFEB , 32'hFFFFFFDD , 32'h00000022 , 32'hFFFFFFED , 32'h0000006E , 32'hFFFFFF5B , 32'h00000004 , 32'h80000000 , 32'h0000003E , 32'h00000022 , 32'hFFFFFFFD , 32'hFFFFFFD2} , 
{32'hFFFFFFFF , 32'hFFFFFFF3 , 32'hFFFFFFFD , 32'hFFFFFFFC , 32'hFFFFFFFF , 32'hFFFFFFF6 , 32'hFFFFFFFC , 32'hFFFFFFFD , 32'h00000002 , 32'hFFFFFFFC , 32'h0000000F , 32'hFFFFFFFA , 32'hFFFFFFF8 , 32'hFFFFFFFD , 32'hFFFFFFFF , 32'h0000000D , 32'hFFFFFFFB , 32'h00000000 , 32'hFFFFFFE3 , 32'h00000013 , 32'h00000000 , 32'h00000005 , 32'h0000001D , 32'hFFFFFFBE , 32'h00000009 , 32'hFFFFFFDA , 32'hFFFFFFDD , 32'hFFFFFFEC , 32'h0000000F , 32'hFFFFFF83 , 32'h00000030 , 32'h0000004E , 32'hFFFFFFC0 , 32'h80000000 , 32'h00000089 , 32'h00000063 , 32'h00000040} , 
{32'h00000002 , 32'hFFFFFFF8 , 32'hFFFFFFFE , 32'hFFFFFFFB , 32'hFFFFFFFE , 32'hFFFFFFFB , 32'h0000000B , 32'h00000009 , 32'hFFFFFFFE , 32'hFFFFFFF3 , 32'h00000005 , 32'hFFFFFFFE , 32'hFFFFFFFD , 32'hFFFFFFF4 , 32'h00000001 , 32'hFFFFFFF5 , 32'hFFFFFFF6 , 32'hFFFFFFFF , 32'h00000001 , 32'h00000000 , 32'h00000016 , 32'h00000013 , 32'hFFFFFFD7 , 32'hFFFFFFF6 , 32'h0000002C , 32'h0000000D , 32'h0000000A , 32'hFFFFFFF3 , 32'h0000002E , 32'h0000003E , 32'hFFFFFF9A , 32'h00000051 , 32'hFFFFFFDC , 32'hFFFFFF75 , 32'h80000000 , 32'h000003E8 , 32'h00000091} , 
{32'h00000002 , 32'hFFFFFFF7 , 32'h00000002 , 32'hFFFFFFFF , 32'h00000000 , 32'h00000000 , 32'h00000001 , 32'h0000000A , 32'hFFFFFFFC , 32'hFFFFFFFE , 32'hFFFFFFFD , 32'hFFFFFFF8 , 32'h0000000D , 32'h0000000E , 32'hFFFFFFFB , 32'h00000003 , 32'hFFFFFFE9 , 32'h00000001 , 32'hFFFFFFFD , 32'h00000005 , 32'h00000001 , 32'hFFFFFFF8 , 32'hFFFFFFD1 , 32'hFFFFFFF1 , 32'hFFFFFFDA , 32'h00000017 , 32'h00000007 , 32'hFFFFFFEF , 32'h00000010 , 32'hFFFFFFBD , 32'hFFFFFFB5 , 32'hFFFFFFA3 , 32'hFFFFFFFD , 32'h00000063 , 32'h000003E8 , 32'h80000000 , 32'h00000029} , 
{32'hFFFFFFFE , 32'hFFFFFFFD , 32'hFFFFFFFD , 32'hFFFFFFFC , 32'h00000007 , 32'hFFFFFFFD , 32'h00000004 , 32'hFFFFFFFA , 32'h00000003 , 32'h00000007 , 32'hFFFFFFFA , 32'hFFFFFFFF , 32'h00000002 , 32'h00000008 , 32'h0000000D , 32'h00000000 , 32'hFFFFFFE6 , 32'h00000000 , 32'hFFFFFFFA , 32'hFFFFFFF7 , 32'h00000008 , 32'h0000000A , 32'hFFFFFFEE , 32'h00000007 , 32'h00000000 , 32'h00000002 , 32'h00000016 , 32'h00000026 , 32'h00000000 , 32'hFFFFFFDD , 32'h00000006 , 32'h00000023 , 32'h0000002C , 32'hFFFFFFBE , 32'hFFFFFF6D , 32'h00000029 , 32'h80000000}
};

logic signed [31:0] VT_1 [37][300] ='{
{32'hFEAEC19C , 32'hD76B1280 , 32'h000009A0 , 32'hF6554840 , 32'hFFFF3F47 , 32'h03C32B60 , 32'hFFFFA3B4 , 32'h0000B288 , 32'hFFFCD535 , 32'hFFFFAC8D , 32'h04BBAA38 , 32'hF5B788B0 , 32'h087D25B0 , 32'hFFFF9BD8 , 32'hFFFD598B , 32'hF64836D0 , 32'hFFFF610B , 32'h00871991 , 32'hFB8CAF70 , 32'h0000897D , 32'hFFFFD067 , 32'h0021E330 , 32'hFBCA91D0 , 32'hFDE049EC , 32'h02B1CC50 , 32'h00003505 , 32'hFE4FE838 , 32'hFF8FE6CC , 32'hFFFEDF21 , 32'h04B0EA90 , 32'hFFFF7DE6 , 32'h00326A03 , 32'h00001384 , 32'hFFFD6401 , 32'hFFFF9EFC , 32'hF3FCFC40 , 32'h031E2408 , 32'h021E3C68 , 32'h00015025 , 32'h0363A9C4 , 32'h0C83F700 , 32'h00008456 , 32'h00026C76 , 32'hFCF8983C , 32'h01504114 , 32'h0E571A00 , 32'hF9622F80 , 32'hFFFF5282 , 32'h04E73710 , 32'hE48C0AC0 , 32'hFF62EEF2 , 32'h00002C75 , 32'h03271960 , 32'h0DB2A850 , 32'h03CDC028 , 32'hFFFFF24B , 32'h035DB090 , 32'hFFFFE75A , 32'h00010CE4 , 32'h00C51917 , 32'hFFD69027 , 32'h06381818 , 32'hE5C818A0 , 32'h0000DC0D , 32'hF4006BC0 , 32'hFFFF764E , 32'hF86FAAF0 , 32'h007F450A , 32'hFFFFDB99 , 32'h000919D1 , 32'h02A3F9C0 , 32'hFAEEF960 , 32'hFFFFE95F , 32'h00027CCC , 32'h00000887 , 32'hF15BFBD0 , 32'hFB596798 , 32'h00006FB4 , 32'hECA3AC60 , 32'h012AC574 , 32'hFFFF207D , 32'hECBE9900 , 32'hF89B9FD0 , 32'h000001D5 , 32'h01AB884C , 32'h10CA0820 , 32'hFA6A6368 , 32'h0000AD3D , 32'hFFFF2900 , 32'h17A9D520 , 32'h0001AFAB , 32'hFB4821B0 , 32'h00004A87 , 32'hFBE2FB20 , 32'hFF4715DF , 32'h0002224A , 32'hFFFE8691 , 32'hFFFFBB45 , 32'h00020326 , 32'hF792D950 , 32'hFE6A8C48 , 32'h00015CC7 , 32'h00C57DD1 , 32'h026C0088 , 32'h0298F664 , 32'h00014EDA , 32'h00481954 , 32'h0000663D , 32'h06FA77B0 , 32'h25D53780 , 32'hFFFF9CC1 , 32'h0220C2A8 , 32'hFFFEFD2F , 32'h0000832A , 32'hF8E09530 , 32'h02A28718 , 32'hFFB58520 , 32'h00002C7A , 32'hFA998AC0 , 32'h0001AA8F , 32'hFFFE4E75 , 32'hF8CD5DD0 , 32'h00027638 , 32'h00004858 , 32'hFFB76585 , 32'hF781C530 , 32'h000033C4 , 32'hFFFF1522 , 32'h00015ACE , 32'hFFFE3E23 , 32'hFFFF8800 , 32'h01133E5C , 32'hFA65FBD8 , 32'h00014771 , 32'hFFFF4D9B , 32'h2D6BB8C0 , 32'h0D643620 , 32'h00018124 , 32'hFFFF2438 , 32'hFFA956D5 , 32'h00000FB6 , 32'hFFFFE0EE , 32'hFEB54EC4 , 32'h0401FAF0 , 32'h0097FD97 , 32'hFD0A3D44 , 32'hFFFF023E , 32'hFFFF190A , 32'h042F1E58 , 32'hFFFFB8FE , 32'hFFFE2CD5 , 32'hFF4548CC , 32'hFFFF5F70 , 32'h00003F95 , 32'h043C1798 , 32'hFFFC28CF , 32'hF425BA10 , 32'hFE4C6568 , 32'h00016715 , 32'h000187D8 , 32'hFFFE28B9 , 32'hF4A22420 , 32'hFF01104F , 32'h09AC04F0 , 32'h04190580 , 32'hFFFF1F1D , 32'hF28EC3B0 , 32'h00005C51 , 32'h0000C8C3 , 32'hEE81B0A0 , 32'h00294F2D , 32'h01B61B20 , 32'hFFFE9E52 , 32'hEFD9B0C0 , 32'hFE6E2F6C , 32'hFE1165B8 , 32'hEC57EBC0 , 32'hFCDC443C , 32'hFE8D0B98 , 32'hFF486ACF , 32'h03507C90 , 32'h000031B0 , 32'hFFFEBA7C , 32'hFFFF1FD8 , 32'hFBA6B1E0 , 32'h04BCD568 , 32'h00FF30C4 , 32'h0128626C , 32'hFA1D19C8 , 32'h02B50C04 , 32'h0001F1EE , 32'hF723DDF0 , 32'hF7357F90 , 32'hFFFDB23A , 32'h002C8633 , 32'hFFFEE865 , 32'h078D0AC0 , 32'h01A1C870 , 32'hFFFE6C3A , 32'h00026ADB , 32'hFFFF14F0 , 32'h0004211D , 32'h00024BA0 , 32'hFFFFC341 , 32'h03AD4F68 , 32'h0144E5D4 , 32'hF8BD4818 , 32'h02760B80 , 32'h0C6559B0 , 32'h0FC8E290 , 32'h00007DC5 , 32'hFFFFF60E , 32'h00025D6F , 32'h000010E4 , 32'hFFFF326C , 32'h00B941B7 , 32'h0094E51A , 32'h0A9F8280 , 32'h0001B23E , 32'hFFFF4BF4 , 32'h0001A502 , 32'hFFFBE58C , 32'hFCC49D78 , 32'h0CCFE5C0 , 32'hFFFF1465 , 32'hFFFE5DAE , 32'hFFFDBAB9 , 32'hEEBB8440 , 32'h026F9698 , 32'h0884B0D0 , 32'hFFFE5BE8 , 32'hFFFE3B5E , 32'h0002692E , 32'hFE799324 , 32'h0233FF40 , 32'h0D42AE40 , 32'hFFFF29AF , 32'hFF497359 , 32'h0001F204 , 32'h0261ABCC , 32'h00013E07 , 32'hFBA70C98 , 32'h0000D4FF , 32'hF31E5AA0 , 32'hFCC22728 , 32'h0AAD4B80 , 32'hFDF5BD78 , 32'hFFFF2C03 , 32'h04A463B8 , 32'hFE6A5830 , 32'h00026C89 , 32'hF88F6498 , 32'h00012C57 , 32'h0045D8DC , 32'hF9D02100 , 32'hFE3332CC , 32'hFFFEDB79 , 32'hFFFE845E , 32'hFF253FCE , 32'h00002E7E , 32'hFE7015B0 , 32'hFFFFDFCD , 32'h006BC89A , 32'hFFFF8D5C , 32'hFA35C888 , 32'hFFFFAC1D , 32'hFFFE178F , 32'h00007528 , 32'hFF70592E , 32'hF9414C98 , 32'hFFFED890 , 32'hFFFD22EE , 32'hFFFF6CAE , 32'h00002311 , 32'hFB1C7EE0 , 32'hFBFBB720 , 32'hFFE7619B , 32'h1CE61260 , 32'h04E3E460 , 32'h00018E78 , 32'h0000ACA2 , 32'h000065E2 , 32'h0423BEE0 , 32'hFFFF3881 , 32'h0002F251 , 32'h033F83E4 , 32'h02D90D68 , 32'h0000BFBF , 32'h1076B4A0 , 32'hFFB02CF4 , 32'h045786C8 , 32'h001ABB95 , 32'h0000A353 , 32'h017E1F78 , 32'hF435FD40 , 32'hFC6BA2E0 , 32'h000075EF , 32'hED0ADC00 , 32'hF8DFF400 , 32'hF3DCB0E0} , 
{32'h058CC0D0 , 32'hEA374CC0 , 32'hFFFFF3BA , 32'h025FF79C , 32'h0001D1B4 , 32'h01C75EE0 , 32'h00034BB7 , 32'h000188AD , 32'hFFFDB7C3 , 32'hFFFF49A0 , 32'h01635990 , 32'hF4635FB0 , 32'hFF85B299 , 32'h0001AC7D , 32'hFFFFECB3 , 32'hEF44C5A0 , 32'hFFFD96B7 , 32'h06CC8C68 , 32'h05EF8C48 , 32'h00025285 , 32'h0000831C , 32'h01941DEC , 32'hFDC8CF58 , 32'hF231D010 , 32'hF2D239C0 , 32'hFFFD0D13 , 32'hFF700878 , 32'hFFC25C61 , 32'h0001D18B , 32'hF4E66630 , 32'hFFFE6A32 , 32'h094799D0 , 32'hFFFF158B , 32'hFFFE3165 , 32'h000194A6 , 32'hF5F6EC50 , 32'hFFCB5290 , 32'h0D2B9C70 , 32'hFFFE50BE , 32'hFE57C1B0 , 32'h007B7911 , 32'hFFFF8EF6 , 32'hFFFFE275 , 32'h047F0E38 , 32'h03668F78 , 32'hFBDDFA88 , 32'hFCE8DDE0 , 32'h00007514 , 32'h0C1A91F0 , 32'hEEC50B60 , 32'hFE855734 , 32'h0002E993 , 32'hFC0C1778 , 32'h0422FF98 , 32'hFF4AD5DC , 32'hFFFF58F2 , 32'hFC415118 , 32'h00025A01 , 32'h00017CD1 , 32'h01A15768 , 32'hFF138D75 , 32'hFFA20282 , 32'h20D1E240 , 32'h0001CFCF , 32'hFAD596C0 , 32'hFFFF55B9 , 32'hFE02C338 , 32'h00B4C29B , 32'hFFFFFE15 , 32'hFA09D168 , 32'hFD5EC74C , 32'h05996C48 , 32'h0002BDF4 , 32'hFFFEE16E , 32'hFFFE0464 , 32'hF7C1CFB0 , 32'h02BC93A8 , 32'hFFFE7685 , 32'hFF5AA767 , 32'h01755AD4 , 32'h00006D80 , 32'hFCC22970 , 32'hFA281CC0 , 32'hFFFE9EB9 , 32'h04CCA008 , 32'hFAF727E8 , 32'h06454118 , 32'hFFFEC449 , 32'hFFFF81FD , 32'hFC6151B8 , 32'h00022C4D , 32'hF80478C0 , 32'hFFFF40C7 , 32'h0A22A480 , 32'hFFF0138D , 32'h00004914 , 32'h00003170 , 32'hFFFDE261 , 32'h0000BCB2 , 32'hF863AC40 , 32'hFF214180 , 32'h00005134 , 32'h02812A7C , 32'h05FF68B0 , 32'hFE4AA144 , 32'hFFFD5C79 , 32'h0062FAC7 , 32'hFFFDB5AB , 32'hFC146BD0 , 32'hD7FE45C0 , 32'hFFFF0B52 , 32'hF5A70670 , 32'h000172D5 , 32'hFFFF127C , 32'h04423370 , 32'hFFF2A666 , 32'hFECF8630 , 32'hFFFC0A8C , 32'h01B581B4 , 32'hFFFF6EB5 , 32'hFFFFAF43 , 32'hFE7D5248 , 32'h0001A69B , 32'hFFFFBC38 , 32'h03AF29A8 , 32'hF9BC2688 , 32'hFFFEE716 , 32'hFFFF2A7F , 32'hFFFF37C7 , 32'hFFFF9803 , 32'h00013D5A , 32'hF48F8840 , 32'h055E1038 , 32'h00001DED , 32'h0000EABE , 32'h05AD7F08 , 32'hFFC667CA , 32'h000072EC , 32'h0001FD5D , 32'h079AE648 , 32'hFFFF227A , 32'hFFFD2870 , 32'h0464D9C8 , 32'hFD7A5470 , 32'h01DB07E8 , 32'hFFA7C628 , 32'hFFFF8E50 , 32'hFFFE2E48 , 32'h00998547 , 32'hFFFFD078 , 32'hFFFFF867 , 32'hFCE92150 , 32'hFFFF6871 , 32'h0000F2FD , 32'hFB3A2768 , 32'h0000113F , 32'h03170D74 , 32'hFFB7A265 , 32'h00002AB6 , 32'hFFFEA889 , 32'h00030D10 , 32'hEBD56500 , 32'hFCE9E8B4 , 32'hF53BD950 , 32'hFAA23198 , 32'h0000C142 , 32'h0AF6E680 , 32'h0001E9B7 , 32'h0001B3E0 , 32'h03965FC8 , 32'hFEDC95E8 , 32'h01CB5784 , 32'h000172C7 , 32'hEE5B73A0 , 32'h01119940 , 32'hFFFE8474 , 32'hFF641FF5 , 32'hFEA83304 , 32'h21456240 , 32'hFF30184E , 32'hFDBE10A8 , 32'h00010F11 , 32'hFFFFCBFB , 32'hFFFF79F3 , 32'hFA6B2C28 , 32'hEA292EA0 , 32'h03D31F70 , 32'hFF63BCA4 , 32'hFCE20E50 , 32'hFACA9370 , 32'h0000B7A0 , 32'hF72731E0 , 32'hFB565568 , 32'hFFFE1CCD , 32'hFF086460 , 32'h000168A8 , 32'hFCD9BD1C , 32'hEA70EAA0 , 32'h0003AA09 , 32'h0000D154 , 32'hFFFF03B9 , 32'hFFFEEF8E , 32'h0000E898 , 32'hFFFEFB26 , 32'h00FF5F07 , 32'h06FEF8D0 , 32'h018BA6A0 , 32'h0A812CD0 , 32'h05BEB068 , 32'hED58F400 , 32'h00012E9D , 32'hFFFDC028 , 32'hFFFEE5EF , 32'h0000EA1C , 32'h00010064 , 32'h01B72264 , 32'h06059CC8 , 32'h0528F258 , 32'h00008FD5 , 32'hFFFEB65F , 32'h00003177 , 32'h0002291E , 32'h0A9ACDC0 , 32'hF295AFB0 , 32'h000095FA , 32'h00020CD0 , 32'h0000270A , 32'hF34B2040 , 32'h09714A40 , 32'hF5F190F0 , 32'hFFFEB4C6 , 32'hFFFF0C7C , 32'hFFFFBB44 , 32'h02697874 , 32'h00B296EC , 32'hF047E330 , 32'h00011780 , 32'h0110CA30 , 32'h00018601 , 32'h07F9D1C8 , 32'h000206A9 , 32'hE8AA4CA0 , 32'h0002B55E , 32'hEB3FAA40 , 32'h0463F530 , 32'h30008080 , 32'h0DD8DF60 , 32'h0001D5E9 , 32'hFE650E10 , 32'hFE2E6C08 , 32'hFFFEAED8 , 32'h094405B0 , 32'h0001FDF5 , 32'hFEFFCBA0 , 32'hFBBD0AF8 , 32'h003801F5 , 32'h00019D1B , 32'h00013075 , 32'h0EF3ED00 , 32'h00015458 , 32'hF82BDF58 , 32'h0000CDDB , 32'h006E39B4 , 32'hFFFFF5F5 , 32'hFEC57878 , 32'hFFFFA40F , 32'h0000BD12 , 32'h00006E9F , 32'hFFFE5FC2 , 32'h0402E938 , 32'hFFFE7B4A , 32'h00005E79 , 32'hFFFF5E7F , 32'h00005CF2 , 32'hF94601A8 , 32'h0AEC2C10 , 32'hEDFB7080 , 32'h09BBCA20 , 32'hF8887D40 , 32'h0000B616 , 32'hFFFFFB30 , 32'hFFFFA957 , 32'h0198C44C , 32'hFFFEAA48 , 32'hFFFED6B6 , 32'hFD191BC4 , 32'h094C3260 , 32'hFFFED277 , 32'hF2503EE0 , 32'h02E6A6A8 , 32'hFF63CF5D , 32'hF2953240 , 32'hFFFF20A7 , 32'h02776F30 , 32'h0251D070 , 32'hFE79773C , 32'hFFFEDDCF , 32'hFC45C578 , 32'h0A587F20 , 32'h0D3B56E0} , 
{32'h066DFC10 , 32'hE5B3EF40 , 32'h000240E5 , 32'hF9164E60 , 32'h0001176C , 32'hFF8E5E1D , 32'h0000B32B , 32'hFFFFB67C , 32'h00027BEE , 32'h000110A0 , 32'hFF8188F3 , 32'hFC069200 , 32'hFD5430A8 , 32'h00005CE3 , 32'h0001C56B , 32'h0B5401D0 , 32'hFFFE821E , 32'hEA5D7DE0 , 32'h0045563F , 32'hFFFF1DD8 , 32'hFFFFE08C , 32'h02C67D9C , 32'h03E39098 , 32'h01B0E534 , 32'hEF9E17E0 , 32'h0000A958 , 32'h046BBEC8 , 32'hFEAC183C , 32'hFFFE6214 , 32'hFE739440 , 32'hFFFFF4CB , 32'hFCB124E8 , 32'h00006EAB , 32'hFFFFEC7F , 32'hFFFDD3AE , 32'hF6A138A0 , 32'hF69F0290 , 32'h07B58958 , 32'hFFFE28FB , 32'hF4ABD140 , 32'h0613BA90 , 32'h00001EEE , 32'hFFFE1BC2 , 32'hFAE3BF58 , 32'h131B6400 , 32'hE9FFDFC0 , 32'hFFFEC594 , 32'hFFFF8663 , 32'hFB9DCE08 , 32'h0169C334 , 32'h009A5D7E , 32'h000149A7 , 32'hFE4AC15C , 32'h010B0B74 , 32'hFD25B680 , 32'h0001CC98 , 32'h003F9313 , 32'h00013593 , 32'h00008AF6 , 32'h02B2BC54 , 32'h00FA6B92 , 32'h0183AEF0 , 32'hF849E8D0 , 32'h0000507D , 32'h097C2810 , 32'hFFFFE8BC , 32'hD931E7C0 , 32'hFD9075CC , 32'h0001D1E7 , 32'h01B4C1E0 , 32'h15532E60 , 32'hF5E960F0 , 32'hFFFFF596 , 32'hFFFFE507 , 32'hFFFE294D , 32'hFCC5C9DC , 32'hFA7AFB80 , 32'h00010503 , 32'hFC9C341C , 32'hFE49D998 , 32'hFFFF4174 , 32'hF1655A40 , 32'hFB3C0E10 , 32'h00007F70 , 32'hFF11D733 , 32'hEF4C18E0 , 32'hFB2B79E0 , 32'hFFFF2928 , 32'hFFFF8794 , 32'h0EC1B780 , 32'hFFFFDE8D , 32'hFD06BB70 , 32'h0000CEAD , 32'hFCE01898 , 32'h000B0D45 , 32'hFFFF831D , 32'hFFFE5C90 , 32'hFFFFC504 , 32'hFFFF76B1 , 32'hFCE5DE14 , 32'h05435CE8 , 32'hFFFDB2BE , 32'hFB1B5410 , 32'hFF07926E , 32'hFFA6D39F , 32'h00015778 , 32'hFFB05073 , 32'h0000B919 , 32'h03EE5CEC , 32'h02C94BDC , 32'hFFFE615D , 32'h05D5F610 , 32'h00032225 , 32'hFFFE6A65 , 32'h0187F960 , 32'hFD8457D8 , 32'h00588DED , 32'h0000C833 , 32'hF9F95BF0 , 32'hFFFF19EF , 32'h00000814 , 32'hFE603E40 , 32'hFFFEFF5D , 32'hFFFF8404 , 32'h0A85CD50 , 32'h0286E008 , 32'h0000CD2C , 32'hFFFF3CD9 , 32'h00021FEB , 32'h000094DF , 32'h00004A7E , 32'hFD5DE770 , 32'h07D33170 , 32'h0000F297 , 32'hFFFDFA10 , 32'hDB31BC40 , 32'hFD77CA0C , 32'hFFFF99F0 , 32'hFFFFA8AD , 32'h02ED03F8 , 32'hFFFF2E05 , 32'h0000A942 , 32'h025FEC90 , 32'h02DF2948 , 32'hFE7EF058 , 32'h020D8EE4 , 32'h0003F9DD , 32'hFFFD60E4 , 32'hFD352C3C , 32'h0002F92A , 32'h00013ECF , 32'h00403351 , 32'h000218C9 , 32'h0001B81B , 32'hFC60494C , 32'h0000DA11 , 32'h0871C3C0 , 32'h00180233 , 32'hFFFCFAD3 , 32'h00005FFE , 32'hFFFF5C3F , 32'hFA2A53B8 , 32'hFF595281 , 32'hFE769E48 , 32'hF51F0BA0 , 32'h00002491 , 32'hF4A22230 , 32'h0002E2B2 , 32'hFFFE73F5 , 32'h007C8FD1 , 32'hFC5C8D7C , 32'hF7E37FA0 , 32'hFFFEB1D5 , 32'h14E9AF20 , 32'hFD13E4DC , 32'hFB7195A0 , 32'h19FBCE40 , 32'hFB7964C0 , 32'hFAE5CFA8 , 32'h00311AA2 , 32'hE5084800 , 32'hFFFF5A7D , 32'h00019C8E , 32'h0000F667 , 32'h04AFFFD8 , 32'hE1B7AB40 , 32'hFFBB0390 , 32'hFF4A32A1 , 32'h02211AC8 , 32'hFA72BA48 , 32'hFFFE0A53 , 32'h000D711D , 32'hFBCF21A0 , 32'h00007E96 , 32'hF50D3A60 , 32'hFFFED6C8 , 32'hFD4935CC , 32'h00AA2CB1 , 32'hFFFFB12C , 32'h0000BDBE , 32'h0001FD1B , 32'h000032BE , 32'hFFFF243D , 32'h00004756 , 32'h02C8F600 , 32'hEAF4BD00 , 32'h039C2E98 , 32'h0DC61940 , 32'h07444600 , 32'hFED10F98 , 32'hFFFEB8C1 , 32'hFFFF0592 , 32'h0000B578 , 32'hFFFD8398 , 32'h00023F22 , 32'hFFEDD644 , 32'h05B9E828 , 32'h04CD60D0 , 32'hFFFF3589 , 32'h00021E0E , 32'h000030E2 , 32'h0001E1A6 , 32'h0974D5F0 , 32'h24F93000 , 32'h000339FF , 32'hFFFF5C33 , 32'hFFFF4C2B , 32'h09C3A190 , 32'h19DF1780 , 32'h0B92D040 , 32'h00001AE0 , 32'hFFFF4818 , 32'h0000D20A , 32'hFAB15DB0 , 32'hFFEF0EF4 , 32'h044A8B98 , 32'h0001DDF1 , 32'h004824A1 , 32'h0002CCA8 , 32'hF88996A0 , 32'h00045985 , 32'h04071C10 , 32'h0002DBD5 , 32'hF41AB650 , 32'hFCF438C4 , 32'hFC33F294 , 32'h09D7D990 , 32'h0001EFC4 , 32'hF5224050 , 32'hFF6AB646 , 32'hFFFF540C , 32'hFEB9069C , 32'hFFFFD2D7 , 32'h00F489CF , 32'hF130FB10 , 32'h059CE0D0 , 32'h00019752 , 32'h000061CC , 32'hFCB36648 , 32'h00012DD3 , 32'h04243250 , 32'hFFFF8CFE , 32'hFDFB2FFC , 32'hFFFFFAA5 , 32'hFFC2FAB9 , 32'h0000ED78 , 32'h0004061B , 32'hFFFCF44D , 32'hFD8BE9A0 , 32'hF5AC51C0 , 32'hFFFD5B96 , 32'h000286AF , 32'hFFFF63A7 , 32'h00002D16 , 32'hF5DEDA60 , 32'hFE5E71C4 , 32'h0CB63E60 , 32'h096C31A0 , 32'h0C0264E0 , 32'hFFFE701D , 32'h000062AC , 32'hFFFF82F9 , 32'h00486F49 , 32'h0000D029 , 32'hFFFF65AE , 32'hFFAEE275 , 32'h06007C88 , 32'hFFFF67FA , 32'hF4770920 , 32'hFF9C4D19 , 32'hFBB10500 , 32'h09D9BEF0 , 32'h0000A017 , 32'h066B8C88 , 32'hFA2FB718 , 32'hFF3B3D60 , 32'h00001939 , 32'h0C48A9C0 , 32'h0379064C , 32'hFCDD08A8} , 
{32'h03449324 , 32'hEF212300 , 32'h000054B1 , 32'hFD9E06B4 , 32'hFFFE5585 , 32'h02166348 , 32'h00009ABC , 32'hFFFF6750 , 32'hFFFE2CEC , 32'h00007204 , 32'hF8592268 , 32'hF3B2A1B0 , 32'hFFA12907 , 32'h00010869 , 32'h00005A12 , 32'hFDBD93F4 , 32'h00016A93 , 32'h009DECF9 , 32'hFE516E44 , 32'hFFFF0FB9 , 32'h00030B37 , 32'h02EB4ED8 , 32'hFF7028D7 , 32'hFECD8AF0 , 32'hFF15E63B , 32'h0001363C , 32'h01AE4D74 , 32'hFD9F3858 , 32'hFFFEF5D1 , 32'h11B2B0C0 , 32'h000219E7 , 32'hF9B53800 , 32'hFFFD3BDA , 32'h0000F84F , 32'hFFFFEC76 , 32'h02AC4E4C , 32'h0F1DC970 , 32'h0B2AC6C0 , 32'h000116EF , 32'h0990BD60 , 32'h01964A18 , 32'h000055BC , 32'h0000A398 , 32'hFA5118D8 , 32'h02C96618 , 32'h09DAE710 , 32'h0DC421B0 , 32'h0002FB14 , 32'h025414D0 , 32'h01E12D84 , 32'h01FB56D0 , 32'h00012CC2 , 32'hFF037378 , 32'h09CBFAF0 , 32'h084AD500 , 32'hFFFFD285 , 32'h004EFED8 , 32'h000026C9 , 32'h00029750 , 32'hFA841D58 , 32'h01D5DE58 , 32'hFEAC33F0 , 32'h045D2C38 , 32'h00004FCB , 32'hF3D43C30 , 32'hFFFF12F0 , 32'h1FCBCFC0 , 32'h003A0697 , 32'h00018ECF , 32'hF439F110 , 32'hF9F1FBC0 , 32'h015F0864 , 32'h0001634D , 32'h00003D06 , 32'hFFFF04A9 , 32'h02B7C228 , 32'hFE403944 , 32'h00003E85 , 32'h03540E00 , 32'h003214CF , 32'h000334B9 , 32'h09ACC290 , 32'h00BE3C42 , 32'hFFFF5AB3 , 32'h03CB9354 , 32'h04B252C0 , 32'h04618710 , 32'hFFFFF28F , 32'hFFFF96DB , 32'hF09B6910 , 32'h00005E3C , 32'h0746D3C8 , 32'h00003A7E , 32'h05E4EAA8 , 32'hFF076E3F , 32'h0000EFAE , 32'h00003780 , 32'hFFFFE1B0 , 32'hFFFF5A74 , 32'hFF571DD9 , 32'h0A12D060 , 32'hFFFDA391 , 32'hFEE663E0 , 32'h101418E0 , 32'h053BAE20 , 32'hFFFF82D8 , 32'h0002028B , 32'hFFFFA417 , 32'hFF65F735 , 32'h04DC1C48 , 32'h00014AEE , 32'hFD87FE3C , 32'h00006C67 , 32'h00024F41 , 32'h0A777890 , 32'h08B00060 , 32'h01FD6124 , 32'h000013C6 , 32'hFC78D0A0 , 32'h0000662B , 32'h00006C7E , 32'hFCF8AEF0 , 32'hFFFF7138 , 32'h00003538 , 32'hF5B99D40 , 32'h0261EE10 , 32'h0001CBE7 , 32'hFFFFDA4B , 32'h0000D885 , 32'hFFFEE578 , 32'hFFFFC3D1 , 32'h0004FC1C , 32'h08EDACB0 , 32'h00010F93 , 32'h0000D173 , 32'h112D17E0 , 32'h011A54D8 , 32'hFFFD7FCA , 32'hFFFF319E , 32'h00242B3E , 32'h0000BF54 , 32'hFFFFF3F6 , 32'hFF9E5EFB , 32'h0B0968F0 , 32'h054F0588 , 32'h00C36B66 , 32'hFFFF35F2 , 32'h0001F7BE , 32'h0106FDAC , 32'h000245D6 , 32'hFFFF00BA , 32'hFF93B905 , 32'h0000917A , 32'hFFFEB684 , 32'hFDCCA4D4 , 32'hFFFF929B , 32'h0DC4BD20 , 32'hFFDFEA8E , 32'h0001B3FD , 32'h0000BF8D , 32'hFFFF1A3C , 32'hF68A0670 , 32'h08561BA0 , 32'h007E1175 , 32'h06B69FF0 , 32'h000139BC , 32'hF39D0CA0 , 32'h00006F5E , 32'hFFFF0E89 , 32'hF688AF20 , 32'h087A41B0 , 32'hFF67ED84 , 32'hFFFE1C9D , 32'h0058BE0A , 32'hFBB8A9D0 , 32'hFC1FEDD0 , 32'h386689C0 , 32'hFE774F44 , 32'hFEAA1624 , 32'h0370FDFC , 32'h008D1FB8 , 32'h00006B48 , 32'h00009F49 , 32'hFFFFCF9F , 32'h0B21DC90 , 32'hF25C79D0 , 32'hFFB39A11 , 32'h029F488C , 32'hFCEDD788 , 32'h030419D4 , 32'hFFFCFFD1 , 32'hFA4A2E68 , 32'hF9009E60 , 32'hFFFE34FE , 32'hFDB0020C , 32'hFFFDE412 , 32'h05B70608 , 32'h0AFF1B60 , 32'hFFFFCF6A , 32'h0001C487 , 32'hFFFF946C , 32'h0000D54D , 32'h00002B70 , 32'h0001DC74 , 32'h055D99A0 , 32'hF7C93770 , 32'hFB1C7340 , 32'h08B20DA0 , 32'hFFD98A83 , 32'h0588D970 , 32'h0000A631 , 32'hFFFF5646 , 32'h000158D2 , 32'h00016577 , 32'hFFFF85DE , 32'hFFAE6A0F , 32'h00277E0A , 32'h045BAF20 , 32'h00016A65 , 32'hFFFF047D , 32'hFFFF1229 , 32'h0000626A , 32'h019F0664 , 32'hEDC51D40 , 32'h0001FF90 , 32'hFFFF327A , 32'h00022A36 , 32'hE586C4C0 , 32'h14869CE0 , 32'h010E0A64 , 32'hFFFF2593 , 32'h000264C5 , 32'h00008FF5 , 32'hFDFF76EC , 32'h0321A104 , 32'hE2F7D940 , 32'h00003930 , 32'hFFF682B0 , 32'hFFFD8C84 , 32'hF6B1E5D0 , 32'hFFFDA86F , 32'h1DAC7F80 , 32'h00013505 , 32'h13218D20 , 32'h117CF920 , 32'h01EC6FB4 , 32'h0E21E6C0 , 32'h0001BF7E , 32'hF9E6BD08 , 32'hFF311BD4 , 32'h0000154C , 32'hFFF5A119 , 32'hFFFF5500 , 32'h01CAE07C , 32'h0947A350 , 32'h08428010 , 32'hFFFE99E9 , 32'hFFFD6A9F , 32'hF5E5C140 , 32'h00021A00 , 32'h0D246820 , 32'h00002DE5 , 32'hFF577943 , 32'h00022F76 , 32'h0AE686E0 , 32'h0000DCCB , 32'h00003AE9 , 32'hFFFD952C , 32'h15B007C0 , 32'hF9B73658 , 32'hFFFED397 , 32'hFFFF3F56 , 32'h000020AB , 32'hFFFEFBB0 , 32'h077629B8 , 32'hF8DD2790 , 32'h1C908FA0 , 32'hFED327A8 , 32'h0A124880 , 32'hFFFEA5BF , 32'hFFFFA4F6 , 32'h00034DA9 , 32'h0220E380 , 32'hFFFF4BBB , 32'h0000970A , 32'h05B4C5A0 , 32'hFDA4107C , 32'h0000CC1B , 32'hFD8D5084 , 32'h01D1C1E8 , 32'h032B8634 , 32'h0415DC58 , 32'h00011CA3 , 32'h0296F7C0 , 32'h01098694 , 32'hFFA14BE0 , 32'hFFFECB87 , 32'hFD0BE50C , 32'hF8EB4400 , 32'h0D58B590} , 
{32'h0724D4A8 , 32'h14BC4520 , 32'hFFFDBBAD , 32'hFE6D0178 , 32'hFFFBF4D9 , 32'h0067A7EA , 32'hFFFE96FC , 32'hFFFF0445 , 32'hFFFDC636 , 32'hFFFF9B84 , 32'hFE2B644C , 32'hFDAA3848 , 32'h02756C60 , 32'hFFFD8F10 , 32'hFFFE7897 , 32'h0867F4A0 , 32'h0000282D , 32'hEB4359C0 , 32'hF69D35C0 , 32'hFFFFE45B , 32'h0000416E , 32'h00343765 , 32'h073395D0 , 32'hFC3791CC , 32'h044BBD10 , 32'h000072E6 , 32'hFE8961E8 , 32'hFDE1FC90 , 32'hFFFE2BF0 , 32'h0A34AD00 , 32'h0000487C , 32'hF2E7BA30 , 32'hFFFDD5E1 , 32'h0000E9FB , 32'h00002E96 , 32'h0702DB90 , 32'hF4072800 , 32'hFA7D6AB0 , 32'h00013670 , 32'h0BADCD40 , 32'h05CD03B0 , 32'h00017304 , 32'h00019148 , 32'h02338C64 , 32'h040DFFF8 , 32'h0CE99280 , 32'hF45B5910 , 32'h0000C89B , 32'hFF7F92AC , 32'h1AB82200 , 32'hFFBA8D0C , 32'h00049A62 , 32'hFDCD08C0 , 32'h01386310 , 32'hFA3ADA80 , 32'hFFFF5844 , 32'hFF9B7DA9 , 32'h00010541 , 32'hFFFFAE98 , 32'h00E93B87 , 32'hFE8799CC , 32'h036149AC , 32'hFC5F43C8 , 32'h0000DDBE , 32'hDF7A2180 , 32'h00014F66 , 32'hE84F2D40 , 32'hFEED4064 , 32'h0001014F , 32'hF4622430 , 32'h00C5D921 , 32'h0D5BBA90 , 32'hFFFEF31A , 32'hFFFD4FB9 , 32'hFFFF3981 , 32'h043D4070 , 32'h038783F0 , 32'h00000034 , 32'h104985C0 , 32'hFFE9F921 , 32'h0001079C , 32'h0AD730B0 , 32'hFD1728B8 , 32'h0001F04A , 32'hFF56BFE9 , 32'hFFB8143D , 32'h002208D5 , 32'h00007E97 , 32'hFFFF3261 , 32'hFFDE1457 , 32'h00002DBB , 32'h066C29C0 , 32'hFFFF1631 , 32'hF2278DA0 , 32'hFED60D14 , 32'hFFFDCE75 , 32'hFFFFA9AA , 32'h000118E8 , 32'h00024CC0 , 32'h078A0138 , 32'h042B1A60 , 32'h000330A4 , 32'hFB80C110 , 32'hF67FB760 , 32'h04E0B8F8 , 32'hFFFF8A11 , 32'h00B86AAD , 32'h0000D327 , 32'h0350FDD8 , 32'h15B7AF40 , 32'hFFFC4FE3 , 32'h04DC6808 , 32'hFFFCAE48 , 32'hFFFF0077 , 32'hF8DF1A98 , 32'h04FC3700 , 32'hFE9CC360 , 32'hFFFFCD28 , 32'hEF3FE100 , 32'h00008B50 , 32'h00020D99 , 32'hFE316DD4 , 32'h0001ECE6 , 32'h0000E8B1 , 32'hF40E9C60 , 32'h0525D418 , 32'h0000DD91 , 32'hFFFED6A8 , 32'hFFFFE206 , 32'hFFFE9DAA , 32'hFFFE3178 , 32'h06E8A148 , 32'h00E86D36 , 32'hFFFEA5AD , 32'hFFFF2683 , 32'h030DFE48 , 32'h08425940 , 32'h00039D05 , 32'hFFFF9DB7 , 32'h0371537C , 32'hFFFC8C59 , 32'hFFFD665A , 32'hFDE8887C , 32'hFD660AD4 , 32'h017C52C0 , 32'hFDE388C8 , 32'hFFFF4576 , 32'h000131DC , 32'hFFFA2880 , 32'hFFFF04EA , 32'h0000F7EF , 32'h00E0B262 , 32'hFFFF6D53 , 32'h0000AEB4 , 32'h01884850 , 32'hFFFF4748 , 32'h041E8F98 , 32'h010A765C , 32'h0001559D , 32'hFFFFC1D8 , 32'hFFFEB1FA , 32'h17434CC0 , 32'h0243A390 , 32'hFD7B4E4C , 32'h02440568 , 32'hFFFFD5ED , 32'hFE61E8B4 , 32'hFFFF8403 , 32'hFFFFBAA6 , 32'h038CF5B4 , 32'h00A6621C , 32'h02291134 , 32'h000112FE , 32'hED76A0E0 , 32'h017FE59C , 32'h0337C0FC , 32'h16404980 , 32'hFB9FF610 , 32'h253A4CC0 , 32'h006AC8A7 , 32'hFB15B010 , 32'hFFFE6BD8 , 32'h0001C426 , 32'h000057A7 , 32'hFF2246BE , 32'h0A160EC0 , 32'hFE370E20 , 32'h0017E0A4 , 32'hFEF23B44 , 32'hFD986E58 , 32'hFFFC89BC , 32'hF9B995C0 , 32'hFFAE3EAE , 32'h000241EE , 32'h082AA840 , 32'h00013EEA , 32'h0C40FA60 , 32'hFF9FC267 , 32'h000160C2 , 32'h0000F87A , 32'hFFFF8CD4 , 32'h0001275B , 32'hFFFFE855 , 32'h00006843 , 32'hFE19E634 , 32'hF939EE70 , 32'h09016860 , 32'hF5904240 , 32'hFC0B66F4 , 32'hFE9BF200 , 32'h0001BC1A , 32'h0001856D , 32'h00015295 , 32'h00015ABD , 32'hFFFE6C3E , 32'h01D73CD0 , 32'h0A380CC0 , 32'hEBA444C0 , 32'hFFFF32F2 , 32'hFFFFDB10 , 32'h00004818 , 32'h000003C4 , 32'h09DF8890 , 32'h1033F7A0 , 32'h0000B8B5 , 32'h00018B87 , 32'h00013EB1 , 32'hF137A8A0 , 32'h0C360F10 , 32'hEAF73B40 , 32'hFFFF0EB5 , 32'h00011699 , 32'h000006E5 , 32'hFD7DA31C , 32'h01991200 , 32'hFFDFA2A2 , 32'hFFFEE86F , 32'h0015CF21 , 32'hFFFE2791 , 32'hFDEC3700 , 32'h0000B91D , 32'hEEFDFD20 , 32'h000249E7 , 32'hEB455960 , 32'h0015AF9E , 32'h0EEF3E50 , 32'hE599EDC0 , 32'h00023939 , 32'h06830C18 , 32'h023ABD70 , 32'h00013BA7 , 32'hF9059F38 , 32'hFFFE7C2E , 32'hFFAE98B8 , 32'h0BDEB150 , 32'h0EA95840 , 32'h000133B4 , 32'hFFFE33D6 , 32'h0807BDB0 , 32'h00016559 , 32'hF8194088 , 32'hFFFFDA6C , 32'hFE7146FC , 32'hFFFE9BE2 , 32'hFD2AE144 , 32'h000093F3 , 32'h0000F90D , 32'hFFFEEC56 , 32'hFD01E868 , 32'hFED77360 , 32'hFFFF5DB9 , 32'hFFFE8D1C , 32'hFFFF8E96 , 32'h00006BE7 , 32'hFAA9C9C0 , 32'hFA4AFDA8 , 32'h03FCE020 , 32'h05B30690 , 32'h01D0A50C , 32'hFFFF2956 , 32'hFFFEC57E , 32'hFFFF61BE , 32'hFF5DA658 , 32'h0000B25B , 32'h00008ABA , 32'hFF130C6C , 32'h182D3380 , 32'hFFFDACF8 , 32'hFFC54912 , 32'h003A4585 , 32'h03222F3C , 32'h0AA361F0 , 32'h00007B3C , 32'hF4D11D30 , 32'h12F0E6C0 , 32'hFCE39070 , 32'hFFFF2674 , 32'hF2F7F5B0 , 32'h11C50AC0 , 32'h0DBB2A00} , 
{32'hFA4D7358 , 32'h12C58AC0 , 32'h00011F05 , 32'hF0179290 , 32'h0000DCFE , 32'hFE7C8184 , 32'hFFFC0D80 , 32'h00016B91 , 32'h00005855 , 32'hFFFFDFAD , 32'h06D87C70 , 32'h15997A60 , 32'hFE07F26C , 32'hFFFEF941 , 32'h000106FA , 32'hF2CF0450 , 32'hFFFD47CE , 32'h18F082E0 , 32'h01B29B68 , 32'hFFFE1EC7 , 32'h0000BED8 , 32'h01E8E11C , 32'hF7777290 , 32'hFA2679F8 , 32'hFEA0BE7C , 32'hFFFE55DE , 32'h0279B8E4 , 32'h032768AC , 32'h00010C81 , 32'h05F55D78 , 32'h0000D39E , 32'hFDB7317C , 32'h00023276 , 32'h0000AF0C , 32'hFFFD96A2 , 32'hFD48C000 , 32'h0F731350 , 32'hF2A46280 , 32'hFFFEC940 , 32'hF41E2CA0 , 32'hFFB4AFBB , 32'h0000F636 , 32'h00021A19 , 32'hFF7DCE3A , 32'hF303B4A0 , 32'hEB520580 , 32'h0CAA3860 , 32'h0000C9AE , 32'hFA510D30 , 32'hF73ACB10 , 32'h00DFABD3 , 32'hFFFFECD3 , 32'h02BCAA84 , 32'h0D02A4A0 , 32'h075D09D8 , 32'h00019888 , 32'hFF7D161C , 32'hFFFDD971 , 32'h0000EE25 , 32'hFB829540 , 32'h01CC3714 , 32'hF9234DF8 , 32'h0E1CD8C0 , 32'hFFFDE998 , 32'hFB793898 , 32'hFFFF6ED8 , 32'hE8A625C0 , 32'hFFE534DE , 32'h00020164 , 32'h00BDDACE , 32'h05F334B0 , 32'h056FFFC8 , 32'h0000EF5C , 32'h00015076 , 32'hFFFF6214 , 32'h055381C8 , 32'hFFA891F8 , 32'h0000573B , 32'h00B335B2 , 32'h00530773 , 32'hFFFEC582 , 32'hEA206280 , 32'hFD579EAC , 32'h0001F40D , 32'h00EA23DB , 32'hF609C420 , 32'h001D3CBE , 32'hFFFD762A , 32'h0000AFF9 , 32'hFF78A2BA , 32'hFFFF6C7A , 32'h07183DB0 , 32'hFFFE4176 , 32'h03657558 , 32'hFFDFDC44 , 32'h000091A2 , 32'hFFFEA555 , 32'hFFFEBCB9 , 32'h0000F00E , 32'hF7F14600 , 32'h000FA415 , 32'hFFFFA775 , 32'hE6F8D480 , 32'hF2547840 , 32'h05A6EE20 , 32'hFFFF5694 , 32'h0047C995 , 32'h000103CC , 32'hFC72FF44 , 32'hFC786398 , 32'hFFFFA72E , 32'h011E15FC , 32'h000091B1 , 32'hFFFF9F6F , 32'h0859D560 , 32'h056CDC80 , 32'hFF3C4EA9 , 32'hFFFEDFEA , 32'h01E699D8 , 32'hFFFFADAF , 32'hFFFCF939 , 32'hFE8197CC , 32'hFFFFB781 , 32'hFFFED6E7 , 32'hFB4528F0 , 32'h004CCA53 , 32'h00011322 , 32'hFFFEFF64 , 32'hFFFFF150 , 32'h0002859C , 32'hFFFF2BD7 , 32'hFE64DB94 , 32'h0438B8A8 , 32'h00007DAC , 32'hFFFEF959 , 32'h14AC66A0 , 32'hFAB374E0 , 32'hFFFDAA1B , 32'hFFFFABA5 , 32'h0B0158C0 , 32'h00023EF0 , 32'hFFFF473C , 32'h01E8E738 , 32'h028975E0 , 32'h053B4328 , 32'h01A1F774 , 32'hFFFD42D4 , 32'h00006D19 , 32'h008CFD38 , 32'h00006F79 , 32'h0002F43F , 32'hFEE7B894 , 32'h00013481 , 32'h0001F382 , 32'hF2114390 , 32'hFFFFDE0B , 32'h0059B954 , 32'h018C798C , 32'hFFFFE5E1 , 32'h0000E7DF , 32'h00005614 , 32'hF3EE85E0 , 32'h06410F10 , 32'hFBFC2F80 , 32'hF7A74450 , 32'hFFFE6E72 , 32'hF4E927A0 , 32'hFFFE819D , 32'hFFFD1B55 , 32'h13324620 , 32'h003E27C8 , 32'h043C0878 , 32'h00010BC9 , 32'h01301BF0 , 32'hFFA11D56 , 32'hFEC98B5C , 32'h07B89CF8 , 32'hFD3A1BB4 , 32'hFC010A00 , 32'h02C27BDC , 32'hFE8D9408 , 32'hFFFF9C1E , 32'hFFFFB55C , 32'h0000AFC5 , 32'hFA4CBE60 , 32'hEF7CD780 , 32'h006238A4 , 32'hFF188DD3 , 32'hFC09D7F8 , 32'h0380AFA8 , 32'hFFFF0213 , 32'hFC3F5C1C , 32'h0A4D6AC0 , 32'hFFFE9201 , 32'hF977BC10 , 32'hFFFE288E , 32'hFD931924 , 32'hEF4CE7E0 , 32'h00001AB6 , 32'h0000769A , 32'hFFFFC4CB , 32'hFFFEC4AB , 32'hFFFFD553 , 32'h00017F69 , 32'hFA93B208 , 32'hEFEC35C0 , 32'h05426B08 , 32'hFE96BD34 , 32'hF94600C8 , 32'h04B6A7B0 , 32'hFFFEAA06 , 32'h00006F74 , 32'h0001CD14 , 32'h00012545 , 32'hFFFCBF49 , 32'hFEE03D6C , 32'hFADF1888 , 32'hFE566F54 , 32'h0001E443 , 32'h00020B74 , 32'hFFFFA444 , 32'hFFFF25C0 , 32'h0414CA50 , 32'h1392DB40 , 32'h0001E433 , 32'hFFFFE151 , 32'h00001F48 , 32'hE30F0C40 , 32'hDB9C6D00 , 32'h116A4C00 , 32'hFFFDE88D , 32'h00008432 , 32'hFFFE51C1 , 32'hFEADC97C , 32'h022A0C00 , 32'h10161EC0 , 32'hFFFFA0B5 , 32'h0068F20D , 32'hFFFD57FE , 32'h1B55D9A0 , 32'h000004DF , 32'h18F7AF60 , 32'h000108A9 , 32'h0B5D1240 , 32'hF49B7930 , 32'hFCBEC43C , 32'hF5516790 , 32'h0001BA36 , 32'hFCF41E10 , 32'h0068D7C8 , 32'h0001D539 , 32'h04A97F80 , 32'h0001F997 , 32'h04468638 , 32'h151ED0C0 , 32'h038462F8 , 32'hFFFFEA4A , 32'h00012519 , 32'hFC1E95E0 , 32'h00020C2A , 32'hF712C340 , 32'h0000A954 , 32'h00404E61 , 32'h000070D6 , 32'h02F6F820 , 32'hFFFEEF44 , 32'hFFFF4115 , 32'hFFFFB67C , 32'h084983A0 , 32'h01B8C570 , 32'hFFFE3CBF , 32'h0000406A , 32'h00001DEF , 32'h0002510A , 32'h05F321C0 , 32'hFACCCFF0 , 32'hFFA6C3BE , 32'h00840E52 , 32'hFC2669E8 , 32'h0000C925 , 32'h00006371 , 32'h000063EA , 32'h0299D73C , 32'h00000111 , 32'hFFFF901B , 32'hFD065244 , 32'h1CC4D8A0 , 32'hFFFFC996 , 32'h033C9F88 , 32'h0458E0F8 , 32'h004EEF7F , 32'h02BE3F78 , 32'h0000AF9C , 32'h0755A960 , 32'h1247A480 , 32'hFF480FAA , 32'h0000D767 , 32'hFBAF23D8 , 32'hFCC922F8 , 32'h0A09F580} , 
{32'hF7D91380 , 32'h0D4C7670 , 32'h00026D04 , 32'h079740D0 , 32'h0000C58D , 32'hFCB2D9AC , 32'h0001BE3F , 32'h0000BA53 , 32'h000032A7 , 32'h0001BB06 , 32'hF8A812D0 , 32'h06953D30 , 32'h011BC604 , 32'h0000D49B , 32'hFFFE7662 , 32'h207D7180 , 32'h0001CE94 , 32'h0BAEBDC0 , 32'hFBB35528 , 32'hFFFE59C6 , 32'hFFFE8290 , 32'h0310EB88 , 32'h11570160 , 32'h0712D990 , 32'hFDBE9F1C , 32'h00014CDD , 32'h02F2F19C , 32'h01110200 , 32'h0002FDE1 , 32'h0E0EC490 , 32'hFFFE97EC , 32'h07BE8C90 , 32'h00008849 , 32'h00009898 , 32'hFFFE6DDB , 32'hF6142320 , 32'hFC223D54 , 32'hFC689B40 , 32'hFFFD1BEB , 32'h13E2C480 , 32'h0C85D890 , 32'h00012C0D , 32'hFFFE4D44 , 32'h00D54F3A , 32'h0991BBE0 , 32'h06CFCA90 , 32'h0CCD5AA0 , 32'hFFFE5480 , 32'hF5C53920 , 32'hF0BC9010 , 32'h0042CD8F , 32'hFFFFC357 , 32'h059D9970 , 32'h04786740 , 32'hFDF2D7B0 , 32'hFFFD75D1 , 32'hFFFC0B5C , 32'hFFFF6D64 , 32'h0000E9E2 , 32'h04997458 , 32'h006F6AB1 , 32'hFF8066E5 , 32'h008D3EDA , 32'h000158FF , 32'hF70BC190 , 32'hFFFE5B0E , 32'h0F742570 , 32'hFD67352C , 32'h0000D90C , 32'h031CB080 , 32'h05C8A580 , 32'hFA0B9F68 , 32'h00016077 , 32'hFFFCC856 , 32'hFFFF36F8 , 32'h041F2118 , 32'hFDAEA6E4 , 32'h00015DF6 , 32'h12996240 , 32'hFE74C614 , 32'h0000176E , 32'hF4B0A770 , 32'hFD0B293C , 32'hFFFF21F0 , 32'h01C5CD50 , 32'h023C7180 , 32'h04DC4C78 , 32'hFFFE78FC , 32'h000109A7 , 32'hF63BCD90 , 32'h0002F509 , 32'hF52445E0 , 32'h0000A9FC , 32'h052957F0 , 32'h0019F211 , 32'hFFFF2C35 , 32'hFFFF0A3C , 32'h00000368 , 32'h00024278 , 32'h04F5ADE8 , 32'h02D05350 , 32'hFFFF5469 , 32'hFD2AD314 , 32'h0D23AEF0 , 32'hFB39C1A8 , 32'h00001100 , 32'h0004DD82 , 32'h0000F388 , 32'h05BB3FC0 , 32'h00836919 , 32'hFFFEB7E3 , 32'h015BF9A8 , 32'h00016514 , 32'h00018DB8 , 32'h053D5658 , 32'h03A0E5D0 , 32'hFD472F60 , 32'hFFFE7881 , 32'hF9076A80 , 32'h00016C06 , 32'hFFFDCED3 , 32'h02ED7F30 , 32'h00001EE8 , 32'hFFFF7A60 , 32'h0D9564A0 , 32'h03ABB658 , 32'h00022842 , 32'hFFFF7C49 , 32'h0001082F , 32'hFFFEAA3B , 32'h0001DC81 , 32'h0A564D10 , 32'h01E58F3C , 32'h00009012 , 32'h0001B103 , 32'hFF206156 , 32'h06465D08 , 32'h000031C9 , 32'hFFFE505E , 32'h077E0C48 , 32'hFFFFABED , 32'h0000C158 , 32'h005EB9E2 , 32'hF20F04F0 , 32'h01817BB8 , 32'h00043E34 , 32'h00027F92 , 32'h0001D202 , 32'hFCF7ABA8 , 32'hFFFF545A , 32'hFFFEB19D , 32'h0352FA5C , 32'h000212EE , 32'h00019925 , 32'hFF26794E , 32'h0002BBE6 , 32'h045A13D0 , 32'h0134AB3C , 32'h0001113B , 32'h000179CA , 32'hFFFE6F9E , 32'h07F99F20 , 32'hFF476C57 , 32'h046A1EB0 , 32'hFFD4E14F , 32'h0000D3DF , 32'h0F919C90 , 32'h00009AB7 , 32'h0001317D , 32'hF9A607A0 , 32'h0292ED10 , 32'hF923D2B0 , 32'h0000373B , 32'h05DE0960 , 32'hFA7EBE68 , 32'h055CD120 , 32'hF0D75800 , 32'hFF674A51 , 32'hF9D7F9E8 , 32'hFF0D728B , 32'hF5F36B80 , 32'h00008325 , 32'h0000ECBA , 32'h0000B564 , 32'h0577D6C8 , 32'hC8948D00 , 32'hFE54BCDC , 32'hFF61B206 , 32'h0A615070 , 32'hF67D42B0 , 32'hFFFD76B3 , 32'h0B71BE90 , 32'hFF6B2C27 , 32'h0001CE28 , 32'h03F65888 , 32'hFFFF2D6A , 32'h0574EE20 , 32'hFD335C48 , 32'h0000DC6F , 32'hFFFF33AD , 32'h0000FC95 , 32'h00039057 , 32'hFFFFFBA9 , 32'h00001F9C , 32'hFBD15DD0 , 32'h0ACB10C0 , 32'hFD75D7B4 , 32'h021736AC , 32'h04390EA0 , 32'h0539EC08 , 32'hFFFF352B , 32'hFFFE04FF , 32'h000343D9 , 32'h0000013B , 32'hFFFE68EB , 32'h040BA940 , 32'h0C0A42C0 , 32'h01EF3A80 , 32'h000036AC , 32'h00005ADE , 32'hFFFF465E , 32'h00021028 , 32'h0095A4E3 , 32'hED4EB1E0 , 32'h0000BFB2 , 32'hFFFEE26C , 32'hFFFFEFBD , 32'hE8E16D80 , 32'hF1438FD0 , 32'hECB023A0 , 32'hFFFED298 , 32'hFFFFBA18 , 32'h000059AE , 32'hFE322B04 , 32'hFF521EBF , 32'hFC384064 , 32'hFFFF563E , 32'hFE707B70 , 32'h00023C26 , 32'h02A873D0 , 32'h000153CC , 32'hFC4BCDF4 , 32'hFFFEADF6 , 32'hE830E260 , 32'hFAC0B370 , 32'hF10EA010 , 32'hEF337B60 , 32'h000008F3 , 32'h02DCDD6C , 32'hFFD962B6 , 32'hFFFBB67B , 32'hFA9BCF98 , 32'h0001990F , 32'h010DC8C4 , 32'hF8C97E40 , 32'h01ECB5C0 , 32'h00002BBF , 32'hFFFEF356 , 32'hFA5E9358 , 32'hFFFCF922 , 32'h002EF3C0 , 32'hFFFE22DA , 32'h009BF43B , 32'hFFFEE206 , 32'h00384A5C , 32'h0000B641 , 32'h0004FE8B , 32'hFFFF3475 , 32'hFD0C8230 , 32'hF1F21A70 , 32'hFFFF0BB8 , 32'hFFFEE885 , 32'hFFFFCEE4 , 32'h00013631 , 32'hFC207034 , 32'h0E0A2A30 , 32'hF8326E00 , 32'h1591C180 , 32'h10341260 , 32'hFFFF1640 , 32'h00020BAB , 32'h0001EFD7 , 32'hFCC2225C , 32'hFFFDD767 , 32'hFFFEE2A5 , 32'h007C449E , 32'hFFA55055 , 32'h0001E823 , 32'h1E532960 , 32'hFFE46EAE , 32'hFB91DD68 , 32'h03A80E38 , 32'h00008483 , 32'h026F6EA4 , 32'h0CE29EF0 , 32'h02BED214 , 32'hFFFFA376 , 32'h18B9A1A0 , 32'hF5DB1610 , 32'hFFF38CDB} , 
{32'h0D309AC0 , 32'h02FA942C , 32'h00009125 , 32'hFB7C9358 , 32'h0000AF45 , 32'hFBB811C0 , 32'h00022FCA , 32'hFFFFE0DE , 32'h00000A43 , 32'h0003317F , 32'h0B94EF30 , 32'hECE7F480 , 32'hF7341750 , 32'h000000EF , 32'hFFFD9391 , 32'h0227225C , 32'hFFFE0A59 , 32'h03A425E4 , 32'hFE92D06C , 32'hFFFFD2F2 , 32'h0000D2BF , 32'h00104D9D , 32'hEE49CEE0 , 32'h02BD7A34 , 32'h05D0C990 , 32'h00006669 , 32'hFF8B1EBB , 32'hFBC87880 , 32'h0001853F , 32'hFA3601D8 , 32'hFFFF040B , 32'hF401B120 , 32'h0000CA45 , 32'h0000B8F3 , 32'hFFFE9CB4 , 32'h0FA8F680 , 32'hF51B7D00 , 32'hF2EAA8C0 , 32'h00001405 , 32'hF5593E50 , 32'hF4771C10 , 32'hFFFFF0C5 , 32'h0000CEE5 , 32'hF9F892F8 , 32'hF1C405F0 , 32'hF5989560 , 32'hF9464DD0 , 32'hFFFFA68A , 32'h00D7DECC , 32'h12FA4F20 , 32'hFF480AEB , 32'hFFFD76CA , 32'hFC6147DC , 32'hF6EF5890 , 32'h01ACF4A0 , 32'h0001104B , 32'hFF8C91D0 , 32'h0000800F , 32'hFFFEFFA0 , 32'h05492718 , 32'h01C2898C , 32'hF80173C8 , 32'h10916C40 , 32'h00024098 , 32'hCDE0F380 , 32'h0000EB9A , 32'hFF046641 , 32'hFF096D14 , 32'h00011261 , 32'hFEC9FE80 , 32'h12844D80 , 32'hFF1AFCB3 , 32'hFFFE8CD4 , 32'hFFFFA5AD , 32'hFFFEE7D4 , 32'hF8AD18F0 , 32'hFC1CF74C , 32'h0000F64F , 32'hFB24DF80 , 32'hFF42479A , 32'h00005762 , 32'hEAF3DE00 , 32'h02FD5A1C , 32'hFFFFC1FE , 32'hFD87212C , 32'hFCE7E880 , 32'h019D0188 , 32'h00005C8C , 32'hFFFFFC2E , 32'h11075C60 , 32'h00020780 , 32'h05EB0D68 , 32'h00026C13 , 32'hFEADA1E0 , 32'h016A3C54 , 32'h0000E578 , 32'hFFFE3B35 , 32'hFFFE2124 , 32'h000218DB , 32'h11624FE0 , 32'hFE8710BC , 32'hFFFED548 , 32'h05DB0C78 , 32'h0ED2C7C0 , 32'h00AC0A53 , 32'hFFFCF8DD , 32'h00352FB7 , 32'h0000E4B9 , 32'h0303B08C , 32'hFCD32AB8 , 32'hFFFF6F73 , 32'h0408A908 , 32'hFFFFE5AD , 32'h0000E9D1 , 32'hFE5BAB78 , 32'h03A01048 , 32'h01BF48A4 , 32'hFFFE880E , 32'hF2B3C030 , 32'hFFFD58D6 , 32'hFFFECE59 , 32'h03763428 , 32'h0000C289 , 32'h0001D6F0 , 32'hDB797CC0 , 32'hFF7D3E6C , 32'h000132F9 , 32'h0000FC1E , 32'h0000F1FE , 32'hFFFF6836 , 32'h00012097 , 32'h00FAB8B2 , 32'hF6D5D7D0 , 32'hFFFFF02C , 32'h0001DEF6 , 32'h05623DF8 , 32'hF5F461B0 , 32'h0001718D , 32'hFFFFBCD4 , 32'h04888468 , 32'h0002344C , 32'h0001AF4E , 32'hFF76141C , 32'h000C5CD2 , 32'h004B22DD , 32'hFFB0D636 , 32'h00033C99 , 32'h0000821F , 32'h003EDBCD , 32'hFFFF41BB , 32'h00002251 , 32'h02C8E1E0 , 32'h0001AF32 , 32'h00038ADF , 32'hF83B16A0 , 32'hFFFE36DF , 32'h0125CA9C , 32'h004E9B25 , 32'hFFFFE3B5 , 32'hFFFE3460 , 32'h00002BBF , 32'h01EB232C , 32'h03C3B6DC , 32'h0373F00C , 32'hFC73FD44 , 32'h0000C01F , 32'hFF6C171D , 32'h00010FB1 , 32'h0001A8B8 , 32'hFB8B24C0 , 32'h02D617A8 , 32'h04794E90 , 32'hFFFEF707 , 32'hF5548B50 , 32'h02AE12C4 , 32'hF9092838 , 32'hF707DC80 , 32'hFC97967C , 32'hFD69464C , 32'hFE1649D4 , 32'h00742F95 , 32'hFFFF70DF , 32'h00036EF0 , 32'h0001C983 , 32'h08451020 , 32'hF7F676E0 , 32'h047A9930 , 32'hFE2D1098 , 32'hFECC5B28 , 32'hFE3DC33C , 32'h0002B759 , 32'hF51A2820 , 32'hF7E0C5A0 , 32'hFFFF9490 , 32'hF8CB8518 , 32'h00003E3C , 32'hF7AD5BF0 , 32'hEE1D4480 , 32'h0001F8DB , 32'h000158C1 , 32'h00043B34 , 32'h00005DDD , 32'hFFFD4374 , 32'h0000355B , 32'hFC29CF1C , 32'h04605B30 , 32'h19220E00 , 32'h042C8AB0 , 32'hF7FC8960 , 32'hF60E1E70 , 32'h0000E984 , 32'hFFFFAAD4 , 32'h000172A8 , 32'h0000F0FD , 32'h00036FE1 , 32'hFDC818A8 , 32'h06BD6B50 , 32'h0BBF8B40 , 32'h000051BA , 32'h00006C5B , 32'h00000570 , 32'hFFFFE7BC , 32'h028FB234 , 32'hF2C4E7B0 , 32'hFFFF00FF , 32'hFFFF0FF9 , 32'h00018A25 , 32'hFC7DC7B4 , 32'h0F243D40 , 32'h176617E0 , 32'h00007E93 , 32'h0000F790 , 32'h00027407 , 32'hFFBDA843 , 32'hFF050881 , 32'hF9736740 , 32'h0002C371 , 32'hFFC18B34 , 32'h0000BC81 , 32'hFBD74130 , 32'h0000484C , 32'hF3DD1CA0 , 32'hFFFFF8B8 , 32'hFE147A6C , 32'hFBF4E060 , 32'hDF5524C0 , 32'h0FEA73E0 , 32'hFFFF8739 , 32'h0A0AC930 , 32'h00F8815E , 32'h0001C048 , 32'hFE11A0EC , 32'hFFFE1D65 , 32'hFE7914C4 , 32'hF31AB6B0 , 32'hF5DE5A50 , 32'h0000E463 , 32'h0001A752 , 32'hFC1C1E4C , 32'h00027945 , 32'h05222B90 , 32'hFFFD84B8 , 32'hFEDBBC8C , 32'hFFFF4985 , 32'hF1B2B110 , 32'h00021836 , 32'h000069C0 , 32'h0000EDFC , 32'h111F9720 , 32'h06DFD588 , 32'h00009852 , 32'hFFFE0310 , 32'h0000F4DA , 32'hFFFF6C18 , 32'h01C35FA8 , 32'h081556B0 , 32'hF7B52450 , 32'hF5948EB0 , 32'h0C234290 , 32'h00003294 , 32'h0002A91B , 32'hFFFF666A , 32'hFD005738 , 32'h0001849C , 32'h00009E12 , 32'hFF7E0313 , 32'hFE049E74 , 32'h00022048 , 32'h10C2B320 , 32'hFCD65D84 , 32'h000A7C96 , 32'hF54A2240 , 32'hFFFEB828 , 32'h01552B44 , 32'hFD6520F4 , 32'h0287BD54 , 32'h00015FE3 , 32'h0D769D00 , 32'hF7194FF0 , 32'hF7FA16F0} , 
{32'h082DCEE0 , 32'h08A750E0 , 32'hFFFEA6BF , 32'hF6C38270 , 32'hFFFF4FE4 , 32'h02040AC8 , 32'h00014097 , 32'hFFFF9C8D , 32'hFFFE45F7 , 32'h00033C9B , 32'h0179C980 , 32'hE8308FA0 , 32'hF9389C30 , 32'hFFFF3BF1 , 32'hFFFEF62B , 32'h1A283B80 , 32'h00014DB6 , 32'h0331836C , 32'h04F758D0 , 32'hFFFF3FB8 , 32'hFFFF86A7 , 32'h00217D4A , 32'h0DDDE370 , 32'h06F675A8 , 32'hFF165DD9 , 32'h0002BB48 , 32'hFEDFC5BC , 32'h000EA277 , 32'hFFFE921C , 32'hE71E7100 , 32'h0001FAE3 , 32'h0145EFB8 , 32'h0003BB7B , 32'h000107E6 , 32'hFFFE65CE , 32'h19777B40 , 32'h0F0A4FD0 , 32'hF06E4F30 , 32'hFFFE54D2 , 32'h06664028 , 32'h0014203C , 32'hFFFE63BC , 32'hFFFDFA8A , 32'h020C1F38 , 32'hECF367C0 , 32'hFDF2C230 , 32'hFF172AE0 , 32'hFFFF250E , 32'h0AF3B660 , 32'h00C64636 , 32'hFF68194D , 32'h00006D25 , 32'hFFE64645 , 32'h13AB7A40 , 32'h0297AA50 , 32'h00012446 , 32'h0049EC44 , 32'hFFFE3684 , 32'hFFFF7AEC , 32'h0172C1EC , 32'hFE883C58 , 32'h00259C23 , 32'hF4BABBC0 , 32'h00003A74 , 32'h03B43104 , 32'h00012536 , 32'hF20A0060 , 32'h02958EB8 , 32'hFFFF60A7 , 32'hE7A92100 , 32'h05C69BA8 , 32'h05411328 , 32'h00007DEC , 32'h00026E49 , 32'hFFFF614C , 32'hFF979B87 , 32'h049D74D8 , 32'h000197BB , 32'hFA402360 , 32'hFEE63ACC , 32'hFFFF27A3 , 32'h0F1FC560 , 32'h02EBE218 , 32'hFFFE4230 , 32'h05ED6440 , 32'h0AF9B4A0 , 32'h003650E9 , 32'h0000BD1B , 32'hFFFF90E7 , 32'h12CD2EC0 , 32'h00002EF2 , 32'hF28A6DC0 , 32'h00016F8F , 32'h09071510 , 32'h0024022C , 32'h0002719E , 32'h0001FE0D , 32'hFFFF494F , 32'h000132C1 , 32'h07348FF0 , 32'h02933224 , 32'hFFFE40FA , 32'h042330E0 , 32'hF7F640D0 , 32'h015AA7AC , 32'h0000A6D8 , 32'hFFFF5B33 , 32'hFFFDA66A , 32'hFC9B33C8 , 32'hEB74D980 , 32'h0000A4F8 , 32'h0D40BF50 , 32'hFFFDB78B , 32'hFFFEE131 , 32'h0A263F30 , 32'h05C10440 , 32'h00ED85C8 , 32'hFFFD5E8B , 32'h06AFC928 , 32'hFFFE2B29 , 32'h00010143 , 32'hFFD830D4 , 32'hFFFF4F9C , 32'h00024D5A , 32'h10C4BFE0 , 32'hEC499C80 , 32'h0000B089 , 32'hFFFCBE98 , 32'h00024B7C , 32'h00017F62 , 32'h00001D3D , 32'h030AA4F4 , 32'h0635BF18 , 32'h0000EF40 , 32'hFFFE7639 , 32'h1696C380 , 32'h00421337 , 32'hFFFE74AF , 32'h00002EE8 , 32'h0118EE10 , 32'h00020E5F , 32'hFFFEEB07 , 32'hFF70FDF4 , 32'h049A82B8 , 32'hFF909038 , 32'hFD98BB7C , 32'hFFFF969E , 32'hFFFE5D31 , 32'hFF035BB1 , 32'hFFFBFEAD , 32'hFFFD4FC7 , 32'h0758C2D0 , 32'hFFFDD6E3 , 32'h0000260F , 32'hFBEF54F0 , 32'hFFFFD947 , 32'h0112EE54 , 32'h01E47874 , 32'hFFFDFC63 , 32'hFFFED635 , 32'h000086F8 , 32'hFDA875F8 , 32'h0544DA38 , 32'hFB94DB48 , 32'h058A88A8 , 32'hFFFF538E , 32'h0B92A250 , 32'h00007E0F , 32'h00010D92 , 32'h149C88C0 , 32'h056A2970 , 32'hF7F3F510 , 32'hFFFCE263 , 32'hFDCAF850 , 32'hFBF59B98 , 32'h00F26CA3 , 32'hF1207720 , 32'h067D8020 , 32'hFD68EEC0 , 32'hFF81B4B7 , 32'hF66B4120 , 32'hFFFFDEE8 , 32'hFFFFD560 , 32'h00017A22 , 32'hFD592DF0 , 32'hF1DD0470 , 32'h09B3F5F0 , 32'hFF80253A , 32'hF6A2B270 , 32'h09669EA0 , 32'hFFFD113B , 32'hF77C0480 , 32'h05AE9C58 , 32'h0001A8D9 , 32'hFFE34035 , 32'h00015ABC , 32'hFCCD306C , 32'h0D8D48F0 , 32'h00011486 , 32'h00048799 , 32'hFFFD89E7 , 32'hFFFEE55F , 32'h0001591B , 32'hFFFEFFAD , 32'hFF92E0D4 , 32'hF85729F8 , 32'h09DEFE00 , 32'hFA9FCC38 , 32'hF4E836E0 , 32'hFD33DE28 , 32'h00000421 , 32'h0001C1F9 , 32'hFFFD16F4 , 32'hFFFE1BDC , 32'hFFFE6E86 , 32'h00D1DD3A , 32'hFC158610 , 32'hFB027D80 , 32'h000104AC , 32'hFFFD3310 , 32'h0001F127 , 32'hFFFEF4D4 , 32'hFD8F4C0C , 32'h084186D0 , 32'hFFFD44F8 , 32'hFFFFB3B9 , 32'h00016C27 , 32'hFF9520BB , 32'h0C9FDE00 , 32'hEA458900 , 32'hFFFE7B1C , 32'h0000B1C7 , 32'h00004BF8 , 32'h0192A8D0 , 32'h01BD4BC0 , 32'h00C483AE , 32'h00011B71 , 32'hFFEC405E , 32'h00023EFE , 32'hEFD05F80 , 32'h00033551 , 32'h056E3BE8 , 32'h000016CA , 32'h0494D2B0 , 32'hFAC69830 , 32'hE93D9B00 , 32'h065DB908 , 32'h00019AEA , 32'h04B47AC0 , 32'h002B2A5C , 32'h00018A20 , 32'h08053A40 , 32'hFFFEDF2C , 32'hFCC9F154 , 32'h0053DDDA , 32'hFC0F4A34 , 32'hFFFDE5AB , 32'h000217F7 , 32'hFD5F9D0C , 32'h0002F442 , 32'h06E6B270 , 32'h00009773 , 32'h0016BF81 , 32'hFFFFA399 , 32'h0D18E680 , 32'hFFFEF6E4 , 32'hFFFD49FD , 32'h0000571D , 32'h0CD04300 , 32'h05708D30 , 32'hFFFF911F , 32'h0000B1AD , 32'hFFFFD49C , 32'hFFFDA2C3 , 32'h0A7A97C0 , 32'hF6F73020 , 32'hF516DE00 , 32'h22AF7D40 , 32'hFBA9D770 , 32'h00010F7D , 32'hFFFEE749 , 32'h0000BAF9 , 32'hFF90995B , 32'h00006E61 , 32'h0000C080 , 32'h03EA953C , 32'hF31B27A0 , 32'hFFFF03EC , 32'hE88CCF20 , 32'hFA29B6A0 , 32'hF23248E0 , 32'h0E042130 , 32'h0000330A , 32'hFECEA95C , 32'hFAEA1A28 , 32'hFF590CD3 , 32'h00010D47 , 32'hF2B0E220 , 32'hFE994564 , 32'h11157EC0} , 
{32'hF6822E40 , 32'h1ED6C0C0 , 32'hFFFF5AFA , 32'hFF4A96BE , 32'hFFFC1444 , 32'h01728A80 , 32'h000228A4 , 32'hFFFF8D3D , 32'hFFFECD8C , 32'hFFFE297B , 32'hF678A190 , 32'hF8EEE528 , 32'hFBC2D910 , 32'h00025A05 , 32'h0003038D , 32'hEE6B80A0 , 32'hFFFEC5CF , 32'hFCB0FDC4 , 32'hFF5F8488 , 32'hFFFCE489 , 32'h0000950E , 32'hFCD1420C , 32'h04DDD0A8 , 32'hF796CAF0 , 32'h07D215A0 , 32'h00027756 , 32'hFF7FBBB5 , 32'h03D6ABD0 , 32'hFFFF23C4 , 32'h027AEDC4 , 32'hFFFE8B57 , 32'hFD692A60 , 32'hFFFEBB4F , 32'hFFFF534E , 32'h00029422 , 32'hF7EBCDE0 , 32'hF8A40420 , 32'h07499468 , 32'h0000F8D7 , 32'h0395B1C4 , 32'hF2D77DD0 , 32'h00013476 , 32'h00005339 , 32'h04720238 , 32'h0370E4B0 , 32'hF56FE840 , 32'hF10D7A00 , 32'h0001A4E8 , 32'hFC81CB18 , 32'hE9781020 , 32'h008EA8E8 , 32'hFFFDE450 , 32'h0039D54F , 32'hF129CA80 , 32'h063CE0C8 , 32'hFFFFF9ED , 32'hFE064F54 , 32'h00036BCB , 32'h0000D1F8 , 32'h00E58BFC , 32'hFDE2A760 , 32'hFB6A1450 , 32'h0BC3AEE0 , 32'hFFFF6D0E , 32'h0EA3B730 , 32'hFFFFECDE , 32'hEB1B82C0 , 32'h014A89F4 , 32'hFFFE4E3D , 32'h04B3DF20 , 32'hF8226FD8 , 32'h11910E20 , 32'hFFFE779F , 32'h000059E3 , 32'hFFFF027E , 32'hF501B9B0 , 32'h00FC28EA , 32'h0000B2C5 , 32'h11B600C0 , 32'hFEFD73D4 , 32'hFFFEB41E , 32'hF5CB3C70 , 32'hFFC15D72 , 32'h00001B72 , 32'hF8079148 , 32'h1C308920 , 32'h04B83D10 , 32'h00000BB2 , 32'h00032666 , 32'hEE577300 , 32'h000157FD , 32'h00770BCD , 32'hFFFF2076 , 32'h00AC0CBD , 32'h007752B9 , 32'h00039B4C , 32'h000299D2 , 32'hFFFF66B1 , 32'h00020E9C , 32'h01FA00D8 , 32'hFB9627B0 , 32'h00005381 , 32'hFB4B71C0 , 32'h01BE2C48 , 32'h034BC4C0 , 32'h00003B17 , 32'h00CB9465 , 32'h00004CC1 , 32'hF6E80850 , 32'h064359B8 , 32'hFFFFAAEA , 32'h0C2E05A0 , 32'hFFFF6675 , 32'hFFFEC08D , 32'hFB3AEE60 , 32'hFFFA1F25 , 32'hFE34261C , 32'hFFFF4E15 , 32'hFD32EF6C , 32'h0000D1CF , 32'h00017AAA , 32'h00A539C0 , 32'h0001FC22 , 32'hFFFBF112 , 32'hED2FED20 , 32'hF4987180 , 32'hFFFF1590 , 32'h00030BB2 , 32'h0002EB4E , 32'hFFFE7665 , 32'hFFFF2051 , 32'hF45CD7B0 , 32'hFB655608 , 32'hFFFF2819 , 32'hFFFEA3F0 , 32'h02E034D8 , 32'hFCF28124 , 32'h0000912B , 32'h0002557D , 32'hFC940658 , 32'h0000578B , 32'h00016988 , 32'hF975DEF8 , 32'hFFAEFBD3 , 32'h00BC28AD , 32'h008FF6DB , 32'h00002AB0 , 32'hFFFF17C6 , 32'h02F9B678 , 32'hFFFF807C , 32'h0001DEE9 , 32'hFE7F7FB8 , 32'h0000DA8A , 32'h0002B459 , 32'h038F3F04 , 32'h000058C7 , 32'hEDEF02A0 , 32'hFEAF49D4 , 32'h0001200B , 32'hFFFF6CA7 , 32'hFFFF38C2 , 32'h09347D50 , 32'h01153778 , 32'hF757CCD0 , 32'h0BAC12A0 , 32'hFFFFE86E , 32'hEA0C5DC0 , 32'h000082B3 , 32'hFFFFFA6D , 32'hF0B1FF70 , 32'h02C1468C , 32'h03FD0720 , 32'hFFFF69D6 , 32'h1BA4CFA0 , 32'h01C663EC , 32'hFE2BF388 , 32'hE7E52EE0 , 32'h1D0D4720 , 32'h03EBEA5C , 32'hFDF3A6D0 , 32'hFCDABF60 , 32'hFFFF4C27 , 32'h000009D2 , 32'h000146AB , 32'hFE756798 , 32'hF35FD6C0 , 32'hFFEF7819 , 32'hFD944CD4 , 32'hFF3778CB , 32'h00F7129F , 32'hFFFFFDFF , 32'h04F473D0 , 32'hFF60C6AB , 32'h00009660 , 32'hEFC88840 , 32'hFFFD18E2 , 32'h0632C790 , 32'h0AFE1C80 , 32'hFFFF1EB7 , 32'h000105B8 , 32'hFFFFB2BB , 32'h0002F84F , 32'hFFFFB7B9 , 32'hFFFE1D13 , 32'hFE9E98F8 , 32'hFCAB5EE0 , 32'h058368E8 , 32'h03358D20 , 32'h01A39608 , 32'h0E126770 , 32'h00019BBD , 32'h0000EFD8 , 32'hFFFEA7A9 , 32'h00002C95 , 32'hFFFDCED5 , 32'h05ACAED8 , 32'h13749600 , 32'h01D53ED8 , 32'h00001373 , 32'h00004A4D , 32'hFFFE6C72 , 32'hFFFF0C1C , 32'h05E90270 , 32'h061DBD80 , 32'hFFFC761D , 32'hFFFDFC72 , 32'hFFFF4942 , 32'hECA42440 , 32'h1D371D60 , 32'h0415AF90 , 32'hFFFE577F , 32'h000197EC , 32'hFFFEAD12 , 32'hFE52F7DC , 32'h015081FC , 32'hFE683E78 , 32'h00010C81 , 32'hFFB82625 , 32'h00029C35 , 32'hE95DBD00 , 32'h00049CEA , 32'h07C44E10 , 32'h00017D51 , 32'h0CC19020 , 32'h02AD3DA0 , 32'h095905A0 , 32'h067A5070 , 32'hFFFF9D24 , 32'hFFC67C06 , 32'hFE097884 , 32'hFFFDAF68 , 32'hFBBECED8 , 32'h00009A99 , 32'h03ABC1B8 , 32'h0B331F00 , 32'hF6B5DDF0 , 32'h00010263 , 32'hFFFEC6BC , 32'h01EECDFC , 32'h00001A39 , 32'h09C23A20 , 32'h000283EC , 32'h01740288 , 32'hFFFDD2F4 , 32'h012594A4 , 32'hFFFDADC3 , 32'hFFFDB7A2 , 32'hFFFEF173 , 32'h00CD2938 , 32'hF2AE64E0 , 32'h0001B596 , 32'hFFFF5620 , 32'h00007876 , 32'h000146D9 , 32'h0E2CB0B0 , 32'hF7EE8ED0 , 32'hF271C940 , 32'h03E45EA0 , 32'h07FBA7D8 , 32'hFFFFC13B , 32'h00008C02 , 32'hFFFFF742 , 32'h00F0A586 , 32'hFFFF87C0 , 32'h00023D40 , 32'h064EA228 , 32'hF58D1500 , 32'h0000CA91 , 32'hF8B36AD0 , 32'hFFC0DA47 , 32'hFE4D94CC , 32'hED4CC240 , 32'hFFFF97D0 , 32'hFD1479B0 , 32'h098E2F80 , 32'h00A57160 , 32'h00018B01 , 32'h07F47A08 , 32'h101F4A60 , 32'h02A786B0} , 
{32'h02B2B1A8 , 32'h18538140 , 32'h000114CD , 32'hF8C56110 , 32'h0001B0CD , 32'h01A2D884 , 32'hFFFB1D58 , 32'hFFFF3F30 , 32'h000057C2 , 32'hFFFBAB33 , 32'h03FC0638 , 32'h0BE864B0 , 32'h04446990 , 32'hFFFF889D , 32'hFFFE8298 , 32'hFA43F120 , 32'hFFFE420C , 32'hFA5BAE30 , 32'hFA6384A8 , 32'hFFFF267B , 32'h0001D2B4 , 32'h03091494 , 32'h0B904D40 , 32'h021AE018 , 32'hFB1E9F70 , 32'h00029003 , 32'h048739A8 , 32'hFEF01CC4 , 32'h0002821A , 32'hF41B40E0 , 32'h000171C7 , 32'h06F689D8 , 32'h00013C98 , 32'hFFFE1158 , 32'hFFFEF66A , 32'hEB8ED500 , 32'hFC6E8EB4 , 32'hF810DAE0 , 32'h0000B084 , 32'h02034A14 , 32'h161CAC80 , 32'h0001C7BD , 32'hFFFF6ACC , 32'h01F4AB74 , 32'h01729BA8 , 32'hEF77DE40 , 32'h11085E20 , 32'h0002C667 , 32'h0BE6B2A0 , 32'h02520A5C , 32'hFF3D1A7E , 32'h0002DFC3 , 32'hFA267228 , 32'h0D2D8550 , 32'hFB560598 , 32'h00017E00 , 32'h02CE0358 , 32'h00022A6F , 32'h000079DC , 32'h05E37018 , 32'h014FB85C , 32'h013C6E60 , 32'hFD53343C , 32'hFFFFD029 , 32'hFF75A275 , 32'hFFFEC53C , 32'h19901920 , 32'h0209FA74 , 32'hFFFF43B5 , 32'hFCAC5DEC , 32'hFB1721B8 , 32'hF1786F90 , 32'hFFFEED04 , 32'hFFFF8D4A , 32'hFFFFE6F6 , 32'h03ADF138 , 32'hFF07D3B6 , 32'hFFFFC67B , 32'h0A352090 , 32'hFDF60698 , 32'h0000E115 , 32'h16D049A0 , 32'hF8E1B6F8 , 32'h00013664 , 32'h040DE5A0 , 32'hF05C56B0 , 32'h0457BA88 , 32'h00000DD8 , 32'hFFFD4BFF , 32'h16B14920 , 32'h000183BF , 32'h08081340 , 32'hFFFF5DFB , 32'hF7E02CD0 , 32'h01099F28 , 32'hFFFE6311 , 32'hFFFFB9AF , 32'h00009642 , 32'hFFFF66DA , 32'hF72F94D0 , 32'h03D377F0 , 32'h000053F9 , 32'h102E4380 , 32'h0ACD61F0 , 32'h0363C808 , 32'h00006A22 , 32'hFF8875D4 , 32'h00006038 , 32'hFFF017FD , 32'h0C1DC230 , 32'h000122E8 , 32'hF9D53B78 , 32'h00031D7A , 32'hFFFF6AF0 , 32'hFF0E1672 , 32'h05E04800 , 32'hFEAFAF58 , 32'hFFFFEBB1 , 32'hF6CFFF40 , 32'hFFFF4E0B , 32'hFFFF048B , 32'hFBDAF410 , 32'hFFFE99FD , 32'h00023C31 , 32'hF5D09C30 , 32'h0CA70820 , 32'hFFFEFF3A , 32'hFFFED4B8 , 32'hFFFE76CB , 32'h000171C5 , 32'h000139B9 , 32'h0052C037 , 32'hFFEAC666 , 32'h0000C8F9 , 32'h00006E4D , 32'h0B1E1550 , 32'hFEEAA840 , 32'hFFFE10C4 , 32'hFFFF6EFA , 32'h01C06274 , 32'h0001095B , 32'h0000B61B , 32'h01C0C540 , 32'h0401CFB8 , 32'h02056EA0 , 32'h02422740 , 32'hFFFE77D0 , 32'hFFFFC937 , 32'hFB6F6FB8 , 32'h0001F77C , 32'hFFFDB3AE , 32'h009AE8CC , 32'h0000722B , 32'hFFFB96F0 , 32'hFE6AA76C , 32'hFFFF33C8 , 32'hFE8EEBEC , 32'h00CB8150 , 32'hFFFE1F04 , 32'h00013D61 , 32'h00006ACE , 32'hFDCD19B0 , 32'hF5A89BB0 , 32'hFFF2FAFE , 32'h088881C0 , 32'h00002369 , 32'hF722E8E0 , 32'hFFFE6267 , 32'h0000E1F2 , 32'h07EF9BB0 , 32'hFDBB5B38 , 32'h00DC4B44 , 32'hFFFF2FBA , 32'h0B1BB520 , 32'h02949328 , 32'h03A101E4 , 32'hF94B07C8 , 32'hFB1C2850 , 32'h004675A4 , 32'hFDC3FE30 , 32'hF82A4AA8 , 32'h000028B7 , 32'hFFFDCB92 , 32'hFFFD79F8 , 32'h035DFAFC , 32'hF0DEBD20 , 32'hFF08339C , 32'hFF731721 , 32'hFCFE1B24 , 32'h017B7E08 , 32'h00003402 , 32'h007D796A , 32'h178BA4A0 , 32'h00001CB8 , 32'h05536170 , 32'hFFFF9567 , 32'h01D6DE58 , 32'h01405D50 , 32'hFFFE29D8 , 32'h00028866 , 32'hFFFCA1B5 , 32'hFFFF5BD6 , 32'h00003176 , 32'h0001C814 , 32'h0250B4A8 , 32'hFBC4EC10 , 32'hF54371A0 , 32'hF76A8BE0 , 32'hF95A90B8 , 32'hFD14CF60 , 32'hFFFE21C3 , 32'h000003C9 , 32'h0000B8C0 , 32'hFFFDC946 , 32'h0000D872 , 32'hFC528F14 , 32'hF56C3B00 , 32'hFB757500 , 32'h0000D758 , 32'h0002B745 , 32'h0000E1F0 , 32'h00000469 , 32'h00F1C678 , 32'hFA825868 , 32'h0000B027 , 32'hFFFE0677 , 32'hFFFF40CB , 32'hF5FBCB20 , 32'h272CA240 , 32'h04AAA3E8 , 32'hFFFE5405 , 32'hFFFF7889 , 32'h00013A2F , 32'h02056E98 , 32'h066D3BD0 , 32'h2E481FC0 , 32'h0001DD80 , 32'hFFFA7219 , 32'hFFFECF53 , 32'h034AE560 , 32'hFFFFC79A , 32'hEB1B2060 , 32'hFFFF6412 , 32'h0EF76200 , 32'hF2866590 , 32'h095A0340 , 32'h1C5E4160 , 32'h0002E10B , 32'h0A0FC270 , 32'hFF8148D8 , 32'h00002108 , 32'hFB8E7780 , 32'hFFFF3266 , 32'h0117A544 , 32'h019D214C , 32'h0087F653 , 32'hFFFF1460 , 32'hFFFEE569 , 32'hFECA7F6C , 32'h000097E4 , 32'h00CD2CCE , 32'h0000B829 , 32'hFF2B45E6 , 32'h0001E465 , 32'h051019C0 , 32'hFFFE7202 , 32'h000020E6 , 32'hFFFFCA87 , 32'hFE937A3C , 32'hF86C3370 , 32'h00012BA1 , 32'hFFFF95F4 , 32'h00009CBC , 32'hFFFEAC6D , 32'hF057D680 , 32'h08369EA0 , 32'hFE1BFE48 , 32'hF1CF1470 , 32'hFC7F8404 , 32'hFFFF949C , 32'hFFFF3A7D , 32'h0001C86A , 32'hFFD2C059 , 32'hFFFF0F37 , 32'h0001B205 , 32'hF75A3EE0 , 32'hFBF81960 , 32'hFFFED99A , 32'hF9C405B0 , 32'hFF8735E7 , 32'h01FB84AC , 32'hF0705A60 , 32'hFFFF092A , 32'h074C4458 , 32'h108D52A0 , 32'h03AC5554 , 32'h000285FB , 32'hF52A1880 , 32'hF03FEA70 , 32'h01FD1FD8} , 
{32'hFA52BAB0 , 32'hFB864388 , 32'hFFFFA61B , 32'h0B6A6960 , 32'hFFFF46D7 , 32'hFFA50854 , 32'hFFFE69BE , 32'hFFFECD00 , 32'h0000D07D , 32'hFFFEF0B3 , 32'hF0BC2930 , 32'h0B792610 , 32'h01D62D64 , 32'hFFFFBE9C , 32'hFFFD43C2 , 32'hF42E0330 , 32'h00007B1A , 32'h12078560 , 32'h00600A13 , 32'h00004559 , 32'hFFFE815A , 32'h00C8161F , 32'h00BAC438 , 32'hF9853008 , 32'hFF3371D3 , 32'h0001A30E , 32'h00F50560 , 32'hFC901CF0 , 32'hFFFE6765 , 32'hFFBB0556 , 32'hFFFED108 , 32'h00B7528C , 32'h00030185 , 32'h0000DE9D , 32'hFFFF5471 , 32'h0954FD00 , 32'hEAC5A5E0 , 32'hFF089D62 , 32'h000188C4 , 32'hF0710E90 , 32'hFA48F928 , 32'hFFFFAAA9 , 32'hFFFFFF19 , 32'h03927C00 , 32'hF606F140 , 32'hFEB043A0 , 32'h08482290 , 32'hFFFF0022 , 32'h0857E430 , 32'h06396AA0 , 32'hFF72D977 , 32'h00012167 , 32'hFF546CB7 , 32'h1548CC60 , 32'h059B3FD8 , 32'h00028583 , 32'h037EE718 , 32'h00000C2E , 32'h0000336D , 32'h038F27F4 , 32'hFCB06D74 , 32'h02E14B84 , 32'hE1693EE0 , 32'hFFFEDB2B , 32'h05B2C188 , 32'h00026E56 , 32'h033C90AC , 32'h0492CFE0 , 32'hFFFE432C , 32'h078529C0 , 32'h082DCE30 , 32'hF3BA4FB0 , 32'h0002B111 , 32'h0001F9AE , 32'h00028A44 , 32'h0563EB40 , 32'hF8EA07E0 , 32'h0000B194 , 32'hF7F63DD0 , 32'hFF89F365 , 32'hFFFE8583 , 32'hF991EC08 , 32'h00AEE06B , 32'h000073E8 , 32'hFD5FA780 , 32'hF7FE8640 , 32'hFF613014 , 32'hFFFDD2CE , 32'hFFFFC897 , 32'h18FF6880 , 32'h00025967 , 32'hFF89F9AD , 32'hFFFFD1B4 , 32'hFF664EFA , 32'h00ABB059 , 32'h000406C0 , 32'hFFFFDE18 , 32'h00002BC0 , 32'hFFFE7895 , 32'hFD724C48 , 32'hFC083ED4 , 32'h00009E53 , 32'hEF3B5AC0 , 32'h13CB7880 , 32'hFC0C2D14 , 32'h00021194 , 32'hFFB2D0A3 , 32'h0000A3C0 , 32'hF62AAB20 , 32'h0710B2A8 , 32'hFFFE217A , 32'hFA421598 , 32'h00013A9C , 32'hFFFF7441 , 32'hF4AB1E00 , 32'h08DA2B20 , 32'h00058BDD , 32'h0001091F , 32'h00C14AFA , 32'hFFFE8593 , 32'hFFFEBF46 , 32'h086DBC80 , 32'h00023E1A , 32'h00005354 , 32'hF3154610 , 32'hF6A29230 , 32'hFFFDE557 , 32'h000254A4 , 32'h0001E37F , 32'hFFFF1673 , 32'h00001FC6 , 32'hFB5BAEE8 , 32'h09CA9A20 , 32'hFFFF4529 , 32'hFFFC68DE , 32'hF6BDD230 , 32'hF2FD4140 , 32'h000266BF , 32'hFFFFCAFC , 32'h04E47AF0 , 32'hFFFFC3C8 , 32'hFFFF0902 , 32'h021E1D10 , 32'hF9EC7538 , 32'h03EC0FC0 , 32'h047C3318 , 32'hFFFC8033 , 32'hFFFEB493 , 32'hFC7B7F0C , 32'h00010B92 , 32'hFFFAF7A3 , 32'hFAAB6F90 , 32'hFFFF219F , 32'hFFFDB2FF , 32'hFF1BF116 , 32'hFFFFC5AA , 32'hFAC59AD8 , 32'hFFD5DBCF , 32'h0002E415 , 32'hFFFDB30D , 32'h0002451A , 32'hF98C5FF0 , 32'hFFF348C4 , 32'hFCBF2F9C , 32'hF8BA4D40 , 32'h0000B3CC , 32'h181537C0 , 32'h0000105B , 32'hFFFF1D93 , 32'h07E51AB8 , 32'h01994148 , 32'hFC5019E0 , 32'hFFFF5DD6 , 32'h19308C00 , 32'hFD20232C , 32'hFC3D9E2C , 32'h053639A8 , 32'h0C0C9E40 , 32'h267B5780 , 32'hFF8C9BDC , 32'h103AACA0 , 32'hFFFFEFE4 , 32'hFFFE6C2D , 32'hFFFFBC83 , 32'hFEEBBF98 , 32'h086D9310 , 32'h02FD5EA0 , 32'h00B247DA , 32'h0E3A8480 , 32'h05142C60 , 32'hFFFF160D , 32'h070E8A20 , 32'hFF9EC79D , 32'hFFFEA37F , 32'hFB29F040 , 32'hFFFFCC14 , 32'h02E12BCC , 32'h106A2920 , 32'h0000EA80 , 32'hFFFF15CE , 32'hFFFEF031 , 32'hFFFE82B2 , 32'hFFFF2061 , 32'h00017273 , 32'hFEEC1EE0 , 32'hF3FD3140 , 32'hED2D8DC0 , 32'h00BB057A , 32'hF9D31690 , 32'h0D273D00 , 32'hFFFEF072 , 32'h0000AE39 , 32'h00006688 , 32'h0001D4F1 , 32'h0002691D , 32'hFD5A056C , 32'hFD72A868 , 32'h07653C10 , 32'h00008F55 , 32'h0001A462 , 32'hFFFF2890 , 32'hFFFF1599 , 32'hF325F260 , 32'hF3DCDF70 , 32'hFFFFE474 , 32'hFFFF3D42 , 32'hFFFE2B05 , 32'hF027EA90 , 32'h17D44F20 , 32'hFE28B57C , 32'h0000A864 , 32'h0000D51A , 32'h00000BD4 , 32'hFBD69AB0 , 32'h04557258 , 32'hEE2E5C40 , 32'hFFFE0BA9 , 32'h014021FC , 32'hFFFD5E7C , 32'h007FD027 , 32'h000140D2 , 32'hFDDC5764 , 32'h0001799E , 32'h00169F8D , 32'hFB48EEB8 , 32'hFEB4DE14 , 32'hE7B47B20 , 32'hFFFEB5D2 , 32'h0249E8C8 , 32'hFF85FDBB , 32'hFFFE6D33 , 32'h00FCBAD0 , 32'hFFFCE002 , 32'h0320C2E0 , 32'h10AA72E0 , 32'h07361260 , 32'h0001B034 , 32'h00019720 , 32'h04562790 , 32'hFFFF48E4 , 32'hF2367270 , 32'h00021E70 , 32'h00221DB3 , 32'hFFFEF193 , 32'hFAE6C518 , 32'h000020EB , 32'h0000CE5E , 32'hFFFFD2AC , 32'h058354F0 , 32'h141FBDE0 , 32'h0001B06A , 32'h0002D4EC , 32'h0000BD11 , 32'hFFFEE8F8 , 32'h07AD5C60 , 32'h05398930 , 32'hE7AD6700 , 32'h01387B6C , 32'h07AC5EE0 , 32'h0000A8CB , 32'hFFFCD33E , 32'h00023D32 , 32'h01D48F80 , 32'h00001AFE , 32'h0001DF22 , 32'h01BAADA4 , 32'h050F5190 , 32'hFFFC1008 , 32'hF909DC30 , 32'h011B6614 , 32'hF7E639E0 , 32'h0A79CD40 , 32'hFFFF30DD , 32'h05BE70D0 , 32'hF42E2210 , 32'h01E5892C , 32'h0003A8DF , 32'h12BC0B00 , 32'hF5FE25D0 , 32'hFA8E6EA0} , 
{32'h0B0664E0 , 32'hE9C2D460 , 32'h00018550 , 32'hFAEB2F30 , 32'h000115C3 , 32'h07A42B50 , 32'hFFFD623E , 32'hFFFF5CF4 , 32'hFFFFDE5D , 32'h00006911 , 32'h049FF378 , 32'h0965EA60 , 32'h025DDED0 , 32'hFFFDFA60 , 32'hFFFB8752 , 32'hF311FDF0 , 32'h00043579 , 32'h0BAF75E0 , 32'hFAE2A170 , 32'hFFFF3491 , 32'h00004F7A , 32'hFE3BA660 , 32'h054475C0 , 32'hF27D24F0 , 32'h0110AF2C , 32'hFFFDFBFA , 32'h039E3CE8 , 32'hFEB66278 , 32'h00010EA8 , 32'h0D114E60 , 32'h00011CA3 , 32'h031E7A8C , 32'hFFFFE841 , 32'hFFFF47EC , 32'hFFFEC1F4 , 32'h006B907D , 32'h0BB798A0 , 32'hF5D413A0 , 32'hFFFDFE41 , 32'h059A1018 , 32'hF8886E68 , 32'hFFFF8277 , 32'hFFFD590C , 32'hFE2008CC , 32'h08BC3730 , 32'h005341FA , 32'h03733E88 , 32'h00025928 , 32'hED27C600 , 32'hF81B43A0 , 32'h01206724 , 32'hFFFCEFE7 , 32'h04E1ACC8 , 32'hF64C2590 , 32'hF73A42E0 , 32'hFFFFC99F , 32'h002BECDE , 32'hFFFFB1A0 , 32'hFFFE4531 , 32'hFC029B90 , 32'h005CB471 , 32'hF37EEFA0 , 32'hFB8CB9F8 , 32'hFFFFC509 , 32'hE0E3F9A0 , 32'h0002BC9F , 32'hF3A8ACD0 , 32'h00CE24D5 , 32'hFFFDF2A8 , 32'h100F8A20 , 32'h0120CCC8 , 32'h02B6B4C0 , 32'h0000132C , 32'h0000D734 , 32'h0000B46C , 32'h053D0250 , 32'h04F41908 , 32'hFFFC777B , 32'hEF9C9940 , 32'h020CF4B4 , 32'hFFFEA219 , 32'h22E8B980 , 32'h055F68C8 , 32'h00005C3B , 32'hFCCA0B58 , 32'hF2A5CC80 , 32'hFDF9A1F8 , 32'h00043D8C , 32'h0000B6C7 , 32'hE3EF86E0 , 32'h00005DEF , 32'hFEFBDCA4 , 32'h00001E6C , 32'hFF17FA87 , 32'h005B0D22 , 32'hFFFE1518 , 32'h00002F3A , 32'h00002CE9 , 32'hFFFF9120 , 32'hF9DD3FE0 , 32'hFAB7E110 , 32'hFFFF9B6F , 32'hF62A4670 , 32'h0BBB1F90 , 32'h035C6704 , 32'hFFFF019A , 32'hFFC89CDD , 32'hFFFF569C , 32'h05858E00 , 32'h008EFAFA , 32'hFFFF79B1 , 32'hEF037700 , 32'h00001F84 , 32'hFFFF4796 , 32'h030B8C68 , 32'hFBAF55E8 , 32'h00ED9AE2 , 32'h0000ABC1 , 32'hFF3716FB , 32'h000060D2 , 32'h00026F95 , 32'h00F20DFA , 32'hFFFF7E54 , 32'h0002AF98 , 32'hED284300 , 32'h0436D8C0 , 32'hFFFE8A65 , 32'hFFFC1F7E , 32'h0001A290 , 32'h00004801 , 32'h0001460B , 32'h03DEC33C , 32'h0BC53760 , 32'hFFFDE4A7 , 32'hFFFD4F8B , 32'hF7ABE820 , 32'hF9196898 , 32'hFFFF3C1D , 32'h00008F17 , 32'hFE0DD484 , 32'h000151E2 , 32'h0000C807 , 32'h0596B4E8 , 32'h07779E78 , 32'hFCFEDFA0 , 32'h00AE9C8E , 32'hFFFEA1AC , 32'hFFFD80E0 , 32'hFBB97CB8 , 32'h00009E1B , 32'h00012BBA , 32'h036A6280 , 32'hFFFFDC3E , 32'hFFFFCEF2 , 32'h0074AECF , 32'h0000AFD6 , 32'hF97F5008 , 32'h01713D80 , 32'hFFFCD211 , 32'h00012730 , 32'hFFFED718 , 32'h05D8A9D0 , 32'h06FD26A8 , 32'h03BABD20 , 32'h10658160 , 32'hFFFE726D , 32'hFA85E080 , 32'h00007489 , 32'h00013C36 , 32'hFFCB33C1 , 32'h00395B82 , 32'hF6F50940 , 32'hFFFE4859 , 32'h0D841A20 , 32'hFCFB82E8 , 32'h02D6A6E8 , 32'hF12EAD70 , 32'hEB93F460 , 32'h22B46C80 , 32'hFFE34715 , 32'h0605D608 , 32'hFFFEBDC0 , 32'h00012C93 , 32'hFFFF48E8 , 32'hFE394818 , 32'hF3C03A40 , 32'hFAED8960 , 32'h00B035B6 , 32'hF5E5D900 , 32'h010F5BB8 , 32'h00010CDB , 32'h06EF6EA0 , 32'h0B174A80 , 32'h0000DED4 , 32'h00549BB9 , 32'h0001D6DE , 32'h00486079 , 32'hF5B82490 , 32'hFFFF472C , 32'h00029D53 , 32'hFFFF3EE1 , 32'hFFFFFD9E , 32'hFFFDDC22 , 32'h0001B6A8 , 32'h02AC4F40 , 32'h088A3FC0 , 32'h0C0A74B0 , 32'h044DB110 , 32'hFFC1B82D , 32'h0606DAD0 , 32'h00017076 , 32'h000015C9 , 32'h0000C2D7 , 32'hFFFFBD6C , 32'h0000782D , 32'hF9718DB0 , 32'h08177200 , 32'hF631CC80 , 32'h0002979C , 32'h000072CC , 32'hFFFE0742 , 32'hFFFEA259 , 32'hFB3189C8 , 32'hF5B2D240 , 32'hFFFFE711 , 32'h0000001A , 32'hFFFDB301 , 32'h0C129770 , 32'hFBCBD8E0 , 32'h0068E469 , 32'hFFFE9F06 , 32'hFFFC59A2 , 32'hFFFF6CBC , 32'h01DF8AD4 , 32'h0080D471 , 32'h117EF3E0 , 32'hFFFE0501 , 32'h004833E2 , 32'hFFFF54FB , 32'hF4404CD0 , 32'h00008E25 , 32'h0D29AFC0 , 32'h0001D80F , 32'h09D47570 , 32'hF7C59C60 , 32'hF4A32020 , 32'hFEE1DA0C , 32'h00000F94 , 32'hFA501838 , 32'h006603FD , 32'h0000EF21 , 32'h017DC8E8 , 32'hFFFF0CDB , 32'hFF2A152F , 32'hFD387E58 , 32'hF35D2EA0 , 32'hFFFFD9C2 , 32'hFFFC85E9 , 32'h0EB13420 , 32'h00015DF0 , 32'h02B24B24 , 32'hFFFFBA0D , 32'hFEECC1A0 , 32'h000170A4 , 32'hFC125648 , 32'hFFFD8FA1 , 32'hFFFC5783 , 32'h00018373 , 32'hF3332550 , 32'hFCB87AE8 , 32'h000140D8 , 32'hFFFF0B8F , 32'hFFFE5FBA , 32'hFFFFD669 , 32'hFEB5BB80 , 32'hF6965F70 , 32'h03A7AD8C , 32'h1FB79D80 , 32'hF9E68650 , 32'h0000F26E , 32'hFFFE8AC7 , 32'hFFFE1A82 , 32'hFC3770E8 , 32'hFFFF1941 , 32'h000017EE , 32'h056F9138 , 32'hF3B92010 , 32'hFFFFBD2D , 32'hE421FA40 , 32'hFCF9DA68 , 32'h02CF7578 , 32'h0ACC9C20 , 32'h0001E1F9 , 32'hFC8E7E1C , 32'h0062F86E , 32'h02A067A4 , 32'h0001B28C , 32'h025B4AA4 , 32'hEC7E7A80 , 32'hF5F74FD0} , 
{32'h1CE285A0 , 32'hFA59A3D0 , 32'h00004C27 , 32'h04357660 , 32'h0001CDCF , 32'h05686AC0 , 32'h000035A3 , 32'hFFFFE69D , 32'hFFFFF2AB , 32'h0001086A , 32'h01288E64 , 32'hFB13A338 , 32'hF21E29A0 , 32'hFFFF347D , 32'hFFFF5112 , 32'hFEE904A4 , 32'hFFFFFE43 , 32'hF87A5148 , 32'hFD5CA768 , 32'hFFFE752F , 32'h00022640 , 32'h005D4A33 , 32'hF8307C90 , 32'h0AA9C060 , 32'hFE252134 , 32'hFFFE5F9E , 32'h0341627C , 32'h023DF8C4 , 32'h00010C63 , 32'hFD888D30 , 32'h00007609 , 32'h0911B0B0 , 32'h00008923 , 32'hFFFD5BB8 , 32'hFFFD5242 , 32'h0A493460 , 32'hFD90BEB4 , 32'hFA75C4C8 , 32'hFFFF6E75 , 32'hEC628D40 , 32'hF2F97B70 , 32'h0001CD50 , 32'hFFFFAF3A , 32'hFEB123AC , 32'hF4A03260 , 32'h00B42A28 , 32'h06BBD7E8 , 32'hFFFD1B4C , 32'h003D29BC , 32'h09DA3700 , 32'hFF4C55E2 , 32'hFFFF420E , 32'h00031C2A , 32'h0187971C , 32'h07DB5510 , 32'hFFFF13B9 , 32'h00880140 , 32'hFFFE55F8 , 32'h0001FEBE , 32'hFE483008 , 32'hFF3466AA , 32'hFE7687D8 , 32'h11D97C60 , 32'hFFFFAD96 , 32'hFC77AF78 , 32'h0000FF76 , 32'h0D36AFA0 , 32'h02D81B00 , 32'h000227A5 , 32'h0C15C9A0 , 32'hFB690720 , 32'h10067800 , 32'h00001C5A , 32'hFFFEB409 , 32'h0000E084 , 32'h10743B80 , 32'h07ED3F30 , 32'hFFFFB8FF , 32'hE960C8C0 , 32'h0273D474 , 32'hFFFF4917 , 32'hF4F9F4C0 , 32'h062A45E8 , 32'h000086D9 , 32'h079C42B0 , 32'hF741A9F0 , 32'hFFEC1FEC , 32'hFFFD1DF7 , 32'h0000A0BC , 32'hF2FC8CB0 , 32'h0001558B , 32'h099D7EB0 , 32'h0000C8B4 , 32'hFB9D8778 , 32'h006CDF66 , 32'h0001A5C6 , 32'h0001DB53 , 32'hFFFCFDF1 , 32'hFFFE7E3D , 32'hFA9EFCA8 , 32'hFEA56D54 , 32'h000053FA , 32'h05599D90 , 32'hFBC43C08 , 32'h04135560 , 32'hFFFF4E53 , 32'hFFD7D367 , 32'h00008E08 , 32'h02801D18 , 32'h157F75A0 , 32'h0000D440 , 32'hFBE34018 , 32'h0000444B , 32'h0002497F , 32'hF9187808 , 32'h03231884 , 32'hFEFE3190 , 32'hFFFF8F24 , 32'hF5601510 , 32'hFFFFADE7 , 32'hFFFF2DAE , 32'hFD10AAA0 , 32'h00016396 , 32'hFFFE7872 , 32'h1C74B4A0 , 32'hF744E610 , 32'hFFFF1F93 , 32'h00018D1D , 32'h000057A8 , 32'hFFFDF230 , 32'h000108ED , 32'hFD3AC260 , 32'hFD6E2054 , 32'hFFFF2CF4 , 32'hFFFF3FEE , 32'h06B4E338 , 32'hEF662F40 , 32'hFFFF394B , 32'h0000BB62 , 32'hF94DF8F8 , 32'h0000CA03 , 32'hFFFFC961 , 32'hFE375E40 , 32'h00E3E82D , 32'h01C9EEF0 , 32'h02892A90 , 32'h00020DBE , 32'hFFFDC32C , 32'hFCD629F4 , 32'hFFFF84B8 , 32'h00004A2A , 32'h03248C84 , 32'hFFFEDA88 , 32'h0001C4EA , 32'h00771649 , 32'h0000D43C , 32'hFE7B56F4 , 32'h00AD62F3 , 32'h0000B4DC , 32'hFFFFC59A , 32'hFFFE3D94 , 32'h178409E0 , 32'h05E65AA8 , 32'hFF5ADD2E , 32'h05D1DAB0 , 32'h00008A64 , 32'h0753BA88 , 32'h00002573 , 32'hFFFC25CE , 32'hFF972C53 , 32'hFA837590 , 32'h032A60AC , 32'hFFFF5489 , 32'h1958B740 , 32'h00B984B7 , 32'h0776D238 , 32'h07ACAAF8 , 32'h0364B9DC , 32'hF094EBF0 , 32'hFEC97928 , 32'h03A83A10 , 32'h0001888D , 32'h0001C997 , 32'h0000A7B1 , 32'hF7AEDC80 , 32'hFCC451D8 , 32'h01A37998 , 32'hFFBFBD1A , 32'hF3D7A990 , 32'hFFA09EB1 , 32'hFFFFEBC5 , 32'hF2A9B230 , 32'h0B38FAE0 , 32'h0000F9BE , 32'hFA4DFB40 , 32'hFFFC99CA , 32'hFDC655F0 , 32'hFAA9DC18 , 32'hFFFDA539 , 32'hFFFF9F9F , 32'hFFFDDBFD , 32'h0001726E , 32'hFFFCFD43 , 32'hFFFE5D49 , 32'h0549BE70 , 32'hF19A2A60 , 32'hF884E178 , 32'hFCF04EA0 , 32'h055F98D0 , 32'hF79B6C70 , 32'hFFFFCD31 , 32'hFFFC8697 , 32'h00000C0F , 32'h00003F4C , 32'h0003008C , 32'hFE75D620 , 32'h1208E520 , 32'h0BEBE890 , 32'h0000F30C , 32'h000067AF , 32'hFFFE879D , 32'h0000817B , 32'h0A32D960 , 32'hF2E7F940 , 32'hFFFF2860 , 32'h00022B68 , 32'h0001823D , 32'h054394F0 , 32'hFBA3F068 , 32'hF6345760 , 32'hFFFF47B8 , 32'h00023B41 , 32'hFFFF4073 , 32'hFA317B28 , 32'h03A27B10 , 32'h06A86500 , 32'h0002A815 , 32'h00CEE22A , 32'h00019F8F , 32'hF7436640 , 32'h00003608 , 32'h030B87D4 , 32'hFFFFF329 , 32'hDF63EF80 , 32'hF9CE1E90 , 32'h04A33938 , 32'h08B8BC90 , 32'hFFFFD456 , 32'hFF275528 , 32'hFFB0C5AC , 32'h0000BF14 , 32'hFA042830 , 32'hFFFE6128 , 32'h04FFC148 , 32'h2A34CD80 , 32'h08838D80 , 32'h000066E6 , 32'h00027D0A , 32'hFAEF69C8 , 32'h00000D64 , 32'hFA2C10F8 , 32'hFFFFEDAB , 32'hFFEAB427 , 32'h00046924 , 32'h07A81F68 , 32'hFFFF5CD1 , 32'hFFFECA3E , 32'hFFFEE6A0 , 32'hE81C7D00 , 32'hF7BAF530 , 32'h000035CF , 32'hFFFF7237 , 32'h0001DF7A , 32'h00009002 , 32'hFA406480 , 32'hFE487698 , 32'hF22C5720 , 32'h07941E08 , 32'h18738F00 , 32'h00003DE3 , 32'hFFFE2C48 , 32'h00013CA4 , 32'h019CC804 , 32'hFFFF835B , 32'h00010ECE , 32'hFC9E7CD4 , 32'hFD284500 , 32'h00001AC5 , 32'h014B248C , 32'hFE572198 , 32'h01155578 , 32'hEF60A7A0 , 32'h00003993 , 32'h06126640 , 32'hEFB74F40 , 32'h01F1E2E8 , 32'hFFFEABDB , 32'hF19E6040 , 32'hF9B9E8B8 , 32'h04F74388} , 
{32'h07C08240 , 32'h08228060 , 32'hFFFF3D64 , 32'hEB4B9980 , 32'hFFFF1A1B , 32'hFE62D140 , 32'h0000C77B , 32'hFFFF3312 , 32'h00003284 , 32'hFFFE9C5E , 32'hF0568D40 , 32'h00BD056B , 32'h09037240 , 32'h0001550E , 32'hFFFC7221 , 32'hFF222DFA , 32'h0000BE60 , 32'hF97D0AB0 , 32'h00C38132 , 32'hFFFDD744 , 32'hFFFF6D6F , 32'h020E09CC , 32'h0127C3E0 , 32'h00B8C801 , 32'h0A8C1A10 , 32'hFFFC8683 , 32'hFBFA7328 , 32'hFE13345C , 32'h000056D4 , 32'h0EA9B2A0 , 32'hFFFF3F9F , 32'h04DCD8C0 , 32'h000094F4 , 32'h00010676 , 32'h00003E66 , 32'h045F08A0 , 32'h060FEB70 , 32'hFD96D574 , 32'hFFFF955D , 32'hF19F25B0 , 32'h11FA48E0 , 32'h00001935 , 32'h00016FFD , 32'hFFF8C66A , 32'hFB1A7630 , 32'h0C1384E0 , 32'hF8F0EE58 , 32'h00016C7E , 32'h0BE3C270 , 32'hFA208330 , 32'hFEE1B458 , 32'h00010249 , 32'hFD9CBEFC , 32'h0CD3CB50 , 32'h022D4F04 , 32'hFFFE156B , 32'hFF831413 , 32'h000193A4 , 32'h00020C74 , 32'h05AC01E8 , 32'h0345B410 , 32'h05618208 , 32'h10C068E0 , 32'h0001A437 , 32'hF0119A90 , 32'hFFFDA25D , 32'hF1CA9E40 , 32'hFF95E3DA , 32'hFFFF7364 , 32'h19326600 , 32'hF50934D0 , 32'hFC4C61D8 , 32'h0004EF9B , 32'h000083AC , 32'hFFFEB635 , 32'h15C83BA0 , 32'hFC9BF264 , 32'hFFFEE63A , 32'hFCA37404 , 32'h0127B77C , 32'hFFFED634 , 32'h0F033C70 , 32'hF9A03FE0 , 32'h0000DA53 , 32'h00992BD7 , 32'h05D06418 , 32'h03674D18 , 32'hFFFB24FE , 32'hFFFCC589 , 32'h027AC7C8 , 32'hFFFF7726 , 32'h0293C014 , 32'h00004F97 , 32'h0879C870 , 32'hFE92CD54 , 32'hFFFDB99C , 32'hFFFF8558 , 32'h000008C4 , 32'h00019157 , 32'hFEE3ABA8 , 32'hFCC06C9C , 32'h0001DA81 , 32'hFA8044C0 , 32'h070ABF08 , 32'hFCE24474 , 32'hFFFE8255 , 32'hFF507D73 , 32'hFFFF515D , 32'h050C80E0 , 32'hF74D8FF0 , 32'hFFFF8DC6 , 32'h029764C8 , 32'hFFFD95F9 , 32'h00008C16 , 32'h0CCAC980 , 32'hFC615248 , 32'h01BC2684 , 32'h000076BA , 32'h062D1530 , 32'h00016B8D , 32'h0000C276 , 32'hF57413B0 , 32'h000102DA , 32'h00012C1C , 32'hF37C5DB0 , 32'h04B5E0B0 , 32'hFFFEBC4C , 32'h00011B08 , 32'hFFFF9B0E , 32'hFFFE13A5 , 32'hFFFE900B , 32'h0521BA80 , 32'hF8378D20 , 32'h0000C167 , 32'h00000EAC , 32'hEBE49680 , 32'hFD446524 , 32'h000064ED , 32'h00005623 , 32'hFD909DD4 , 32'h0001CAED , 32'hFFFF9090 , 32'hFC631B8C , 32'hFA129E60 , 32'hFE0EE780 , 32'hFDE0EED4 , 32'hFFFEE81E , 32'hFFFFEFCB , 32'h02ABCA98 , 32'hFFFE6C71 , 32'hFFFC8FC9 , 32'hFECB235C , 32'hFFFF3ED7 , 32'hFFFE47E4 , 32'hF5950E30 , 32'h00010EF6 , 32'hF6B01E60 , 32'h00E1D2F9 , 32'hFFFF20F2 , 32'hFFFFF238 , 32'hFFFF8CEA , 32'hF278E160 , 32'hF3282D50 , 32'h0232F868 , 32'hFA0E3098 , 32'h00008428 , 32'hD8F3C000 , 32'h0000E43C , 32'hFFFD77D3 , 32'h09751B10 , 32'hFC0EF09C , 32'hFFCEC0A2 , 32'h00025FC5 , 32'hEA9E7C60 , 32'hFE36C678 , 32'h09A4F810 , 32'hF97EA928 , 32'h0856A490 , 32'hF222EBF0 , 32'hFF0728D9 , 32'h136320A0 , 32'h0001BDD1 , 32'h00005975 , 32'hFFFFC9DC , 32'hF5FD3A90 , 32'hEF05BBC0 , 32'hFF526B68 , 32'h0111AFC8 , 32'hFD83DBC8 , 32'hFD8D3D90 , 32'hFFFEDE5E , 32'hEECFC2C0 , 32'hEE92C9C0 , 32'hFFFF2D06 , 32'hF462CA70 , 32'h0001A4B4 , 32'hFFE8A2D6 , 32'h19DA5E60 , 32'hFFFF18CA , 32'h0000FD03 , 32'hFFFEDCAE , 32'h00010352 , 32'h000027A8 , 32'hFFFF2B48 , 32'h018209BC , 32'h01F0617C , 32'hF10E0CE0 , 32'hFE932FEC , 32'hEBBE0C00 , 32'hFC2FE6C0 , 32'h0000081D , 32'hFFFF111C , 32'h0002552F , 32'hFFFEBD82 , 32'h0002EDE5 , 32'hFF032BFF , 32'hEDB289E0 , 32'h06C6BFC8 , 32'hFFFE0D5F , 32'hFFFF305B , 32'hFFFC1095 , 32'h00017648 , 32'hF4859ED0 , 32'h01E16BDC , 32'h00000A6A , 32'h0001C491 , 32'h00004A18 , 32'h16C093C0 , 32'h0FAC3CF0 , 32'hFA3B0758 , 32'h00010FE1 , 32'hFFFEEFE1 , 32'h00000F24 , 32'h01379DE8 , 32'h00514B28 , 32'hEFA50D80 , 32'h0001663F , 32'h0066D4B8 , 32'hFFFDD94C , 32'h0DE04910 , 32'hFFFE7F4C , 32'h043EF418 , 32'hFFFF9329 , 32'hF643BBA0 , 32'h03B82500 , 32'hF9B678A0 , 32'hF5CD4BD0 , 32'hFFFDED29 , 32'h04190750 , 32'hFFA6A913 , 32'h00020F85 , 32'h06A6D430 , 32'h00007CCD , 32'hFEB0BA30 , 32'h08EF9400 , 32'h0EA35AA0 , 32'h00022667 , 32'h0000CA43 , 32'h011A10E4 , 32'h0001B273 , 32'hE5455240 , 32'hFFFBE11B , 32'h023BEEF8 , 32'hFFFFFF00 , 32'h034B62F4 , 32'hFFFEAC31 , 32'h00010E64 , 32'hFFFD3DC7 , 32'hF822C378 , 32'hEA97DD80 , 32'h0002C907 , 32'hFFFFEA07 , 32'h000041C0 , 32'h000052A8 , 32'hFB678A30 , 32'hFE6C8E50 , 32'hF71941F0 , 32'h0690F7B8 , 32'h03F85580 , 32'hFFFFBBA9 , 32'hFFFEFFB3 , 32'h00003F48 , 32'h00946FA3 , 32'hFFFFD0C0 , 32'hFFFF897C , 32'hF9EF9230 , 32'hF31061B0 , 32'hFFFEEF74 , 32'h03E19FB8 , 32'hFBC9B730 , 32'h07315000 , 32'hFC24BFB0 , 32'h00005F09 , 32'hF8B600D8 , 32'h011A5C00 , 32'hFCBDFEAC , 32'hFFFEEBBE , 32'h04A8F0B8 , 32'hF9E1B020 , 32'h015ACAE8} , 
{32'hEBC5E840 , 32'hEB400D00 , 32'hFFFE7A7A , 32'hF641D3D0 , 32'h0000CABD , 32'h090392F0 , 32'hFFFF8477 , 32'h00002A22 , 32'hFFFF47AC , 32'h00036CA1 , 32'h02461DFC , 32'h0CF95AD0 , 32'hFFF72EAD , 32'h0001DCD9 , 32'hFFFF60ED , 32'h215CB2C0 , 32'h0000AE6B , 32'hFB0835B8 , 32'hF837EFD8 , 32'h00018801 , 32'hFFFF6F9F , 32'h01B8ABE8 , 32'h056455C8 , 32'h0CB62D20 , 32'h0A264890 , 32'hFFFE4002 , 32'hFFA1DCBE , 32'h00B251FB , 32'hFFFF5C0F , 32'hEEBD0440 , 32'hFFFE59F0 , 32'hF85B8C98 , 32'hFFFD377E , 32'hFFFEFE6D , 32'hFFFF1A35 , 32'h00E1A338 , 32'hEA2EBEE0 , 32'h04445548 , 32'h0000C6F3 , 32'h07B1E5D0 , 32'h076D54C0 , 32'h000242BD , 32'h00007D5B , 32'hFBD5E958 , 32'hFE3ECF24 , 32'h0A752240 , 32'hF46F9410 , 32'hFFFD6127 , 32'hFE84EEA8 , 32'h05DEC838 , 32'hFFB30A32 , 32'hFFFE532B , 32'h007A6EB8 , 32'h02AE627C , 32'hFF2AB52E , 32'h00012620 , 32'hFF17FE36 , 32'h0001D85C , 32'hFFFE72FE , 32'h00C5F408 , 32'hFEF93E24 , 32'hFC463F68 , 32'h0DB117E0 , 32'h0003A0DD , 32'h09051720 , 32'hFFFE7887 , 32'hE3936A40 , 32'hFFE05A0A , 32'h0000BDF5 , 32'h14A4A7A0 , 32'h0F5D4790 , 32'h08CF46D0 , 32'h00003418 , 32'h0000EEE6 , 32'h0001D113 , 32'hF9D32450 , 32'h047E04D0 , 32'h0000532C , 32'hFC2ABB68 , 32'hFD3F7E58 , 32'hFFFCFA47 , 32'h01C46918 , 32'hFF662607 , 32'hFFFE2A13 , 32'h0AA3EE20 , 32'hF091D510 , 32'hF9657510 , 32'hFFFF5BA3 , 32'hFFFFD211 , 32'h0969E960 , 32'hFFFE0FFC , 32'hF82BFDD0 , 32'hFFFF1DAC , 32'hFF1B454B , 32'hFF4B1DEC , 32'h0000993F , 32'h00008B02 , 32'h0000D4FE , 32'hFFFFACDD , 32'hF3109820 , 32'hFCEAFBF8 , 32'h00000B79 , 32'hF079B050 , 32'h0830C4C0 , 32'h03423C64 , 32'h00023706 , 32'h002D19FB , 32'hFFFFB515 , 32'h05E55A20 , 32'hFAAF0990 , 32'hFFFEEFF4 , 32'h05964688 , 32'h00004A3B , 32'hFFFEBC77 , 32'hF6A075D0 , 32'hF4DFEF20 , 32'hFEECE048 , 32'hFFFF867C , 32'h01B7AC40 , 32'h00012FC4 , 32'hFFFCD075 , 32'hFEC27AB4 , 32'hFFFF5330 , 32'hFFFF4E18 , 32'hFB7D2D90 , 32'h01A58CF4 , 32'h00002C1C , 32'hFFFF75CD , 32'hFFFF224D , 32'h0001DC98 , 32'h00005243 , 32'h09201950 , 32'h04A0AEA0 , 32'hFFFE9B71 , 32'hFFFEBDF9 , 32'h036B43B4 , 32'hF7193820 , 32'hFFFFBDB0 , 32'h00015711 , 32'h0E557A60 , 32'h00000ED9 , 32'hFFFCFAC1 , 32'h098F0CF0 , 32'h006FD1EC , 32'h02BC00E8 , 32'h000E2B00 , 32'h00032B6E , 32'hFFFE40B4 , 32'h047DAB98 , 32'hFFFEA971 , 32'hFFFFDAB1 , 32'h01418368 , 32'h00030E96 , 32'h00014F39 , 32'hF5361DA0 , 32'h0001FF9E , 32'hFFAF3C5C , 32'h00CD7ECC , 32'hFFFE4B0D , 32'h0000AD63 , 32'hFFFF3F0F , 32'h13EDCE00 , 32'h00B9F274 , 32'h034DCF18 , 32'h11304B40 , 32'hFFFF432E , 32'hFC16F028 , 32'h0000A183 , 32'h000086FF , 32'h07D79958 , 32'hFACE5A10 , 32'h01FA2E98 , 32'hFFFF75B5 , 32'hFE415518 , 32'hFE8D4C54 , 32'hE9AE94E0 , 32'h006471A1 , 32'h06B545D0 , 32'hFFCACC85 , 32'hFF2E36F2 , 32'h090A4150 , 32'h0000B92F , 32'h0001E7CC , 32'hFFFF4490 , 32'h07119260 , 32'h00E268FC , 32'h034D6BDC , 32'h0019E929 , 32'h02F613F4 , 32'hFB717C20 , 32'h0000A512 , 32'hEB056480 , 32'hFCE759FC , 32'hFFFE1BE3 , 32'h16D04A00 , 32'hFFFE124A , 32'hFD1641EC , 32'hFBB647C0 , 32'h0000FC3F , 32'hFFFF51D5 , 32'h0000094D , 32'hFFFF780E , 32'hFFFCA06B , 32'h00014B3F , 32'h02331720 , 32'h116A23E0 , 32'hF355FE70 , 32'hFB45BF18 , 32'h0AFB0740 , 32'hFAAB24A8 , 32'h000295F9 , 32'hFFFFDFA9 , 32'h0000021B , 32'hFFFD930A , 32'h0000F13A , 32'hFB9475E0 , 32'h06429DC0 , 32'hF80FE298 , 32'h000060F3 , 32'hFFFFCD75 , 32'h0001A9EB , 32'h00006042 , 32'h059F82C0 , 32'hE1D7BAA0 , 32'h0000B781 , 32'hFFFC2438 , 32'hFFFD9D37 , 32'hF5475530 , 32'h0CBCE3B0 , 32'hFCB82230 , 32'h0000BFE6 , 32'hFFFDFC8C , 32'hFFFE91F0 , 32'h01DB5F64 , 32'h015786F4 , 32'hFC8F2F04 , 32'hFFFFBC2C , 32'h000CC993 , 32'h000021D1 , 32'h16958880 , 32'hFFFFBE74 , 32'h0C4037B0 , 32'h00001F63 , 32'h1D16EE60 , 32'hFDBAA874 , 32'h06EED920 , 32'h08AA3EF0 , 32'h00006805 , 32'hF1C8F680 , 32'h016517FC , 32'h0000BE0B , 32'hFF80F6DB , 32'h000047B9 , 32'h03C6EB70 , 32'h0ADE0FB0 , 32'hFB0388F0 , 32'hFFFF2116 , 32'h0000470B , 32'hEEC174A0 , 32'h00004D35 , 32'h0E5313A0 , 32'h00031112 , 32'hFF6B6B99 , 32'hFFFF8EC3 , 32'h133C2240 , 32'hFFFFB8CC , 32'hFFFFA343 , 32'h00025FE3 , 32'hF2DB4FE0 , 32'hF828FE78 , 32'hFFFDB4E9 , 32'hFFFEFE7E , 32'h00002711 , 32'h000007A9 , 32'h0B4196B0 , 32'hFB7B2688 , 32'hF7400830 , 32'hF9F23348 , 32'hF745C5E0 , 32'h0001D864 , 32'h0000D746 , 32'h00003520 , 32'hFD730E20 , 32'hFFFE6BBF , 32'hFFFE5D80 , 32'h01176CDC , 32'h02CD8544 , 32'h00019446 , 32'h0A80BD30 , 32'hF5BCD6E0 , 32'hFDDCACAC , 32'hFC4A66B8 , 32'hFFFD6E21 , 32'hFCC5B270 , 32'hFC2B2EB0 , 32'hFEF02080 , 32'h0001B66A , 32'hF820CC40 , 32'h08E9C940 , 32'hF6214790} , 
{32'h083F79F0 , 32'h0152A108 , 32'h00001534 , 32'h06724F98 , 32'hFFFFF642 , 32'hFA8EC260 , 32'h0001803D , 32'h0001482E , 32'h00006082 , 32'h000012BA , 32'hF3682560 , 32'h0DCB3950 , 32'hFCDDB958 , 32'h00003D80 , 32'h00004A75 , 32'hF57DBD30 , 32'h0000B405 , 32'hFE7308CC , 32'h084F85F0 , 32'hFFFE0CA6 , 32'h0000AFD4 , 32'h00626A05 , 32'h04F17130 , 32'h03C9A36C , 32'hF9DAE040 , 32'h0001F02A , 32'hFD08F6F8 , 32'h01BB14F0 , 32'h0000548E , 32'hFD8D57BC , 32'h00001331 , 32'hF3952C10 , 32'h0000B1EF , 32'hFFFEB96E , 32'h000083A1 , 32'h0E5B2430 , 32'h17C2CEC0 , 32'hFEAFABE8 , 32'h00000147 , 32'h0994ECC0 , 32'hF1AEAD80 , 32'h0001EDCD , 32'h0000AD1D , 32'h0114C624 , 32'hFEEA97E8 , 32'hFC922B30 , 32'hFE41C528 , 32'h00017CEE , 32'h02A3B964 , 32'hEAFA0E80 , 32'hFFF62540 , 32'h0000E863 , 32'h02803C34 , 32'hF8BA2CA0 , 32'h044E3F28 , 32'h00001017 , 32'h03024028 , 32'hFFFF2063 , 32'hFFFDF838 , 32'hF98F8F88 , 32'hFE2F7A5C , 32'hFD5B04CC , 32'hF96B08D8 , 32'hFFFF3243 , 32'hF32E9460 , 32'h00006A1C , 32'hE6838F40 , 32'h00C785CA , 32'h00031494 , 32'hFAB4E690 , 32'hE448E5E0 , 32'h06AB2B48 , 32'h0000750C , 32'hFFFE46FB , 32'hFFFEC50E , 32'hEF8EC1C0 , 32'h03411A44 , 32'hFFFFEECB , 32'h108E27C0 , 32'h006229E3 , 32'hFFFA777F , 32'h0AB56F70 , 32'h02FA77AC , 32'h00026C44 , 32'h024B26FC , 32'hE70D1280 , 32'hFB4D59A8 , 32'hFFFF1A35 , 32'h0001A8B8 , 32'hF42263D0 , 32'h00008057 , 32'hFC66D3D8 , 32'hFFFF75FB , 32'h017F2208 , 32'h00446973 , 32'h0001267C , 32'hFFFEA394 , 32'hFFFEFC27 , 32'hFFFF8006 , 32'h04BEDE70 , 32'hFB020528 , 32'hFFFE0794 , 32'hF6E47340 , 32'h0343931C , 32'hFD612538 , 32'hFFFD18F5 , 32'hFF95ED08 , 32'hFFFD54F3 , 32'h02902CBC , 32'h279A18C0 , 32'h00005CD5 , 32'h06A69718 , 32'h00002C66 , 32'hFFFE1043 , 32'hF80EE478 , 32'h06D9E1D0 , 32'h010D6B40 , 32'h0001873E , 32'h0B2C02C0 , 32'h00011D73 , 32'h0000AE71 , 32'h0338E9B4 , 32'h0001E20D , 32'h00018D92 , 32'h0788CE50 , 32'h00F8EE0D , 32'h0000E989 , 32'hFFFD8FF4 , 32'hFFFF9A19 , 32'h0000804C , 32'hFFFFB3BB , 32'hFC8B702C , 32'hF8CB16D8 , 32'h0001872C , 32'hFFFE9AB2 , 32'hEBBD0DC0 , 32'hF9268C98 , 32'h0000D0DD , 32'h00001AE0 , 32'h0C8BF890 , 32'hFFFF60D1 , 32'h0001429D , 32'h04A7DDE0 , 32'h02E1FB90 , 32'hFC010108 , 32'h014E15AC , 32'hFFFEA069 , 32'hFFFCAB37 , 32'hFEB1E2DC , 32'hFFFE1082 , 32'h00022FBF , 32'hFF2DB29E , 32'h00023007 , 32'h00005779 , 32'hFA699188 , 32'h000456BE , 32'hFE5C34E4 , 32'h00A66888 , 32'hFFFF8BD2 , 32'hFFFFA3A2 , 32'hFFFD7F94 , 32'hF6781BB0 , 32'h02944A58 , 32'h05D99868 , 32'h01246B28 , 32'hFFFDE726 , 32'h0CAD8710 , 32'h00013023 , 32'hFFFEBEAB , 32'h0EFB9740 , 32'h0134BE54 , 32'hFAF4D2B8 , 32'h0000F2AE , 32'hDBEAE1C0 , 32'hFFD4532F , 32'hF9BA4450 , 32'hF1531B20 , 32'h08A65620 , 32'hEAA660E0 , 32'h0254AB4C , 32'hFE6222A8 , 32'h000057DA , 32'hFFFEC505 , 32'hFFFE8AD4 , 32'h0637A818 , 32'hFAF06440 , 32'hFFA9CEDB , 32'hFF115DCB , 32'h08AB7AF0 , 32'h06B60ED8 , 32'hFFFF5ADF , 32'h0BBACC50 , 32'h04465808 , 32'hFFFFB2ED , 32'h025F4678 , 32'hFFFF1B3D , 32'h0ACD96D0 , 32'h023EAB4C , 32'hFFFE1B07 , 32'h0001B6AF , 32'h00018D83 , 32'h0000F55E , 32'hFFFF4396 , 32'h0000B988 , 32'hFDAB9BC0 , 32'hFE0016AC , 32'hF90D3E38 , 32'h034ECFD4 , 32'h014A0758 , 32'hFB4AAA78 , 32'hFFFE4802 , 32'h000134D8 , 32'h0000432F , 32'h00018DEB , 32'hFFFF4DF5 , 32'hFB5EBE40 , 32'h088F52C0 , 32'h120A0700 , 32'h00011B96 , 32'h000209D1 , 32'hFFFEA95C , 32'h00020F09 , 32'h024380DC , 32'hF2F6B740 , 32'h000019C4 , 32'h00013E8B , 32'h0000F148 , 32'hF6439C10 , 32'h0C8842F0 , 32'hF39FF800 , 32'h000043A8 , 32'h00020F68 , 32'hFFFF649C , 32'hFC2B785C , 32'hFFEC5A73 , 32'hFB7C5DD0 , 32'h0000C467 , 32'hFF4B929A , 32'hFFFEC66B , 32'hFBFECAD0 , 32'hFFFFF2BB , 32'h067AE620 , 32'hFFFFEDB2 , 32'hFEF21E98 , 32'h049AA0A0 , 32'hFBF2EEA8 , 32'h11BAB480 , 32'h0000EFCF , 32'h016794E4 , 32'h00B936C8 , 32'hFFFE3212 , 32'h062719B0 , 32'h000181F6 , 32'hFDA58D24 , 32'hF1B9CDC0 , 32'h15D0DD60 , 32'hFFFFEBA0 , 32'h00001A99 , 32'hF800C1F0 , 32'hFFFEEEAE , 32'h020C3600 , 32'hFFFFB797 , 32'h026687A0 , 32'hFFFF19C4 , 32'h04BC58E0 , 32'hFFFE6580 , 32'h000093BB , 32'hFFFFD95C , 32'hFA6744B8 , 32'h152E1DA0 , 32'hFFFF9B12 , 32'h0002A8C9 , 32'hFFFEFDB2 , 32'hFFFE0AC1 , 32'hFA7CA5E8 , 32'h0DB2E620 , 32'hFAE43100 , 32'hF26DAAA0 , 32'h096209E0 , 32'hFFFD1FA3 , 32'hFFFDDF7E , 32'h0000CAED , 32'h056B9EE0 , 32'h00010A21 , 32'hFFFF9505 , 32'h0210CDCC , 32'h16DDEB20 , 32'hFFFCA81E , 32'hF1FEEBA0 , 32'h04826520 , 32'hFC1D456C , 32'hF9D0E8E0 , 32'hFFFF22A3 , 32'h016397B8 , 32'hFA265400 , 32'hFF60DEAA , 32'h00043A1E , 32'hF3F42CE0 , 32'hF354A050 , 32'hF4B4AF70} , 
{32'h1233A680 , 32'h03C0A2CC , 32'hFFFDAE99 , 32'hFDB13EA0 , 32'hFFFE6628 , 32'h06B55158 , 32'hFFFEA58A , 32'hFFFDC2A4 , 32'h00019A86 , 32'h00009ABE , 32'h060F5330 , 32'hF94738E0 , 32'hFAEB7190 , 32'h000090B6 , 32'h0000E397 , 32'h0763CEF0 , 32'hFFFFFA94 , 32'h0892F140 , 32'hFC794610 , 32'hFFFF8125 , 32'hFFFD633D , 32'hFFE44718 , 32'hF8222A00 , 32'h086B51F0 , 32'h07EAE868 , 32'h0000435F , 32'h0083DEB7 , 32'hFFD480C9 , 32'h000001D8 , 32'h150057E0 , 32'hFFFE2673 , 32'h01F55FCC , 32'hFFFE6645 , 32'h00002AC9 , 32'h000273F6 , 32'hF10A8300 , 32'hE97CBD00 , 32'hEE0E1E40 , 32'hFFFF28D4 , 32'h08B64430 , 32'hF12C3700 , 32'h00002081 , 32'hFFFF99A9 , 32'h05BF8D60 , 32'h19264DA0 , 32'hE9689F60 , 32'h0121BE80 , 32'h0000835A , 32'h076030C0 , 32'h062CEE80 , 32'hFF3409C3 , 32'hFFFF0BB6 , 32'hFB5CC1E8 , 32'h016D1464 , 32'hF7C9CF90 , 32'h00022A5E , 32'h00515E1F , 32'hFFFF23AB , 32'hFFFF8621 , 32'h02EE90D0 , 32'hFE4C5E28 , 32'h09E67E80 , 32'hF6498D90 , 32'hFFFEFBF3 , 32'h0BEEFC80 , 32'h00001188 , 32'hEBF93740 , 32'h0085856E , 32'hFFFE2142 , 32'hFCF438C0 , 32'hE6F5A360 , 32'hF376AF90 , 32'hFFFFD9E0 , 32'h0000C888 , 32'hFFFF3937 , 32'h07A6FB58 , 32'hFAF817F8 , 32'hFFFEBF21 , 32'hF8879508 , 32'h02990F7C , 32'h00005A3F , 32'h123A94C0 , 32'h01CB53C4 , 32'h00007347 , 32'h07072AF0 , 32'h03548A08 , 32'h050623F0 , 32'hFFFFBED1 , 32'hFFFFFA17 , 32'h05AA1ED0 , 32'hFFFEB3F2 , 32'h011394BC , 32'hFFFF75A9 , 32'hF6EF9830 , 32'h004C708E , 32'h0000E0C6 , 32'hFFFF8CAA , 32'hFFFE386C , 32'hFFFFC78D , 32'hF438CB40 , 32'hFFEB6307 , 32'h00020FAC , 32'hF674E0F0 , 32'h02FC4720 , 32'h01D67F2C , 32'hFFFF354D , 32'h002CEF91 , 32'h00017E5D , 32'h065D25C0 , 32'hF3D40F40 , 32'hFFFF513D , 32'h0A6EF8D0 , 32'h0000ACF0 , 32'h000112DE , 32'hFACE7D20 , 32'hFA367028 , 32'h0112A44C , 32'hFFFE4FA9 , 32'h063E3528 , 32'h00008428 , 32'h0001A760 , 32'h036EA8C4 , 32'h00021E1B , 32'hFFFDE5FE , 32'hF8C1E798 , 32'hF8E021B0 , 32'hFFFDF087 , 32'h0002F8C9 , 32'hFFFDF0F3 , 32'hFFFD72EC , 32'h00012280 , 32'h034D1984 , 32'hF7DEC720 , 32'hFFFEE079 , 32'hFFFF2B2C , 32'h0A60B330 , 32'hFD025934 , 32'hFFFFC8E8 , 32'h00005C27 , 32'h0BA30950 , 32'h000000B9 , 32'hFFFCB98A , 32'h01B04538 , 32'h0336528C , 32'hFF540D19 , 32'hFE13E634 , 32'h0000277B , 32'hFFFFF065 , 32'h0045AE95 , 32'hFFFED2EB , 32'hFFFEE37B , 32'hFDBC9D7C , 32'h000041A4 , 32'h00029822 , 32'h0A62F0C0 , 32'hFFFF484B , 32'hFA59FED8 , 32'h0119F0E0 , 32'hFFFFFCE0 , 32'h00001DF0 , 32'hFFFF213C , 32'hFC7C5ACC , 32'h023541EC , 32'h038A1718 , 32'h03A783E0 , 32'h000036D3 , 32'hF6F59A80 , 32'hFFFD8D55 , 32'h00019BB0 , 32'hFB3DCA88 , 32'h029BF3F8 , 32'h000EB73A , 32'h00013254 , 32'h04F3B3D8 , 32'h00A004D6 , 32'h00C72FEE , 32'h03A68908 , 32'hF944D850 , 32'hD9B90100 , 32'h008D89E5 , 32'hFC9C5474 , 32'h0001BD55 , 32'h000092EC , 32'hFFFF66FD , 32'hFE6DFFA8 , 32'h12ED6560 , 32'hFC7EE608 , 32'hFF3D7548 , 32'h01FB9AC4 , 32'hFA48BC78 , 32'h0003E153 , 32'h080CE6B0 , 32'hFA4DBEE8 , 32'hFFFF6F15 , 32'hF1D4AEB0 , 32'h000109E7 , 32'hFB6AC600 , 32'hF5E3CDC0 , 32'h000159A1 , 32'h00005891 , 32'h000076F4 , 32'hFFFDC30C , 32'h0002EF2C , 32'hFFFEA601 , 32'h0AD1D530 , 32'hFB6A3AF8 , 32'h1DFD7CE0 , 32'h0014C49A , 32'hFB2F0CE8 , 32'hFBB30150 , 32'h00010D9E , 32'h000087C0 , 32'hFFFFACA1 , 32'h000130D2 , 32'hFFFEE7B3 , 32'hFE9D9C48 , 32'hF6A5D9A0 , 32'hF487A7F0 , 32'h0000C995 , 32'h0001D174 , 32'hFFFFE5AD , 32'hFFFF04C3 , 32'hFF73D531 , 32'hEC9DAD20 , 32'hFFFD0EE5 , 32'hFFFF2640 , 32'hFFFC8DF4 , 32'hEF82CA80 , 32'hFC1C0D60 , 32'hF6538C00 , 32'h000150C8 , 32'hFFFF4AC9 , 32'hFFFECC10 , 32'h045409B0 , 32'hF9B160D0 , 32'hEA389EE0 , 32'h0000E168 , 32'hFF1D8B57 , 32'h00002AA4 , 32'h02F74D50 , 32'hFFFDB559 , 32'hEB683080 , 32'h0001F958 , 32'h034538C4 , 32'hFE1C20B0 , 32'h144BCD60 , 32'hF212E960 , 32'hFFFE1BC4 , 32'hF9A65190 , 32'hFF56D745 , 32'hFFFF6812 , 32'hFB0B8AD8 , 32'h0001D2DD , 32'h02A25754 , 32'h06BE1238 , 32'h009AEFB6 , 32'hFFFF7138 , 32'hFFFF2242 , 32'hF19E32E0 , 32'hFFFEFB7C , 32'h0F25D5C0 , 32'hFFFF99FE , 32'hFFF4FBF7 , 32'hFFFF91C0 , 32'hFEB1868C , 32'h00017FEC , 32'h00002BD7 , 32'hFFFF4270 , 32'h07CAACA0 , 32'hFBA59970 , 32'h0001386D , 32'h00008741 , 32'hFFFFF482 , 32'hFFFE66BB , 32'hEFEDAD00 , 32'h04AA5850 , 32'hF61D2980 , 32'h0D52DB90 , 32'h02F5EFB0 , 32'hFFFFEF61 , 32'h000133A1 , 32'hFFFEA8EF , 32'hFF9C35C1 , 32'h00014A43 , 32'h000227D3 , 32'hFA2EFF78 , 32'h0BAE2320 , 32'hFFFFCC49 , 32'hF0DC75D0 , 32'h01BABCB4 , 32'h060FD698 , 32'h032C8978 , 32'h0001C1AA , 32'hFEE528D4 , 32'hF86FDC08 , 32'hFF79F50F , 32'h000038A3 , 32'h0BABF300 , 32'hE260DC40 , 32'h0266DF60} , 
{32'h01851698 , 32'h064AE4E8 , 32'h00015FDB , 32'h05F4D770 , 32'hFFFF9442 , 32'h02485A58 , 32'hFFFE10CD , 32'h000040B7 , 32'h000111AE , 32'hFFFEB627 , 32'hF99778E0 , 32'hFF0F978C , 32'h081E48D0 , 32'h0000DE34 , 32'hFFFFD0A4 , 32'hFF999E2D , 32'h0000BD1A , 32'h066060B0 , 32'hFE7EF8D0 , 32'hFFFEBC2B , 32'hFFFFA377 , 32'hFC76421C , 32'h00674008 , 32'h086BF4B0 , 32'h11571D80 , 32'h0000667B , 32'h005E3300 , 32'h00693F18 , 32'hFFFE8776 , 32'h0B80A8B0 , 32'h0002ED52 , 32'h139BA840 , 32'hFFFC5241 , 32'hFFFFDAB4 , 32'hFFFF06C9 , 32'hF6846930 , 32'h18D6C200 , 32'hE73D24C0 , 32'h00001152 , 32'hEACDDE20 , 32'hFF0F9509 , 32'h00000A20 , 32'h0000111C , 32'h043DFCA8 , 32'h15844980 , 32'hF3A7DC20 , 32'hF4C8DEB0 , 32'hFFFCFDC7 , 32'hFF88AE20 , 32'hF17B3240 , 32'h0054591D , 32'h0000C973 , 32'h012BA6C8 , 32'h0AF480B0 , 32'hF4F06D80 , 32'hFFFE12B0 , 32'h00F064DC , 32'hFFFFFDE6 , 32'h000167D3 , 32'hFD7D5CA0 , 32'hFECEFDF4 , 32'hF93D9EE0 , 32'hF192EA10 , 32'hFFFFDDBB , 32'hF7ED2E50 , 32'hFFFF2159 , 32'hF6FDBFF0 , 32'h0035EAAE , 32'h0000B270 , 32'h012B5310 , 32'hF96663C8 , 32'hFA606F20 , 32'h0001FA92 , 32'h00013C45 , 32'h00005556 , 32'hFF138EE3 , 32'h049D3A60 , 32'h000125A1 , 32'h02E2CD7C , 32'h01B35034 , 32'hFFFECFAA , 32'hFCC8C3D0 , 32'hF6B22240 , 32'h00008C07 , 32'h0FC84A80 , 32'hFC87F880 , 32'h05B26288 , 32'h000238A3 , 32'h0000191D , 32'h08185E70 , 32'hFFFE9CFB , 32'h09DC8B10 , 32'h0000625F , 32'h0807F1C0 , 32'hFF8C5E3C , 32'hFFFED507 , 32'h0000DC11 , 32'h00000136 , 32'h00016240 , 32'hF9A2CBC0 , 32'hFEED7A0C , 32'hFFFEF55D , 32'hFD8EAE08 , 32'h06B8CAD8 , 32'h0129A7FC , 32'h00006CB9 , 32'h0030610A , 32'hFFFE0258 , 32'h103EE1A0 , 32'h06BAEE38 , 32'h00001394 , 32'hF32909C0 , 32'h000108EB , 32'h0001C969 , 32'h041B4618 , 32'h025591A4 , 32'hFD561C20 , 32'h00027A3F , 32'h0134DBF8 , 32'h000081B4 , 32'h0001FF1B , 32'h00CC7F91 , 32'hFFFE5955 , 32'hFFFEBF4D , 32'h0BB2E670 , 32'h0290C754 , 32'hFFFF24D8 , 32'hFFFE34EF , 32'h0001EF7B , 32'h0000BCA8 , 32'hFFFF43F1 , 32'h0865B220 , 32'h04A9B310 , 32'h00000DC9 , 32'hFFFEC1C1 , 32'hF8D7AF38 , 32'hF721AF60 , 32'hFFFF0B78 , 32'h000264D2 , 32'h0086342B , 32'h0000B6FC , 32'hFFFFD248 , 32'hFED8003C , 32'h008E0FF9 , 32'h015D6784 , 32'hFC6379D8 , 32'hFFFFCE5D , 32'hFFFDACA8 , 32'hFE1448EC , 32'h0001C221 , 32'hFFFFD89D , 32'h01CD42BC , 32'hFFFF6447 , 32'h000077C7 , 32'h035E2C0C , 32'h00010AF4 , 32'h021D3C28 , 32'hFFC62512 , 32'hFFFD8CFF , 32'h0002E439 , 32'h00003D84 , 32'hF9E57B78 , 32'h035A60D0 , 32'h06A1DB90 , 32'h06283A98 , 32'h0001073E , 32'h14EC2E40 , 32'h0000C973 , 32'h00007489 , 32'hF2D9CD90 , 32'hFFF70699 , 32'hFF29C93A , 32'h000040D9 , 32'hFFE22825 , 32'h02433B18 , 32'h0A7AB2E0 , 32'h01AFF92C , 32'hF2C26170 , 32'hF2042650 , 32'h01B792F4 , 32'hFFC9AFD8 , 32'hFFFFD41F , 32'h00002D36 , 32'h0000FD6A , 32'hF6E25D00 , 32'h0311DBD4 , 32'hFCA11000 , 32'hFF08543C , 32'hFE46C868 , 32'h04481710 , 32'hFFFDF9D4 , 32'h02C8248C , 32'h02AD3040 , 32'hFFFF43C2 , 32'h21310A80 , 32'h00003936 , 32'hFDA59F90 , 32'hFB8EDE98 , 32'h0000F5CA , 32'h0000643B , 32'hFFFF88C8 , 32'hFFFFD3C8 , 32'hFFFE1949 , 32'h00004E95 , 32'hFA3F5760 , 32'h0DC4A020 , 32'h13EE9BE0 , 32'h0A17E950 , 32'h002BFF23 , 32'hFB4AED18 , 32'h00006423 , 32'h00002FA0 , 32'h00009FEF , 32'hFFFEF6DE , 32'h0001F663 , 32'h01CA1A90 , 32'h02A0BBDC , 32'hF94C05C8 , 32'h0002F2C8 , 32'hFFFF8F80 , 32'hFFFD653A , 32'hFFFFE94E , 32'h0163B0D4 , 32'hFBBE04D8 , 32'hFFFE49F1 , 32'h00007830 , 32'h00016736 , 32'h0B614E80 , 32'h1AB54F20 , 32'h114518C0 , 32'h00002B79 , 32'h0001DF86 , 32'hFFFCD594 , 32'h05C2AE00 , 32'h03F91B1C , 32'hFE9E4F00 , 32'h00006F00 , 32'h0145CE04 , 32'h000086DB , 32'hFCF1C57C , 32'h0001958A , 32'hFE445208 , 32'h0001DB94 , 32'hF66C3A90 , 32'h038847A8 , 32'h09E8CEA0 , 32'h0B6D8F00 , 32'hFFFFB851 , 32'h02F10D40 , 32'hFF5FCC2E , 32'h00008256 , 32'h08559C50 , 32'hFFFF1E6B , 32'h03D14AFC , 32'h17690260 , 32'h01ADAEC8 , 32'hFFFFE9CB , 32'h00004B7E , 32'hF7923220 , 32'hFFFF3387 , 32'hF7291E60 , 32'h00002841 , 32'h00EA6330 , 32'hFFFEA1CB , 32'hF8E91B78 , 32'hFFFDD272 , 32'hFFFF76B9 , 32'hFFFFF421 , 32'h0C1739F0 , 32'h057AD9A8 , 32'hFFFEB923 , 32'hFFFF856C , 32'hFFFF3B6B , 32'hFFFEF8DC , 32'h2DF24DC0 , 32'hF76F1520 , 32'hFE6E91C0 , 32'hFCEA2D34 , 32'hFBC9DDF0 , 32'h0000087E , 32'h00003630 , 32'h00016B7C , 32'h022BC324 , 32'hFFFEA938 , 32'h00010BDA , 32'h026429C4 , 32'hFB3E8250 , 32'hFFFF732E , 32'h0F455660 , 32'h012B74F8 , 32'h00E1747B , 32'h0DA0C490 , 32'h00004B54 , 32'hFA9A38C8 , 32'h052B2310 , 32'h00740DE3 , 32'h000094CA , 32'h08465430 , 32'h250EA840 , 32'h08CCE670} , 
{32'h0039F1C9 , 32'h03E50064 , 32'h0000101F , 32'hFBA0F160 , 32'h0002AEF4 , 32'h00B76A3A , 32'hFFFDCD20 , 32'h00004046 , 32'hFFFD3076 , 32'h0003953F , 32'h05A80E98 , 32'h080628F0 , 32'h089B0140 , 32'h000152E9 , 32'h00007565 , 32'hF844D100 , 32'hFFFFD47B , 32'h04919F40 , 32'h03E37AB4 , 32'hFFFF1D19 , 32'hFFFFE991 , 32'h01C2E28C , 32'h0C2A8180 , 32'hFE270F0C , 32'hED847100 , 32'hFFFFD9ED , 32'h01111168 , 32'h03F568F0 , 32'h0001C46E , 32'hEC8CB600 , 32'h00009F7F , 32'h09413850 , 32'hFFFFF7BD , 32'h0002F07E , 32'h00007454 , 32'hFCBFB820 , 32'hE448AD40 , 32'h040B7AE0 , 32'h00014E9B , 32'hFB05B420 , 32'h01FB2D3C , 32'h000042B9 , 32'hFFFF404A , 32'hFED6C2B8 , 32'hFDDB7AF4 , 32'hEFAE3200 , 32'hFEF6A0EC , 32'h00010CCC , 32'hFE22C0BC , 32'hFCAD78C4 , 32'h01D96550 , 32'hFFFE8C88 , 32'h068AE868 , 32'hFA5E1A20 , 32'h0F058B40 , 32'h00013FFA , 32'h010C0C14 , 32'hFFFFCEF6 , 32'h0001EEC7 , 32'hFF128188 , 32'h01CD2934 , 32'hFCE7AF38 , 32'hEDD625A0 , 32'hFFFF5B52 , 32'hF4C36120 , 32'h0000F8CF , 32'h05593520 , 32'hFFFFC1C3 , 32'h00023E8A , 32'hF51BF280 , 32'hFEB0D5E4 , 32'hFD3CAF20 , 32'h00006701 , 32'h00002A17 , 32'hFFFECA4F , 32'h04E2F590 , 32'h02BD8EBC , 32'h0000FD69 , 32'h1136C220 , 32'hFEF2F000 , 32'h0001698B , 32'h1D223540 , 32'hF5DE0C80 , 32'hFFFC4409 , 32'h009E4126 , 32'hFAFFFBD0 , 32'h01BBEDD0 , 32'h000079A9 , 32'h0000F6F5 , 32'hFAE28470 , 32'hFFFEEE83 , 32'h04EDDFC0 , 32'hFFFFBE51 , 32'hFF4B342D , 32'h002D50DF , 32'h0000C6AB , 32'h00001A35 , 32'hFFFF9B45 , 32'h0002A480 , 32'h00A6F5A6 , 32'hFE27CA90 , 32'h0003D19F , 32'hEF7AECA0 , 32'hF2BD2250 , 32'h055BF3C0 , 32'h00004BA6 , 32'hFF6DB25A , 32'h00014898 , 32'hF9456A50 , 32'h061A1238 , 32'hFFFEAFC5 , 32'h01D69908 , 32'h0000D2DF , 32'hFFFE1FC9 , 32'hF8435C50 , 32'hF9E97340 , 32'h00FEA380 , 32'hFFFEDD00 , 32'hFF871279 , 32'hFFFF6160 , 32'h00005F47 , 32'hFE2858FC , 32'hFFFF8399 , 32'hFFFFEB26 , 32'h05BC1280 , 32'h112BFA60 , 32'h00000BF8 , 32'hFFFF98D6 , 32'hFFFE3111 , 32'h0001503E , 32'hFFFF853B , 32'hF51A5DA0 , 32'hFD230A0C , 32'h0000178F , 32'h00015346 , 32'h1D7D5F20 , 32'h07804548 , 32'hFFFD8BEA , 32'h00015876 , 32'h049E7F38 , 32'hFFFFDD0D , 32'hFFFE70FC , 32'hFF06C7EC , 32'hFC9744E8 , 32'h01504768 , 32'hFE7FA25C , 32'hFFFED9C4 , 32'hFFFF91B9 , 32'hFF0A22F0 , 32'hFFFEFCCE , 32'h000178CC , 32'hFB1D47E8 , 32'hFFFEC149 , 32'h00006E05 , 32'hEEC4D860 , 32'h0000C7B6 , 32'hFFD97DCF , 32'h0127B61C , 32'hFFFE8BA8 , 32'h0001622E , 32'h00019B25 , 32'h06ED0A80 , 32'hF8289C90 , 32'hF8F27688 , 32'h02400588 , 32'h000141CF , 32'h098127C0 , 32'h0000CC50 , 32'h0002555C , 32'hF8FE9C28 , 32'hFC3770B4 , 32'hFBC3AD00 , 32'hFFFF075B , 32'hEEC1D660 , 32'hFC5F86A8 , 32'h099836B0 , 32'h09D9C230 , 32'h15F7F020 , 32'hFF628527 , 32'h01114510 , 32'hF37CF350 , 32'hFFFE3A1A , 32'h0000D7E2 , 32'h00011287 , 32'hF93A3530 , 32'h1123ADA0 , 32'h05A3B698 , 32'hFECAE1E4 , 32'hFF7272B8 , 32'hFACF8290 , 32'h00008FB0 , 32'hF1C80380 , 32'hFC0A3E10 , 32'hFFFF7C01 , 32'hFBEE3428 , 32'hFFFFB799 , 32'hFD0D0294 , 32'hF9813618 , 32'h00002A42 , 32'hFFFF87E1 , 32'hFFFEF8F1 , 32'h00006589 , 32'h00012238 , 32'h00003D7A , 32'h03769550 , 32'h033FF008 , 32'h0A819A30 , 32'h000A98A3 , 32'h075A57C0 , 32'h011AFE20 , 32'hFFFEFAEB , 32'hFFFE968A , 32'hFFFF0762 , 32'h00027089 , 32'hFFFFD3F2 , 32'hFC973EC0 , 32'hFF0FD7AB , 32'h09C03E40 , 32'h0000740B , 32'hFFFFE9AA , 32'h00005339 , 32'hFFFF2B54 , 32'h0385D450 , 32'h0A4EE350 , 32'hFFFFAC44 , 32'h000218A3 , 32'hFFFF0643 , 32'h153A9C80 , 32'h02EEF758 , 32'hF4835490 , 32'h0000DBC5 , 32'hFFFF4CD6 , 32'hFFFF7C30 , 32'hF2FC5CA0 , 32'hFE28BF14 , 32'hEE39E180 , 32'h000083F7 , 32'h01307FAC , 32'hFFFF6423 , 32'h04110A38 , 32'hFFFEE11B , 32'h17459740 , 32'h0002427D , 32'hFA06B890 , 32'hFEFDE8DC , 32'hFB04F0F0 , 32'h1FA99220 , 32'hFFFFD7C8 , 32'hF5033E60 , 32'hFFF4DA6C , 32'h0000631B , 32'h06945EA8 , 32'hFFFFD65A , 32'h00E65C59 , 32'h11ED9C60 , 32'hFA6C4A98 , 32'hFFFDA46B , 32'hFFFEFBE4 , 32'h053AF190 , 32'hFFFD5F9F , 32'hF728BCD0 , 32'hFFFEDD78 , 32'h015E8FD8 , 32'hFFFF94BE , 32'hF5CB9530 , 32'h00004022 , 32'hFFFE23BB , 32'h000133CE , 32'hFA599888 , 32'hFD0F2360 , 32'hFFFFE222 , 32'hFFFE39F7 , 32'hFFFDBD33 , 32'hFFFF5723 , 32'hFE1D87A4 , 32'h0066D85A , 32'h01B474F0 , 32'h133D5880 , 32'hF4CAFFF0 , 32'h0000E3E1 , 32'hFFFEC93C , 32'h00007586 , 32'hFEB02210 , 32'hFFFDD2B3 , 32'hFFFD1A53 , 32'h01D0613C , 32'hFD929854 , 32'h00001718 , 32'h11EC8760 , 32'h0133A398 , 32'h002B3CEF , 32'hFD66F2F0 , 32'hFFFD9B2A , 32'h03B5E620 , 32'h08F188A0 , 32'hFDFFB448 , 32'h00007688 , 32'h2BAB6380 , 32'hFA7768F0 , 32'hECDF4C20} , 
{32'hF9E27210 , 32'h04CE5780 , 32'h0001E232 , 32'hE4B13E80 , 32'h000040B2 , 32'hFB1F3AD0 , 32'h00010ADD , 32'h0001042F , 32'h000181CE , 32'h00003ABC , 32'hF63EF950 , 32'h0C8F63A0 , 32'hF9CDDDD0 , 32'hFFFF3D84 , 32'hFFFEDAF9 , 32'h00B52672 , 32'h0000694C , 32'h242CC1C0 , 32'h00AAD52A , 32'h000333D6 , 32'hFFFFEBAB , 32'h052146D8 , 32'hFE5C7968 , 32'hFEC190BC , 32'hF8F796D8 , 32'h00014D9A , 32'h024533F8 , 32'hFE97398C , 32'h0001E90E , 32'hFAC65178 , 32'hFFFFD896 , 32'h06775F28 , 32'h00009694 , 32'h0001BB9C , 32'hFFFEC9D0 , 32'h0ADDD8A0 , 32'hFB4DC160 , 32'hF62F4B70 , 32'hFFFF8B40 , 32'h0A6DCB80 , 32'hFDEEDB98 , 32'h0000E3E4 , 32'hFFFFE99F , 32'h00C4BE77 , 32'h01A0E03C , 32'h12582420 , 32'h0316E1AC , 32'h0000D716 , 32'h037B3DDC , 32'h071AA960 , 32'h001AF671 , 32'h00036F95 , 32'h010AAC78 , 32'h039FC84C , 32'hF8C26E88 , 32'h00017A02 , 32'h00F1A572 , 32'hFFFEB020 , 32'hFFFFEEF7 , 32'hFB8B2DA0 , 32'h00745652 , 32'hFBD0FC70 , 32'hFBDC9958 , 32'h00006039 , 32'hF87384A0 , 32'h000009AB , 32'hE6B59F20 , 32'h0212732C , 32'h00000B76 , 32'h00B7ED96 , 32'hF6DB8D00 , 32'hFEF7F14C , 32'h000171D8 , 32'hFFFFBDBD , 32'hFFFF2070 , 32'hEE90BA60 , 32'hFE1253A0 , 32'h0003E5C1 , 32'h09330320 , 32'h01A2E98C , 32'h00001A06 , 32'hF0C12E70 , 32'h042641B8 , 32'h00000F47 , 32'h0129E1F8 , 32'h097BDD50 , 32'h00D72B1D , 32'h0002E352 , 32'h0000B370 , 32'hF5E89800 , 32'h00005E89 , 32'h01A943FC , 32'h0000C90E , 32'hFC930D98 , 32'h00B20AC1 , 32'hFFFDF32B , 32'h0001C4BE , 32'h0000857D , 32'hFFFEE215 , 32'h061B34A8 , 32'h05D516E8 , 32'hFFFF4163 , 32'h077754B0 , 32'hFF6FD330 , 32'h031D393C , 32'h00011ACF , 32'h000A2D7A , 32'h0000438B , 32'hFEC3CD7C , 32'h0020FD81 , 32'h000165B5 , 32'h03455398 , 32'hFFFFB526 , 32'hFFFF65A2 , 32'hF9C0B2B0 , 32'h099754A0 , 32'h01B4C9C4 , 32'h0001F173 , 32'h02CD1440 , 32'hFFFE795D , 32'hFFFFC834 , 32'h009B7E62 , 32'hFFFED7CF , 32'h00012737 , 32'h1EBA7160 , 32'h1312F4E0 , 32'hFFFF688F , 32'hFFFFFB90 , 32'hFFFCCD72 , 32'h00022A34 , 32'hFFFFF849 , 32'h005475E6 , 32'h063852C0 , 32'hFFFF5EE8 , 32'h0000764F , 32'hFFE45ACB , 32'h02BC003C , 32'hFFFF078C , 32'hFFFF849F , 32'h072C59E0 , 32'h00015EE2 , 32'h0001E827 , 32'hFF2FD53B , 32'hFB5D1080 , 32'h01243F58 , 32'hFF6637E0 , 32'hFFFF8FE7 , 32'hFFFF5D3E , 32'hFCA4CA34 , 32'h0001DF26 , 32'h000140B6 , 32'hFEE89E30 , 32'hFFFD8818 , 32'hFFFC2B9D , 32'hFF6F8795 , 32'h00032F15 , 32'h0D6D9400 , 32'hFF24957B , 32'hFFFFF63E , 32'h0000B794 , 32'hFFFEF486 , 32'h0320F7B0 , 32'hFF205A86 , 32'h03079E44 , 32'h0BD0C850 , 32'hFFFFE5B7 , 32'hD6F23780 , 32'hFFFF951B , 32'h00006B26 , 32'h09F67D20 , 32'h08C0E520 , 32'hFFFF54A7 , 32'hFFFF8B9C , 32'h1E036500 , 32'h0019589A , 32'h09B5A9F0 , 32'h0B612330 , 32'hF5225320 , 32'h03478CB0 , 32'hFDD5D594 , 32'h03EAB3DC , 32'h0003D1EC , 32'hFFFE2F83 , 32'hFFFFF46E , 32'h06A45B08 , 32'h1AC80EA0 , 32'h021779F0 , 32'hFFF06C29 , 32'h01260188 , 32'h0567F300 , 32'h0000481E , 32'hF5FF8EC0 , 32'h0EC91E50 , 32'h0000631B , 32'h0DB271B0 , 32'h00024C29 , 32'h03E82644 , 32'hFCE695E0 , 32'hFFFFC0E5 , 32'h00020346 , 32'h0001660B , 32'hFFFE8B8D , 32'h000031DE , 32'h00024E00 , 32'hFBE9D9E0 , 32'hFDF7AED4 , 32'h00F24EBF , 32'hFE534718 , 32'h0096E387 , 32'hFE385EC4 , 32'hFFFF283A , 32'h0002F79C , 32'h00007FA8 , 32'h0000ED28 , 32'h000168F3 , 32'h03F02F24 , 32'h03E4CE60 , 32'h241C2240 , 32'hFFFF8110 , 32'h00007A1E , 32'hFFFF6310 , 32'h00029B07 , 32'hF91648A0 , 32'hF1131620 , 32'hFFFFEE23 , 32'hFFFE4ED7 , 32'h0001C225 , 32'hFAB8CE38 , 32'h059F2288 , 32'hF55925A0 , 32'h000259CF , 32'h00002347 , 32'hFFFFB40A , 32'h006E2BFA , 32'hFFF2FE22 , 32'hFF960BEC , 32'hFFFFE73A , 32'hFE0013D8 , 32'hFFFCD6E9 , 32'h093BB7A0 , 32'hFFFF327F , 32'hF4923C00 , 32'hFFFF1CD3 , 32'hEC37A1C0 , 32'hFF104766 , 32'h066250C8 , 32'h07DB1A98 , 32'hFFFF8DB4 , 32'h05C469A8 , 32'h001068E4 , 32'hFFFE8C42 , 32'h09A4ABD0 , 32'h00004416 , 32'hFBF99858 , 32'hEA918440 , 32'hED97B1C0 , 32'hFFFFF9BA , 32'h0000BAE3 , 32'h0113F698 , 32'hFFFE39F8 , 32'hF19572C0 , 32'hFFFEA933 , 32'hFEF2EC80 , 32'h0002D68D , 32'hF87F33C8 , 32'h0000C5F0 , 32'h0000DB7E , 32'h000132F3 , 32'h0DE3D1C0 , 32'hFFC46AC5 , 32'h00024868 , 32'hFFFFD61A , 32'h0001A71B , 32'hFFFFA25F , 32'hFAC05918 , 32'hFB97CBB8 , 32'h09C27640 , 32'hFAC57488 , 32'hFFFFC056 , 32'hFFFF4E59 , 32'h0000A9EC , 32'h0000C288 , 32'hFD140FE8 , 32'hFFFF1CEF , 32'h00017938 , 32'hFF77A77A , 32'hECFB1720 , 32'hFFFEAB01 , 32'hF91DA450 , 32'hFCB67DD8 , 32'hFC67D374 , 32'hFE80F138 , 32'h0000C401 , 32'h0528C7E0 , 32'hFDAF26E0 , 32'h020E2F50 , 32'hFFFF9844 , 32'h0C12DD50 , 32'h0241975C , 32'h03FA0988} , 
{32'h0190FA00 , 32'h08034580 , 32'h00005725 , 32'hF84155F0 , 32'h0000EEA5 , 32'hFBC454C0 , 32'h000259CF , 32'h0001BF1C , 32'h000255E7 , 32'h0000ECA0 , 32'h06F326B0 , 32'hF3A6E3B0 , 32'hFBA78F78 , 32'hFFFEF8A2 , 32'hFFFF8E93 , 32'hE60AA660 , 32'h0001259A , 32'hE10CA5A0 , 32'h0B97D5D0 , 32'hFFFF5B0A , 32'hFFFDB894 , 32'h01227AD4 , 32'hF8D083D0 , 32'hFA96B8F0 , 32'hEB21D340 , 32'hFFFF56D3 , 32'h00983C1A , 32'h0016967C , 32'hFFFFC887 , 32'hF4ECEED0 , 32'hFFFE0943 , 32'hFCE6F47C , 32'hFFFDC6B0 , 32'hFFFF6C41 , 32'hFFFDBE6B , 32'h0629B320 , 32'h140B4060 , 32'h07D955B0 , 32'h00024BF0 , 32'h047C9568 , 32'hF7FCB400 , 32'h0001D68B , 32'h000063DD , 32'hFF494821 , 32'h11D741E0 , 32'hF57CCDA0 , 32'hFD95DFD0 , 32'h00002477 , 32'hF52B1EF0 , 32'hFD25CFF8 , 32'h00AB77E0 , 32'hFFFF1845 , 32'h03FA22A0 , 32'hF38DDC20 , 32'hFEB28658 , 32'hFFFFD083 , 32'h00CDF7C9 , 32'hFFFFBC55 , 32'h000143D4 , 32'h030ECA40 , 32'hFE41282C , 32'hFC21D190 , 32'hEB343860 , 32'h0000DF26 , 32'hF37AA180 , 32'hFFFE7BA5 , 32'hF25F98B0 , 32'hFEA8C9C8 , 32'h0002266A , 32'h23225240 , 32'hFFA18C47 , 32'hF6F88CC0 , 32'h00006607 , 32'hFFFFF041 , 32'h000090AB , 32'hFF6C0672 , 32'h01372660 , 32'h0001039B , 32'h0CCD99B0 , 32'hFE9D4324 , 32'h0001169B , 32'h043BDEC0 , 32'h0816B5B0 , 32'h0000AA75 , 32'hFFEAD8B6 , 32'h0219322C , 32'hFEEF971C , 32'h0000C778 , 32'hFFFF04B0 , 32'h1CCCF3C0 , 32'h00019910 , 32'h00678E78 , 32'hFFFDBA2C , 32'h02B56890 , 32'h003BA326 , 32'h0001FEB2 , 32'h0001FCCC , 32'hFFFEBDEA , 32'hFFFFACCA , 32'h04EBE6F8 , 32'h0134A7DC , 32'h0000CE9D , 32'h070F1788 , 32'h118A6240 , 32'h04D04090 , 32'h0000625D , 32'h0010F6E6 , 32'hFFFE77E7 , 32'hFA36B7D0 , 32'h01EAF358 , 32'h00004FD7 , 32'h23B2D200 , 32'hFFFF6DAA , 32'h00014A7C , 32'h08469990 , 32'h00968FC4 , 32'hFD05AA3C , 32'h000008A5 , 32'h0A8F8970 , 32'h0000DBCE , 32'h0001B9C8 , 32'h01E86E24 , 32'h0001301A , 32'h0002069F , 32'h03C82444 , 32'hF4EDFD10 , 32'hFFFFDF6C , 32'hFFFCA3FE , 32'h000002EA , 32'hFFFDDAAB , 32'h00013C0B , 32'hF6CE2EE0 , 32'h04E6C540 , 32'hFFFEFF6A , 32'h000123E2 , 32'h0F00ED60 , 32'h0219CB10 , 32'h0000064E , 32'h00017012 , 32'hFCA460DC , 32'hFFFDB375 , 32'h000053A5 , 32'hFFDBF98F , 32'hFC7A9CB0 , 32'h00CBB56C , 32'hFF6D78AC , 32'hFFFFD8B1 , 32'hFFFFBBAF , 32'hFB601E20 , 32'hFFFFBE85 , 32'h0000EAF4 , 32'h02962E3C , 32'hFFFE9CB2 , 32'h000135CE , 32'h0A950E10 , 32'h0000CC67 , 32'h08069CC0 , 32'hFF558552 , 32'h0001248C , 32'h00013C9D , 32'h00000669 , 32'hF88595B0 , 32'h08FBE2D0 , 32'hFA859D78 , 32'h01E43F9C , 32'hFFFEBD53 , 32'hFE99FC68 , 32'hFFFE6150 , 32'h0001A6A3 , 32'h0B8CB330 , 32'hFD2C3AC0 , 32'h03A9ECC8 , 32'hFFFF088B , 32'h0AEED520 , 32'h012F3A6C , 32'h0276E530 , 32'h064C0DD0 , 32'h073034E8 , 32'h073E8160 , 32'hFFC86473 , 32'h0C450550 , 32'hFFFF20FB , 32'hFFFF698C , 32'hFFFF900E , 32'h07590858 , 32'hF56959F0 , 32'h0181D4D4 , 32'hFFD6592E , 32'h014A6E64 , 32'hFEE9C900 , 32'hFFFFA900 , 32'hFF9992A5 , 32'hFE8B83E8 , 32'hFFFE19A3 , 32'h093CA2B0 , 32'hFFFCE6E3 , 32'hF47AE830 , 32'hFB49E830 , 32'h0000B716 , 32'hFFFEB3B6 , 32'h0001CCB0 , 32'hFFFF488C , 32'hFFFD9853 , 32'hFFFF3B32 , 32'hF677AA80 , 32'h0FFD44E0 , 32'h03030E38 , 32'h01D1F5A4 , 32'h11E6B8E0 , 32'hEC73FF00 , 32'h0000442D , 32'hFFFE3B84 , 32'hFFFE545B , 32'hFFFF98DA , 32'hFFFF90AA , 32'hFE3E91D0 , 32'hFA791428 , 32'hF7954120 , 32'h000007CF , 32'h00009C6E , 32'h0000F530 , 32'h00000494 , 32'hF7F75340 , 32'hF6138260 , 32'h0000124A , 32'hFFFF1794 , 32'hFFFF412E , 32'hFC68B4C0 , 32'hEC02E340 , 32'hECA3DE40 , 32'h000232BA , 32'hFFFE384A , 32'h00013655 , 32'hFABF28C8 , 32'hFBD440D0 , 32'h01016334 , 32'h00028DA8 , 32'hFF56FC2E , 32'h00047CD6 , 32'h0684F078 , 32'hFFFE9FA8 , 32'hFE3A1088 , 32'hFFFBE179 , 32'hFB2D07A0 , 32'h005BCD9F , 32'h0690C108 , 32'hF9A41218 , 32'h00004000 , 32'h01FF3C74 , 32'hFD4020CC , 32'h00020B91 , 32'hFD748018 , 32'h0002583B , 32'h02C6144C , 32'h13CFFDC0 , 32'h08BBAC70 , 32'hFFFE860C , 32'h00010F20 , 32'h0F0E8F20 , 32'hFFFCB2E9 , 32'h064DD320 , 32'hFFFEAF6F , 32'hFF24DA74 , 32'h00014473 , 32'h04634BF0 , 32'hFFFEE488 , 32'hFFFD7078 , 32'h000028C2 , 32'h01941000 , 32'hF4CB3DD0 , 32'h000093E4 , 32'hFFFD6158 , 32'hFFFCFCB8 , 32'hFFFFDA41 , 32'h036A3F64 , 32'hFA394B10 , 32'h0A65CF90 , 32'hE9232E00 , 32'h0378E3A0 , 32'h00005B6F , 32'h0000D910 , 32'h0002100C , 32'h02F45E54 , 32'h0000E369 , 32'h0001B85D , 32'hFB618510 , 32'hE804CA40 , 32'hFFFF9A0F , 32'h0BAC6FF0 , 32'hFEF7B5D4 , 32'hF515EFC0 , 32'h0ED32700 , 32'hFFFF0092 , 32'h09F05060 , 32'h02EE9FFC , 32'h01307B4C , 32'hFFFFBAF0 , 32'h0182B578 , 32'hF2723540 , 32'hFDFBF564} , 
{32'h02C91B58 , 32'hFA90B440 , 32'h000131E8 , 32'hFD7235C4 , 32'h00007F06 , 32'h014A490C , 32'hFFFE3BF6 , 32'h000089A1 , 32'hFFFE8FC9 , 32'h00013220 , 32'hFBADC170 , 32'h0EB5DBA0 , 32'hFD7B5C7C , 32'hFFFE8CA6 , 32'hFFFF9355 , 32'hF6769B20 , 32'h0000DD65 , 32'h0F547780 , 32'hFE31CF50 , 32'h0000D8CE , 32'hFFFEE8EE , 32'h04634068 , 32'hFB67D4A8 , 32'hFE3532EC , 32'hF7359A30 , 32'h0001043B , 32'h01E99CE4 , 32'hFDF116B4 , 32'h000024C7 , 32'hFAA45BA0 , 32'h00002515 , 32'hECFCC580 , 32'h0000B27F , 32'hFFFFE3D0 , 32'h00008175 , 32'h0B354030 , 32'hF695C050 , 32'h00568F59 , 32'hFFFDDDC6 , 32'h09481580 , 32'h06D4C270 , 32'h00002CFE , 32'h0001FBE3 , 32'h001C7CEC , 32'h09EEDDA0 , 32'hED07BCC0 , 32'h09158EF0 , 32'h0001D58E , 32'hF7FC16B0 , 32'h00C115E1 , 32'hFFB31436 , 32'hFFFFAA55 , 32'h0216BD68 , 32'hEEE19BA0 , 32'hFB90D290 , 32'h0001AFFE , 32'hFE4E6320 , 32'hFFFC83B4 , 32'h0002EC27 , 32'h03F23C58 , 32'hFF1AD976 , 32'hF71E4CB0 , 32'h1A4272E0 , 32'hFFFFC5FB , 32'hFAD91DE0 , 32'h000160C9 , 32'hF8720CA0 , 32'h02248D78 , 32'h00031F8B , 32'hE2BDF880 , 32'hFB467448 , 32'hF82DBCC8 , 32'hFFFF8569 , 32'h00005687 , 32'hFFFFF077 , 32'hFEE6FE24 , 32'h01EF3C30 , 32'hFFFFF20C , 32'hF39078A0 , 32'h002019B5 , 32'h0000434A , 32'hF945AC70 , 32'h00B280E6 , 32'h000085ED , 32'h059D2438 , 32'h0307B4E0 , 32'h05D7E940 , 32'hFFFFCAF5 , 32'hFFFF348C , 32'hFBDD4398 , 32'hFFFFA5D8 , 32'h01B95CEC , 32'h00019344 , 32'h021FE9D4 , 32'h00072CCF , 32'h000011B6 , 32'h00001B7E , 32'hFFFEB558 , 32'hFFFEAD2C , 32'hF2DC9550 , 32'hFAF70FE0 , 32'h00003306 , 32'hF16B91A0 , 32'h0F27F510 , 32'hFFE73446 , 32'hFFFF57DF , 32'hFF202E30 , 32'h000043EE , 32'h02DDD0CC , 32'h02671D6C , 32'hFFFF45C0 , 32'hFEB2E648 , 32'hFFFFBD02 , 32'h00007CD7 , 32'hFE1F7C14 , 32'hFC2BB900 , 32'hFED35494 , 32'h000062E9 , 32'hFA5433B0 , 32'hFFFF62F6 , 32'hFFFF4095 , 32'h05A46108 , 32'h0001CC56 , 32'h000296F0 , 32'hE1E12320 , 32'hF7DF9DF0 , 32'hFFFF2DF9 , 32'hFFFF4155 , 32'h000135BD , 32'hFFFFE515 , 32'hFFFE976F , 32'hFD917094 , 32'h04E1C220 , 32'h000012F7 , 32'h0000D337 , 32'h1C394880 , 32'h08EC8DF0 , 32'hFFFD4E3D , 32'h00008651 , 32'h0DBF3090 , 32'h0000C9CE , 32'h00011740 , 32'hFE31EAB8 , 32'h000B48C4 , 32'h006F585B , 32'h005E131B , 32'h00035454 , 32'h00013637 , 32'hF9C64520 , 32'h00007E74 , 32'hFFFFB8A4 , 32'h020AD6EC , 32'hFFFE2462 , 32'h0002C442 , 32'h000E9418 , 32'hFFFEC68F , 32'hFFA4FC89 , 32'hFFB1151A , 32'h0003A5E3 , 32'h000025B6 , 32'h00014C70 , 32'h07CAF510 , 32'h09CB93B0 , 32'h00D219B0 , 32'h0ABBC3C0 , 32'hFFFD8B9F , 32'h0A002430 , 32'h0000F42C , 32'hFFFDD7AC , 32'h006B31C4 , 32'hFFB353BA , 32'h0247D3D4 , 32'hFFFE0E96 , 32'hFD148C04 , 32'h009B423B , 32'hFBDCD6D0 , 32'h07ACDCF0 , 32'hFC850B74 , 32'hEE45E540 , 32'h0094DC9B , 32'hFFEF114B , 32'hFFFEFD18 , 32'hFFFF3E27 , 32'h0000C44E , 32'h01DE0480 , 32'hF2A68C90 , 32'hFD0448C4 , 32'h0048154F , 32'h084CCB20 , 32'hFA5674E0 , 32'h0001FB47 , 32'h01AC6F40 , 32'h0A1BAD70 , 32'hFFFEDF90 , 32'h0FA74B90 , 32'h00009001 , 32'hF8FCA280 , 32'h2EF25B40 , 32'hFFFD90D8 , 32'h00001E6A , 32'hFFFE6BEC , 32'hFFFE31C7 , 32'h00025DAC , 32'h00025437 , 32'h06B21AA8 , 32'hF6331D20 , 32'hF481D490 , 32'h024B4990 , 32'h015623E0 , 32'hFDF02EA4 , 32'h000035DD , 32'hFFFFF6F4 , 32'h000151B7 , 32'h0000AE23 , 32'h00002B91 , 32'h021DECD0 , 32'h0C8C12F0 , 32'h0D12B060 , 32'hFFFE211D , 32'h000319FB , 32'h00001211 , 32'hFFFD070F , 32'hFEDF3B50 , 32'h0F31C050 , 32'h0000BED8 , 32'hFFFC1243 , 32'h0001C089 , 32'h248AEF40 , 32'hF8A5FE70 , 32'hF4D0D7D0 , 32'h0002A2B1 , 32'hFFFF50A1 , 32'h0000666C , 32'hFFDC1D5C , 32'h00C67001 , 32'h091BAB50 , 32'hFFFE687D , 32'h00518FB6 , 32'hFFFC89C7 , 32'h016B8EB8 , 32'hFFFECD45 , 32'hF0266450 , 32'h000080B7 , 32'hFFC60FEB , 32'hFC0A27E4 , 32'h121F43C0 , 32'hEC832400 , 32'hFFFDBA36 , 32'h044C7558 , 32'hFE038530 , 32'hFFFEE21C , 32'h0417D180 , 32'h0000AE89 , 32'hFE5B3114 , 32'hFDA3D628 , 32'h09191030 , 32'h0000BE5A , 32'hFFFF91B2 , 32'hF8046E90 , 32'h0002E7B0 , 32'h00C69B1C , 32'h0001003A , 32'hFEDA93E8 , 32'h00014865 , 32'h013E20B8 , 32'hFFFECCE8 , 32'h0001DAB4 , 32'h00029CAE , 32'hFABBB0C8 , 32'h090FB130 , 32'h000060BA , 32'h00014552 , 32'hFFFFEA42 , 32'h0002A400 , 32'h09FF1E30 , 32'h11BE97C0 , 32'h061992D0 , 32'hFAFBECB8 , 32'hFF0470BE , 32'h00000086 , 32'hFFFFAB06 , 32'h00000D1A , 32'hFE9DE5E4 , 32'hFFFD695E , 32'h00011F12 , 32'hFECBBA6C , 32'hE3A87C20 , 32'hFFFF52DF , 32'h03AED228 , 32'h02C2DC80 , 32'hFC7AA62C , 32'h09824580 , 32'h0000D381 , 32'h01F8D504 , 32'hF9568C10 , 32'hFE018F14 , 32'h00023908 , 32'h028EBAB4 , 32'h08F08900 , 32'h064A4068} , 
{32'hFFC86155 , 32'h06A523B8 , 32'hFFFEB4D3 , 32'h0F0A6E40 , 32'h00006EB4 , 32'h0148A134 , 32'h0000EADA , 32'h0000450C , 32'h0000051F , 32'hFFFE41A0 , 32'hFB88DCF8 , 32'h09441DA0 , 32'hF8267BC0 , 32'h0000F63F , 32'hFFFF9511 , 32'h058E7820 , 32'h0000C99E , 32'hF3AEECE0 , 32'hFF580804 , 32'hFFFE8F97 , 32'h0000FE6B , 32'hFE2C8AB8 , 32'hFA209B90 , 32'hFFA43696 , 32'hF5942EF0 , 32'hFFFECF30 , 32'h014B458C , 32'hFFD07FEF , 32'hFFFF8C83 , 32'h080097B0 , 32'h000157F5 , 32'hF71D2600 , 32'hFFFF37CC , 32'hFFFF5185 , 32'hFFFFC24E , 32'h0BABC000 , 32'hFDA6A820 , 32'hF0F882D0 , 32'hFFFEAA28 , 32'h1F114EA0 , 32'hF3312C30 , 32'hFFFE3545 , 32'hFFFDE75C , 32'h040FAFF0 , 32'hFB6B63D0 , 32'h02CC8F80 , 32'hF8976068 , 32'hFFFFC2A0 , 32'h01F63C60 , 32'h04C02AA0 , 32'h00F0E1F3 , 32'h000156F5 , 32'hFD402A50 , 32'h16AB4560 , 32'h015A4A50 , 32'hFFFECA3E , 32'h008AB3CE , 32'hFFFFD0DC , 32'hFFFED326 , 32'hFD8A79F0 , 32'h01522AFC , 32'h034C5404 , 32'hF904D188 , 32'hFFFF41A9 , 32'hE3FAF1E0 , 32'hFFFEFB4C , 32'h01068E94 , 32'hFF80FD17 , 32'hFFFD7934 , 32'h14A818A0 , 32'hF71BE490 , 32'hF1C34700 , 32'h0000E470 , 32'h0000C6CF , 32'hFFFFBDD0 , 32'hFF3B0476 , 32'h01FAE7D0 , 32'hFFFEB151 , 32'hFC649FB8 , 32'h0055CE47 , 32'h00010E2F , 32'hE8105540 , 32'h0C2DC580 , 32'hFFFF61EA , 32'h0955F780 , 32'h0E4A92A0 , 32'hF71E36B0 , 32'hFFFDE2E2 , 32'hFFFE537E , 32'h12D09F40 , 32'h00010FCC , 32'hFD23A1A0 , 32'hFFFECDF6 , 32'hF9B44310 , 32'hFFA0011D , 32'h00046A1B , 32'h000118EA , 32'hFFFEC503 , 32'hFFFEDFD2 , 32'hFBCCA8D0 , 32'hFE663C98 , 32'h0002FFE8 , 32'h045B51E8 , 32'hF6DF71E0 , 32'hFF4C3846 , 32'hFFFE4E43 , 32'hFF887941 , 32'h00020CFF , 32'hFDD2A7D8 , 32'h0153F694 , 32'h0001A0A3 , 32'hE96D8E80 , 32'hFFFEF872 , 32'h00001770 , 32'hFD9A1CE8 , 32'h0117AF48 , 32'h027C581C , 32'hFFFDA377 , 32'h01A91918 , 32'hFFFF3C7E , 32'hFFFF1171 , 32'hF9FFAA50 , 32'hFFFFB7B6 , 32'hFFFE3E93 , 32'hFA4FD520 , 32'h01CEBA58 , 32'hFFFFAF3B , 32'h00047250 , 32'h0001412E , 32'hFFFFC054 , 32'h0000D242 , 32'hFD7628B0 , 32'h081D30C0 , 32'h0000F66F , 32'h0001355E , 32'hF6401C00 , 32'h03AB2674 , 32'h0000AB40 , 32'h000078F2 , 32'hFD33FBF4 , 32'h0000FBE3 , 32'h00010CBA , 32'hFF27E1BC , 32'hFAB9C268 , 32'hFF5CC9CC , 32'hFFA46D37 , 32'hFFFFC762 , 32'hFFFDCC36 , 32'hFF6BDFAA , 32'hFFFEDEA4 , 32'hFFFF35FC , 32'hF7743E60 , 32'h0000C3E6 , 32'h00003CEA , 32'hFB970610 , 32'h0000AB7A , 32'hF938FAA0 , 32'h01317244 , 32'hFFFCF6E3 , 32'hFFFE1B77 , 32'h00008133 , 32'hF46B8B40 , 32'h03C91060 , 32'hF8EFD748 , 32'hF426BCB0 , 32'hFFFFED9B , 32'h08471AA0 , 32'h0000EA9F , 32'hFFFDFA35 , 32'hF5AA0240 , 32'hFB28E978 , 32'hFC081648 , 32'hFFFE34BC , 32'hFFA9E76E , 32'hFD360B38 , 32'hFD8828F0 , 32'h03DB6C04 , 32'hFB34B6A0 , 32'h04FFCE70 , 32'h00486B37 , 32'hFB2E1110 , 32'h00014A02 , 32'h0000A287 , 32'h000139DE , 32'hFC9310A0 , 32'h041E5C70 , 32'h0164A638 , 32'h013671F8 , 32'hFF0FCAF6 , 32'h02DC0F34 , 32'hFFFC3E92 , 32'h09CC0780 , 32'h04E93748 , 32'hFFFFE55A , 32'hF05264A0 , 32'hFFFEB7C3 , 32'hF847CF18 , 32'h0C4984A0 , 32'h00024FAF , 32'hFFFFFD6A , 32'h0002274E , 32'h000152D6 , 32'h0000C2B6 , 32'h0000F37F , 32'h03BA556C , 32'hFFEEB507 , 32'h0FE90CF0 , 32'hF87CAF90 , 32'hF8883AE0 , 32'h002C215B , 32'hFFFD81A2 , 32'h0001B316 , 32'h0000D06A , 32'h00004E5C , 32'h00000249 , 32'h02944814 , 32'hEFC56980 , 32'h1599AB00 , 32'hFFFF2B8C , 32'hFFFED422 , 32'hFFFF3AC4 , 32'h000026EB , 32'hFDA02DD0 , 32'hF6AC2E00 , 32'hFFFFFD7F , 32'hFFFE561A , 32'hFFFE523E , 32'h14F1F6C0 , 32'hF4041A70 , 32'hEF7FD300 , 32'h00011C6D , 32'hFFFFC1EF , 32'h0001BA1B , 32'hFF504DF0 , 32'hFF172106 , 32'h0C5DD240 , 32'hFFFF2A79 , 32'hFEA14A90 , 32'h000184D8 , 32'hF5D62160 , 32'hFFFFF2C3 , 32'h172F07A0 , 32'hFFFF2E5E , 32'h155E6A80 , 32'hEF705F20 , 32'h2187D840 , 32'h12C0AF80 , 32'hFFFF89AE , 32'hF08D0FF0 , 32'hFF176CF3 , 32'h00014ACE , 32'h03B6BD08 , 32'h00014D8A , 32'hFDC164DC , 32'hF2E9E810 , 32'hFB98E440 , 32'h000017D6 , 32'hFFFECF9D , 32'hFF640590 , 32'h0000882B , 32'h0AFAEBF0 , 32'hFFFDF479 , 32'hFF5C1E43 , 32'hFFFC340D , 32'h18F8FF80 , 32'h0000FE82 , 32'hFFFFEE88 , 32'hFFFCFC8A , 32'hF713BFD0 , 32'hF548B0E0 , 32'h00029879 , 32'h000071A5 , 32'h00004941 , 32'h0000E95E , 32'hFE690D9C , 32'hFBAD4168 , 32'hF6A92C70 , 32'h08116190 , 32'h0C5826E0 , 32'hFFFFBC5D , 32'hFFFF48BD , 32'h0000E487 , 32'h01A78CD4 , 32'hFFFFFEE6 , 32'hFFFFC71B , 32'hFB060F48 , 32'h06FD7DB0 , 32'h00010110 , 32'h0AB185F0 , 32'h02E0AB1C , 32'h01B24924 , 32'hF88EB7F0 , 32'h000015C8 , 32'h00497BE8 , 32'h0D607500 , 32'h03BC8C4C , 32'hFFFE21A1 , 32'h0A547F20 , 32'h131AE620 , 32'h0DCA92E0} , 
{32'h04F03ED8 , 32'h0DD8BBD0 , 32'h00015F34 , 32'h0A307440 , 32'hFFFEDDA3 , 32'hFCBC20B8 , 32'hFFFFD68D , 32'h0000AAD9 , 32'hFFFDD0E3 , 32'h00013A73 , 32'hF1A6F970 , 32'h09043120 , 32'h0171FB8C , 32'hFFFFFBC7 , 32'h00011657 , 32'hFE7313D4 , 32'h000113F5 , 32'hED679F80 , 32'hFC16FA78 , 32'h000009D0 , 32'h00005996 , 32'h031B8390 , 32'hF89AE600 , 32'h000F25C0 , 32'h09D47750 , 32'hFFFDD025 , 32'hFD437214 , 32'hFF3BD8C2 , 32'hFFFFB116 , 32'h09AC6110 , 32'h00020B33 , 32'h02630120 , 32'hFFFF9B7C , 32'h00018576 , 32'hFFFEED5E , 32'hF1851190 , 32'hFE85827C , 32'hF3211E30 , 32'hFFFE2633 , 32'hF2602F70 , 32'hECFDE860 , 32'hFFFFB68C , 32'hFFFDC33A , 32'h007480C8 , 32'h02F344A4 , 32'hEC4658C0 , 32'h04F157F0 , 32'h0003CCC8 , 32'hF0581D30 , 32'h08086AE0 , 32'h00114DB4 , 32'h0001E3FA , 32'hFED47100 , 32'hFE216D10 , 32'hFAADA0C8 , 32'hFFFF16DA , 32'hFFBD2189 , 32'h0000B0B7 , 32'hFFFEDED0 , 32'hFFAAB3A2 , 32'hFF45C989 , 32'h04D7ED68 , 32'hFD153214 , 32'hFFFF61E5 , 32'h1EE5AEC0 , 32'hFFFF725E , 32'h03FDF024 , 32'h0128AC9C , 32'hFFFED07B , 32'h0B1C0590 , 32'hFA98F4A0 , 32'h07491750 , 32'h0000004B , 32'h00013475 , 32'h0000B638 , 32'hC8FB9180 , 32'hFDA708B0 , 32'h00023888 , 32'hF7D122A0 , 32'h006512A8 , 32'h000060B3 , 32'h0149A578 , 32'hFB3A2550 , 32'h00008D8C , 32'hFC7C22C8 , 32'h0D083520 , 32'hF0D3D800 , 32'h0000EEF1 , 32'h0000DD49 , 32'h035D7F9C , 32'hFFFFD474 , 32'h0185ABBC , 32'hFFFF554D , 32'h04152B48 , 32'hFE8AFA74 , 32'h00015A3A , 32'h00018380 , 32'h0001D11F , 32'h00009758 , 32'h01DBF16C , 32'h02A2E7C0 , 32'h00014D8B , 32'hF963FA58 , 32'h0B2C3B00 , 32'hFD077288 , 32'hFFFFCA35 , 32'hFF3E36F6 , 32'hFFFEDCD3 , 32'h013646AC , 32'hF4479EC0 , 32'hFFFE60E2 , 32'h062BD538 , 32'h0000EEFE , 32'h00024FE8 , 32'h06EC81D0 , 32'hFC518774 , 32'hFFA54213 , 32'h00026B6B , 32'h0B0DA860 , 32'hFFFF41DE , 32'hFFFE2D6F , 32'h02163ACC , 32'h000153BF , 32'h0002962A , 32'h091AFBC0 , 32'h08D6E6B0 , 32'hFFFFDD44 , 32'h0000A9D8 , 32'hFFFFBE0E , 32'hFFFDED6C , 32'hFFFE9B1B , 32'h0442C268 , 32'h0D5545B0 , 32'h00019F87 , 32'h00017592 , 32'h130917A0 , 32'h02B0E470 , 32'hFFFFA63D , 32'h00017240 , 32'hFBA462D8 , 32'h0000A2F4 , 32'h00012AE6 , 32'hFA9060E0 , 32'h003E4C9B , 32'hFE67D260 , 32'hFF7DE5CD , 32'hFFFFE851 , 32'hFFFF6ACC , 32'h02FFF3F4 , 32'hFFFFC8C0 , 32'hFFFFB12C , 32'h02C5DF70 , 32'hFFFF215D , 32'hFFFEB730 , 32'hEF08A3E0 , 32'h0000A6BA , 32'h075711B0 , 32'h0015EEBA , 32'hFFFFD153 , 32'h000159D3 , 32'hFFFFC1CE , 32'h069423D0 , 32'h03D32644 , 32'hFF455700 , 32'h04D23AE8 , 32'hFFFE8F37 , 32'h020F8CA4 , 32'hFFFE7607 , 32'hFFFF40BD , 32'h0A577F00 , 32'hFF665766 , 32'hFCA8D594 , 32'h0002077A , 32'hE8CC17E0 , 32'hFC6D8F98 , 32'hF85648A8 , 32'h117D0B00 , 32'hF1ED6590 , 32'h0D31B710 , 32'h01795890 , 32'h03F711B0 , 32'h0001D513 , 32'hFFFE8E50 , 32'hFFFDB232 , 32'h001F1B3B , 32'hF9B4A040 , 32'h010C7F84 , 32'h01922C88 , 32'h098B0FF0 , 32'h01043090 , 32'hFFFDBA4E , 32'hF61C90B0 , 32'hFEF6C480 , 32'h0002064D , 32'hF11DC310 , 32'hFFFFBB51 , 32'h0F83FC90 , 32'h05BA80F8 , 32'hFFFF7FB8 , 32'hFFFFE9A4 , 32'h0000D48B , 32'h0000FC0A , 32'h00001FB6 , 32'hFFFE6F22 , 32'hF83A83D8 , 32'hFF438631 , 32'h003C37B3 , 32'hFD6B2A7C , 32'hF56B7E20 , 32'hFD86C3F0 , 32'h0000E90C , 32'h000273FA , 32'h00000B3C , 32'h0000666C , 32'hFFFFAB1C , 32'h0482CF18 , 32'h074F8F00 , 32'h05AC9E48 , 32'hFFFFC2EE , 32'hFFFEF297 , 32'h00019191 , 32'hFFFF1B98 , 32'hFB561450 , 32'hF0BFB740 , 32'h0001F6AA , 32'h0000F263 , 32'hFFFD751D , 32'h1713A760 , 32'h0E82E540 , 32'h03979F20 , 32'hFFFEAFB4 , 32'h0001097D , 32'hFFFE8651 , 32'h0010A114 , 32'h021A8A10 , 32'h02BA7194 , 32'h0001FD86 , 32'h00523735 , 32'h0000FE50 , 32'h01E5E6CC , 32'h0002A84E , 32'h08896460 , 32'hFFFCA038 , 32'hF6E844F0 , 32'hF3EF7540 , 32'hFA0F0188 , 32'hF6D6AB70 , 32'hFFFF5921 , 32'hFE5E2ECC , 32'hFF8FAED6 , 32'hFFFEEEC0 , 32'h096F4EA0 , 32'h00003E88 , 32'h00E6224A , 32'h01694978 , 32'hE5465200 , 32'h0000D304 , 32'hFFFEB629 , 32'h0548C7B8 , 32'hFFFE6ADE , 32'hFC37B81C , 32'h0000B7D7 , 32'hFFF1D110 , 32'hFFFD635D , 32'hF9F89F58 , 32'h00012448 , 32'h0001AEAE , 32'h00019B03 , 32'hFE2F09D8 , 32'h04455D10 , 32'hFFFFCE15 , 32'h000278AC , 32'hFFFF39DF , 32'h000284C2 , 32'hF77D65B0 , 32'h0A538410 , 32'h06120A80 , 32'h0C876410 , 32'h14C61400 , 32'hFFFD4412 , 32'hFFFE17A0 , 32'h0001C229 , 32'hFB1A7130 , 32'hFFFE4CB6 , 32'hFFFFF4BC , 32'hFF9664A9 , 32'h028C31A4 , 32'hFFFF80B0 , 32'h0CBD6CE0 , 32'h02C5E258 , 32'h0277AD00 , 32'hFD7F1710 , 32'hFFFDFC02 , 32'hF6B63C30 , 32'h10616DC0 , 32'hFF3CDB10 , 32'h00018A72 , 32'hE8A3AB60 , 32'hF4A87400 , 32'hF9A353D0} , 
{32'h17019F00 , 32'hFEB95A98 , 32'h0002B7C1 , 32'hF19CD600 , 32'h00012A3B , 32'hFD848D30 , 32'h000157F7 , 32'h00015666 , 32'hFFFFA6C3 , 32'hFFFF8483 , 32'h0869B120 , 32'h0C8ADDA0 , 32'hF96ED338 , 32'hFFFEC3D9 , 32'hFFFE2A68 , 32'hF8763E08 , 32'h0001BC3B , 32'h18854440 , 32'hFD47CA70 , 32'hFFFD7229 , 32'h000245D8 , 32'h01DC0D7C , 32'h05C94040 , 32'hFD002DE4 , 32'h07B9A3B0 , 32'hFFFFB4BA , 32'hFD937D84 , 32'hFEF83B5C , 32'h00012B0A , 32'h027E3368 , 32'hFFFF4F62 , 32'hF7BDEB60 , 32'h0002EB02 , 32'hFFFE83F1 , 32'h00001E7F , 32'h028EB6F4 , 32'h058DED00 , 32'hF1A32830 , 32'hFFFF0517 , 32'hFFCA4359 , 32'hFBD6F3C0 , 32'h0000981F , 32'h0000E062 , 32'h01E69124 , 32'h0BEB79E0 , 32'hF7435C70 , 32'hF254CF20 , 32'h0002CB59 , 32'hF5E40CF0 , 32'h01A25CEC , 32'h000AAD8E , 32'hFFFE7003 , 32'hFE151784 , 32'h0237D470 , 32'h070C66A8 , 32'hFFFF2814 , 32'h00CE6962 , 32'hFFFEACC5 , 32'h000046EB , 32'hFB427E58 , 32'h04183E30 , 32'h02B394E0 , 32'hF7AC66C0 , 32'hFFFF62A9 , 32'h2458E000 , 32'h00020368 , 32'h084C8070 , 32'hFF4DD611 , 32'hFFFE2CCA , 32'hEF22D1A0 , 32'hF714BCF0 , 32'hFFCC76BE , 32'h000023B7 , 32'h00005763 , 32'h0000A0BF , 32'h22DFF380 , 32'hFE70DA4C , 32'hFFFF72C8 , 32'hF4A2AA00 , 32'h007156B3 , 32'h0000ACF0 , 32'hFA09EFD8 , 32'h082FDE10 , 32'hFFFFFDE9 , 32'h0001710D , 32'h06069B88 , 32'h06093950 , 32'h00016114 , 32'h00034C90 , 32'h0BC75E80 , 32'h000042CA , 32'hFD546238 , 32'h000073B5 , 32'h0AAF1450 , 32'hFEBD7520 , 32'hFFFEEEF0 , 32'h000247F8 , 32'hFFFF3267 , 32'h0000F121 , 32'hFFF16621 , 32'hFECD8838 , 32'hFFFDD3E9 , 32'hEC9CA400 , 32'h08EBC8C0 , 32'hF87C03D0 , 32'hFFFDA26C , 32'h003285C5 , 32'h0000A1BB , 32'hFA0DF118 , 32'h118FC860 , 32'h00008F40 , 32'h01C53814 , 32'hFFFFD580 , 32'h00019359 , 32'hFAAF9CD0 , 32'hF4C5C650 , 32'h01D6C320 , 32'h0001A881 , 32'hF57F5690 , 32'h000141AB , 32'hFFFBE9F2 , 32'hF7C06C90 , 32'h000014EF , 32'h0002033D , 32'h1194E540 , 32'hEF212060 , 32'h00012E1C , 32'h00009C19 , 32'h00008247 , 32'h00009F83 , 32'hFFFE7128 , 32'h0070BDA1 , 32'h0AF06AC0 , 32'h0000BE94 , 32'h0000C1C1 , 32'hFA93E2D0 , 32'h00C1E775 , 32'hFFFF603B , 32'hFFFEAA12 , 32'h02856808 , 32'hFFFEBB8A , 32'h00020C7D , 32'hFFDB3FA0 , 32'h0395FB34 , 32'hFD1BF71C , 32'hFDB116F4 , 32'hFFFCA2E5 , 32'h00001CB8 , 32'h05FFB1F8 , 32'hFFFF075E , 32'h000054F8 , 32'h03C43534 , 32'hFFFFD01B , 32'hFFFEECB6 , 32'h04D21778 , 32'hFFFFBA07 , 32'hFF585248 , 32'h010797E0 , 32'h00012EEF , 32'h00010F60 , 32'hFFFE32F7 , 32'h04E4D368 , 32'h013D86CC , 32'hFEA3D1EC , 32'hFD37049C , 32'hFFFEFB30 , 32'hF09E5880 , 32'hFFFF2742 , 32'h00015318 , 32'h000AF9BF , 32'hFFA5EACF , 32'hFC1596D8 , 32'h00026009 , 32'hDEF049C0 , 32'hFDC3E050 , 32'hF8A59A00 , 32'hFF376190 , 32'h0919CCF0 , 32'h1E9C6980 , 32'h02D764F0 , 32'hF266A360 , 32'hFFFF9639 , 32'hFFFFD76D , 32'h00020B9E , 32'h03B3CCA8 , 32'hFA7CB738 , 32'h00C78DF5 , 32'h029C5F14 , 32'hF6A8B510 , 32'hFAD115B8 , 32'hFFFD4536 , 32'hF09F9C40 , 32'h06E4A350 , 32'h0000F0D9 , 32'hFF556047 , 32'hFFFFF2DF , 32'hF5721540 , 32'h05367088 , 32'hFFFD1C2B , 32'hFFFF3F83 , 32'hFFFF5B5E , 32'hFFFF4182 , 32'hFFFFE1A6 , 32'hFFFFDD54 , 32'h068E2C08 , 32'h01A27B70 , 32'h01F2497C , 32'hF648B7D0 , 32'hF5069FB0 , 32'hF2433FB0 , 32'hFFFF3D29 , 32'h0000F3A6 , 32'hFFFFBD8A , 32'hFFFEC152 , 32'h0001BE0D , 32'hFA7D7000 , 32'h07620BF8 , 32'hF305A3E0 , 32'h00004498 , 32'hFFFF10B6 , 32'hFFFFF6A2 , 32'hFFFF47F5 , 32'h031CAD40 , 32'hEA45A5A0 , 32'h0000B74A , 32'hFFFF50E6 , 32'h00008BDB , 32'hFC9FE524 , 32'hFAD2F540 , 32'h0982D6A0 , 32'h000023BA , 32'h00012287 , 32'hFFFFD408 , 32'h003F836C , 32'h03B4FC40 , 32'h015A4FF4 , 32'hFFFFD12A , 32'h0037999E , 32'hFFFF5093 , 32'hF73C66B0 , 32'hFFFDF352 , 32'hFED2E890 , 32'hFFFE9270 , 32'hFB22EC00 , 32'hF36D9A60 , 32'hFCCD941C , 32'h05C82278 , 32'hFFFF6CB3 , 32'h00A9AEC2 , 32'h01075D98 , 32'hFFFF0CBC , 32'h0093EEF1 , 32'h00023496 , 32'hFB6E3EC8 , 32'hE7DCEB00 , 32'h070048B8 , 32'hFFFFE589 , 32'hFFFEF9B1 , 32'h13FE9AC0 , 32'hFFFEBBCC , 32'h0A4CE9F0 , 32'h000090A4 , 32'h00AD0580 , 32'hFFFF362E , 32'hFFD3F606 , 32'hFFFEC9F8 , 32'h00001344 , 32'hFFFF1D52 , 32'h0285A200 , 32'hEBEF64C0 , 32'hFFFDD93F , 32'hFFFF64AE , 32'h00011226 , 32'hFFFDB0E0 , 32'h01FF5E0C , 32'hF0B5A630 , 32'h0611F270 , 32'hEA2A1D00 , 32'h0E6A5120 , 32'hFFFD8623 , 32'hFFFF42EF , 32'h0001190A , 32'hFFE0E59F , 32'h00004B10 , 32'h00025376 , 32'h004A855E , 32'hFD7228F0 , 32'h0001E812 , 32'h0AA51D40 , 32'hFD455DC4 , 32'hFB743770 , 32'hF97B88E0 , 32'h00019C07 , 32'hFD495C54 , 32'hFE290E34 , 32'h00136C25 , 32'h00025D8D , 32'h0EAE5270 , 32'h0A871B20 , 32'hF93BF2F8} , 
{32'hF01673F0 , 32'hF4B16C30 , 32'h00027B2C , 32'h010F6D58 , 32'hFFFF019A , 32'hFD30A368 , 32'hFFFE33C5 , 32'hFFFE7701 , 32'hFFFF7C11 , 32'hFFFFF195 , 32'h0D46B0E0 , 32'h1B91C9E0 , 32'hFC593310 , 32'h0000427D , 32'h000012B2 , 32'hF69F2B20 , 32'hFFFEFBB2 , 32'hFEA49644 , 32'h091A23C0 , 32'hFFFEA2E1 , 32'h00014931 , 32'h00BC45FE , 32'h08EA6540 , 32'h0049F982 , 32'hF20CBF20 , 32'h0000FF21 , 32'h008C8C6E , 32'h014FE8FC , 32'h00000662 , 32'h14AE8CA0 , 32'hFFFFA341 , 32'hFDFA085C , 32'hFFFF307E , 32'hFFFF52AB , 32'h000149F6 , 32'h07E659A0 , 32'h03CB06E4 , 32'hF3B1EB90 , 32'h0002C572 , 32'h0670AA30 , 32'h118C1C00 , 32'hFFFFDA67 , 32'hFFFFD19D , 32'hFF1BB018 , 32'h0CF42050 , 32'hFC156A50 , 32'h09E6FF10 , 32'h00001222 , 32'h055F3980 , 32'h0297CA60 , 32'hFF4E28C3 , 32'hFFFFDAA0 , 32'hFDA6FFCC , 32'h065CC950 , 32'hF2494150 , 32'hFFFDD6BE , 32'hFF6146D9 , 32'h000087B9 , 32'hFFFFC725 , 32'hFAEA6350 , 32'h00790D2C , 32'h03A2FA88 , 32'h0317C908 , 32'h000107D6 , 32'h0205FBB8 , 32'h0001FAAE , 32'hF59CA270 , 32'hFE8CA7B8 , 32'h00004297 , 32'h00C8BB41 , 32'h052AE7A8 , 32'hFEEBB0FC , 32'h00003682 , 32'hFFFDAF4F , 32'hFFFFC63D , 32'h0DCAB420 , 32'h01705FD4 , 32'hFFFE7416 , 32'hE6313F40 , 32'h0122CC60 , 32'h000073A0 , 32'h02D8AF38 , 32'hFF1642A1 , 32'h000026E2 , 32'hF86A2DC0 , 32'h0118747C , 32'h03704768 , 32'hFFFFCB26 , 32'hFFFF7518 , 32'hE2711840 , 32'hFFFFB114 , 32'h01FAF5B4 , 32'h00008EBD , 32'hF8438498 , 32'h000EE30F , 32'hFFFFF8F4 , 32'h0001ADDD , 32'h0000E53D , 32'hFFFE7DD6 , 32'h068A8678 , 32'h007F3A46 , 32'h000150C9 , 32'h04E5D0B8 , 32'hF2379ED0 , 32'h03C21F14 , 32'hFFFFB4BC , 32'h0041C363 , 32'h00008C6A , 32'hFBC9C5C0 , 32'hF9FFC8D0 , 32'h0000B085 , 32'h092D3420 , 32'hFFFF9FA6 , 32'hFFFE02E5 , 32'h0104AEBC , 32'h0023CAB5 , 32'hFF69E4C2 , 32'hFFFF5B66 , 32'hFF3B7342 , 32'hFFFDF882 , 32'hFFFFA4EF , 32'h00F870C3 , 32'hFFFF4F4C , 32'hFFFFD850 , 32'h064B1148 , 32'hF1F53720 , 32'hFFFDAB06 , 32'hFFFE59F9 , 32'hFFFF8A51 , 32'h0000A7AF , 32'hFFFFA17E , 32'hFC883948 , 32'h05A5E2B8 , 32'hFFFFAFAF , 32'hFFFFAC62 , 32'h16011200 , 32'h07D03ED0 , 32'h0000427A , 32'h00006068 , 32'hFA6275F8 , 32'h00008F53 , 32'h00004E75 , 32'h01A1393C , 32'hF6343200 , 32'h017C5D14 , 32'h016815D4 , 32'hFFFECF58 , 32'hFFFDF9FC , 32'hF936AD48 , 32'hFFFFCD66 , 32'hFFFE84DD , 32'h01363A00 , 32'h0000DAB6 , 32'hFFFF29FE , 32'hFE2BD358 , 32'h0003EF4C , 32'hFDD70BDC , 32'hFF2BF262 , 32'hFFFF42F7 , 32'h0000C473 , 32'hFFFF5833 , 32'hF9A53C08 , 32'h00FBCDCC , 32'hFD735C34 , 32'hFA130E80 , 32'hFFFF5507 , 32'h0F823230 , 32'h000163F9 , 32'hFFFFEEE3 , 32'h17949E40 , 32'hF9A1D3A0 , 32'h05721970 , 32'hFFFE9294 , 32'h055BFB28 , 32'h04D69C10 , 32'h07F3ABD8 , 32'hF6ACE9F0 , 32'hF4991C90 , 32'h03F44A98 , 32'h000392EE , 32'hFC058128 , 32'h00005F96 , 32'h000157CA , 32'hFFFF3846 , 32'hFAF1C960 , 32'h05CF4748 , 32'hFE06E3F4 , 32'hFFF03EEA , 32'hF69BD1A0 , 32'h048C0EE0 , 32'h0000AF7E , 32'h0B276E00 , 32'hF992AF78 , 32'hFFFE7044 , 32'hE8A6BEC0 , 32'hFFFE9335 , 32'hF724CE90 , 32'hF9488F18 , 32'h00014BF3 , 32'hFFFEC0A4 , 32'h0002761E , 32'hFFFF929C , 32'h00000FD7 , 32'hFFFF1576 , 32'hF9602FC8 , 32'h0C1E6520 , 32'h12A97AE0 , 32'h096D64F0 , 32'h05142D80 , 32'h0AA11F30 , 32'hFFFDB900 , 32'h0000B5AE , 32'h00006331 , 32'h0002303A , 32'hFFFFACE1 , 32'h01C74B70 , 32'h02078718 , 32'h077576B8 , 32'hFFFE5E88 , 32'h0001998A , 32'h00004425 , 32'hFFFF0911 , 32'h05037A98 , 32'h066FF5E0 , 32'h00005C99 , 32'hFFFFD107 , 32'hFFFFE37F , 32'h0008E293 , 32'h2AF34980 , 32'hF11011C0 , 32'hFFFF313B , 32'hFFFFADC9 , 32'hFFFEABD1 , 32'h029CE210 , 32'h0248C994 , 32'hF02F8D30 , 32'h00003423 , 32'hFE82F3E4 , 32'h000209B1 , 32'hFF61FFC4 , 32'h00007501 , 32'hF6F60970 , 32'hFFFEFD96 , 32'h0E6E3BB0 , 32'h082C04D0 , 32'hEF3C9640 , 32'hFBF8C568 , 32'hFFFDD5D6 , 32'h04E9E250 , 32'h001D74F5 , 32'h0000985B , 32'h0805A260 , 32'h0000A6DE , 32'h00E63DA4 , 32'hFDCCFE44 , 32'hFAD33918 , 32'h0000696A , 32'hFFFEAC01 , 32'hFFF9AA45 , 32'hFFFE9376 , 32'hFB95E708 , 32'h000068AB , 32'hFD6A703C , 32'h0001367F , 32'h0AE03D40 , 32'h00016581 , 32'hFFFE3F05 , 32'hFFFF62A3 , 32'hF2D71F80 , 32'hF9AF0248 , 32'h0000FBCB , 32'h00002AAF , 32'h0001CF38 , 32'h00000563 , 32'hF969D6D0 , 32'hF72AB230 , 32'h015D882C , 32'hE4DC1840 , 32'h05771310 , 32'hFFFEF2B5 , 32'h0000DFB7 , 32'hFFFFCAFE , 32'hFF64448E , 32'hFFFFB7D1 , 32'h0000C1DB , 32'h00913B9C , 32'h05C6FB90 , 32'hFFFF70AE , 32'h25FCF640 , 32'hFE938E50 , 32'hF40096D0 , 32'hF9793650 , 32'h0001213C , 32'hFBCA2160 , 32'hF4916480 , 32'h01240690 , 32'hFFFFAF63 , 32'hF480F570 , 32'h00D1B4F5 , 32'h04249080} , 
{32'hF5D4E4B0 , 32'h0FD1EF80 , 32'h00000090 , 32'hF92AD518 , 32'hFFFF8175 , 32'hFD7083EC , 32'h0000CAD0 , 32'hFFFF9534 , 32'h00020645 , 32'hFFFBE4A8 , 32'hFD878174 , 32'hFCC10130 , 32'hEF226980 , 32'h0001ABFE , 32'h000061C3 , 32'h1737F9C0 , 32'hFFFEBB7F , 32'hF6769AF0 , 32'hFFCDC765 , 32'h00020D81 , 32'hFFFF5808 , 32'hFE3434CC , 32'h06932728 , 32'h070D2308 , 32'h008EB947 , 32'h0002EDB9 , 32'hFFFDEFFB , 32'h027FE84C , 32'hFFFF7274 , 32'h08017190 , 32'h00016E86 , 32'h00004080 , 32'h00030792 , 32'hFFFF689E , 32'h0000A444 , 32'h0C4F1770 , 32'h06E0FA50 , 32'h169B8500 , 32'hFFFF8C9A , 32'hEF49F6A0 , 32'hDD3DBFC0 , 32'h00007157 , 32'h00014004 , 32'h0247DF0C , 32'h101B5780 , 32'hFA8738A0 , 32'h068F1FD8 , 32'hFFFF535F , 32'h0375AE88 , 32'h00DD3418 , 32'h0109DD68 , 32'h0001994C , 32'h00912879 , 32'hFDDCC1A8 , 32'h04E45168 , 32'hFFFD56E8 , 32'h012C7684 , 32'h0000029E , 32'hFFFDF83E , 32'hFEEE02B8 , 32'h0049AE4B , 32'h00D4B36E , 32'hF3CBA460 , 32'hFFFFF4F6 , 32'hF19DCAD0 , 32'h00027DE0 , 32'hF42392D0 , 32'h0742A6C8 , 32'hFFFF45A1 , 32'hF11AF8F0 , 32'hF9D18000 , 32'hFA9D94D0 , 32'h0001737A , 32'h0002E154 , 32'hFFFE8056 , 32'h0A1477A0 , 32'h0045DD6C , 32'hFFFF7FF7 , 32'h0D5E7C50 , 32'h012155D8 , 32'hFFFECACC , 32'hF376BEA0 , 32'h09A75490 , 32'h000256EE , 32'h0116E864 , 32'hF0A61130 , 32'h01299968 , 32'hFFFF5436 , 32'h000214E8 , 32'hF5C953E0 , 32'h00012360 , 32'h02F04880 , 32'hFFFF6F7A , 32'h05EB8D60 , 32'h0021B773 , 32'hFFFD028F , 32'h000002ED , 32'h00003DF6 , 32'hFFFE6F54 , 32'hF8740508 , 32'hFD170760 , 32'h000147E3 , 32'hFB8F3950 , 32'h0061BA37 , 32'hFCEF6CE8 , 32'h00001395 , 32'hFFDF4FC1 , 32'hFFFC12BD , 32'h0680F1B8 , 32'hED839A80 , 32'hFFFE1FC7 , 32'hF46E5340 , 32'h00004265 , 32'h00009F4D , 32'hF7AB9DC0 , 32'h031AFBD0 , 32'h01FD72B4 , 32'h00018321 , 32'h03381C58 , 32'hFFFF5BD3 , 32'h000089F9 , 32'hFC6B02F0 , 32'h00009ABA , 32'hFFFFAB7B , 32'hF45A6110 , 32'hF97253D8 , 32'hFFFF40B1 , 32'h0002FC48 , 32'h00007F55 , 32'hFFFEDF04 , 32'hFFFEDA2C , 32'h0355AA4C , 32'h06F691A8 , 32'hFFFE0325 , 32'hFFFEDED2 , 32'h100AEDC0 , 32'hF78D9110 , 32'h0000D216 , 32'hFFFFB4F6 , 32'hF05F92D0 , 32'hFFFFE567 , 32'hFFFE1CD7 , 32'hFEFA5448 , 32'hF8D295D8 , 32'hFDB0F230 , 32'h01F68044 , 32'h0000E8D2 , 32'h00001C01 , 32'hFC69DB24 , 32'hFFFF8BB7 , 32'hFFFFE8E2 , 32'hFB25AA18 , 32'hFFFE5873 , 32'hFFFDD605 , 32'h0C8837A0 , 32'h00017F66 , 32'hFC0453AC , 32'hFBDA0768 , 32'h0001A966 , 32'hFFFDD59B , 32'hFFFEF6A5 , 32'hF9819F60 , 32'h053E49C8 , 32'h00C75C11 , 32'hF9A49DC8 , 32'h0000844D , 32'hF9C3FAA0 , 32'h00002D49 , 32'hFFFFDC16 , 32'hF990E540 , 32'hFD46FB0C , 32'hFC19FF60 , 32'hFFFFB65B , 32'hECAE69A0 , 32'h00AE1A13 , 32'hFDC3298C , 32'h05AD4990 , 32'h063C31D0 , 32'h0550CAE0 , 32'h0301F678 , 32'hEF0E6E40 , 32'hFFFF426B , 32'hFFFDF5AE , 32'hFFFFFCBB , 32'hF4EC8940 , 32'h004C5B88 , 32'hFA104210 , 32'hFCAC5740 , 32'hEF6B47E0 , 32'h02A6D808 , 32'h0002CEB8 , 32'h0D74B1D0 , 32'h0E07C2C0 , 32'h0000E860 , 32'h09FBE310 , 32'hFFFFFE72 , 32'h06CD5CD0 , 32'hF4820A10 , 32'h00001886 , 32'hFFFF027A , 32'h00017780 , 32'hFFFD4603 , 32'h00017551 , 32'h0000181D , 32'hFAC8F168 , 32'hFC697B78 , 32'hD24D3080 , 32'h01F894AC , 32'hFBD59D48 , 32'hF9F80D98 , 32'hFFFED551 , 32'h0000793F , 32'h0000BD00 , 32'hFFFFEB68 , 32'hFFFF2166 , 32'hFAA7D5B0 , 32'hF8CF6BA0 , 32'hFD24E1B4 , 32'h00004E59 , 32'h00002BF4 , 32'hFFFEB61F , 32'hFFFDD94A , 32'hF8A3EB28 , 32'h05047FF0 , 32'h00000B17 , 32'h0001ED9F , 32'h0000BCB0 , 32'hFCD7BFA0 , 32'h0420A710 , 32'h044578B0 , 32'hFFFDB630 , 32'hFFFD69D3 , 32'h000168FB , 32'h012D5F14 , 32'hFEB318B8 , 32'h01AB0BD8 , 32'hFFFF91CD , 32'hFFFF21E3 , 32'h00024DF2 , 32'hF4A3FDD0 , 32'hFFFD1F7F , 32'hF9C9B138 , 32'hFFFEDE9F , 32'h048080B0 , 32'h00C71975 , 32'h0B933D20 , 32'h02E68A3C , 32'h0000A981 , 32'h02B8D240 , 32'hFE970138 , 32'hFFFD038D , 32'h0077E933 , 32'h00002E1D , 32'hFEB38DB4 , 32'hFD995D24 , 32'hD91C7680 , 32'h00006078 , 32'h000072EE , 32'hF1D14D80 , 32'h0000EBA2 , 32'hEFC64760 , 32'hFFFEB2C1 , 32'h01503934 , 32'h0000068C , 32'hFD1CEE14 , 32'hFFFDD64A , 32'hFFFF112D , 32'hFFFEF38A , 32'hF5BE8E70 , 32'hF2E053C0 , 32'hFFFFF3DA , 32'h0002C111 , 32'hFFFE5758 , 32'hFFFECE42 , 32'hF6211280 , 32'hEF051D00 , 32'hF9AAC470 , 32'hFD2D91D4 , 32'hFF774AD5 , 32'h0000B7E8 , 32'h00005E1D , 32'h000019C8 , 32'hFDCB52C4 , 32'h00014104 , 32'h0004B24F , 32'h00C4429D , 32'hFB071608 , 32'hFFFD0209 , 32'h11AA3980 , 32'h00686B59 , 32'h016CFA34 , 32'h0CDC5310 , 32'hFFFE9821 , 32'hFBE76338 , 32'hEBDBB660 , 32'h0393B9EC , 32'hFFFF1FA9 , 32'hFEF4DB2C , 32'hF175D730 , 32'hFB853A80} , 
{32'hFCE5F05C , 32'hF5852DA0 , 32'hFFFFEBBF , 32'hFAD03F78 , 32'h0000A5BB , 32'h0145EB48 , 32'h00004F54 , 32'h00008489 , 32'h00008365 , 32'hFFFD5C57 , 32'h01D39EC8 , 32'hF9334C40 , 32'h026AA194 , 32'h0002D6DB , 32'hFFFFA07B , 32'hEF4EAC60 , 32'h000020E7 , 32'hD78E82C0 , 32'hF9D9F438 , 32'hFFFE04AF , 32'hFFFE68DD , 32'hFA5DE710 , 32'h0EEC5830 , 32'hFF8F0C1E , 32'hF4A749D0 , 32'hFFFEA57C , 32'hFFFAB8A3 , 32'hFF751B5C , 32'h0000DB18 , 32'h0E6D8570 , 32'hFFFEF008 , 32'hFC97EAE0 , 32'hFFFF2185 , 32'h0000F510 , 32'h00024BB3 , 32'h14B15F40 , 32'hF85AB208 , 32'hEBC0E640 , 32'h000091BA , 32'h019BF4D0 , 32'h0AC5EC00 , 32'h00013F81 , 32'h0001F113 , 32'h02C5D8E0 , 32'hEE0026C0 , 32'h0F23E080 , 32'hFE55D568 , 32'hFFFEA66B , 32'h0CBFFBF0 , 32'hF0EDD330 , 32'hFFD0CAF0 , 32'h00030505 , 32'hFFAB71A4 , 32'hF27F2DB0 , 32'hF6F4FB50 , 32'hFFFEA25E , 32'hFD51C830 , 32'h000014B6 , 32'hFFFE9A21 , 32'h01DFEA30 , 32'h0011A660 , 32'h00626020 , 32'h02C9EF44 , 32'h0001ABC9 , 32'h0E369DD0 , 32'h0000A5AE , 32'hF56E6430 , 32'hFD5D54D0 , 32'hFFFD3032 , 32'hF33BFD60 , 32'hED0B8AA0 , 32'h08710160 , 32'hFFFDC51E , 32'hFFFF7D86 , 32'hFFFF399C , 32'h0457D9D0 , 32'h0216A460 , 32'h00016A51 , 32'hEBAFA960 , 32'h036DE848 , 32'hFFFF2D27 , 32'hF4882400 , 32'hFF8864BC , 32'h000216E1 , 32'h018DB7C0 , 32'hE6049D20 , 32'hFBB32AF0 , 32'hFFFE5C4A , 32'h00023797 , 32'h0E691690 , 32'hFFFD737F , 32'h024AC7C4 , 32'hFFFF2404 , 32'hF7964920 , 32'h00BDE46A , 32'hFFFEA91B , 32'hFFFDBC0E , 32'hFFFE3855 , 32'h00005AE5 , 32'h05E30DE0 , 32'h05508050 , 32'hFFFF1484 , 32'hFB811C20 , 32'hF8D43C50 , 32'h0784D8B8 , 32'hFFFECBBE , 32'hFFDB7DF0 , 32'h0000BE57 , 32'hFDD3F0BC , 32'hF4EAA8B0 , 32'hFFFEA318 , 32'hF48668F0 , 32'hFFFE4951 , 32'h00018BC1 , 32'h0DE488C0 , 32'hFE868368 , 32'h02BE4A80 , 32'hFFFD99D8 , 32'hFA9F37F0 , 32'h0000725E , 32'h000083C0 , 32'h0A064C70 , 32'hFFFFDE47 , 32'hFFFC7221 , 32'h05850998 , 32'h1111B860 , 32'hFFFE9956 , 32'h000027EE , 32'h000171F9 , 32'hFFFFEEFB , 32'hFFFF738C , 32'hFCCC8078 , 32'h069642D0 , 32'hFFFFC353 , 32'h0003AF12 , 32'h03A44314 , 32'h0873FD60 , 32'h000021F0 , 32'h0002BCF2 , 32'hF35E71E0 , 32'hFFFF510D , 32'hFFFE74A0 , 32'h033AA044 , 32'h007B1413 , 32'h022CC168 , 32'h019CAD30 , 32'h000165FA , 32'h00004B08 , 32'hFFE9064C , 32'h0001BC7E , 32'hFFFED2F1 , 32'h02CA95C0 , 32'hFFFEDE76 , 32'h00007811 , 32'h068C83F0 , 32'hFFFF2B62 , 32'hF5603BC0 , 32'h009514D3 , 32'hFFFF9E71 , 32'h00008542 , 32'hFFFFC779 , 32'h0D2FB2A0 , 32'hF4175BC0 , 32'h039BC844 , 32'h14A69E80 , 32'hFFFEC2E8 , 32'hFADEA0E0 , 32'hFFFF53CB , 32'hFFFF5A6C , 32'hF20F6B10 , 32'h08DF6F10 , 32'hFD795D9C , 32'hFFFF40DC , 32'hF8EDAE98 , 32'hFB109F28 , 32'hFFFB6EC7 , 32'hFC36157C , 32'hF5DD6220 , 32'hF89C5E90 , 32'hFFD3794E , 32'h02494108 , 32'h00020F46 , 32'hFFFE3674 , 32'h00001938 , 32'hF987DBB0 , 32'hF3027B10 , 32'hFF4574CC , 32'hFF2AFC82 , 32'h032E399C , 32'hF8BAE410 , 32'hFFFFA8D8 , 32'h0EA98370 , 32'h08223F70 , 32'hFFFDE400 , 32'hF235BF00 , 32'hFFFEE758 , 32'h0BF581A0 , 32'hFCD285E8 , 32'h00010CBC , 32'hFFFE5ED0 , 32'hFFFFF356 , 32'h00002689 , 32'hFFFD1A49 , 32'hFFFEA617 , 32'h007B8B84 , 32'hFCCE265C , 32'hF7406840 , 32'hF7EC7AF0 , 32'hFCA03400 , 32'hF35930C0 , 32'h000039CF , 32'h0001993A , 32'h00019BFD , 32'hFFFF32BC , 32'h0000EB7B , 32'hF9D9D830 , 32'h03C2EDDC , 32'hF3C40840 , 32'hFFFBB278 , 32'hFFFF690C , 32'h0000AADF , 32'h000075F0 , 32'hFB49ABD8 , 32'hFBE16118 , 32'hFFFF4F2F , 32'hFFFF308C , 32'hFFFDDF3A , 32'hF36EC880 , 32'h0021D90F , 32'hF27C8040 , 32'hFFFE3A7B , 32'h00015A41 , 32'hFFFF261B , 32'h01C326A0 , 32'hFCFE19C4 , 32'h00D64E86 , 32'h00012C96 , 32'hFF36F5B8 , 32'hFFFE8513 , 32'h0E34B8B0 , 32'hFFFFDFD0 , 32'h0BB5C650 , 32'hFFFF2275 , 32'h04A6B380 , 32'hF4F631D0 , 32'h02DE2364 , 32'hFCEDEFD0 , 32'h00022EAC , 32'h01DFA5B0 , 32'hFE2F0334 , 32'h00008B77 , 32'hF5D131B0 , 32'h00006FFE , 32'hFE0F3E2C , 32'h03417EFC , 32'hEE78CD20 , 32'hFFFF7996 , 32'h0000A683 , 32'h06D94930 , 32'hFFFF313E , 32'hF749F860 , 32'h000396DA , 32'hFE989294 , 32'h0001E80A , 32'hF8011688 , 32'h0000549D , 32'hFFFFFDB2 , 32'hFFFEF9DA , 32'h17172B80 , 32'h1A31A5E0 , 32'h0002D012 , 32'h0001B418 , 32'h0000566D , 32'h00027247 , 32'h0F453660 , 32'hFCA509B0 , 32'h0834F9F0 , 32'hF76E15A0 , 32'h08A8EDD0 , 32'hFFFF4A18 , 32'h0000D8A5 , 32'h0001E15E , 32'hF8DE8618 , 32'hFFFE39A1 , 32'hFFFED441 , 32'hF98A8838 , 32'hF8B39E18 , 32'hFFFE1AD8 , 32'h01A154C8 , 32'h04110B60 , 32'h02024668 , 32'hF487C6F0 , 32'hFFFDAC75 , 32'h06053BA8 , 32'hF88D7380 , 32'h0097F391 , 32'hFFFDB844 , 32'h1F4A68A0 , 32'h01A5A6E8 , 32'h03509080} , 
{32'hF59A9830 , 32'hF92DE0D8 , 32'hFFFCE6AC , 32'h00FF9F24 , 32'hFFFEC177 , 32'hFE21D0D8 , 32'h00004913 , 32'hFFFDE5C9 , 32'h000019B3 , 32'hFFFFF874 , 32'hFD08E750 , 32'hF0958CB0 , 32'h06A7DE98 , 32'hFFFF23DB , 32'h0003A49A , 32'h0EFBBA70 , 32'hFFFFE4C8 , 32'h19AD3A00 , 32'hF8D96DC8 , 32'h00004E90 , 32'hFFFC4939 , 32'hFF5B906B , 32'hFD9A93B0 , 32'h076D9240 , 32'hFD6C4B8C , 32'hFFFFAA71 , 32'hFFBB16E3 , 32'hFFCCD951 , 32'h00019A23 , 32'h0E29FB40 , 32'h0000167A , 32'hF75A8CA0 , 32'h0000ADDD , 32'h00024723 , 32'hFFFBF290 , 32'h01095114 , 32'h04C210B8 , 32'h047DD8F0 , 32'h0000BE9D , 32'h049FD038 , 32'hF98F8DE8 , 32'h0001A0EE , 32'hFFFFFDCE , 32'hFF436EDE , 32'h114BBD40 , 32'hE8016F80 , 32'hFD971C6C , 32'hFFFF1854 , 32'hFD007A2C , 32'h0B5BBAC0 , 32'hFFEB07AE , 32'hFFFFECDC , 32'hFA76A480 , 32'hF83854C0 , 32'hF838AEB8 , 32'h00006EF2 , 32'h00CC88CB , 32'h000119D5 , 32'hFFFF60CC , 32'hFBCBE4B0 , 32'hFDF9D61C , 32'h051C7F88 , 32'h0369B5D0 , 32'h0001A872 , 32'h034DF248 , 32'hFFFC1F40 , 32'hF3CE5030 , 32'hFF8E9A48 , 32'h0004F122 , 32'h21A59380 , 32'hFB27C1C8 , 32'h068A43F0 , 32'h0000F2B5 , 32'hFFFEE39E , 32'hFFFE5CEC , 32'h09691FE0 , 32'h03CD5EE0 , 32'h0000EE7A , 32'hF9D2C768 , 32'hFEDEADFC , 32'hFFFFFF24 , 32'h07D58E40 , 32'h03E3416C , 32'h00002C86 , 32'hFAB33C40 , 32'h0FF7A2B0 , 32'hFFB6DC6A , 32'h0001BA13 , 32'hFFFC7469 , 32'h03C0E1EC , 32'hFFFF0B5F , 32'h0FF012A0 , 32'hFFFE017D , 32'hF9484278 , 32'h0025EBE9 , 32'h00010238 , 32'hFFFE1587 , 32'h0000ADDA , 32'h0000C395 , 32'h08ADC540 , 32'hFDDC8284 , 32'hFFFFAD46 , 32'h120A5940 , 32'h0021EB8A , 32'h0014F250 , 32'h00011396 , 32'h000B5508 , 32'h000122B9 , 32'h04717D50 , 32'h03C412B8 , 32'hFFFFA539 , 32'hFF9DE69E , 32'h0000A1D8 , 32'hFFFF912F , 32'hFE7D3AA8 , 32'hFFAF804D , 32'hFE785084 , 32'h0000CB30 , 32'h05010F40 , 32'h00004455 , 32'hFFFEBA29 , 32'h06601D70 , 32'h0001159A , 32'h0002173E , 32'h04B42018 , 32'hFD4337F0 , 32'h00008142 , 32'hFFFE6E61 , 32'h00015482 , 32'h00017D5F , 32'hFFFFD3EC , 32'hFEB83964 , 32'h0BB5C030 , 32'h00001F9A , 32'hFFFF6E9C , 32'h094EE700 , 32'h020C53EC , 32'hFFFEEF4D , 32'hFFFD86B5 , 32'h0C5E74E0 , 32'h00030936 , 32'h0000A9C7 , 32'h01E6B1F0 , 32'h01EED324 , 32'h027768FC , 32'h05989A28 , 32'hFFFFFD57 , 32'h00037381 , 32'hFE2F389C , 32'hFFFFC762 , 32'hFFFF6C1F , 32'hFB35E8F8 , 32'h0003D808 , 32'h0001C429 , 32'h07362500 , 32'h00011FAA , 32'h038B764C , 32'h006F38F7 , 32'h0002EE72 , 32'h00022F72 , 32'hFFFF0FFD , 32'h089F7A70 , 32'hFD4E3CFC , 32'hFEF2773C , 32'hF56A60E0 , 32'hFFFD9488 , 32'h099E8D80 , 32'hFFFF9232 , 32'hFFFF0608 , 32'hFD42C2B8 , 32'h04787F38 , 32'hFF1B372F , 32'hFFFF989E , 32'hEF8A9DA0 , 32'hFC179794 , 32'h028FA4BC , 32'h08D618B0 , 32'hE8F91620 , 32'h06444978 , 32'hFE987BEC , 32'h11AC1120 , 32'hFFFF67F9 , 32'hFFFEF413 , 32'hFFFE2C2C , 32'h0290CCA8 , 32'hFDE88160 , 32'hFE04B540 , 32'h05009250 , 32'h05268180 , 32'hFBD2C768 , 32'hFFFE075B , 32'h031816A0 , 32'hFEB66608 , 32'hFFFEB60A , 32'hDFE2E980 , 32'hFFFED236 , 32'hFF879A09 , 32'h0DC45730 , 32'hFFFDD6FA , 32'hFFFFAD08 , 32'h00005350 , 32'h00006FB5 , 32'hFFFF4AF0 , 32'hFFFEFCCA , 32'hFD369E44 , 32'h04E682D8 , 32'hD927D9C0 , 32'hF913D6B8 , 32'hFDD8057C , 32'h0D721CB0 , 32'h0001288B , 32'h0000E3DD , 32'hFFFD7275 , 32'h000288D9 , 32'hFFFFB1DA , 32'hFD074D24 , 32'h0541DB98 , 32'hF80CEE00 , 32'h00012D84 , 32'h00006D44 , 32'hFFFF3EEC , 32'h0000A357 , 32'h03B88150 , 32'h10D826A0 , 32'h0002F21D , 32'h00004114 , 32'hFFFF0F29 , 32'hF33B5B40 , 32'hF2942C10 , 32'hF0E3DDF0 , 32'hFFFE115B , 32'hFFFDFF3D , 32'h0000720D , 32'hFFEFE135 , 32'hFF55AAEB , 32'h075588B0 , 32'hFFFD0D05 , 32'h001D0D0B , 32'hFFFFCB5E , 32'h07A245B8 , 32'h00015A41 , 32'hEE27E800 , 32'hFFFEC318 , 32'hFE1F5D8C , 32'h0088D6FD , 32'hEFCC8F60 , 32'h3176B6C0 , 32'hFFFF8CBF , 32'h06FB4C78 , 32'hFF58B600 , 32'hFFFDAD54 , 32'hFC91F828 , 32'hFFFE5A99 , 32'h02DFE524 , 32'h08D18AD0 , 32'h02DF4A1C , 32'h0002DABD , 32'h00002602 , 32'hFC5FE470 , 32'hFFFEC080 , 32'hFCC1D308 , 32'h0000ECCE , 32'hFF012B3B , 32'hFFFEF6A2 , 32'hFB155A60 , 32'hFFFF90AD , 32'h0000018D , 32'h00001203 , 32'h09880FD0 , 32'h074413C8 , 32'hFFFF04E0 , 32'hFFFF550E , 32'hFFFF7A03 , 32'h0000FA68 , 32'h0C7C93C0 , 32'h03973544 , 32'hFA930EC8 , 32'h03B8822C , 32'hF8DAB1D8 , 32'h0002713E , 32'hFFFF018F , 32'h000287D8 , 32'hFAD84DE0 , 32'hFFFF0C67 , 32'hFFFE22B4 , 32'hFF4DC853 , 32'h02DB9F20 , 32'h0000A399 , 32'hF47340D0 , 32'hFF047F77 , 32'hFE00A6CC , 32'hF57FA440 , 32'h000041D8 , 32'hFBDCC400 , 32'h00D47EDF , 32'hFD5052EC , 32'h0000C7B0 , 32'h0C186670 , 32'h0F72ED00 , 32'hFCFCCAA8} , 
{32'hF7AAD550 , 32'hF7874800 , 32'hFFFF76FB , 32'h01976DF4 , 32'hFFFFAD07 , 32'hFF87AD72 , 32'hFFFF8737 , 32'hFFFF8603 , 32'h000035EC , 32'h000294C4 , 32'hFF6F08FC , 32'hF1E00980 , 32'h02E99830 , 32'h000192F6 , 32'h00011DC0 , 32'hE6F68A60 , 32'h00000243 , 32'h0C7FE4B0 , 32'h0108C280 , 32'hFFFE3BE5 , 32'h00007812 , 32'hFE5B6634 , 32'hF3FF0D30 , 32'hF9FF00C0 , 32'hFC6A1A80 , 32'hFFFF6302 , 32'h00A464D0 , 32'hFF448227 , 32'hFFFFD03D , 32'h07F130C8 , 32'hFFFFDA26 , 32'h0230EEEC , 32'h00018A20 , 32'h0000FB66 , 32'hFFFFC6BB , 32'h0E440390 , 32'hFE3A6DA8 , 32'h01454B88 , 32'hFFFFFA29 , 32'h049B43A0 , 32'hFB2E0778 , 32'h00015483 , 32'hFFFFFEDB , 32'h04BC4D70 , 32'h0C385210 , 32'h19E11D80 , 32'h00455489 , 32'hFFFECA99 , 32'hF6963080 , 32'hFF85C054 , 32'h008ACF75 , 32'hFFFCBFF8 , 32'hFE90E340 , 32'h03923B78 , 32'hF7D26830 , 32'hFFFEF746 , 32'hFD81E7B0 , 32'hFFFE5386 , 32'h0001A5C6 , 32'hFD01A048 , 32'hFF3CD270 , 32'h02280184 , 32'h179C8060 , 32'hFFFD1A4C , 32'h0D9D0C50 , 32'hFFFC20B3 , 32'hF59EDB90 , 32'hFDA196E0 , 32'h00033B61 , 32'h00F14F29 , 32'h12E67BE0 , 32'h0189BBB0 , 32'h00014827 , 32'hFFFFA705 , 32'hFFFF87DC , 32'h11CC81C0 , 32'h00CC9730 , 32'hFFFC24CA , 32'h2EF88080 , 32'hFD12DE44 , 32'hFFFDE1C4 , 32'hEF0C5580 , 32'hFFB0B491 , 32'h0000297C , 32'h04557D68 , 32'hF7B8E510 , 32'h09848000 , 32'hFFFF5F39 , 32'hFFFFB5DC , 32'h09A9C1F0 , 32'hFFFF28B5 , 32'hFBF9C1D8 , 32'h00011542 , 32'h00FA5469 , 32'h00376387 , 32'h0000AAFF , 32'hFFFF687D , 32'hFFFEC4A2 , 32'h00027CC5 , 32'h01D49314 , 32'h022CE0E0 , 32'h0000C6DC , 32'hF6A4BF10 , 32'h05B432C0 , 32'hFFF377BE , 32'h00009C53 , 32'h002B92B5 , 32'h00014E86 , 32'h0BBA6F00 , 32'hF7C477A0 , 32'hFFFF9245 , 32'h030FF208 , 32'h0001EAAA , 32'h00011368 , 32'hF8D3C008 , 32'hFA5D8310 , 32'hFA6E13B0 , 32'hFFFE3B6D , 32'hFD49FD34 , 32'hFFFDB1DF , 32'h00022DC8 , 32'h0131D9A0 , 32'h00023978 , 32'h00009C9F , 32'h162296E0 , 32'hF18AABF0 , 32'hFFFFB76C , 32'hFFFE4267 , 32'h00018578 , 32'h0002030A , 32'h000091FB , 32'hFABEC808 , 32'hF2D34BB0 , 32'hFFFFA7ED , 32'hFFFFE6CF , 32'hFFB0CFC4 , 32'hFEBC4F1C , 32'hFFFFE006 , 32'h0000437D , 32'h06E5CB00 , 32'h0000C698 , 32'hFFFF7BE6 , 32'h020C0494 , 32'hF98DF658 , 32'hFEAA1B04 , 32'hFD837018 , 32'h00001335 , 32'h00004D26 , 32'hFD7129B4 , 32'hFFFF7217 , 32'h000062A3 , 32'hFF095577 , 32'h0000AACA , 32'h00000EBF , 32'h0FDAE790 , 32'h0000248D , 32'h02A91548 , 32'h0211CD54 , 32'h0000C107 , 32'hFFFE6AC5 , 32'h00017892 , 32'hFF42FE69 , 32'h0276DCFC , 32'h05CA7E48 , 32'h09C9C980 , 32'hFFFFF7F0 , 32'h133E6AE0 , 32'h0000ED0B , 32'hFFFDBD82 , 32'hF9B67010 , 32'h03F38710 , 32'h05AC75E0 , 32'hFFFF8E73 , 32'hEE9B67E0 , 32'h08DA9310 , 32'hF40D7480 , 32'h0A3C2860 , 32'hF3B01290 , 32'hF78A9850 , 32'h01416AAC , 32'h07CC73A0 , 32'hFFFF40B2 , 32'h00014DB6 , 32'hFFFF81FF , 32'h01DD4FB4 , 32'h14DE91C0 , 32'hFD0D51FC , 32'hFE362868 , 32'hF7199730 , 32'hFA3013F0 , 32'h000226D3 , 32'h0432CB80 , 32'hFD33B5E0 , 32'h00001AEA , 32'hF1AB2D10 , 32'hFFFD2A6C , 32'hFB52DBE8 , 32'hFD4CECE0 , 32'hFFFD0C5D , 32'hFFFFBAAE , 32'hFFFF5F6D , 32'h0003DA00 , 32'hFFFF68AF , 32'h000127D7 , 32'hFFAE9DDB , 32'hFED15E34 , 32'hF86A12D0 , 32'hFFBCD26C , 32'hFC272654 , 32'hFE88E268 , 32'hFFFFC58E , 32'hFFFED9FD , 32'h00014CE1 , 32'hFFFF5857 , 32'h000227CC , 32'hFE773264 , 32'hFE28D30C , 32'h0732C438 , 32'hFFFFEB96 , 32'h0000AF55 , 32'hFFFF1A48 , 32'h00009826 , 32'h02C006D8 , 32'hFCE6BDD0 , 32'h000123D7 , 32'hFFFD4BDD , 32'hFFFFD0AC , 32'h0BF4D660 , 32'h1E37D020 , 32'h0380E864 , 32'hFFFEF648 , 32'h0001301F , 32'hFFFEC517 , 32'h05A721E0 , 32'hFEF5616C , 32'h1C8C82E0 , 32'hFFFEB435 , 32'h0057ABD3 , 32'h0000D3F9 , 32'hF5CD68E0 , 32'h0000CFA5 , 32'h095710B0 , 32'h0002AFCB , 32'h06E44B18 , 32'hF13266B0 , 32'hF3309E20 , 32'hF4009570 , 32'h0000DB71 , 32'h01281958 , 32'hFF66127C , 32'hFFFCF9BC , 32'hFE8CB678 , 32'hFFFF92A5 , 32'hFE331534 , 32'h0A457DD0 , 32'h04A33F10 , 32'h0000B85B , 32'hFFFEBCAD , 32'h05F49300 , 32'h00010BBC , 32'h02CCF694 , 32'hFFFE5DC5 , 32'h0339FAF4 , 32'h00001296 , 32'h088FC6C0 , 32'h000192EB , 32'h00008AD6 , 32'hFFFFD382 , 32'h0083CCA6 , 32'h014E1EC4 , 32'hFFFF72EC , 32'h0001CC57 , 32'h0000B248 , 32'h0000A984 , 32'hFA259060 , 32'h01C1F0B4 , 32'h04D46DB0 , 32'h16003440 , 32'hF630F3D0 , 32'h000005AF , 32'hFFFFE144 , 32'h00004102 , 32'h01CFBB08 , 32'h0000F1D3 , 32'hFFFFE22A , 32'hFF7461E6 , 32'hFA8DAB70 , 32'h00023696 , 32'h04D72188 , 32'hFFA3718A , 32'h0A0321D0 , 32'hFA9E7340 , 32'hFFFF8639 , 32'hFF9515EF , 32'h1784BE60 , 32'hFECF8FC4 , 32'hFFFD8064 , 32'h07CFEB28 , 32'hE595B5E0 , 32'h081482C0} , 
{32'hD2B1AF40 , 32'hF65C0EB0 , 32'h00015FCF , 32'hFBBD6060 , 32'h00007060 , 32'hFE7DF808 , 32'h0001E249 , 32'hFFFF2993 , 32'hFFFF1795 , 32'h0001646D , 32'hFE2B78D4 , 32'hF41D90E0 , 32'h07F5EEB0 , 32'h0001C5CB , 32'hFFFDBA6D , 32'hFF49C23B , 32'h0000E871 , 32'hFCCD7704 , 32'hFEE69FD4 , 32'hFFFDE62B , 32'h000227B3 , 32'hFE819684 , 32'hFE01A804 , 32'h0084A5AF , 32'h01453088 , 32'h0000A60C , 32'hFD70AC54 , 32'hFFE79F21 , 32'h00009A8F , 32'hF9486968 , 32'h0000DE78 , 32'h03EB92FC , 32'h0000A5C3 , 32'hFFFF909F , 32'hFFFF6C25 , 32'hEE6910E0 , 32'h0CB3B960 , 32'hF84823C8 , 32'h00017679 , 32'h0CFD7700 , 32'h00BA50A8 , 32'h00006119 , 32'h0000B795 , 32'hFC3FFDE8 , 32'hF9E4C0C0 , 32'hD9B92000 , 32'hFF1C0DBC , 32'h0000705F , 32'hF6C86180 , 32'h0867CCC0 , 32'h00C3AF25 , 32'h0003908A , 32'h01D51574 , 32'hF49C5470 , 32'h08857EA0 , 32'hFFFF3149 , 32'h0024BA1D , 32'h0003630A , 32'hFFFD91D7 , 32'hFEF57190 , 32'h03C50D50 , 32'hFBDDB598 , 32'hFD611458 , 32'hFFFD4DF6 , 32'hF2B7D8E0 , 32'h0000EB18 , 32'h198850E0 , 32'h0194451C , 32'h000025B8 , 32'hFBD83E50 , 32'hF05AB8C0 , 32'h06A4DCC8 , 32'hFFFED948 , 32'h0001894B , 32'h0000C074 , 32'h06DE75D8 , 32'h00A740AF , 32'h00015FC9 , 32'hE9BFA220 , 32'h019886E8 , 32'h00014720 , 32'hD5EBC640 , 32'hFBCA2868 , 32'hFFFF4D50 , 32'h05E7F8E0 , 32'h00306BA1 , 32'hFE0910E8 , 32'h000238EE , 32'h0000E40F , 32'h0393D388 , 32'hFFFF9943 , 32'hFD4FD940 , 32'h00005C3E , 32'h0714BFA8 , 32'hFF6A66F9 , 32'hFFFE92C0 , 32'h0001151B , 32'hFFFF515B , 32'h00010874 , 32'hFB28CA70 , 32'h01DAC13C , 32'hFFFEE600 , 32'hF78D2170 , 32'hF292DE80 , 32'hFB1FAF78 , 32'h0000A46A , 32'h0054AE82 , 32'h000102F5 , 32'h0318A428 , 32'h0BFAD750 , 32'h00015078 , 32'h0AE4F640 , 32'h000249D3 , 32'hFFFF827A , 32'hFD370BA4 , 32'hFF38B44C , 32'h00E65400 , 32'h00017328 , 32'h01D12348 , 32'h0002938A , 32'hFFFE3A5D , 32'hFE1977CC , 32'hFFFF640D , 32'hFFFE65DC , 32'hFF925D5A , 32'hF8A1BAE0 , 32'h0002740B , 32'h0000A3B4 , 32'h0001BBAC , 32'hFFFE5774 , 32'hFFFEE170 , 32'hFFEF570B , 32'h07219288 , 32'hFFFF77BA , 32'hFFFE6D84 , 32'hF27A9E60 , 32'hFDF48E74 , 32'hFFFF6235 , 32'h0002D5C1 , 32'hFCB21FF8 , 32'h0001E639 , 32'h00020A9F , 32'h01D03DD4 , 32'hEC3AC920 , 32'hFC6B7E38 , 32'hFFB366A1 , 32'hFFFF56CC , 32'hFFFECF91 , 32'h020E2318 , 32'hFFFFB2C5 , 32'hFFFCB6E4 , 32'h0319AE68 , 32'hFFFFF45A , 32'h00016906 , 32'hFD5051F4 , 32'hFFFFE35E , 32'h071E0628 , 32'h025ABA90 , 32'h0001AD4E , 32'hFFFE448B , 32'h00000F95 , 32'h0BD9E400 , 32'hFFAA5DF1 , 32'hFFEBB052 , 32'hFF89D1CA , 32'hFFFF3A5F , 32'hF96D41B0 , 32'hFFFC8599 , 32'h00001FB1 , 32'hFDE765FC , 32'hFD4546B4 , 32'h00089A0B , 32'hFFFF260A , 32'hF9593B80 , 32'hFF815996 , 32'h04BBF9C8 , 32'h08C4C020 , 32'h06E868D0 , 32'hF7EC93E0 , 32'h00BE0C4B , 32'h08C8E9C0 , 32'hFFFECD07 , 32'hFFFF9813 , 32'h00013026 , 32'hFC2D139C , 32'hFF33900E , 32'h01DAE1EC , 32'h0105A850 , 32'hFB5D7B60 , 32'h00FE5EFD , 32'h00001EC8 , 32'hF41F4480 , 32'h09CB8600 , 32'h0001A482 , 32'hFD7D4C34 , 32'h00002D87 , 32'h0309960C , 32'hEE600300 , 32'h000039E0 , 32'hFFFEDB5D , 32'h00005DB9 , 32'h000110B1 , 32'hFFFEA526 , 32'hFFFEA27F , 32'hF1BDE740 , 32'h0BF7D8E0 , 32'h0350704C , 32'hF655E440 , 32'hF4C7A380 , 32'hFD2FF8A8 , 32'hFFFFC988 , 32'hFFFFDDA9 , 32'hFFFDC54B , 32'hFFFFB9FE , 32'h00026F4C , 32'hFD964C40 , 32'h043A0DD0 , 32'hFD482A00 , 32'hFFFFD774 , 32'hFFFEE237 , 32'h00013D92 , 32'h0000A511 , 32'hFE8E7384 , 32'hF90CC2C8 , 32'h00010770 , 32'hFFFEF41F , 32'h0000CC27 , 32'h04764DB8 , 32'h13CB4680 , 32'hE7F787C0 , 32'hFFFE0F15 , 32'h0001730E , 32'hFFFEC7BC , 32'hFBA3FB08 , 32'h00C1AA4B , 32'hFC358A8C , 32'h00014F0B , 32'h00A11D43 , 32'hFFFC1FAC , 32'hF1906C40 , 32'h00004E73 , 32'hFAD7CCE8 , 32'h00002D04 , 32'h06BC5B88 , 32'hFD6A6158 , 32'h023C607C , 32'hEDCE5F40 , 32'h0000B63F , 32'hFED99DB8 , 32'h00746E5F , 32'hFFFF3F60 , 32'hFF12AEE2 , 32'h00013E40 , 32'hFD25F9D4 , 32'hFAD7C558 , 32'h0A996740 , 32'hFFFD39A3 , 32'h000049F2 , 32'hF6732BD0 , 32'hFFFF78E7 , 32'hEB0AE560 , 32'h000003A7 , 32'hFED19AEC , 32'h000095A3 , 32'h00DC882D , 32'h0000E62B , 32'hFFFF5E28 , 32'hFFFF2FDA , 32'hFC72151C , 32'hFD5D7BDC , 32'h00004E52 , 32'h00029578 , 32'h00003416 , 32'h0000A262 , 32'h001911E7 , 32'hF94E9AA0 , 32'h097A72E0 , 32'h07EDA238 , 32'hE35F31C0 , 32'h0000B2DC , 32'hFFFFDD8C , 32'h0000E335 , 32'h01945B14 , 32'h000145A1 , 32'h0001065D , 32'hFFF64D7B , 32'hFEBD8D78 , 32'h00020553 , 32'hE560A840 , 32'hFF94F84E , 32'hFB31D120 , 32'hFC5B290C , 32'hFFFF12D2 , 32'hFD07D584 , 32'h081756A0 , 32'hFE1CD6FC , 32'h00020138 , 32'h0508B340 , 32'hF14F19E0 , 32'hF5702E50} , 
{32'h17E4B280 , 32'h0CF71230 , 32'hFFFF7707 , 32'h07D3CE18 , 32'hFFFED64C , 32'hFF89A8B8 , 32'hFFFF7AF8 , 32'hFFFEBC3B , 32'h0001097B , 32'h000055A2 , 32'h0D8560B0 , 32'hFF14774D , 32'h0673D400 , 32'h0000CF88 , 32'h00026DB8 , 32'h06D35B50 , 32'hFFFEFCD3 , 32'h15F982E0 , 32'hFFD73B76 , 32'hFFFED8AA , 32'h0001BB2F , 32'hFDDB4A90 , 32'hF5A20270 , 32'h05AA5768 , 32'hFBA815F8 , 32'hFFFEC2F4 , 32'hFF46E6DE , 32'hFE088B10 , 32'h0001EF18 , 32'hF8128EC0 , 32'hFFFF3409 , 32'hFBB9F6D8 , 32'hFFFF7D1D , 32'h0000EAF3 , 32'h00030BD1 , 32'hF9BC0AF0 , 32'h0ADC84A0 , 32'h130D6960 , 32'hFFFEE01A , 32'hFBAF0F88 , 32'h0F69BEF0 , 32'h0001C16C , 32'h0000FA2C , 32'hFE496BF0 , 32'hF9E8B528 , 32'h0D595C80 , 32'hFD8C0C78 , 32'h00029777 , 32'hF6EC92D0 , 32'h08FCBF80 , 32'h00154204 , 32'h0000B1F4 , 32'h002C2FD7 , 32'hE8151720 , 32'hFF102155 , 32'h0000A011 , 32'hFB9EFBE0 , 32'h00005938 , 32'hFFFEC682 , 32'hFFEBAE4D , 32'h02031BC8 , 32'hFFF5C7B4 , 32'hFFB1DC53 , 32'h0000A4DF , 32'hF87A7BF0 , 32'h00010F87 , 32'hFE0BAA40 , 32'hFCA3F85C , 32'hFFFF57AF , 32'h062581A0 , 32'hF2DF1AA0 , 32'h034716CC , 32'h00019D0F , 32'hFFFFEEA6 , 32'hFFFDDBF3 , 32'h0BB31B20 , 32'hF9121900 , 32'hFFFD63B1 , 32'hE85F3700 , 32'h0167F7A8 , 32'hFFFF6D0F , 32'h0C1DB7B0 , 32'hFC0F9C80 , 32'h0001EA69 , 32'h03E9CCDC , 32'h12FC70E0 , 32'h027B03A8 , 32'hFFFFC796 , 32'h00009644 , 32'h0DC57020 , 32'h0002EA39 , 32'h0665F6B0 , 32'hFFFEF171 , 32'hFD3C0138 , 32'h0025BBE7 , 32'h0000114A , 32'h000083DE , 32'h00019133 , 32'h0000253F , 32'hFE286438 , 32'hFD0ED744 , 32'hFFFFE6C8 , 32'hF8F5C820 , 32'hF192AAE0 , 32'hFD450560 , 32'h0000162A , 32'h009B38CF , 32'h00014615 , 32'hFE614EF4 , 32'hECEABD20 , 32'hFFFCE0F6 , 32'h165FFDE0 , 32'h00014430 , 32'hFFFFDF2A , 32'h11718D00 , 32'hFBCE48D8 , 32'h024FFCD4 , 32'h00019F9D , 32'h09412790 , 32'hFFFFB904 , 32'h00016043 , 32'h095C5300 , 32'hFFFFA81F , 32'h00012A90 , 32'hFC17832C , 32'hF2658800 , 32'h000087FD , 32'h00020D28 , 32'h0001247B , 32'h00024909 , 32'hFFFD9ABC , 32'h01DF00BC , 32'h04B51C40 , 32'h00029CD5 , 32'hFFFF8514 , 32'hF07D82A0 , 32'h028B29FC , 32'h00000574 , 32'h00006ABA , 32'hFABFC320 , 32'h0000BA50 , 32'h00013DEA , 32'hFD6D8D8C , 32'h07101350 , 32'hFD734FCC , 32'h017669A0 , 32'h00000E0B , 32'hFFFEC7A8 , 32'hFDBC18F4 , 32'hFFFF5E15 , 32'h000171EB , 32'h019C8648 , 32'hFFFDCEEE , 32'h000139D9 , 32'hECFA3B00 , 32'hFFFA8AB2 , 32'h01311098 , 32'hFE124E8C , 32'hFFFF3EFF , 32'h000093A9 , 32'hFFFEA2DC , 32'h08599B40 , 32'hFB8AA5D0 , 32'hFF7B8542 , 32'hFB20C720 , 32'hFFFEFB8D , 32'h06236140 , 32'hFFFDB5BA , 32'hFFFFEEF9 , 32'h00FF7A10 , 32'h04CCF2D8 , 32'h0095611C , 32'hFFFFB4FA , 32'hFFE4DC48 , 32'hFFC56C8C , 32'hFB61CF30 , 32'hFD89CC20 , 32'hF3F0BFB0 , 32'hF926E348 , 32'hFF6D8BD3 , 32'hFCAC7A58 , 32'hFFFE7034 , 32'h000010AE , 32'hFFFF20A4 , 32'h00FE2A91 , 32'hFFC44B4B , 32'h040D7C80 , 32'h032F0BA8 , 32'hFEC0B8C4 , 32'h00B58C6B , 32'hFFFB5470 , 32'h0C54FC60 , 32'h06C097F0 , 32'h000034E8 , 32'h14A4F4C0 , 32'hFFFF13B9 , 32'hF7A12BF0 , 32'hF70224B0 , 32'h000148DF , 32'hFFFE07F0 , 32'h0000D6C0 , 32'h00009874 , 32'h00002A05 , 32'hFFFF6FDF , 32'h047E2D58 , 32'h0C5B7A20 , 32'hEA53AE80 , 32'hF3FAFB30 , 32'h082ADC30 , 32'h06E362E0 , 32'h00000F67 , 32'h0001318C , 32'hFFFF1B06 , 32'h00006797 , 32'hFFFFC566 , 32'h03D11B80 , 32'h0002DF45 , 32'h17DC3EA0 , 32'hFFFE91F6 , 32'h00014358 , 32'h00013DAD , 32'h000112B1 , 32'h01DAC530 , 32'h05C4E1F8 , 32'h00002BEA , 32'h000309D0 , 32'hFFFFDF96 , 32'hF550C100 , 32'h19D843E0 , 32'hFA82EB78 , 32'hFFFD8C1D , 32'hFFFDE972 , 32'h00001310 , 32'hFF4893C8 , 32'hF887A8C8 , 32'h162650E0 , 32'hFFFF986A , 32'hFF3F8929 , 32'h000147DE , 32'hEF4BB820 , 32'h0000B3BA , 32'h1744AD40 , 32'h00008DA5 , 32'hFED20ECC , 32'h06CAE770 , 32'h1BD99120 , 32'hF0F77A80 , 32'hFFFE1318 , 32'h00566E65 , 32'h01197B34 , 32'hFFFE60C1 , 32'h077B67B8 , 32'hFFFDAF84 , 32'h02BFE7B4 , 32'h050F38A0 , 32'hFD151AD0 , 32'hFFFF7F39 , 32'hFFFEE24E , 32'hFFFA26A9 , 32'h0000EF1E , 32'h05EB7C20 , 32'hFFFD89B1 , 32'h00C7A1D6 , 32'h0001618E , 32'hF507BBE0 , 32'h0001D453 , 32'h0000EBA1 , 32'h0000A5CD , 32'h12D8C7C0 , 32'h0A92C8C0 , 32'hFFFEBFD7 , 32'hFFFFF85F , 32'h0001C87E , 32'hFFFE96F4 , 32'hF80E30D0 , 32'hF8566050 , 32'h081E8410 , 32'h070B1490 , 32'h0D9F65F0 , 32'hFFFE2EC2 , 32'h00019BFA , 32'h00002C50 , 32'hFD96E9EC , 32'h0001DFC0 , 32'h000197D8 , 32'hFC6E05FC , 32'h13D6AD40 , 32'h000156A3 , 32'h0E1FB7D0 , 32'hFCC2E7F4 , 32'hFC91D14C , 32'hFAB3A190 , 32'hFFFF8D76 , 32'hF923F1F8 , 32'h01502E94 , 32'h01A59BF8 , 32'h0002F413 , 32'h0C258DD0 , 32'hFC45D844 , 32'hEB38A760} , 
{32'hEBA33EE0 , 32'hF6063130 , 32'h00006A4A , 32'hF69057C0 , 32'h00010E75 , 32'h0101A644 , 32'h0002C806 , 32'hFFFCA747 , 32'h000051F1 , 32'hFFFF934F , 32'hFF1DCA0B , 32'hF9654188 , 32'hF619A400 , 32'hFFFBE7C4 , 32'hFFFDE102 , 32'hF86DE1B8 , 32'hFFFDA966 , 32'h07B49210 , 32'hF8BAA0B0 , 32'h0000C271 , 32'hFFFFAC31 , 32'h01DB8C3C , 32'hF597CD90 , 32'hFA322E98 , 32'h0CF8AD70 , 32'h000024FF , 32'h01D8C398 , 32'h00543A56 , 32'hFFFEE77A , 32'h0AE6DAF0 , 32'h0001BAD0 , 32'h0A59DD10 , 32'hFFFFFF6D , 32'h00003FC7 , 32'hFFFF755A , 32'h03432758 , 32'h082ACE30 , 32'h04DA6498 , 32'hFFFFF9FE , 32'hFEC20098 , 32'hFF9645A3 , 32'h0000A8A0 , 32'hFFFFA8AF , 32'hFDC8FF98 , 32'h02AD0E84 , 32'h12794680 , 32'h01FE5978 , 32'h0001753B , 32'hFCCA3508 , 32'h07C9EB30 , 32'hFF22E516 , 32'hFFFBBC3A , 32'hFAED96C0 , 32'hFE2FE8F4 , 32'hFE88CBBC , 32'h00004BC1 , 32'h02A8D820 , 32'h0002A0B5 , 32'h00008F00 , 32'h0403A448 , 32'h00BC5D8F , 32'h028C169C , 32'hF5BADB00 , 32'hFFFEF8D8 , 32'h09185A60 , 32'h0000A81D , 32'hF5F4ABC0 , 32'h0207E4C0 , 32'hFFFFE1B3 , 32'hD4E11B40 , 32'hFC38CC40 , 32'h01386A58 , 32'hFFFF25C6 , 32'h0003DCEB , 32'hFFFD42C7 , 32'hF0F00320 , 32'h0351FD68 , 32'h00015591 , 32'hFFEE7DEB , 32'h00CD6B6F , 32'h000064CB , 32'h0456F0A8 , 32'h06FC5600 , 32'h00009BB7 , 32'hF95BF720 , 32'hFE82BCF0 , 32'h001F4E0C , 32'h0001D15A , 32'h00005259 , 32'h0B9705D0 , 32'hFFFBF94E , 32'h040C5C10 , 32'h0000DBAD , 32'hFE71A190 , 32'h00303BB8 , 32'hFFFD902A , 32'hFFFF14C6 , 32'hFFFF25E6 , 32'h0000BE3C , 32'h03005F58 , 32'hFCBB7E6C , 32'h0000DCAE , 32'hF572D4C0 , 32'hDFD20E80 , 32'h019100D8 , 32'h0000B0C9 , 32'hFF78A4AE , 32'hFFFFEDBD , 32'h02279CA0 , 32'h0C1ABA10 , 32'h0000E864 , 32'h0A74B3F0 , 32'hFFFFD6D7 , 32'h0001839D , 32'h0B4E2A10 , 32'hFF9C1C4F , 32'h02A19FCC , 32'h0000E014 , 32'h03168250 , 32'h0000C0B8 , 32'h000337CE , 32'h009FC490 , 32'h00007C9C , 32'hFFFD430B , 32'hEF2764C0 , 32'hFD80BF68 , 32'h0001BE4A , 32'hFFFEA8B4 , 32'h00000E30 , 32'hFFFE1CAB , 32'hFFFECFCB , 32'h0084AA23 , 32'hFBECE910 , 32'h00014186 , 32'h0002556E , 32'hEADB51E0 , 32'hF20CC310 , 32'hFFFEBD89 , 32'h00000426 , 32'h05C2E3B0 , 32'hFFFFD04E , 32'hFFFD49F4 , 32'h01DA24A8 , 32'hFCA45700 , 32'hFF8FE4F0 , 32'h03993A88 , 32'h000026F7 , 32'h000099E9 , 32'h00303A3E , 32'h000107E2 , 32'h0002F558 , 32'h01C93E58 , 32'h0000DC74 , 32'h0000A35C , 32'hF2AD7F20 , 32'h00014462 , 32'hFE942520 , 32'h01AAA144 , 32'hFFFD88BE , 32'h000194BE , 32'h0001DA02 , 32'hFD57DF24 , 32'h01D0E2DC , 32'h021976BC , 32'hFE5EA390 , 32'hFFFDCB6C , 32'hF4793710 , 32'hFFFE0BAE , 32'hFFFED369 , 32'h00BC0AA5 , 32'h0335F040 , 32'hF8E71C20 , 32'hFFFFF5AF , 32'h16C512C0 , 32'hFD3B5360 , 32'h07837250 , 32'h0538C7C8 , 32'hF1D506D0 , 32'h07813548 , 32'h01DF1A3C , 32'hED167BC0 , 32'hFFFF9DCD , 32'h00011361 , 32'h00005492 , 32'h03EDC828 , 32'hEFBD0F60 , 32'hFDB8AAA4 , 32'h00BDED48 , 32'h04054B98 , 32'h0084BE53 , 32'h0003A2B5 , 32'hFC4AADA4 , 32'hFD40B34C , 32'h00002C45 , 32'hE9481360 , 32'hFFFFA2CB , 32'h00B4F3F2 , 32'h0F6AB270 , 32'hFFFEABE2 , 32'hFFFF061F , 32'hFFFFECA2 , 32'h000050A1 , 32'h0000D227 , 32'h000105E8 , 32'h01C0B5E4 , 32'h17E8F4C0 , 32'hFB1D8EB0 , 32'hFF3A3AFA , 32'h01BD6AF8 , 32'hED36F980 , 32'h00003CF7 , 32'hFFFF978D , 32'hFFFFC63C , 32'h0001B314 , 32'hFFFF20F2 , 32'h00322D97 , 32'hF5896910 , 32'h00B876C2 , 32'hFFFFE31A , 32'h00009C76 , 32'hFFFEDFA2 , 32'h00012287 , 32'h03F1D040 , 32'hEB6C0100 , 32'hFFFFA41F , 32'hFFFCE0FD , 32'h0002A6D7 , 32'h078944E0 , 32'hF1369670 , 32'hFA9B8508 , 32'h00006F55 , 32'hFFFF9109 , 32'h00002B1A , 32'h017AFDC8 , 32'h00CD5DD2 , 32'h00F1EFA6 , 32'h00004989 , 32'h002A5EEF , 32'hFFFE36A9 , 32'hED2FA9A0 , 32'hFFFFBB1A , 32'hF6148FD0 , 32'h00012CA6 , 32'h018A2734 , 32'hFEEA246C , 32'h03623F20 , 32'h1684B920 , 32'h0002896B , 32'h030499B8 , 32'hFE60D850 , 32'h000051D3 , 32'hFE14ACEC , 32'hFFFFBC13 , 32'h04729CF8 , 32'h1BD8C240 , 32'h075AF628 , 32'h0000FE20 , 32'hFFFEC689 , 32'h0A790CD0 , 32'h000001FB , 32'h02F94798 , 32'h00006245 , 32'h0141A1C4 , 32'h0000D522 , 32'hFB071C98 , 32'hFFFF982A , 32'h00002F77 , 32'hFFFEFC2D , 32'hFDCD909C , 32'h07E5E550 , 32'h00001E41 , 32'hFFFFDC7C , 32'h00019B78 , 32'hFFFF9EB9 , 32'hFB5B7080 , 32'h0B922A20 , 32'hF0D49D60 , 32'h039B197C , 32'hE87DF600 , 32'hFFFE5B81 , 32'hFFFE28B3 , 32'hFFFFAC42 , 32'hFE5976C8 , 32'hFFFE735E , 32'hFFFE1AA3 , 32'hFD984A00 , 32'h00E895C2 , 32'hFFFF7641 , 32'h22F39B80 , 32'hFE1BFEDC , 32'h08609410 , 32'h04FE1F38 , 32'hFFFE8258 , 32'h04775D70 , 32'h029DF174 , 32'hFFD96AB5 , 32'hFFFD81D2 , 32'hF40BC310 , 32'hFAFC68A8 , 32'hFA671A28} , 
{32'h029DA078 , 32'h068FC000 , 32'h00017A93 , 32'h07715940 , 32'h000099A8 , 32'hFCB3BCC0 , 32'hFFFE581D , 32'hFFFF02B9 , 32'hFFFE2BED , 32'h0001412A , 32'hF3DE6610 , 32'h02303F88 , 32'hFDEAED80 , 32'hFFFE1127 , 32'h0000DAE9 , 32'hF7630270 , 32'h0001EB36 , 32'h01C318F0 , 32'h05AD9448 , 32'hFFFF9DB9 , 32'h0000DEBE , 32'hFE5FC1B4 , 32'h148E1E00 , 32'hFC3653E0 , 32'h004B5D73 , 32'h00006B1C , 32'h0102DC40 , 32'h015B28DC , 32'h000217CC , 32'hF6C0D7A0 , 32'hFFFF7D6C , 32'h01C6FE3C , 32'h00037619 , 32'h0000B31F , 32'h0001D83D , 32'hD325F080 , 32'h0D9A4420 , 32'hFC48253C , 32'hFFFF2D34 , 32'h033FF918 , 32'h01C1D024 , 32'hFFFECC17 , 32'h0000A4E0 , 32'h024BBCB0 , 32'h20CF5000 , 32'h1AFBF3E0 , 32'hF9E613C0 , 32'hFFFE34F9 , 32'h0081F2F9 , 32'h0C328F30 , 32'h00391EEA , 32'h00029E4C , 32'h0512B720 , 32'h010D6A68 , 32'h03CABA78 , 32'hFFFEE1A3 , 32'hFE1F41D0 , 32'hFFFC2449 , 32'h0000D3CC , 32'hFDD734D4 , 32'h015CA074 , 32'hFB48F388 , 32'h05084960 , 32'h00001DE6 , 32'hE03160E0 , 32'h00022424 , 32'hFA2D3E18 , 32'h0045A48D , 32'hFFFF1B2D , 32'hF2FEEF80 , 32'h0128AC04 , 32'hEEF4C780 , 32'h0001288B , 32'hFFFEB552 , 32'hFFFDF707 , 32'hF3513B60 , 32'h00B99875 , 32'hFFFF338C , 32'hE20B1C80 , 32'h00ECAFA0 , 32'h00012441 , 32'hF2A71C20 , 32'hF0271C70 , 32'hFFFE2B31 , 32'h011AB650 , 32'h00E0FA51 , 32'hFF2C5B9D , 32'h000031FC , 32'h00020CCF , 32'h051E69E8 , 32'hFFFDF787 , 32'h03FBFDCC , 32'h000073EB , 32'h03D50528 , 32'h006379DC , 32'hFFFDC595 , 32'hFFFEEFCF , 32'h00014FEE , 32'h00021AC3 , 32'h0A6EC4E0 , 32'hFCC009D0 , 32'hFFFFDE57 , 32'hF5FECC80 , 32'h0DCC0010 , 32'hF8365440 , 32'hFFFE4382 , 32'hFFA210AE , 32'hFFFFD339 , 32'hFC66FED8 , 32'hF0D1D590 , 32'hFFFF2625 , 32'hFEFD8610 , 32'h00027CE8 , 32'h0002917B , 32'h022369D0 , 32'hFDA5D948 , 32'h02ADAC54 , 32'hFFFF9296 , 32'hFEB2C130 , 32'hFFFE8136 , 32'hFFFEDB7F , 32'h01070140 , 32'hFFFE3C05 , 32'hFFFFDE12 , 32'h080FC750 , 32'h0308EE80 , 32'h0000DB8D , 32'h0000EB90 , 32'h0001B5DE , 32'h00002857 , 32'h00001C59 , 32'hFBC12570 , 32'hF5FD2590 , 32'h0001EB32 , 32'h00012F92 , 32'h09A26F00 , 32'hFE9A91F8 , 32'hFFFE28FF , 32'h000087BB , 32'h037E1150 , 32'hFFFD7D50 , 32'h000001CB , 32'hFD2349B0 , 32'hFAEBFBB8 , 32'hFE7F12B4 , 32'h026E72F0 , 32'hFFFEBECD , 32'h0000FF07 , 32'h016A05A4 , 32'hFFFD059B , 32'h000064D6 , 32'hFD72D210 , 32'hFFFE3788 , 32'h00014B01 , 32'h00B92A6A , 32'hFFFE8460 , 32'h037EA1FC , 32'h02A881D0 , 32'h00009D69 , 32'hFFFF3D17 , 32'hFFFF0481 , 32'h034958DC , 32'hFC0F0274 , 32'hFF33F4D7 , 32'h013AB248 , 32'h00010490 , 32'hF9D81FD0 , 32'hFFFFCC5F , 32'h0003CC96 , 32'h06B75E30 , 32'hFED3B5CC , 32'h00C0B1F1 , 32'h0001F824 , 32'hFFB9D8B2 , 32'h00EE39DF , 32'hF20866D0 , 32'hF599AB80 , 32'h040F8F00 , 32'hFD7F7560 , 32'h01201278 , 32'hE9E04CA0 , 32'hFFFD6B28 , 32'h000096A9 , 32'h000127A0 , 32'hF5892560 , 32'h150731A0 , 32'hFD9D0E08 , 32'hFD0B1BBC , 32'h0672BBE8 , 32'hFE9EC038 , 32'hFFFC5CD5 , 32'h094DF9A0 , 32'h01835F98 , 32'h0000B960 , 32'hEED533E0 , 32'hFFFF0FC1 , 32'h013061C0 , 32'hFBC0E6C8 , 32'h0003DD9C , 32'hFFFD071D , 32'h00007E3F , 32'hFFFFED28 , 32'h00000015 , 32'h0000695E , 32'h06BFBFD0 , 32'hE78D3840 , 32'hE469A280 , 32'hFF5C117E , 32'h099F3E60 , 32'hEECFEA40 , 32'h0000E081 , 32'h00001C00 , 32'hFFFF611E , 32'h0000119D , 32'h0002723A , 32'h04948C20 , 32'hF6BD3B50 , 32'hFB0A4730 , 32'hFFFF797F , 32'h00010B5C , 32'hFFFFFD83 , 32'h0001B256 , 32'h07E0E9B8 , 32'hF2A665A0 , 32'h00004D41 , 32'h00029158 , 32'hFFFF5F4F , 32'h0415CF70 , 32'hFC5EFB94 , 32'hF7F03890 , 32'hFFFE875D , 32'h0002BA72 , 32'hFFFFA81E , 32'h015890F8 , 32'h011646B4 , 32'hFC65B8F0 , 32'hFFFE523A , 32'h0136266C , 32'h00008C79 , 32'hFCBDA8BC , 32'h000279E0 , 32'h09704830 , 32'h0000C0A7 , 32'h017D9128 , 32'hFF467A08 , 32'hE1C24720 , 32'hFB74D3E0 , 32'hFFFF7663 , 32'h092D52E0 , 32'hFF78D9A7 , 32'h00007662 , 32'hFBC06408 , 32'hFFFF03C2 , 32'h031BDFDC , 32'h115EFB80 , 32'h02EDB184 , 32'hFFFD7C0B , 32'hFFFFAEE7 , 32'h06968FD0 , 32'hFFFE7F26 , 32'h10D34AC0 , 32'hFFFDD0AB , 32'h01B6F69C , 32'h0000771B , 32'h09B7DE00 , 32'h0002FFDE , 32'h0002A930 , 32'h00007B70 , 32'hFCC625C8 , 32'hFB122098 , 32'h0000F719 , 32'h0002B484 , 32'hFFFEABCC , 32'h0000C1A1 , 32'h02D8B324 , 32'h05374AE8 , 32'h0020D970 , 32'hF9455B38 , 32'hFE13ED58 , 32'hFFFD1931 , 32'hFFFD4FF6 , 32'h00004341 , 32'h0024759E , 32'h00006B6B , 32'hFFFC843A , 32'h01561560 , 32'h02AC5908 , 32'hFFFBCB8D , 32'hEF277840 , 32'h022E9270 , 32'hFC9B7E2C , 32'hFB934268 , 32'hFFFF10B8 , 32'h04B15860 , 32'h04245FF0 , 32'hFDA318D0 , 32'hFFFFF8DF , 32'h053E3F00 , 32'h12D5B860 , 32'hFC745CD0} , 
{32'hFEDF6CE4 , 32'h09EBB050 , 32'h0000D66E , 32'h04993208 , 32'hFFFDDB71 , 32'h02B4E8D4 , 32'hFFFD830C , 32'hFFFEE498 , 32'hFFFF40D7 , 32'hFFFF1D9F , 32'hF73C9BD0 , 32'hF6412260 , 32'h059AE0E8 , 32'h0001E27C , 32'h000255BA , 32'hFCEFAAA4 , 32'h000284D8 , 32'hF858EA90 , 32'h01741740 , 32'h000186E7 , 32'h00008BA3 , 32'hFA5AA6F8 , 32'h00DAEE65 , 32'hFD5DA990 , 32'h016DEC14 , 32'hFFFF977C , 32'h0055AE88 , 32'h01166F18 , 32'hFFFFBA5E , 32'hFBCBA248 , 32'hFFFFA177 , 32'hF9251BD0 , 32'h0002360D , 32'h00002FC3 , 32'hFFFF25C8 , 32'h015EEED4 , 32'h03A28CB4 , 32'hFB8FB538 , 32'h0002244F , 32'h000CF683 , 32'h0F5C0560 , 32'hFFFF6D58 , 32'h0000DE6B , 32'h059270A0 , 32'h021F9940 , 32'hF385ADE0 , 32'h14764F80 , 32'hFFFD94CD , 32'h0055A1E6 , 32'hFEF4FB0C , 32'h00981EA5 , 32'hFFFD99E0 , 32'h02FED3C0 , 32'h03C92474 , 32'h0A444E40 , 32'hFFFF40D7 , 32'hFEED99EC , 32'hFFFEA5A5 , 32'h00009E7C , 32'hFA9F04F8 , 32'h052447A8 , 32'hF7A44420 , 32'h0A17E940 , 32'hFFFFF0AC , 32'hF6EF05B0 , 32'hFFFD2EA0 , 32'hF0B146F0 , 32'hFBCE3A68 , 32'hFFFEE18B , 32'hFA63BBA8 , 32'h06C50DF8 , 32'hFDB36BC0 , 32'hFFFFE982 , 32'hFFFE6022 , 32'h00007968 , 32'hFB22ACF0 , 32'hFFC4351F , 32'hFFFEB635 , 32'hE27088C0 , 32'h00754592 , 32'h0001DB47 , 32'hEFD89120 , 32'hFE2E7468 , 32'hFFFFDA2C , 32'h037EC2FC , 32'h03E0925C , 32'hF8DD8D08 , 32'hFFFF0658 , 32'h000046D1 , 32'hF3221340 , 32'h00018747 , 32'h02655594 , 32'hFFFF2F3A , 32'h0886A4A0 , 32'h00835E6C , 32'h0001851D , 32'hFFFF6D72 , 32'h0000A97D , 32'h00014A32 , 32'h006A758E , 32'h0229AC2C , 32'hFFFFC32D , 32'hFF8BAB06 , 32'h0D27DEB0 , 32'hF9510960 , 32'hFFFFA021 , 32'hFEC67380 , 32'h0001B334 , 32'hF9B52628 , 32'hEE3A3700 , 32'hFFFF59E8 , 32'h05F3FC48 , 32'hFFFE1C9B , 32'h0000A96A , 32'hF9A5EE90 , 32'h043AE0B8 , 32'h009C2015 , 32'hFFFF507D , 32'hF632BEE0 , 32'hFFFF82D4 , 32'hFFFEC5A2 , 32'h028176A0 , 32'h0000BB5F , 32'h0000D0C7 , 32'h10261160 , 32'h04858D50 , 32'h00004CE5 , 32'h0002CA1B , 32'h000015C3 , 32'h0000A9EA , 32'hFFFE30C9 , 32'hFEFC81D8 , 32'h02F648E0 , 32'h00004DD3 , 32'hFFFEB944 , 32'hEB08CAC0 , 32'hFCD514F8 , 32'h0001AC9C , 32'hFFFF8A2A , 32'h03EAAAD4 , 32'h00012E7F , 32'hFFFF7CD4 , 32'hFE98CD3C , 32'hFE69F8A4 , 32'h013FB034 , 32'hFDB8B1A8 , 32'hFFFF7E53 , 32'h000040AC , 32'hFE26EB90 , 32'hFFFD39D1 , 32'hFFFF439E , 32'hFE606244 , 32'hFFFE7C37 , 32'hFFFE184C , 32'h1245FD60 , 32'hFFFC895A , 32'hF51CF6F0 , 32'h0010D521 , 32'h00010610 , 32'hFFFF7A76 , 32'hFFFF6C3C , 32'h042CF9B8 , 32'hFA09F178 , 32'hFB0EA510 , 32'hF81B3160 , 32'hFFFFD64C , 32'hF7461E90 , 32'h0000A2CA , 32'hFFFF81D0 , 32'h000A00E7 , 32'hFFE9D078 , 32'h00695C30 , 32'hFFFECB98 , 32'hFE5FF380 , 32'h004BB499 , 32'h04BEADC0 , 32'hFE625944 , 32'h11D0D380 , 32'h0ED05060 , 32'h00E6B36A , 32'hFC57F328 , 32'hFFFE050E , 32'h0001A8CE , 32'h00009F6C , 32'hFF45632D , 32'h1FA13300 , 32'hFE4B85A0 , 32'hFFD0F197 , 32'h01820000 , 32'hFC7E3008 , 32'hFFFFF589 , 32'h0CBD4B80 , 32'h06B68360 , 32'hFFFE218A , 32'h17916CC0 , 32'hFFFFE893 , 32'h06CDF708 , 32'h1F264420 , 32'h000136FA , 32'h000034AA , 32'hFFFFB73C , 32'h0000844F , 32'hFFFF44B2 , 32'h00002FC6 , 32'h01AF8054 , 32'h171C0440 , 32'h04C4E838 , 32'hFF1DC76F , 32'hFD783A1C , 32'h0B72A0F0 , 32'hFFFEC833 , 32'h000013C8 , 32'hFFFFC631 , 32'hFFFFE357 , 32'h00002630 , 32'hF901DD08 , 32'h0B8E5030 , 32'hE595EDE0 , 32'h000222A3 , 32'hFFFED6B6 , 32'h00009E87 , 32'hFFFE72EE , 32'h06B44310 , 32'h052F3660 , 32'h0002BB70 , 32'h0000DE23 , 32'hFFFC5F8F , 32'h0163E4BC , 32'hFC96D734 , 32'h04985CB8 , 32'hFFFEF1E6 , 32'h0003488C , 32'h000000DF , 32'hFF7D8449 , 32'hFF59BB68 , 32'h00AA6CB9 , 32'hFFFFF565 , 32'hFF4B6204 , 32'h0000AC67 , 32'h099700D0 , 32'hFFFF53E9 , 32'h07A15768 , 32'hFFFFAC65 , 32'hFA6FEBF0 , 32'h04DE36F8 , 32'h06858158 , 32'h1F8ABB80 , 32'hFFFFFE8B , 32'h006713C2 , 32'h01603BBC , 32'h0001D060 , 32'hF8762830 , 32'hFFFF22A9 , 32'h018A816C , 32'hFE52FF6C , 32'h0B0FDA60 , 32'hFFFEECF6 , 32'h000152BB , 32'h010DBAC8 , 32'hFFFEC4A5 , 32'h0766A430 , 32'hFFFF2C46 , 32'hFFF8849B , 32'hFFFE8A98 , 32'h013817F0 , 32'h00002387 , 32'hFFFE608B , 32'h00006FC6 , 32'h0E1A39A0 , 32'h01B40EA8 , 32'hFFFED425 , 32'h00006A06 , 32'h00006D5C , 32'h0002D9EA , 32'h00881FB9 , 32'h07739398 , 32'h00153BA5 , 32'h0EDA4450 , 32'h03FB3788 , 32'h000163D6 , 32'hFFFEC8C5 , 32'hFFFEC675 , 32'h03D40DEC , 32'h00039680 , 32'h0000003B , 32'h01D21C64 , 32'h07867CE0 , 32'h0002858E , 32'h1B76F5C0 , 32'h02720F6C , 32'h01A4CD2C , 32'hFDD49F68 , 32'h0001FF5E , 32'h00528DCC , 32'h045CB3E8 , 32'h019A283C , 32'hFFFE9AF2 , 32'hF9B4C370 , 32'hCF99C680 , 32'h0F1728E0} , 
{32'hE8F8DC20 , 32'h0BFA0240 , 32'hFFFE3B69 , 32'h00908E90 , 32'h0000A5FE , 32'h00BC7DBC , 32'hFFFE8351 , 32'h000144AD , 32'h000071AC , 32'hFFFFCEE0 , 32'h013E3924 , 32'h0641BB80 , 32'hFB2ADCC8 , 32'hFFFF2D85 , 32'hFFFE7D4F , 32'h06D26510 , 32'hFFFFB898 , 32'hFF981BDD , 32'hFD5D39B8 , 32'hFFFFA290 , 32'h0000CB6C , 32'h024B4A80 , 32'hF770E450 , 32'h037C2888 , 32'h0C401670 , 32'h00005952 , 32'hFF6AB808 , 32'h01A041DC , 32'hFFFF080A , 32'h041D67F8 , 32'h00011467 , 32'hFD4B5F5C , 32'hFFFE8E4D , 32'h0001DFC7 , 32'h0000169A , 32'hF51D8950 , 32'h050A1FE8 , 32'hF2B8EB00 , 32'h0000EFB2 , 32'hFC3606FC , 32'hF8474770 , 32'hFFFF4A24 , 32'hFFFEFEF9 , 32'h02FDB1F0 , 32'h0D322160 , 32'h31F35180 , 32'h0A6EF970 , 32'h000081EB , 32'h0297A1EC , 32'h037BFD8C , 32'hFF642388 , 32'hFFFD703A , 32'hFCCC1D84 , 32'hFC2F0630 , 32'hF8F4BD38 , 32'h0001A6E3 , 32'h0204F7B8 , 32'hFFFF0EF1 , 32'h0001C8D5 , 32'h011651A8 , 32'hFEA32220 , 32'h020A2D70 , 32'hF8972F68 , 32'hFFFFE4AA , 32'h0B1B01D0 , 32'h0000073C , 32'h0393D344 , 32'h0231BEC4 , 32'hFFFF4E73 , 32'h0FBEF9D0 , 32'h0583B100 , 32'h030C5D90 , 32'h0002B3F3 , 32'hFFFEC0CC , 32'h000337E0 , 32'h07BDA050 , 32'hFF8804A7 , 32'h0000B6A8 , 32'hF6ADC2B0 , 32'h006E3346 , 32'hFFFF12ED , 32'hEAF104E0 , 32'hFF54676A , 32'hFFFE76E5 , 32'h029E4D5C , 32'h013794D8 , 32'h01C1C934 , 32'h0000FEF0 , 32'h00024885 , 32'hF9C62148 , 32'hFFFFF271 , 32'h07116788 , 32'h0000A605 , 32'hFA860FB0 , 32'h0021C366 , 32'h00015D61 , 32'hFFFEF9EB , 32'hFFFEBDBF , 32'hFFFE224F , 32'h033F689C , 32'h004CA437 , 32'hFFFEFB56 , 32'h0171042C , 32'hF7568330 , 32'h01A5AF30 , 32'h000167F1 , 32'hFF47C98D , 32'hFFFFF480 , 32'hFED0AD30 , 32'h0AC3C190 , 32'hFFFE8EB0 , 32'h1279F760 , 32'hFFFDD028 , 32'h0000870B , 32'h06F95E08 , 32'hF9486618 , 32'hFEA30778 , 32'h0000C61E , 32'h04BD81B8 , 32'hFFFF42D5 , 32'hFFFFCA26 , 32'h052D2470 , 32'hFFFECFF3 , 32'h0001C9C6 , 32'hFCB3EC98 , 32'h0069D3CE , 32'h00019268 , 32'hFFFEE902 , 32'hFFFBA509 , 32'h000171B9 , 32'hFFFEC18E , 32'h08CBC1B0 , 32'h060C7C68 , 32'hFFFFA593 , 32'h00026B41 , 32'h0B7E90A0 , 32'hFC8390DC , 32'h00014944 , 32'hFFFE95ED , 32'hFCBB3764 , 32'h0000521B , 32'hFFFF538F , 32'hFDCCA7CC , 32'hFAA0D558 , 32'hFFE04AD5 , 32'hFED8C764 , 32'hFFFF3FC8 , 32'hFFFFE7EF , 32'hFF3E1AA2 , 32'h00022F23 , 32'h0000695D , 32'h0715C920 , 32'h000016DA , 32'h000134AB , 32'hF8C965B0 , 32'h0001EB92 , 32'hFE4D528C , 32'hFE108BA8 , 32'hFFFE176F , 32'h00007761 , 32'hFFFFEE0E , 32'h06A71B90 , 32'hF9159CD0 , 32'h0207CFC0 , 32'h024AA24C , 32'hFFFED3AF , 32'h0D4A98C0 , 32'hFFFF5932 , 32'hFFFF0CF1 , 32'hFF53B8FC , 32'h003EBC6F , 32'hFB4EF2C0 , 32'h00017B95 , 32'hEAA7DB20 , 32'hFBD179B8 , 32'hFF4A8F1D , 32'hFB692C98 , 32'hFD206F78 , 32'h0FD0BF30 , 32'hFFE58E50 , 32'hFEF19398 , 32'h00004E53 , 32'h00018462 , 32'h00019870 , 32'hFFEF7B7E , 32'hE8A9B020 , 32'h02054864 , 32'h015C2688 , 32'h03B7C604 , 32'hFC983C28 , 32'hFFFF1BDC , 32'h00771E8D , 32'h0154CD24 , 32'hFFFE1A24 , 32'h1AF7E580 , 32'hFFFF58E1 , 32'hF88EB088 , 32'h07DE06A8 , 32'hFFFEA9BC , 32'hFFFF0C45 , 32'hFFFF2605 , 32'h0000681A , 32'h00007A41 , 32'hFFFFAC0D , 32'h01EAEDE0 , 32'hDF100080 , 32'h19FDD600 , 32'hFFA4A48C , 32'h03C6CFE8 , 32'hFA4D2588 , 32'h00010808 , 32'h00004F4D , 32'h00000BE5 , 32'h00008F18 , 32'h000015C5 , 32'hF9A36B60 , 32'h011E1D34 , 32'h0C8047F0 , 32'h00004DA9 , 32'h00003713 , 32'h0000EFBB , 32'hFFFFADF5 , 32'h0078E0C9 , 32'h19CD46C0 , 32'h0001A623 , 32'hFFFEE8D7 , 32'h0001F102 , 32'h0A588D10 , 32'hFEC92D78 , 32'h08C02E90 , 32'h00011015 , 32'hFFFF4DAC , 32'hFFFFA1B0 , 32'h0385288C , 32'hFC3CC400 , 32'hEE251CC0 , 32'h0000DB4D , 32'h00A83534 , 32'hFFFDF1F3 , 32'hFF41F269 , 32'h000090A9 , 32'hF89290A8 , 32'h000040F3 , 32'h09B94EE0 , 32'h078DABF0 , 32'h101773A0 , 32'h1A768240 , 32'hFFFE8623 , 32'h013619F0 , 32'hFFE9313C , 32'hFFFFA719 , 32'h06CD8320 , 32'h0000BCAF , 32'h028C53B4 , 32'h0DBBD210 , 32'hFD8E3474 , 32'h00005323 , 32'hFFFD5E38 , 32'h07B10AD8 , 32'hFFFE71DD , 32'h05E9DBB8 , 32'h00014F0F , 32'h005AFDE9 , 32'hFFFF70CE , 32'hFBE05028 , 32'hFFFE59F3 , 32'h00007B9C , 32'hFFFEE2A0 , 32'h0147460C , 32'hFB689B38 , 32'h00019770 , 32'hFFFFA86E , 32'h000017B5 , 32'hFFFBFDE1 , 32'hFB2141F0 , 32'h060CCF88 , 32'hF7B24650 , 32'hF4BB2C70 , 32'hFB33B788 , 32'h00014D3F , 32'h00008562 , 32'h00003FEA , 32'hFD3ACF7C , 32'hFFFEA3D0 , 32'hFFFDEC7A , 32'hFC7C67C8 , 32'hFB649B38 , 32'hFFFFB778 , 32'hE48B79A0 , 32'hFE623FFC , 32'h01A963AC , 32'hFBE3FB30 , 32'hFFFEA7E9 , 32'hFC6ECFA4 , 32'hFCA3D370 , 32'h0154E10C , 32'h00020032 , 32'h0D6B8D00 , 32'hDDAC28C0 , 32'hFF35CA21}
};

logic signed [31:0] VT_2 [100][100] ='{
{32'h02D33D1C , 32'hFBDECF08 , 32'h03C11398 , 32'h00004324 , 32'hFFFFEA8B , 32'hFD4B2D1C , 32'hEF1A9340 , 32'hFBA0C710 , 32'h0000CAF5 , 32'hF47EE460 , 32'hFF1A0D52 , 32'hF1348020 , 32'hE69778E0 , 32'h076EF6A0 , 32'h0F43A650 , 32'hF5DC22C0 , 32'hE804D920 , 32'hF63C72A0 , 32'h03C5A2F8 , 32'h0000C796 , 32'hF7548A90 , 32'hF0C05D20 , 32'hF9C5EB68 , 32'h0002262E , 32'hE40BBFE0 , 32'hF28EC2E0 , 32'hF63E1C00 , 32'h0127BCFC , 32'h04A52C58 , 32'h160FCAA0 , 32'hE92E7FA0 , 32'h0B0DDE60 , 32'hFD8D0510 , 32'hE0A58A40 , 32'hFFFFD6F8 , 32'h025AFA24 , 32'hFB6BD288 , 32'h09069570 , 32'h00EFCAB6 , 32'h0012A364 , 32'hEED818C0 , 32'h00C2B8A3 , 32'hFE6B38BC , 32'hFE38D9E0 , 32'h043369D0 , 32'hFF3741B7 , 32'h0A82D1A0 , 32'h01AB379C , 32'hE615B140 , 32'h0D34D230 , 32'hFE8374D0 , 32'hE86A45A0 , 32'h0AA27C50 , 32'h09522680 , 32'hF8097F88 , 32'h0DE339E0 , 32'h0FDE07C0 , 32'h12EBECA0 , 32'h0A6C4210 , 32'h16E367E0 , 32'h057012B8 , 32'h091E8090 , 32'hE86C8600 , 32'h0B0D9F70 , 32'hFBAB0350 , 32'h1AD6E3C0 , 32'hFFFED0AF , 32'hF3E9DDA0 , 32'h02130224 , 32'hFF7DA3BF , 32'hFEA2A3CC , 32'hFF3336DE , 32'hFDA6C6EC , 32'hFA394100 , 32'hFBDE9740 , 32'hFA292258 , 32'hFC2E7EE4 , 32'h0B0E0160 , 32'h1C852800 , 32'hFBEC9E08 , 32'h149BE8E0 , 32'h18E38CA0 , 32'h0666FFE8 , 32'hFFFF8634 , 32'hF5AB8EF0 , 32'hFFAEBC1E , 32'hEE4C7700 , 32'hE803B860 , 32'h0C3FEB50 , 32'h0000A6D0 , 32'hEC4BAD80 , 32'hFAE53758 , 32'h000949B7 , 32'hE97D66E0 , 32'hFFFFE1D9 , 32'h11C01000 , 32'h0B578B60 , 32'h09F64890 , 32'hF9845B18 , 32'hEEDC4000} , 
{32'h0D870E60 , 32'hEF38E560 , 32'h0131F7D0 , 32'hFFFFA297 , 32'hFFFFC33B , 32'h173B3AC0 , 32'h016B7C3C , 32'hF693EF10 , 32'h00006E67 , 32'hD3000E40 , 32'h10521FE0 , 32'h038CE3B0 , 32'hE8503800 , 32'hF8C9EA10 , 32'h0E766F30 , 32'h14462CA0 , 32'hF3BAA470 , 32'h0236C7EC , 32'h06A8C110 , 32'hFFFFEAF1 , 32'hFB65CFD0 , 32'h0C211240 , 32'hFC107600 , 32'hFFFF5C9F , 32'h0769CE28 , 32'hF2779D30 , 32'h05BC9B38 , 32'h02D2CCC0 , 32'h00E26E79 , 32'h0DCF5380 , 32'hFA36D258 , 32'hEE05FE00 , 32'hFC30F9B4 , 32'h085B6E80 , 32'h00009341 , 32'hFFCA32A9 , 32'h059E8740 , 32'hEA6A22C0 , 32'h02D7CBA0 , 32'hF2440820 , 32'hEF525F40 , 32'h004D7828 , 32'hFCE05980 , 32'h0DC01F10 , 32'h18FC92E0 , 32'hFC4C9894 , 32'h06463468 , 32'hF75A0790 , 32'hFCF749B0 , 32'hFB5B5128 , 32'h07026A78 , 32'h0D1F4CE0 , 32'hE6DBE9C0 , 32'h05C30DE8 , 32'h13F6E380 , 32'h037BFBC4 , 32'h26731840 , 32'hF439E2F0 , 32'hEE7C0980 , 32'h12145020 , 32'hF623F510 , 32'h07DD5258 , 32'h08E66A60 , 32'h0DCA5830 , 32'h03A4C45C , 32'hF1CABDD0 , 32'h0001222E , 32'hFC49FA10 , 32'hF9EECE40 , 32'hFB0DC8D0 , 32'hFE344360 , 32'hEF556BE0 , 32'hFCA4BE54 , 32'h0A31F6C0 , 32'hEF19EF20 , 32'h09BAD6C0 , 32'hF2AB44A0 , 32'hEC578AC0 , 32'h0FF0A0F0 , 32'hF537E3B0 , 32'h0532FC18 , 32'hFEABA9B8 , 32'hFECDF260 , 32'h00006AC8 , 32'hFDE0B8F8 , 32'h09F3DE00 , 32'h09B873F0 , 32'h1069C520 , 32'h0B69CF50 , 32'hFFFEB1AD , 32'h0AF3C100 , 32'hFE5E99A4 , 32'hFBB71A40 , 32'h169D6000 , 32'h000083E4 , 32'h06DF2B88 , 32'hFD3E9EA0 , 32'hE6FEA9E0 , 32'h17238180 , 32'hFABCBED0} , 
{32'h09ECF500 , 32'h12C71240 , 32'h02630FD8 , 32'hFFFFCFD3 , 32'h0000793D , 32'hECC3DD20 , 32'hF1975620 , 32'hE0E86640 , 32'hFFFFC4BE , 32'h00984EF0 , 32'h029E7BA8 , 32'hF84D4EE8 , 32'h128E5E20 , 32'hF1E92950 , 32'h0C370F40 , 32'hFC99D63C , 32'hF96C7C60 , 32'hFA645E98 , 32'h05AAD120 , 32'hFFFF8637 , 32'h04730D58 , 32'h0C9B0A40 , 32'h163F9240 , 32'h0001F520 , 32'h0F926BE0 , 32'hF49C4ED0 , 32'hFC9E9048 , 32'hFA536C18 , 32'hFC4473F4 , 32'hFFFFD597 , 32'hF4766170 , 32'h1690D360 , 32'h030EBE30 , 32'h0E8195A0 , 32'h00015111 , 32'h0C3BFFC0 , 32'h02F80218 , 32'h115D8440 , 32'h099E62C0 , 32'h09E45FC0 , 32'h00CCAD69 , 32'hFFED7912 , 32'hF5AAFB10 , 32'h216D4A80 , 32'hECEC7340 , 32'hFAF03378 , 32'h11882FA0 , 32'hFA46C2E8 , 32'hEB5EE960 , 32'h02EB4EC0 , 32'h14DFE680 , 32'h0C27D9E0 , 32'hFF67C046 , 32'hEF9C3660 , 32'h01EA9E90 , 32'hF5F329A0 , 32'hF99D6C28 , 32'hEF768C00 , 32'hF561BE80 , 32'hF58C6D00 , 32'h04E084A0 , 32'h070987D8 , 32'h0E777910 , 32'h03E581B0 , 32'h0C7B1230 , 32'h0E068870 , 32'h00019874 , 32'hF7FF44A0 , 32'hFF09468F , 32'hF492DE40 , 32'h09250E70 , 32'hF1677A90 , 32'h0165C65C , 32'h0FAB7230 , 32'h00BF604C , 32'h01461E2C , 32'h066872F0 , 32'hEE4CBC60 , 32'h16FEF9E0 , 32'h1F0EAC80 , 32'hF1C26CB0 , 32'h12B0C980 , 32'hF0153A10 , 32'hFFFF494F , 32'hF5BB1550 , 32'hFA6EF388 , 32'h092F6B60 , 32'h19D92B60 , 32'h110C0780 , 32'hFFFF3E07 , 32'h07ACDF48 , 32'hFF26BF4A , 32'hEC78C9C0 , 32'hF0689510 , 32'hFFFFA129 , 32'h08046A20 , 32'h18CDA7E0 , 32'h0C475E20 , 32'hEFF986C0 , 32'h037A0454} , 
{32'hE9EAA040 , 32'hF5BA60F0 , 32'h03B7B898 , 32'h0000D17A , 32'h00005804 , 32'hF41BDC40 , 32'hFBAF7898 , 32'h0B7B7D80 , 32'h0000683C , 32'hFED3839C , 32'hF25440F0 , 32'hF8E8F1B0 , 32'hF30906A0 , 32'h0B7037F0 , 32'hEE66FD00 , 32'h0AE63D80 , 32'hF3CC8900 , 32'hE77BAE60 , 32'hECBA5C80 , 32'hFFFE9BAA , 32'hFC848830 , 32'h12EB5EE0 , 32'h0166FD74 , 32'hFFFFAE02 , 32'hED70E840 , 32'hFEC6FC60 , 32'hFF9636BE , 32'hFE6434C0 , 32'h0CCFAF00 , 32'h03078670 , 32'hF1A0B200 , 32'h02B01444 , 32'h00D00C86 , 32'h19904440 , 32'hFFFFCF17 , 32'hEE086AE0 , 32'hFAFA10B8 , 32'h08AA6240 , 32'h01F06E24 , 32'h0638D840 , 32'h140CA920 , 32'hFFA120D4 , 32'hFDC2A340 , 32'h2272D840 , 32'hE39E5820 , 32'h017B89B0 , 32'hE1EA5C00 , 32'hEB39F480 , 32'h04197BE0 , 32'h06211C70 , 32'h1170EE80 , 32'h0CC1C250 , 32'hEDA1ED40 , 32'h000590EE , 32'h0F6C5A90 , 32'h06593A88 , 32'hF8B84CC8 , 32'hE6BFDC60 , 32'h0EA270D0 , 32'h03133204 , 32'hFC91A838 , 32'h0F33BC90 , 32'hF9BECE08 , 32'hFBD49F90 , 32'hEC3CB9A0 , 32'h075558E0 , 32'h0000E37F , 32'hEE883EE0 , 32'hFF91D9A6 , 32'hEE005B60 , 32'h0AF35E50 , 32'hF4544140 , 32'h130F30A0 , 32'hFAFFBBD8 , 32'hFDF200C8 , 32'h120BA0C0 , 32'h16DDA040 , 32'h00C7A5E6 , 32'h0676A530 , 32'hFA779078 , 32'h0C7BBE10 , 32'hED14D9A0 , 32'h12EB77A0 , 32'h00000CB5 , 32'h08CE3DF0 , 32'h16C26420 , 32'hFA8BBB60 , 32'hEE994D80 , 32'h03F31F24 , 32'hFFFF9355 , 32'hFBC793A0 , 32'h01E9E420 , 32'h007BA223 , 32'hFF244BDA , 32'hFFFF9948 , 32'h0026D1CF , 32'hEA1E6240 , 32'h02D396D8 , 32'h02AD46BC , 32'hF5B298F0} , 
{32'h196E63C0 , 32'hEFE95060 , 32'h0E3916A0 , 32'h0000FB83 , 32'hFFFF51DB , 32'hFE49B658 , 32'hF718B6C0 , 32'hF5E4CF00 , 32'h0000E374 , 32'hFD156694 , 32'h043AD1E0 , 32'h0C1FA060 , 32'hF6ED4600 , 32'hF44FD770 , 32'h033C9EE0 , 32'hF9DD1F08 , 32'hF4DC80A0 , 32'hF4A9F590 , 32'h041EFF88 , 32'h000013F7 , 32'hFBBC4828 , 32'hE71DD020 , 32'h00A4F348 , 32'hFFFDE713 , 32'h0EB77B00 , 32'h06C53A70 , 32'hFD701F48 , 32'hFA8DD4A8 , 32'h013BDAF8 , 32'h1D850840 , 32'hF2BC8210 , 32'h0E454F90 , 32'hFA34E0D8 , 32'hF2D71000 , 32'h00004059 , 32'h072CCBF0 , 32'h04FE5530 , 32'hFD8E1220 , 32'hFFD5CBD6 , 32'h0E604910 , 32'hFDCF91A8 , 32'h010F3808 , 32'h0008A459 , 32'hF91D4D50 , 32'hE9A00400 , 32'h079C1AB0 , 32'h126F2920 , 32'hF9F90D98 , 32'h051A73D8 , 32'hF4AAA370 , 32'h0923A420 , 32'h11EC4660 , 32'hFE4FC894 , 32'h0BA63A60 , 32'h0D6371D0 , 32'hF4DB1D70 , 32'hF6EE85F0 , 32'hFA53DDA0 , 32'hF92ECEA0 , 32'hF2D6E1A0 , 32'hF08F09D0 , 32'h1109D5E0 , 32'hFB645788 , 32'h0095D0C5 , 32'h10583DA0 , 32'hF202AE80 , 32'hFFFFFF71 , 32'h14AEA7C0 , 32'hFC4FD10C , 32'h17092DA0 , 32'h052EB5A8 , 32'h05FB3530 , 32'h1531A6A0 , 32'hF59B2750 , 32'h160D3280 , 32'h002D77DC , 32'hFE144AB4 , 32'h0F5E33B0 , 32'hF0F741A0 , 32'hFC0788CC , 32'hFBCA87E0 , 32'hF005B480 , 32'hF52A5250 , 32'h0000AA45 , 32'h16DCC220 , 32'h0FE2D320 , 32'h1F654540 , 32'hFECED660 , 32'hEA803FA0 , 32'hFFFF71C9 , 32'hF3ECF3B0 , 32'h019BDBFC , 32'hFE8E1B9C , 32'hE30B32C0 , 32'hFFFFFDE9 , 32'h1933D420 , 32'hE90CF3C0 , 32'hF47A6A00 , 32'hFCDACB54 , 32'hE2202DC0} , 
{32'hFE797FD0 , 32'hF0E1D290 , 32'h1427C9A0 , 32'hFFFEFD0D , 32'hFFFF7354 , 32'hFF58DDD0 , 32'hF3220EE0 , 32'hFDBD8004 , 32'h0000CF4B , 32'h077F9030 , 32'h0D623F30 , 32'h192802C0 , 32'hF8648B80 , 32'hFBFBA4F8 , 32'hEED52320 , 32'hECFF0920 , 32'h0399B3A4 , 32'hF887F340 , 32'hDF365780 , 32'hFFFFA8C4 , 32'h1552DD80 , 32'h062DD9E8 , 32'hFA979EE0 , 32'hFFFFCC68 , 32'hEE0DD8E0 , 32'hFBD1CC78 , 32'hEE591B80 , 32'hFBF7C658 , 32'hF16192D0 , 32'h1F7431C0 , 32'h1764DE00 , 32'hF41C2BA0 , 32'hF73BC940 , 32'h0AC80580 , 32'hFFFFA96C , 32'hF520DA30 , 32'h0688E428 , 32'hEE6A4440 , 32'hF5C94E40 , 32'hF894FD20 , 32'h115D9B40 , 32'h00FE1E6A , 32'hFF273147 , 32'hF231FB30 , 32'hFC7903A4 , 32'h0F95A370 , 32'hEA3A7C80 , 32'hF85C6EE0 , 32'h14C12880 , 32'h172D55A0 , 32'h14671D60 , 32'h0A873540 , 32'hF6BDDC50 , 32'hF3D58610 , 32'hEAB105A0 , 32'hF52B7600 , 32'h07D790F0 , 32'h0C51A000 , 32'hFB5D8518 , 32'h106BEF00 , 32'hFA3FC978 , 32'h09C9E980 , 32'h0CE939C0 , 32'h08BC0430 , 32'h05B997F0 , 32'h0DA86FB0 , 32'hFFFFFC49 , 32'hFE13E988 , 32'h02CE8BB4 , 32'h072CCA70 , 32'hF8685A50 , 32'h045CBFE8 , 32'hFDA67520 , 32'h04F32058 , 32'hFAC847F8 , 32'hF0305850 , 32'h05BC48B8 , 32'hEC2A6B00 , 32'h02183508 , 32'h0381E46C , 32'hF83C2890 , 32'h17E12420 , 32'h03F836A4 , 32'h0000993D , 32'h0C564790 , 32'hE665EC60 , 32'hFC8FD810 , 32'h1E8AD6A0 , 32'hFF5CFF54 , 32'h0000E3B8 , 32'hEA1AE340 , 32'h00C00476 , 32'h09BD1470 , 32'hF4F15FE0 , 32'h0003124D , 32'h0064B86E , 32'h0A9CF710 , 32'hFFAFC335 , 32'hFBF61618 , 32'hF44369B0} , 
{32'h0949D0F0 , 32'hF5C6D5F0 , 32'hF6B9D370 , 32'h00001215 , 32'h00006BAA , 32'hEDC05B80 , 32'h041DFFA0 , 32'hE1C578E0 , 32'hFFFFEE08 , 32'h0D96C620 , 32'h0AF56350 , 32'hF94DCCC0 , 32'h114B6AA0 , 32'h097F1980 , 32'hF7DB2530 , 32'hF38EA250 , 32'hEC94D820 , 32'h024A3410 , 32'h08B1C630 , 32'hFFFEF076 , 32'h216B0BC0 , 32'h09D0F930 , 32'hE9267280 , 32'h0000951B , 32'hFE8D7650 , 32'h14473540 , 32'h0A720510 , 32'h12C91BE0 , 32'hF210DFE0 , 32'h0B382D60 , 32'h1968B5C0 , 32'h0D923DD0 , 32'hFADE4710 , 32'h00FD2BCE , 32'h0000485D , 32'h0742E9D8 , 32'hF6F52460 , 32'hE735F0A0 , 32'hF8C46830 , 32'h023269A8 , 32'hFBDA3F30 , 32'h000E45EA , 32'h037751DC , 32'h01253854 , 32'hECDEA860 , 32'hD9489540 , 32'h06AD7518 , 32'h17B3B420 , 32'hF18CAA30 , 32'hFD5EB674 , 32'h07AA21C0 , 32'hEEF58680 , 32'hF2365370 , 32'hFAA76378 , 32'h05E716A0 , 32'h0B4B88C0 , 32'hFEDCF978 , 32'hF1A28BC0 , 32'h049DC928 , 32'h0AFA19E0 , 32'hEBC72720 , 32'h0620C8B0 , 32'hF4C349C0 , 32'hF7EEB330 , 32'hFB5573D0 , 32'hF442EDD0 , 32'h00002A20 , 32'h1771EB60 , 32'hF64818A0 , 32'hEF6490A0 , 32'hF96445F8 , 32'hFB456390 , 32'h066879A0 , 32'h02D2B1FC , 32'hF6C78940 , 32'h0AF58940 , 32'h0919ABD0 , 32'h079AE9E8 , 32'hFF685025 , 32'h0D369450 , 32'h17195B00 , 32'h12A695E0 , 32'h06F31DA0 , 32'hFFFF7C9D , 32'h0D6AFA60 , 32'hF6CC6A10 , 32'hF501E930 , 32'hF4CBF080 , 32'hF98D9658 , 32'h0001AC5A , 32'h0FB78D00 , 32'h01D9A2D8 , 32'h136A8E80 , 32'h0F6CA140 , 32'hFFFE8455 , 32'h07E3E480 , 32'hFE02F65C , 32'hF0958FB0 , 32'hFBAA3ED8 , 32'hFCAF1A70} , 
{32'hFAFAF9C0 , 32'hFE1C9640 , 32'h0DA484F0 , 32'h00004AA8 , 32'h0000AE40 , 32'hFCDA5434 , 32'hFD581318 , 32'hF6E7AD90 , 32'h0000385F , 32'hEFC09180 , 32'hF2AB1390 , 32'hF1CE0B60 , 32'hEFF0AD00 , 32'hF3972C50 , 32'h12C31860 , 32'hFCC9D7FC , 32'hF8EE7E40 , 32'h021F7EF4 , 32'hF5976A00 , 32'hFFFFC5F9 , 32'h04A29390 , 32'h11CF67A0 , 32'hF09158A0 , 32'h0000F77E , 32'h0095EFFC , 32'h08CFF480 , 32'h05DFC5A8 , 32'hF35E8700 , 32'hECDAD660 , 32'hF906B440 , 32'h0B367E30 , 32'hEFBDE140 , 32'h1F76DA40 , 32'hFB2C7188 , 32'h00015918 , 32'h07A576F8 , 32'hFB0F7C38 , 32'h03A8E020 , 32'hF43CE6F0 , 32'hDD954500 , 32'h0548CE48 , 32'hFFCBBB8A , 32'hFEE0EAF4 , 32'h0EA53410 , 32'hFB6F8C48 , 32'h0712A208 , 32'hF8428980 , 32'h0CF28BB0 , 32'h018A1730 , 32'h0ABA3280 , 32'h0D850960 , 32'h09F2FE70 , 32'h0A252760 , 32'hFDB021D4 , 32'hECD896A0 , 32'h0A873040 , 32'hDEC81A40 , 32'h04152230 , 32'h0FF0A4E0 , 32'h04DEB8F0 , 32'hF966AAB0 , 32'hF612F210 , 32'h0ECA71B0 , 32'hF8949EF0 , 32'hF03C2C90 , 32'hE5475B80 , 32'h00004760 , 32'hF71807A0 , 32'hF4C2C700 , 32'h0C2412F0 , 32'h0DB54C50 , 32'h07C8A000 , 32'hEF2CED80 , 32'h001A142E , 32'h0C229150 , 32'hF2616C80 , 32'h0507B850 , 32'h03C7A268 , 32'hF8796AE0 , 32'h02541B68 , 32'h1360E6E0 , 32'hFCBCC0A8 , 32'hEF8759E0 , 32'h0000AF1A , 32'hED4F4B80 , 32'h07FFA798 , 32'h037EF528 , 32'hF2F6FBF0 , 32'hFB99DFC8 , 32'h00022845 , 32'hFBC59190 , 32'h0602FBD8 , 32'hE6658980 , 32'hF59FAEA0 , 32'h0000572B , 32'h1BE8F620 , 32'h100DA0A0 , 32'hD7A48780 , 32'hFD9D354C , 32'h04668390} , 
{32'h0B734140 , 32'h182D2A40 , 32'hF97DD3F8 , 32'h0001985C , 32'hFFFFA020 , 32'hFC206558 , 32'hFA6C9BB0 , 32'h1D7FCDC0 , 32'hFFFE8B24 , 32'hECAAACE0 , 32'h018C00DC , 32'hF0A26180 , 32'hDF7A9840 , 32'h0769B2E0 , 32'hF75B23D0 , 32'h07309150 , 32'hFC3678E8 , 32'hDDDA3E00 , 32'h0EC5B6E0 , 32'hFFFF3425 , 32'hFA9249A8 , 32'hF9307948 , 32'h036FE26C , 32'h00011139 , 32'h19B7CD00 , 32'h0CE422F0 , 32'h0393C694 , 32'h09A1CF20 , 32'hF1FD7320 , 32'hE8412CC0 , 32'hF4201660 , 32'h11405840 , 32'hD97130C0 , 32'hFA0606F0 , 32'h00010211 , 32'hF9F84650 , 32'hFDDA6C98 , 32'hFB142F80 , 32'h04780590 , 32'hFCE31D84 , 32'h0AEAC520 , 32'hFF5A2009 , 32'hF996FCA8 , 32'h0387B470 , 32'hFDDBFE24 , 32'h09C58570 , 32'hF426C530 , 32'h09890C40 , 32'h09C88720 , 32'h0B75AED0 , 32'h1154AF60 , 32'h08050D90 , 32'hF70468E0 , 32'hF504E4B0 , 32'hF84A0A48 , 32'h0B12A150 , 32'hFDCF9BE4 , 32'h0524C0D0 , 32'hF8CFBFF0 , 32'hF6E21210 , 32'hF007CB20 , 32'h02C4276C , 32'hF0E3D890 , 32'hFA2C4878 , 32'h104852E0 , 32'hF81D2CC8 , 32'h00000155 , 32'hEA66D660 , 32'h04822A20 , 32'hFEFA7E7C , 32'hFE33DD00 , 32'h03FB4170 , 32'h0CA69C10 , 32'hFE2ED0BC , 32'hF4B18130 , 32'hF63FE920 , 32'hF936A978 , 32'h190B0A60 , 32'hECA267E0 , 32'h11B44EE0 , 32'h0340032C , 32'h15F88260 , 32'h09964170 , 32'h0000F859 , 32'h06DC3408 , 32'hF7783E10 , 32'h04558D80 , 32'h079359B8 , 32'hF0B37DF0 , 32'hFFFE9991 , 32'hFFAAA734 , 32'hF6D9A320 , 32'h0B905E30 , 32'h0C2BC280 , 32'hFFFF1656 , 32'h013CCAC0 , 32'h22ECD2C0 , 32'hF540D340 , 32'h07CB1B08 , 32'h0994E690} , 
{32'hF91F0210 , 32'hF9104360 , 32'hE66E5EA0 , 32'hFFFE787D , 32'hFFFEF83D , 32'h144F3780 , 32'h08211710 , 32'hDED9E840 , 32'hFFFE6377 , 32'hE4EC02A0 , 32'hF14AAC40 , 32'hF863A1C8 , 32'hE81B1660 , 32'h008CF813 , 32'hF3B96920 , 32'hF339DF90 , 32'h25382F80 , 32'h01C7CF18 , 32'hFACA1D48 , 32'h0001DEF7 , 32'hF37F8070 , 32'hF5D336D0 , 32'h07503E28 , 32'h000058CE , 32'h03CAFD4C , 32'hFA71D0B0 , 32'h03B4C2D4 , 32'hF91FFAA0 , 32'h03C9FB78 , 32'hF3F83050 , 32'hF48B6350 , 32'h09311B20 , 32'hEC52CD40 , 32'h016C0B90 , 32'hFFFEF4C7 , 32'hF2F64830 , 32'h051DC2F0 , 32'h022C3958 , 32'hEF2098E0 , 32'hF1000720 , 32'h00E2EAA4 , 32'h0011CEB2 , 32'h03D9623C , 32'h0761BB48 , 32'hF6703120 , 32'hEEB752C0 , 32'hF9DE82C8 , 32'hFAFD6388 , 32'h05EF7410 , 32'hE22AA360 , 32'h0C22B480 , 32'hEA33D440 , 32'hF3367B70 , 32'h0467B348 , 32'h051F8E70 , 32'hF5B22650 , 32'hF4D5E0C0 , 32'hF7C7E0D0 , 32'hF431E290 , 32'hFA8510C8 , 32'h047B8FA8 , 32'hFBA61D28 , 32'h00D3744B , 32'h05710438 , 32'hED2ADF80 , 32'hEF935BC0 , 32'h00017BB4 , 32'h0DFE7D10 , 32'h010CBE24 , 32'h0B404EA0 , 32'h080CC8C0 , 32'hF6309AC0 , 32'h020514BC , 32'h01D4CC80 , 32'hFADB6768 , 32'hFAF8E488 , 32'h0341C35C , 32'hE93B6CE0 , 32'h006FE6EB , 32'hFAB38698 , 32'hEB0DEF40 , 32'h073A3A70 , 32'hFC7DE334 , 32'hFFFE9EED , 32'h03322828 , 32'hE16A3780 , 32'hE90B3040 , 32'hE8B66C20 , 32'hFD03E548 , 32'hFFFF8B2D , 32'hF58F65F0 , 32'hFCD233E0 , 32'h1033D900 , 32'hE60779C0 , 32'h0000EEB8 , 32'hFB258888 , 32'h086052B0 , 32'hF59F7D10 , 32'hEA48D940 , 32'hF879C2B0} , 
{32'h24305100 , 32'hF59F6410 , 32'hFEC474E8 , 32'h000038D1 , 32'hFFFF137B , 32'h07BB6850 , 32'hFDE25A5C , 32'h11D2CC80 , 32'h0000203C , 32'h07A323F0 , 32'hFF4371D6 , 32'h0AE81D50 , 32'hF4997870 , 32'h05B536A0 , 32'h035BE178 , 32'h03AC4A4C , 32'hFFE4BA46 , 32'hF9546580 , 32'hF799D720 , 32'hFFFFFA04 , 32'h21994100 , 32'h009337F3 , 32'h112F8920 , 32'h0000D103 , 32'hF3D09040 , 32'hFD7CFAE8 , 32'hF805F1C8 , 32'hF691FA70 , 32'h151C6DE0 , 32'hF009D650 , 32'h26B78940 , 32'hDD69C8C0 , 32'hE50C16E0 , 32'hDC85FA00 , 32'h000117F6 , 32'h0AD9C670 , 32'h01B5C010 , 32'h04A29F78 , 32'h00DD4623 , 32'hF8B39F40 , 32'hF5798770 , 32'h000058AE , 32'hFB6A39C0 , 32'h0F205D60 , 32'h023F38F0 , 32'h06153760 , 32'h0FEA8410 , 32'h004A4D19 , 32'h011D0634 , 32'hFB9C3910 , 32'h0C44A240 , 32'hF8FA9FB8 , 32'hF87E9250 , 32'hEEDA19E0 , 32'h0D97ADE0 , 32'h0421D2D8 , 32'hF41489A0 , 32'hE51248E0 , 32'hF56EC5E0 , 32'h00F4C308 , 32'h00968C31 , 32'hF0C382D0 , 32'h03882BDC , 32'hFC7FE9D4 , 32'h00004A91 , 32'h002BAE38 , 32'hFFFCEB67 , 32'h0478EE30 , 32'h00CE2B0D , 32'hFD290A3C , 32'h07AB50B8 , 32'hF294B650 , 32'h028C3990 , 32'h0450AEC0 , 32'h033DA214 , 32'hFE7A2D58 , 32'h002D2B90 , 32'hFEBBA88C , 32'h06081DD0 , 32'h070CA0B0 , 32'h10AD2920 , 32'hE9CC27A0 , 32'h13127860 , 32'hFFFD561F , 32'hFCACCC08 , 32'hF11784A0 , 32'h0EF73260 , 32'hEA9DB000 , 32'h004682F4 , 32'h000215E6 , 32'hF6285880 , 32'h02570A74 , 32'hF516F600 , 32'hEFA2D400 , 32'hFFFE7B66 , 32'h020A55E4 , 32'h0AFB8600 , 32'h1D1A1D20 , 32'h069B67C8 , 32'h0D77CD40} , 
{32'h1542AA60 , 32'hF766B230 , 32'hF796C970 , 32'hFFFE4A28 , 32'h00035AC5 , 32'hF65D06A0 , 32'h0771EFE8 , 32'h082ED960 , 32'h0001B258 , 32'h034423CC , 32'hF45E9730 , 32'hFC705B28 , 32'h0880D160 , 32'h09AF1E70 , 32'hF64FCAB0 , 32'hF7D41010 , 32'h0A745560 , 32'h0AB9F710 , 32'hE24755C0 , 32'h0001AC0E , 32'hE7CA3680 , 32'hFC9A7F6C , 32'h07DA2E78 , 32'hFFFE2200 , 32'h134688C0 , 32'h08CBA3E0 , 32'h030CA654 , 32'hFF086608 , 32'hEE8AD440 , 32'h05B43068 , 32'hDE5DC3C0 , 32'hFCCE5300 , 32'h13552B60 , 32'hD64418C0 , 32'hFFFF16BF , 32'h148D5FA0 , 32'hFD02E9C4 , 32'hF31B1590 , 32'hF97A15A8 , 32'hFA0B0D60 , 32'h0B3D7AA0 , 32'hFF18E3AD , 32'h00645FCB , 32'h0CA5ABB0 , 32'hFFBCFD58 , 32'hF6B9DD00 , 32'h1C085F00 , 32'h01210048 , 32'h152C31A0 , 32'h11675180 , 32'h089920B0 , 32'h0313DADC , 32'hE8F728C0 , 32'hFB3352F8 , 32'hEF73F1E0 , 32'hF991D9F8 , 32'hEB176D00 , 32'h00C96018 , 32'h0F75B3F0 , 32'hFC465338 , 32'h00533DBC , 32'h09F4F750 , 32'h01A1D098 , 32'h09EF3A20 , 32'h099EE420 , 32'h0C6C5FA0 , 32'hFFFC57E0 , 32'h084D32F0 , 32'h03697B0C , 32'h000858E0 , 32'h012171BC , 32'h07DE8B58 , 32'h0B9CD290 , 32'hFE0BC960 , 32'hF241D5D0 , 32'hFF96322C , 32'h118198E0 , 32'hEC851CA0 , 32'h16D8A2E0 , 32'hDFF94840 , 32'h08C55FA0 , 32'hF4C96F60 , 32'h0C254720 , 32'h00023ABB , 32'hFCEF21CC , 32'hFEAB2A94 , 32'h04159460 , 32'h02F95EE4 , 32'h01B51E68 , 32'hFFFD132C , 32'h0D5B0CC0 , 32'h0243AE44 , 32'h0DF8F180 , 32'h1CD83720 , 32'hFFFE9C45 , 32'hFBD46490 , 32'h0F4B6A90 , 32'h0586D468 , 32'h00C693DE , 32'hFF282D51} , 
{32'hF025B550 , 32'hF31B9DC0 , 32'h060F2540 , 32'h0002E5C9 , 32'hFFFF8383 , 32'h02AD0F2C , 32'hFD13B3C4 , 32'hEE1F1940 , 32'h0002BFF1 , 32'hFC7122E8 , 32'hEF2750C0 , 32'h099E26C0 , 32'h0A05F1D0 , 32'hF34200B0 , 32'h022D8194 , 32'hF1429EC0 , 32'hEFE76980 , 32'h06833B58 , 32'h0B903620 , 32'h00000D69 , 32'hF42CE8C0 , 32'hF739ADE0 , 32'h0B382390 , 32'hFFFEF727 , 32'h0B1C7120 , 32'hFAD10E90 , 32'hF6C51F70 , 32'h09122520 , 32'hF9559B80 , 32'hF9016EA8 , 32'h076841E0 , 32'hE5A08480 , 32'hEBBD64C0 , 32'hF6289610 , 32'h000084FF , 32'h12241F80 , 32'h114E2F80 , 32'h3AFAC800 , 32'h128FB940 , 32'hFA33C6C8 , 32'h1D6B6680 , 32'hFF5D7943 , 32'hFCA289D0 , 32'hFAACF0F8 , 32'h107802C0 , 32'hF4C89F90 , 32'hF00D15D0 , 32'h10210B00 , 32'hEA5EE040 , 32'h1533AA60 , 32'h050410B8 , 32'h07798AA8 , 32'hDAB07940 , 32'hF85B4578 , 32'hF5366800 , 32'h0025076B , 32'hFEBA5FA8 , 32'h07FDCD58 , 32'hF8E425D0 , 32'h0677C420 , 32'hED0B7B40 , 32'h03DDF0E0 , 32'h0B8DD8A0 , 32'hFEBD21C0 , 32'hFC46BF68 , 32'h08D0B900 , 32'hFFFDA7FA , 32'h06470518 , 32'hF63A6500 , 32'hFAE79750 , 32'hEF884AC0 , 32'hF52C95A0 , 32'h09759D70 , 32'hFB867218 , 32'hFE6DCEC8 , 32'hFE56149C , 32'hFC495D60 , 32'h05401CA8 , 32'hEFE9C2A0 , 32'hF8402E78 , 32'hF6004CB0 , 32'h054779F0 , 32'hF0BE1E90 , 32'hFFFF3295 , 32'hFBAB9CF0 , 32'h024AE894 , 32'h05CCEA88 , 32'hE8B302E0 , 32'h00D44CE5 , 32'hFFFE091E , 32'hFEE8A754 , 32'hFA7962A0 , 32'h0AD5D880 , 32'h0DF93BA0 , 32'h00003CA7 , 32'hFD0FB3B4 , 32'hF258AE80 , 32'h03E0EB70 , 32'h030C4D5C , 32'hF61FDB80} , 
{32'h0FF97950 , 32'hF2F8DCA0 , 32'hEF952760 , 32'hFFFF8552 , 32'hFFFE934F , 32'hFA222FD8 , 32'hF0D4E060 , 32'hE7452860 , 32'h0000DAFB , 32'h0E5ACC00 , 32'h08334980 , 32'h0F9F3DF0 , 32'h16D3F200 , 32'h0145DA88 , 32'h003A72BB , 32'h04FF3960 , 32'h0D368F30 , 32'hFB2100B0 , 32'hF9C41318 , 32'hFFFFD75D , 32'h0E41D4D0 , 32'h0631BAD0 , 32'h010BF3DC , 32'h00023F50 , 32'h02B14C9C , 32'h10AC59E0 , 32'h04DAD3E0 , 32'hF9D24038 , 32'hF4344CC0 , 32'hF89C8B78 , 32'hDF4ABD00 , 32'hFAE4B7B0 , 32'hE4C7D3C0 , 32'h1A3589E0 , 32'h00022995 , 32'hF2091C90 , 32'h068928F8 , 32'h008C3258 , 32'hFDAEE344 , 32'hF1A11010 , 32'hE80DCEE0 , 32'hFEDC6078 , 32'h03FF3894 , 32'hF12085D0 , 32'h0671FDA0 , 32'h09D4A320 , 32'h00131799 , 32'hEDA48120 , 32'hE7C7B5A0 , 32'h07C5E578 , 32'h11C2B6A0 , 32'h24D0E340 , 32'h15BF3C00 , 32'h0EA08A90 , 32'h06800588 , 32'h014CFABC , 32'hF5C49F50 , 32'hFEB032CC , 32'h0316EB28 , 32'h0F0C5050 , 32'hFC112B9C , 32'hF7C63D40 , 32'h03E3B88C , 32'h012E32B8 , 32'h05435448 , 32'h0D34B5B0 , 32'hFFFE3F95 , 32'hF692C570 , 32'h03048F40 , 32'h0DB14AF0 , 32'h030E6360 , 32'h06D96418 , 32'h04012730 , 32'h01BE3608 , 32'h0B8FFCF0 , 32'hF1BB1580 , 32'h07203808 , 32'h1756BC40 , 32'h0A9D3110 , 32'hEC121BC0 , 32'h00AE0B81 , 32'h001EE2EB , 32'h07A46478 , 32'h0001D22B , 32'hF4568300 , 32'hE9442680 , 32'hFEE2BBA0 , 32'hDD5EE2C0 , 32'h033EAB54 , 32'h000190A5 , 32'h0C042FE0 , 32'hFE474774 , 32'hFC473590 , 32'h0C9F46B0 , 32'hFFFC1595 , 32'hF22FB1C0 , 32'h03A04890 , 32'hF6EA4770 , 32'h14FF19A0 , 32'hFF7BD9D4} , 
{32'hE9511720 , 32'hF9298CF0 , 32'hFB1B87C8 , 32'h00005385 , 32'h00017F9C , 32'hF3B3CA10 , 32'h0C1051C0 , 32'hFFED6F2E , 32'hFFFED011 , 32'h113A7300 , 32'h05066218 , 32'h089CF800 , 32'h1A3FAA00 , 32'h00F466F8 , 32'h04A74918 , 32'h15B76E40 , 32'h085D5740 , 32'h0104CB2C , 32'h06DF43D0 , 32'hFFFF93F8 , 32'hFB3ABB88 , 32'h09056130 , 32'h1701D460 , 32'h00002E36 , 32'hF30DAFD0 , 32'h064CE178 , 32'hFCB29CF8 , 32'hF9A02968 , 32'h08B24420 , 32'h1AB02B60 , 32'h0E134B00 , 32'hFB7345D0 , 32'h103FA440 , 32'hF09FAC70 , 32'h0002DF72 , 32'h0043BFEE , 32'hEFBE5A20 , 32'hFE292A80 , 32'h0337FB80 , 32'h05580488 , 32'h06CFF788 , 32'h01FE2654 , 32'h0146FA88 , 32'hFB2CA8F8 , 32'h0CC25A60 , 32'h048C3068 , 32'hFA387EE8 , 32'hEACCC320 , 32'hFC0F4E98 , 32'hFE2160E4 , 32'hFBB64890 , 32'h040D7C88 , 32'hE4975680 , 32'hFC2710E4 , 32'h06B63B18 , 32'h03B07508 , 32'hFDEC426C , 32'hFAED6048 , 32'hE7835340 , 32'hDFB21A00 , 32'hFD1BF9C4 , 32'h045DAEF8 , 32'hF7396B00 , 32'h0877CBF0 , 32'h01C52224 , 32'hE5B7DB00 , 32'hFFFEEEE2 , 32'hF83AF588 , 32'hFF7244BA , 32'h12CA6CE0 , 32'hFECA2A14 , 32'h0A309C90 , 32'h043B0350 , 32'h034CAC80 , 32'hF7EC8B80 , 32'h08BD6A60 , 32'hF265A180 , 32'h16E82DE0 , 32'h13D12FC0 , 32'h08923380 , 32'hF5939BB0 , 32'h0B1836E0 , 32'h0D631730 , 32'hFFFE0F03 , 32'hF728A220 , 32'h0BC19050 , 32'hF38D69A0 , 32'hEB25C2A0 , 32'hFEF0EBD8 , 32'h00001949 , 32'hF1123020 , 32'h03D44280 , 32'h02E2D578 , 32'hFE2E3E40 , 32'hFFFDB923 , 32'hFA71C1D8 , 32'h313BC080 , 32'hE912AFA0 , 32'h05DD3988 , 32'hE7C45940} , 
{32'h05912C90 , 32'h1A1C6860 , 32'hF4330D00 , 32'hFFFE7E78 , 32'h00013129 , 32'h004BB525 , 32'hFF60C718 , 32'hFDE205AC , 32'hFFFF6D04 , 32'h117AA7C0 , 32'h0D4B0E60 , 32'hFFB0070A , 32'hF6DB4C40 , 32'hFBF4D400 , 32'hF786E510 , 32'hE45BF7A0 , 32'h14E01720 , 32'h0D01B540 , 32'hFB973830 , 32'h0002E0CE , 32'h03FE4C7C , 32'h1A5E52C0 , 32'h01177D14 , 32'h0001B573 , 32'hF33310B0 , 32'h011C6A28 , 32'hF621D4C0 , 32'h021B2F28 , 32'h05FE3020 , 32'h05F54EF0 , 32'hED151720 , 32'h09DD4E40 , 32'hFF11398A , 32'hEB03FC40 , 32'hFFFCCED2 , 32'hF52BC970 , 32'h0122D6A0 , 32'h14AB3DE0 , 32'h093AC110 , 32'h0DBACF50 , 32'hF9EEF268 , 32'hFFA8AC43 , 32'h04FEBC18 , 32'hFE0C8C2C , 32'h07369E38 , 32'h1ED56D80 , 32'h055E7570 , 32'h0BB2BD90 , 32'hFC0C6920 , 32'h20937D00 , 32'h1162BAA0 , 32'hD89A6940 , 32'h0172DCDC , 32'hEE003F60 , 32'h107CEF60 , 32'hFA2813A0 , 32'h0D670C50 , 32'hF3B39BE0 , 32'hFCC4FEEC , 32'h0C877CD0 , 32'hE9E805C0 , 32'h01CB14D0 , 32'h046138B8 , 32'h0AC60D90 , 32'h08393720 , 32'hF5747A10 , 32'h00028323 , 32'hF99B3680 , 32'hFEEEFC60 , 32'hFB317950 , 32'hFC26B994 , 32'h016122EC , 32'h00AB49FC , 32'h065A8D40 , 32'h0A42B4D0 , 32'h121E6FC0 , 32'h03DFECDC , 32'h04604318 , 32'hFF48E099 , 32'hFBD1B608 , 32'hF73AFBA0 , 32'hE827C960 , 32'hF9632780 , 32'h00007C36 , 32'h03C66210 , 32'h055415E8 , 32'hFB752728 , 32'h03EE2A00 , 32'hFEE18988 , 32'h000073F1 , 32'h0341BD40 , 32'h025F862C , 32'h01528654 , 32'hF52FD3F0 , 32'h0001F431 , 32'hF31F03D0 , 32'hF52E5720 , 32'hCE84E840 , 32'h03E6E008 , 32'h12EB1880} , 
{32'hF359BF20 , 32'h15EA65E0 , 32'h062E3258 , 32'h00011548 , 32'h00000380 , 32'hEE4E9900 , 32'hEBDB5200 , 32'hFBF7F278 , 32'hFFFF58C3 , 32'hF77FCDD0 , 32'hFEA45E88 , 32'h180DCDE0 , 32'h00C5A049 , 32'h125322A0 , 32'h03DB06A4 , 32'h14345220 , 32'hF094B200 , 32'h00F4F55B , 32'h1F8DBB20 , 32'h0003A7AC , 32'h004B3223 , 32'hF9869050 , 32'h04AC4070 , 32'hFFFEE444 , 32'h05E50918 , 32'hFD6F841C , 32'hF44D8CE0 , 32'hFD0CF89C , 32'hFBE39800 , 32'h0F013260 , 32'h05588E18 , 32'hFB0C8A88 , 32'h07FD3BB8 , 32'h0B452150 , 32'h00006219 , 32'hED9FC0E0 , 32'hF62FB2F0 , 32'h05085198 , 32'h0B8E26A0 , 32'hF6332390 , 32'hEB6F9EC0 , 32'h006DE9A1 , 32'h04130C00 , 32'h04535F10 , 32'hFDD55318 , 32'hE9D497A0 , 32'hF5C7CCD0 , 32'h05333340 , 32'h0D575D40 , 32'h0D5510D0 , 32'h0971E120 , 32'hF6EACAE0 , 32'hF7C392C0 , 32'hF02B7CD0 , 32'h03E0A2B0 , 32'hE9BB7A00 , 32'h13583AA0 , 32'hF1AB1B70 , 32'h185C2E40 , 32'h054C32A8 , 32'hFE143B6C , 32'hF8D1A9A8 , 32'hE3003F80 , 32'hF8D8E2F0 , 32'hFC7B9A64 , 32'h055277C8 , 32'h0004B371 , 32'h0D756E30 , 32'hFE318C24 , 32'h04222060 , 32'h0AB4BC50 , 32'h0970CC70 , 32'hF1A30B90 , 32'h04B2E450 , 32'h06E6A678 , 32'hF6333850 , 32'h08A1C7E0 , 32'hFA9E1530 , 32'hF6BCD5D0 , 32'hD6BBE080 , 32'hEEFDBAA0 , 32'hE065AD00 , 32'hF2F5C960 , 32'h00023F40 , 32'h0355AFA8 , 32'hF153CF80 , 32'h09612AE0 , 32'hFCE76B10 , 32'hF5C5D9B0 , 32'hFFFD699B , 32'hFFD9E278 , 32'h00C98ADA , 32'h081D0C60 , 32'hFE220638 , 32'hFFFF5D96 , 32'h0E333EC0 , 32'h22D5E940 , 32'h0859E5C0 , 32'hF8A2B560 , 32'h0A111D90} , 
{32'h02633858 , 32'hFC9D0EE8 , 32'h001B6A30 , 32'hFFFE0D4B , 32'h0001D81E , 32'h06A71B70 , 32'h099823A0 , 32'h070542A8 , 32'h00003769 , 32'h2491D180 , 32'hFA0B7378 , 32'hE0EF15A0 , 32'hF7807F80 , 32'hE1419660 , 32'h18F91220 , 32'h0A063FC0 , 32'h08C7D650 , 32'h08A488A0 , 32'hFBBD0B68 , 32'hFFFFAF7E , 32'h1F03C120 , 32'hFCB52D90 , 32'hEED076C0 , 32'h00024DB8 , 32'h2DE2EB80 , 32'hF2AA72B0 , 32'hF063D1F0 , 32'hFFA9630A , 32'h17A10AA0 , 32'hFCB324CC , 32'hFCEE4234 , 32'hFCE72608 , 32'hFBB6A320 , 32'h0E31CB00 , 32'h00000C64 , 32'hED779280 , 32'hF8DEE218 , 32'hF4776800 , 32'h03C64D20 , 32'hFF0C2274 , 32'h286C4500 , 32'h00600E74 , 32'hFF926666 , 32'h011D5700 , 32'h04DA5880 , 32'hEFC3E160 , 32'h0AFA8690 , 32'hF3209840 , 32'hF848ACD8 , 32'hF1984970 , 32'hF8558490 , 32'hFBB192F0 , 32'hF52DD3F0 , 32'hFB8367E0 , 32'h080A86F0 , 32'hFA14A710 , 32'h0FAC4C80 , 32'h121E7180 , 32'h1024C1E0 , 32'h0B3C0310 , 32'hF55BE9A0 , 32'h034D5928 , 32'h08097A00 , 32'hFACBEF48 , 32'h0683EDB0 , 32'h1218A700 , 32'hFFFB6687 , 32'hF5EF1340 , 32'hF86749C0 , 32'hFC3CC970 , 32'hF61DB220 , 32'h09E8A480 , 32'h0BFF5980 , 32'h042A31C8 , 32'h031B164C , 32'hF67F42B0 , 32'hFD203BA0 , 32'h01827F18 , 32'h09E22050 , 32'hEDBF3BC0 , 32'h06D15B20 , 32'hF2C0EE40 , 32'h01175ADC , 32'hFFFD9258 , 32'h0682A348 , 32'h013999A8 , 32'hFC426CB0 , 32'hF879A320 , 32'h01E3138C , 32'h00014C10 , 32'hF538C480 , 32'hFB18C920 , 32'h050B6ED0 , 32'hEF876520 , 32'h000406C4 , 32'h0810CC00 , 32'h121DDD00 , 32'hF35A7F70 , 32'hFBCB1BC0 , 32'h0557D198} , 
{32'hFCC4079C , 32'hFA3BDDA8 , 32'hFDC09EDC , 32'hFFFE0C4D , 32'hFFFEC3D9 , 32'hF5026ED0 , 32'hF59639C0 , 32'h00D408A8 , 32'h0002240A , 32'hFC65836C , 32'h03DA6250 , 32'hE51D7FA0 , 32'hE1076060 , 32'h0AE26E50 , 32'hEFB3F920 , 32'h08F4C3B0 , 32'hFDE1E4A4 , 32'hE6188C80 , 32'hFA5B7DC0 , 32'h0000C613 , 32'h10C9CF80 , 32'h009D440B , 32'h0D286490 , 32'h00028E06 , 32'hFB308950 , 32'hF3703D00 , 32'hF9FCBB68 , 32'h065507B8 , 32'h0088AC1C , 32'hE7C54E80 , 32'h16CE9D20 , 32'h01265F3C , 32'h1BB2D7A0 , 32'hEE1306A0 , 32'hFFFF9657 , 32'hFCEBE568 , 32'hF835F2B0 , 32'h0E417E80 , 32'hFC524EAC , 32'h05A0E800 , 32'hEB687780 , 32'h00C99202 , 32'h06827748 , 32'hE8D1C840 , 32'h034A66C8 , 32'hF5E1C650 , 32'h05535AA8 , 32'hFD3F6004 , 32'hF9C57180 , 32'h0C65F230 , 32'hE32C38C0 , 32'h1F9A6080 , 32'hFB293470 , 32'h0F1F3520 , 32'h099FA120 , 32'hFC7983E0 , 32'hFE82C034 , 32'hF7D493F0 , 32'h0B86A200 , 32'hF1BC3360 , 32'hF4B9E740 , 32'hFDB782CC , 32'h1372E0C0 , 32'h093CEA10 , 32'hF602BC30 , 32'h195EC340 , 32'h00018864 , 32'h116DE3E0 , 32'h04580568 , 32'h046CCA50 , 32'h02650D40 , 32'h09C2F230 , 32'h0C990950 , 32'h046EC1D0 , 32'h0BB8BE60 , 32'h08B12790 , 32'h03FCAD1C , 32'hF6E32550 , 32'h02ABBDB4 , 32'hF67B6C30 , 32'hEEDD87A0 , 32'h16AB6860 , 32'hF5A44C00 , 32'h00055DE1 , 32'h1C368EC0 , 32'hFD98DFC4 , 32'h0ADF87C0 , 32'hFD42995C , 32'h1473FFC0 , 32'h000293E3 , 32'h110D7920 , 32'h065BEBF8 , 32'h076D8F28 , 32'hF734EE20 , 32'hFFFE0CFB , 32'hF1836A60 , 32'h0790A7C0 , 32'hE724B500 , 32'h01ECDBD8 , 32'h0894BCE0} , 
{32'h04022010 , 32'hFCA9B0B4 , 32'h09595120 , 32'hFFFFDC8C , 32'hFFFDB310 , 32'h0EB5C310 , 32'h01E7DBD0 , 32'hF88B7850 , 32'h0000B780 , 32'hFE0DEB5C , 32'h09FF15E0 , 32'hF21CDA90 , 32'hF97728A8 , 32'hFB5951E0 , 32'h04EB2CF0 , 32'h052B7F20 , 32'h0EF053E0 , 32'h0BB297B0 , 32'h06F33468 , 32'hFFFF6B04 , 32'hF2D047F0 , 32'h1A92F220 , 32'h1CB1D240 , 32'hFFFEFC4C , 32'h1DF2D420 , 32'hF93018A8 , 32'h004C431B , 32'hFD67E2F0 , 32'hECC49740 , 32'h104EACC0 , 32'h139C71E0 , 32'h013538A8 , 32'h0B090F50 , 32'h014C3AF8 , 32'hFFFDFD52 , 32'hFFBC7B19 , 32'hFCBED614 , 32'h04C6A6B0 , 32'hF7453CC0 , 32'hF6618E90 , 32'hFDF2D874 , 32'hFEDAEE84 , 32'h0B1FCDB0 , 32'h051E0D10 , 32'hEF9F78E0 , 32'h0912DD30 , 32'hF4A536C0 , 32'h2472F500 , 32'h013CC894 , 32'h1427BCC0 , 32'h12EFD300 , 32'h0109E9A8 , 32'hFEC35C78 , 32'h1C24D1A0 , 32'h0D50E450 , 32'h071F13A8 , 32'h1CA68E40 , 32'h14DCBAC0 , 32'hFDD0E8FC , 32'h06826280 , 32'h16DE82E0 , 32'hFEBF1B18 , 32'h063E2AB8 , 32'h08668210 , 32'hF37A1410 , 32'hFF973668 , 32'h0003ACCA , 32'hFF3CDE76 , 32'h01C08124 , 32'h0FAD3D80 , 32'h01574E98 , 32'h0B555FF0 , 32'h130400A0 , 32'h044995F8 , 32'h0E8D57F0 , 32'hFDB231BC , 32'h0258AD0C , 32'h14E2A360 , 32'h0DE57910 , 32'h12D60DA0 , 32'hFCD6C23C , 32'hF1C3BDF0 , 32'h1A4C1D00 , 32'hFFFE13D3 , 32'h1B4B5660 , 32'hFE1DAEF4 , 32'hF81A21B0 , 32'hF28E7CD0 , 32'hF99A2DF8 , 32'h0000FB97 , 32'h0DF77D50 , 32'h0AEA46C0 , 32'h0090B5C3 , 32'h04CA73A0 , 32'h0000AB89 , 32'h01C6B79C , 32'hFDFFA2B0 , 32'h1D07B5C0 , 32'hF2C8E410 , 32'h07C8CD68} , 
{32'hEA44FFA0 , 32'h0F1B6840 , 32'h09E669C0 , 32'h000096B0 , 32'hFFFF03D4 , 32'h00EC96AE , 32'hFD81018C , 32'h063A73F8 , 32'hFFFF59AE , 32'h2662E5C0 , 32'h05E14868 , 32'h06BF35B8 , 32'hDE869F40 , 32'h05EFB7E8 , 32'hFC25ED08 , 32'h0286C040 , 32'h1311ABE0 , 32'hEE824E80 , 32'h0853D5C0 , 32'hFFFC6B1E , 32'hEAB7EA20 , 32'h18CBBD00 , 32'hF2323120 , 32'hFFFD8EB4 , 32'hF43E9380 , 32'hFAEA5C20 , 32'hF6498440 , 32'hFF865FDB , 32'hFEB81CE4 , 32'h05C87E48 , 32'hF5BD4D60 , 32'hF905E148 , 32'hEFB5A2C0 , 32'hFA15F540 , 32'h0000C034 , 32'h05793B48 , 32'h06753418 , 32'hF8722C60 , 32'h043F2128 , 32'hF0B5A1E0 , 32'hEE662380 , 32'h0082ABFC , 32'hF8793B18 , 32'h04A772E0 , 32'hE2AF4240 , 32'hECB8E6A0 , 32'h171D2080 , 32'h15C924E0 , 32'h027676F8 , 32'hF9CB08D0 , 32'hEDBB47E0 , 32'h275CA400 , 32'hFDFC0FB4 , 32'hEA215380 , 32'hFA0056F0 , 32'hF491EFA0 , 32'h0B874BD0 , 32'h0FD60710 , 32'hFC724C2C , 32'hF9067950 , 32'hF64BFB20 , 32'h02C61638 , 32'h09CC4960 , 32'hF7BFFD40 , 32'h0CDA6690 , 32'hF6899F70 , 32'hFFFE956E , 32'h0A8F4330 , 32'hF74F4000 , 32'h047E9528 , 32'hE9E01560 , 32'h017F3D50 , 32'hFBDDC100 , 32'h058F9C18 , 32'hFE17AD80 , 32'h0D09F810 , 32'hFA602060 , 32'hF4E692E0 , 32'h02F5B998 , 32'h0C551870 , 32'hF82454B0 , 32'hF280A1A0 , 32'h04AA6D48 , 32'hFFFFDEBF , 32'hE5555B40 , 32'hF69BFE40 , 32'hEDBE8F40 , 32'hEE7A0C60 , 32'h059343F0 , 32'hFFFE6233 , 32'h02EDD974 , 32'hFE14D0B0 , 32'hFB478170 , 32'h038D8F58 , 32'hFFFE8DA3 , 32'h0FA29340 , 32'hF467C740 , 32'h04A6B520 , 32'h03912CA4 , 32'hF7132D70} , 
{32'h06D0C790 , 32'h049598B8 , 32'h16BCC620 , 32'h00004368 , 32'h00027E1E , 32'hFC4A838C , 32'hF99E6628 , 32'hF4C67A30 , 32'h000090E0 , 32'h02422B08 , 32'hF4156FC0 , 32'h0AA3EE90 , 32'h0A476960 , 32'hF2C93AC0 , 32'hE42CBF60 , 32'h00878AE4 , 32'hE50DB620 , 32'h085A6030 , 32'hD5B53C00 , 32'h00040C97 , 32'hE31741A0 , 32'h035DB7F8 , 32'hF2E23900 , 32'h0000E122 , 32'h0205C5EC , 32'hFD385B64 , 32'hF2A54BC0 , 32'h09927E30 , 32'h146D4200 , 32'hDCC20D80 , 32'hF514AA80 , 32'hF305C9E0 , 32'h17A86740 , 32'hF31EFE50 , 32'hFFFEC8F7 , 32'hE1ADB7E0 , 32'h0B07C2A0 , 32'hF69CB7A0 , 32'h03491820 , 32'hFB7D17D0 , 32'hF8FA0580 , 32'hFFDCD35B , 32'hFFDADF3D , 32'h034FF68C , 32'hF84B4930 , 32'hFB7BE060 , 32'h036D1B5C , 32'h0420D410 , 32'hEEE80AA0 , 32'hF7F37210 , 32'h07E9B218 , 32'hFE837624 , 32'h05995238 , 32'hEFC72740 , 32'h0B3570F0 , 32'hF851A6D8 , 32'h161E1FA0 , 32'h09483FB0 , 32'hEA78CD60 , 32'hF93D9598 , 32'h1406EB40 , 32'hF7A0E640 , 32'h03FDD8E4 , 32'hFA4BF498 , 32'h01B42294 , 32'hF97FE108 , 32'hFFFDA614 , 32'h08ABD1D0 , 32'hF9C74398 , 32'hFAF2A000 , 32'h0BE6B6F0 , 32'h0459D1F0 , 32'h04788310 , 32'h03007B30 , 32'hEC9D6380 , 32'h0742E630 , 32'hFB0C6F28 , 32'h23BBB800 , 32'hF8A91848 , 32'h0285E0EC , 32'h06579DA0 , 32'h025AF638 , 32'hF1C416A0 , 32'hFFFE9745 , 32'h1902A480 , 32'hE9CF1060 , 32'hFF83AE91 , 32'hFE119E4C , 32'h03B19358 , 32'h00010D41 , 32'hF81410F8 , 32'h0072ED68 , 32'hFDE51544 , 32'h07EAC828 , 32'hFFFF7E16 , 32'h09AD06F0 , 32'h0AC9D0C0 , 32'hFE19D058 , 32'h036B8DC0 , 32'hFD222F54} , 
{32'hFDD1C334 , 32'hFBBD9560 , 32'h0141B9F4 , 32'hFFFFBD77 , 32'h0001D516 , 32'hF5342FD0 , 32'hF9F835B0 , 32'hF810F9E8 , 32'hFFFF5CB6 , 32'h0487E6B8 , 32'h0ED91D10 , 32'h0514F510 , 32'h191C1EE0 , 32'h039EE8DC , 32'h047EDBF0 , 32'h0650E670 , 32'hF4E7D2E0 , 32'hEF1E0B00 , 32'h2371BB80 , 32'hFFFDFA59 , 32'h00B2182B , 32'hF40B64E0 , 32'hFF733BA3 , 32'h0004B997 , 32'hFBA6C010 , 32'hF3D0A2B0 , 32'hF4FD6620 , 32'hFA667578 , 32'h13A48680 , 32'hF408ABC0 , 32'hDCDC8140 , 32'hE1A5F2C0 , 32'hFD1650BC , 32'hF4C7A740 , 32'hFFFEEF19 , 32'h18CAA5C0 , 32'h0B752250 , 32'hF8E719D0 , 32'hEFE2DDC0 , 32'hF78D8D70 , 32'h02AED97C , 32'h00235E5B , 32'h007D3AAF , 32'h059B8728 , 32'hDE92EB40 , 32'hF7E7DDD0 , 32'hEBD3B360 , 32'h0C635A60 , 32'h1539C660 , 32'h05587FA0 , 32'hF643EB50 , 32'hFBA7E660 , 32'hF29E8920 , 32'h12945980 , 32'h08532230 , 32'h161F4D40 , 32'hF8A64EB0 , 32'h0FA8B430 , 32'hF9E26908 , 32'h0B7EEFD0 , 32'h09045BD0 , 32'hF6158000 , 32'h142C3200 , 32'h01E4E60C , 32'h05CF05B0 , 32'h0053B849 , 32'h00004CBC , 32'hFF78EF57 , 32'hFF343286 , 32'hFAEDFFA8 , 32'h0385D5E0 , 32'h0010439F , 32'hFFE92E21 , 32'hFABF0C30 , 32'h07DDDC08 , 32'h08D836B0 , 32'hFD6C18DC , 32'hFC4CC44C , 32'h03004358 , 32'hFCE56EFC , 32'h0E7D1D30 , 32'hF7FB33F0 , 32'hFB188AB0 , 32'hFFF9C47C , 32'h1187FA40 , 32'hF5E8AB50 , 32'hE6306360 , 32'h19F33BE0 , 32'hF46DBBB0 , 32'h0001B000 , 32'hFD7C73C4 , 32'h03D59984 , 32'hFA631468 , 32'hE701CA00 , 32'h00054131 , 32'hE56BCE20 , 32'h0B2B8F00 , 32'hEFC13680 , 32'h11965C60 , 32'h0648A528} , 
{32'h106DDDA0 , 32'h10887440 , 32'h140609E0 , 32'h000326B3 , 32'h00035207 , 32'hEA88C360 , 32'hE7D20220 , 32'hFEC98A58 , 32'h00049D73 , 32'hEE0A6B20 , 32'hFF5DCC94 , 32'h0F0EEC30 , 32'hF143FD90 , 32'hF25ED450 , 32'hFBF40658 , 32'hFF437CBD , 32'h0AF09F40 , 32'h046DCBA8 , 32'hFE50AACC , 32'h0000AF03 , 32'h0685E7A8 , 32'h09345260 , 32'hEC7F35C0 , 32'hFFFEF445 , 32'h077ED558 , 32'hF9CB1930 , 32'hF6FD4470 , 32'h0C489A80 , 32'h047DB758 , 32'hEF2A9A60 , 32'h0DD8C070 , 32'hFA91DE30 , 32'hF9ABB8E8 , 32'h0337EDF8 , 32'h00015A15 , 32'hF0C03680 , 32'hFFEC8A6F , 32'h065030F0 , 32'hF8852180 , 32'h1504F1E0 , 32'hF9FB8158 , 32'hFF79EE42 , 32'h00E52D81 , 32'h02AAAC7C , 32'hF0251BF0 , 32'hE0A4E000 , 32'hFC26D308 , 32'hFD959710 , 32'hEA02C060 , 32'h0A648810 , 32'h013E4D0C , 32'hF1952120 , 32'hF99BF9E8 , 32'h1EAC2C20 , 32'hEE2A0D40 , 32'h00C49760 , 32'hE7C92000 , 32'hFF1DC329 , 32'hEAE34040 , 32'hF5BEF8F0 , 32'hFDBCBC58 , 32'hF8380228 , 32'h034B062C , 32'hFF8F2D5B , 32'h0EC67BE0 , 32'hED5B33A0 , 32'h0000C112 , 32'hF7A4BB10 , 32'hF3784C60 , 32'h18EB5900 , 32'hF475E4E0 , 32'h08213AE0 , 32'hEFAA86E0 , 32'hFB7D4120 , 32'h00A34C90 , 32'hF95F8AF0 , 32'hFE921950 , 32'h06427990 , 32'h186EA840 , 32'hE9308140 , 32'hF903E870 , 32'hF7DC28E0 , 32'h1E39FBC0 , 32'h000356D6 , 32'hF2686540 , 32'h1DB55FC0 , 32'hFA76A648 , 32'h12949F00 , 32'h0DD3C300 , 32'h0000E100 , 32'hF83974E8 , 32'hFE2711E0 , 32'h10172940 , 32'h03A732EC , 32'h0000B112 , 32'hF1805C20 , 32'hF6971B30 , 32'h0661D1C8 , 32'hF973C8D0 , 32'h01303C10} , 
{32'hF423E300 , 32'h01FE0C98 , 32'h01670108 , 32'hFFFC8215 , 32'h00017126 , 32'h11801460 , 32'hFFFFCF77 , 32'hF142E8D0 , 32'h0000EC94 , 32'h11B24000 , 32'h0290B2E4 , 32'hF5E4EF30 , 32'hF19FDDE0 , 32'hF62D04E0 , 32'hFEBED440 , 32'h0E9F3B70 , 32'h0019F6C1 , 32'h0BC046B0 , 32'h090A5980 , 32'hFFFAA0D4 , 32'h0EED3E90 , 32'hFBE28B80 , 32'hEAAAD900 , 32'h00025C5A , 32'h0EC691F0 , 32'h090CE950 , 32'hEF283320 , 32'h028F04C8 , 32'h0284F340 , 32'h059FBEE0 , 32'hF500E580 , 32'hF87A4AB8 , 32'h0B32EC30 , 32'h00800FA4 , 32'h0000104D , 32'hFFB37E46 , 32'hFF9E9D98 , 32'h05BDD7D0 , 32'h0C7DAE80 , 32'hFD983318 , 32'hE99104C0 , 32'h009D521D , 32'hF7DF0080 , 32'h0EDDD6A0 , 32'h09BE18E0 , 32'hF42BBF50 , 32'h0AD1C140 , 32'hFD035A80 , 32'h1DFC6560 , 32'h19FA53C0 , 32'h15051840 , 32'h03CF9D4C , 32'h10F79D80 , 32'hF6409FC0 , 32'hF37903E0 , 32'h02F512AC , 32'h04F594D0 , 32'hEF747200 , 32'hEF6B2AA0 , 32'hDF5EF380 , 32'h0D24F210 , 32'h06585070 , 32'h0B6DDB40 , 32'h0AD76610 , 32'hFDA8C318 , 32'hFCDDD0A0 , 32'h0000ADB1 , 32'hFC0ADB64 , 32'hFC7C5308 , 32'hEE7AC4C0 , 32'h0CDCF500 , 32'hF7158A40 , 32'hF7D00270 , 32'hFAAA9E78 , 32'h0E203B90 , 32'h02A3F5EC , 32'hF9990510 , 32'hFD83DAAC , 32'hFFEAFEA6 , 32'hED2D2C40 , 32'h06FB40F8 , 32'h2D93B580 , 32'h0576D1C0 , 32'hFFFF36C6 , 32'h07F89D88 , 32'h0D5549F0 , 32'hFDE4943C , 32'hEEF166C0 , 32'hD942F180 , 32'hFFFE6D43 , 32'hED119120 , 32'h06673920 , 32'h05B06F00 , 32'h0134A338 , 32'h00006A9E , 32'hEB96C800 , 32'hEFEAA4E0 , 32'h0F20C430 , 32'h04F06DB8 , 32'h06FE2E60} , 
{32'h012741E8 , 32'hFBE48188 , 32'h131C4AC0 , 32'h0004B683 , 32'hFFFFAF3B , 32'h02B24E88 , 32'hF94D9E40 , 32'hFCCBFFE4 , 32'hFFFCEA40 , 32'h0E065F90 , 32'h09E4E2F0 , 32'hF02DECB0 , 32'hF339B0D0 , 32'h060B9E10 , 32'hF79A01F0 , 32'h18828680 , 32'hF9F9F538 , 32'hF87DC648 , 32'h00C36E65 , 32'hFFFED736 , 32'h2A1EB380 , 32'hF9528F90 , 32'h01AB896C , 32'h00029ED9 , 32'h0C7E1D90 , 32'h02B45BF8 , 32'h09D86D40 , 32'hF33C11F0 , 32'hFAD607A8 , 32'h04AE3148 , 32'hF14DF520 , 32'h0B127F30 , 32'h024D2B64 , 32'hE37A91A0 , 32'h00003F6F , 32'hF7416190 , 32'h0343F2AC , 32'h0B5F03B0 , 32'hF1AB4D90 , 32'hFBBA5000 , 32'h072F9278 , 32'h02FC60D0 , 32'h00E0A53B , 32'h0FEC00A0 , 32'h0A9D6540 , 32'h0CBBECF0 , 32'hDCBD53C0 , 32'hFFEE6C5F , 32'hFBDEFFB0 , 32'hF8646420 , 32'hF87E6290 , 32'hEBF8B720 , 32'hFB5B0710 , 32'hFA2D8EE0 , 32'hFE330CD8 , 32'hFC2B01DC , 32'h02B35710 , 32'hEFAA3B20 , 32'hF7F14CB0 , 32'hFDB81C18 , 32'h1AA32540 , 32'h1011F040 , 32'h0C3A4CD0 , 32'h000D4A06 , 32'h1AE000E0 , 32'h0AAA40B0 , 32'hFFFEB2F8 , 32'h1151B660 , 32'hF9F51D88 , 32'h1C910520 , 32'h1181AC60 , 32'h049BA120 , 32'hF51ECE80 , 32'h05E04EB8 , 32'hFBA2DA48 , 32'h03DE09F8 , 32'h0109AB8C , 32'h07D7B110 , 32'hF007C110 , 32'hFF281BCB , 32'hFB89C800 , 32'hFB2A15C0 , 32'hF0C82B00 , 32'hFFFF196E , 32'hE4CD13A0 , 32'hF7792430 , 32'hE4AB5620 , 32'h04763628 , 32'h064B6938 , 32'h00023415 , 32'h1754CC40 , 32'hFFABC254 , 32'h0191F858 , 32'h171654C0 , 32'hFFFDD6DA , 32'h06A6CEB0 , 32'hEF11DA40 , 32'h05A28478 , 32'hFE883D9C , 32'hEA22DC00} , 
{32'h07382DD8 , 32'hF5982010 , 32'hF3F68B30 , 32'hFFFB2206 , 32'h0001FF1A , 32'h170666E0 , 32'hF72E1850 , 32'h014DA2F4 , 32'hFFFF1DF1 , 32'h132AF2E0 , 32'h0A8C5FE0 , 32'h068CA468 , 32'h022F6564 , 32'h12C348A0 , 32'hF439D980 , 32'hE5DE8480 , 32'hFBA581B8 , 32'hD08CA500 , 32'hFE91952C , 32'hFFFCEC09 , 32'h0A146C60 , 32'h08F0E330 , 32'hFEFA51EC , 32'h00018502 , 32'h12BD0740 , 32'hEFC66740 , 32'h0CBC7FB0 , 32'h0C2B9820 , 32'hFEE920FC , 32'h05A27320 , 32'hF7CF1120 , 32'hE99EC7C0 , 32'h1328FD80 , 32'hF910ED70 , 32'h0002EAC2 , 32'hF5E4E000 , 32'hFD1D2818 , 32'h12452D20 , 32'h0F853D50 , 32'hFFEF6926 , 32'h0997E330 , 32'h005C4330 , 32'hF9855118 , 32'hF2902590 , 32'hEAAB5D80 , 32'hFF56F8CD , 32'hFFCFC22F , 32'hF0B1FB60 , 32'hF1027C30 , 32'hF0B736B0 , 32'h09C4CAC0 , 32'hED56E4E0 , 32'h16B66D80 , 32'h1124F220 , 32'hEFF75680 , 32'hF935E228 , 32'h16C5AC40 , 32'h022ED114 , 32'h0C67D580 , 32'hF9DB3D30 , 32'h08E56AE0 , 32'h00BDB9BE , 32'h065CDA18 , 32'h0D382B90 , 32'hF41ABF40 , 32'hDD5F88C0 , 32'h00013737 , 32'hFD453398 , 32'hFC819640 , 32'hFDF34E90 , 32'hEFD316C0 , 32'hF3619E40 , 32'hF8A6F208 , 32'hFE009530 , 32'hF4B1A5B0 , 32'hF940F808 , 32'h0736FCD8 , 32'hF231F6D0 , 32'hF94DB9F8 , 32'hFE9D3AC8 , 32'h039E1950 , 32'hFE88879C , 32'hF9D13338 , 32'h000564EE , 32'hF8156A40 , 32'h10FE1760 , 32'h109925A0 , 32'hFDC3F244 , 32'hF07EF800 , 32'h0002C06B , 32'h13B2D260 , 32'hFD6F0590 , 32'hFD38D308 , 32'h051A1930 , 32'h0002AC88 , 32'hF7742BF0 , 32'h1AD42240 , 32'h09959F30 , 32'h031580E4 , 32'hF5C50DF0} , 
{32'hD95B84C0 , 32'h006B9A50 , 32'h0758A080 , 32'h00014295 , 32'hFFFBD61D , 32'hFE4020F8 , 32'h06D76F70 , 32'h049F1AE0 , 32'hFFFCC17F , 32'h02D08450 , 32'hF5DBBD10 , 32'hF6112950 , 32'h0810D3C0 , 32'hFEBE8F1C , 32'h0EF486A0 , 32'hE49DEAE0 , 32'hF0290ED0 , 32'hFAE14DE0 , 32'h0395F284 , 32'hFFFD0F40 , 32'h02BE6F3C , 32'hF5C4C040 , 32'h07391EE8 , 32'h0000B889 , 32'h06E700B8 , 32'h0917DEB0 , 32'h089AA160 , 32'h0767C000 , 32'h00C8BC6F , 32'h01D28B8C , 32'hF72ED3E0 , 32'hE3D4C5C0 , 32'hFE4FD2C4 , 32'hF71378C0 , 32'hFFFE9722 , 32'hEBE15B60 , 32'hFFBCC246 , 32'hE1388560 , 32'h0A6EE320 , 32'h168BD400 , 32'hEB3B0500 , 32'hFFFB0156 , 32'hFCD4F630 , 32'h0CE7B9F0 , 32'h0D9519A0 , 32'h18D96480 , 32'hEFD794A0 , 32'h10123660 , 32'hED019B20 , 32'hF68A6F40 , 32'h10A521A0 , 32'h042D7D78 , 32'h0232DAE8 , 32'hFB28EBF0 , 32'h0202AC4C , 32'h08944BB0 , 32'hEDFD2F40 , 32'h086B1FA0 , 32'hF7844690 , 32'hEDEAD700 , 32'h009D0013 , 32'h01219488 , 32'h0D2920C0 , 32'h00159B42 , 32'h02582E90 , 32'hFC7669B0 , 32'h0001D364 , 32'h042CF630 , 32'h0BF81F90 , 32'hFB6CC508 , 32'hF9AA49E0 , 32'hF8AF7EB8 , 32'h012804A8 , 32'h0834AB50 , 32'h0E82BBB0 , 32'hFB239FE0 , 32'hF9D56A70 , 32'hF214E910 , 32'h055E2150 , 32'hED467260 , 32'hF74B2A50 , 32'h0223E860 , 32'h186E0020 , 32'hFFFCFD9B , 32'h01EB60BC , 32'hF96EFD20 , 32'h025FA77C , 32'h04F2F3E0 , 32'h0854A2D0 , 32'hFFFD70BF , 32'h22C7E800 , 32'hFAED9E88 , 32'h20DC2C40 , 32'hE7DBC880 , 32'h0002E972 , 32'h20713C80 , 32'hFCECE5B8 , 32'h037FDEB8 , 32'h0623E090 , 32'h093E6120} , 
{32'h06CF1198 , 32'hFA1AE5A8 , 32'hF5E980F0 , 32'h00001C0B , 32'h000349B1 , 32'h1AE8F7C0 , 32'h022EA364 , 32'h08879F70 , 32'h0003BA21 , 32'h035078EC , 32'hF2325420 , 32'hFDA81718 , 32'h063C4290 , 32'hF7BF0070 , 32'h03DF5DA0 , 32'hECA6C1E0 , 32'h0ADE2100 , 32'hEB52E8C0 , 32'h0975BA80 , 32'hFFFEDB41 , 32'hEC8CF6A0 , 32'hFE4D644C , 32'hE5772F80 , 32'hFFFF97D2 , 32'h074EEFE0 , 32'hF2C847C0 , 32'hFE00FE74 , 32'h01D4C6E0 , 32'hF1307DB0 , 32'h068C1F60 , 32'h1E150FE0 , 32'h0C5369C0 , 32'h20AF2A80 , 32'h0171AC60 , 32'h00014358 , 32'h0B4DAE40 , 32'hFC78BC54 , 32'h032AA35C , 32'hEB89EA20 , 32'h100D1300 , 32'hFC734778 , 32'hFD773D08 , 32'hEC5C5220 , 32'hFE3F6784 , 32'hE7B18480 , 32'hFFF9181A , 32'hF999E6C0 , 32'hED2BD140 , 32'hF31F6BF0 , 32'h0C0E62D0 , 32'h00CB86A6 , 32'h07C89290 , 32'hFFCCF9AA , 32'hEFADA6A0 , 32'h0771B7B8 , 32'h141E52C0 , 32'hFB40CE10 , 32'hEF9F8C60 , 32'hE53FEFC0 , 32'h11FDDD20 , 32'h0714BA80 , 32'h02D405AC , 32'hF36E7890 , 32'hFB92CF50 , 32'h0B397280 , 32'h184FEC80 , 32'h000077A3 , 32'hFEEE8000 , 32'hFEA5D38C , 32'hF6E0B1C0 , 32'h0B7CB220 , 32'hF0204C10 , 32'h0B56BE50 , 32'hF5858FD0 , 32'h05C97F38 , 32'hFB9DD410 , 32'hDE43DCC0 , 32'h0901F980 , 32'hF4F4AB90 , 32'hE41731A0 , 32'hEEED9140 , 32'hF44A8A00 , 32'h0BE0C870 , 32'hFFFD4BB6 , 32'hF06E7B70 , 32'hEBA61920 , 32'hF151D4B0 , 32'h031B6118 , 32'hF662C7C0 , 32'h0005C847 , 32'h073B7698 , 32'h04FD6FE0 , 32'hF883FAE0 , 32'h055161E0 , 32'hFFFC9095 , 32'h031C2A2C , 32'h06008FF8 , 32'hF7F1D4F0 , 32'h056BCE80 , 32'h04AE4390} , 
{32'h19A4B800 , 32'hF65BFC80 , 32'h0369D424 , 32'hFFFE2A27 , 32'hFFFE58E9 , 32'h0E4B0410 , 32'hF8ED5480 , 32'hFF9DEE8A , 32'h0001A74B , 32'h05680740 , 32'hFDBDD67C , 32'hFCB39858 , 32'hFDEC5254 , 32'hE54D8B60 , 32'hDFC69440 , 32'h03F1A178 , 32'hEE544640 , 32'hFAC8C6E0 , 32'h22B32CC0 , 32'hFFFE1CDD , 32'hFD58F060 , 32'h010568BC , 32'h00092856 , 32'hFFFF8EED , 32'hF3514500 , 32'h03429438 , 32'hEE75EDE0 , 32'h04550138 , 32'hE4C35C20 , 32'hF662A850 , 32'h07CD8038 , 32'h044ED070 , 32'hF6A634D0 , 32'h0D001C10 , 32'hFFFC9BFF , 32'h06C8C520 , 32'h07F79BB8 , 32'hDA2A64C0 , 32'h135B1520 , 32'hF9981FE0 , 32'h03B66000 , 32'h0008F23E , 32'h05BBC698 , 32'h133FE8E0 , 32'hF05A7F40 , 32'h1D9BED80 , 32'h012BCA40 , 32'hF7D55210 , 32'hF6416DE0 , 32'h09D1FA80 , 32'hED62F060 , 32'hE328B8C0 , 32'h017C5000 , 32'hFA6A1CB0 , 32'hFF90A310 , 32'hF845BCE0 , 32'hEFB81020 , 32'h15733F40 , 32'h00BAAB17 , 32'hEDC2E360 , 32'h08CE8C70 , 32'h0279A734 , 32'h0C6427F0 , 32'h0018D10E , 32'hE2A0C180 , 32'h11308D20 , 32'h0002D287 , 32'h01DA98E8 , 32'h01BE7FB4 , 32'h00C5BD07 , 32'h01A7460C , 32'h021D7D04 , 32'hFCB1CEA8 , 32'h0BC567E0 , 32'h059D8548 , 32'h08B30AA0 , 32'hF9ABD358 , 32'hF5E87A70 , 32'h0D91C730 , 32'hFD114B70 , 32'hEEE408C0 , 32'hF3289F30 , 32'hF1A81C90 , 32'h0000992E , 32'hFB30ABF0 , 32'h0BA4CFF0 , 32'h08E1BEA0 , 32'hE9A22F40 , 32'h01D28CD4 , 32'hFFFF1C31 , 32'hF6C61820 , 32'hFB795AF8 , 32'h0EA8F920 , 32'h112D39A0 , 32'h00022F23 , 32'hFB81DDF8 , 32'h08305CA0 , 32'hF8DB5070 , 32'h03B6CCE4 , 32'hF76CE7B0} , 
{32'hFA5E4230 , 32'hF74EA130 , 32'h01EAFC20 , 32'h0001B9FD , 32'h0000B212 , 32'hF2F0AA90 , 32'h0444B5E0 , 32'hFBE0DBA0 , 32'h00008E6B , 32'hF7E03B00 , 32'h01A7E2E0 , 32'hF9985878 , 32'h0E6EC570 , 32'h015F1AEC , 32'hED0D7B40 , 32'hE7B013C0 , 32'hEB1BC160 , 32'h0008A211 , 32'h060D4790 , 32'hFFFF25CE , 32'hFEC95B74 , 32'h1F973660 , 32'h0153FBA4 , 32'hFFFDB787 , 32'h170ADA20 , 32'hF7DB1F40 , 32'hFE717588 , 32'h07AC9440 , 32'h0EC4E960 , 32'hF19F0910 , 32'h1211E100 , 32'h03D09D28 , 32'hED60DAA0 , 32'hF0E17800 , 32'h00010F55 , 32'hF9F2CD08 , 32'hFBEB0818 , 32'h0FBF9780 , 32'hF25AE070 , 32'h00483B04 , 32'hF60F14F0 , 32'hFFD4814B , 32'h0040FC87 , 32'h10A2CB80 , 32'h0C650480 , 32'h08AD33E0 , 32'hFBE644E0 , 32'hE53460C0 , 32'h18483720 , 32'hF935B430 , 32'hEEA1CBC0 , 32'h0BA03E40 , 32'h088F1450 , 32'h048575B0 , 32'hF66AB450 , 32'hF2A31500 , 32'hFBD90CF8 , 32'h1ACC6360 , 32'hF19CDD10 , 32'h0CDA6C20 , 32'h00B89CE3 , 32'h0C1B2730 , 32'hDA117900 , 32'hFBC81F68 , 32'h1ABFDFC0 , 32'hFC664E8C , 32'hFFFE0841 , 32'hF2BBEBE0 , 32'hFF54F4FB , 32'hFC4E9FB0 , 32'h035F2048 , 32'h03A7D0CC , 32'hEBF51EA0 , 32'h0C00EC70 , 32'h1BD65880 , 32'h068026D8 , 32'hFA290D80 , 32'hE4D785C0 , 32'h12687520 , 32'h00A02EAC , 32'h09EC9140 , 32'hFC6F560C , 32'hFBF95950 , 32'h00006DED , 32'h132D3880 , 32'hFB218300 , 32'hFB4E82D0 , 32'hEC38ED00 , 32'hEDDAF900 , 32'h0002E77E , 32'h0ADB9A70 , 32'h049A56D0 , 32'hF77914D0 , 32'h0A02BE00 , 32'h00047AE6 , 32'h032A1D00 , 32'hFBEE9DD8 , 32'hF6856A50 , 32'hF3B9DFF0 , 32'hF67A58D0} , 
{32'h0D301140 , 32'hEA8002A0 , 32'h1758A640 , 32'hFFFF8AF6 , 32'hFFFD26C9 , 32'hFF401C62 , 32'h0F857840 , 32'hFABD4738 , 32'h0001FA9F , 32'h17B59F00 , 32'hFBE9F878 , 32'hEA125880 , 32'h0344AD38 , 32'hF7A80520 , 32'h0C39B2C0 , 32'h039CB120 , 32'hFC5D29D0 , 32'hF0BAD320 , 32'hE98D7120 , 32'hFFFF3E0D , 32'h0150C66C , 32'hFCF009E4 , 32'h12327320 , 32'h000240A6 , 32'h00B0203C , 32'h1991AB00 , 32'h0FC19230 , 32'h07F61D88 , 32'h034956B0 , 32'hF7CD9870 , 32'hFC5ECE94 , 32'h00E0B2A1 , 32'hF19CCC20 , 32'h16F0CE80 , 32'hFFFF7653 , 32'h0496B980 , 32'hFBECA7B8 , 32'h1A266F00 , 32'h02725CB4 , 32'hEAA7F0E0 , 32'hE3B53300 , 32'hFED34CEC , 32'hFAD54BB8 , 32'hFCABF470 , 32'hFBDB7FE8 , 32'hFD18C440 , 32'hFA1E6338 , 32'h03E0174C , 32'h10627BE0 , 32'h18D73980 , 32'hFE19E61C , 32'hF365FAF0 , 32'h0B7A0700 , 32'h033C3424 , 32'hFA8F8260 , 32'h12258B40 , 32'h086C1C50 , 32'hF62AF640 , 32'hF10DDD00 , 32'hEA1A1360 , 32'h040A5BA0 , 32'hF9A94988 , 32'hE115F240 , 32'hF588D3F0 , 32'hEE065480 , 32'hFED9D0F0 , 32'hFFFF0AF6 , 32'h027C6FA8 , 32'hFA1C3E10 , 32'hFF03EAC5 , 32'hEB3F59E0 , 32'h0EF26CC0 , 32'h0B8569A0 , 32'hF2A0D120 , 32'hEE314EA0 , 32'hFF9A2941 , 32'hE37B15C0 , 32'hEBAD5E40 , 32'h10A65A80 , 32'hF90EBBE0 , 32'hFF42FBBE , 32'hEB111600 , 32'hF1B58ED0 , 32'hFFFF1B1E , 32'hFF10F31F , 32'hF9BB7E58 , 32'hFE3C537C , 32'h18533F40 , 32'h0A7FD910 , 32'h00008E9B , 32'hFD1FA3E8 , 32'hF5F1A5B0 , 32'h0A7503E0 , 32'hF98A3A50 , 32'h000257AE , 32'h08983EA0 , 32'hFEB03684 , 32'hF5940FE0 , 32'hFC60F614 , 32'hF8280FD8} , 
{32'h10F363E0 , 32'h064EDF68 , 32'h0655FE70 , 32'hFFFFEF26 , 32'hFFFF1EEE , 32'h0A3F7910 , 32'h282F2C40 , 32'hEB6DA980 , 32'hFFFB101C , 32'hF7B655A0 , 32'hF84D45E8 , 32'hE7A509C0 , 32'h003D10E7 , 32'h01D51660 , 32'h1FCE7440 , 32'h11087260 , 32'hFE0CCBDC , 32'hFB294798 , 32'h0D39D470 , 32'hFFFC294A , 32'hF4D23C60 , 32'h042203B8 , 32'hF7FEF520 , 32'hFFFCF7E6 , 32'hEBD41D00 , 32'h03A6C3F8 , 32'hF8012AC0 , 32'hF83BC340 , 32'h04417250 , 32'h141E0080 , 32'h01739E30 , 32'hF249F840 , 32'hF13DEEC0 , 32'hED0CE6E0 , 32'h00049237 , 32'hDA5D5980 , 32'hEBD5D260 , 32'h0EB9F2E0 , 32'h16D2F220 , 32'h0702C1D0 , 32'h023898B4 , 32'hFEAEA9A8 , 32'hFF52D3DB , 32'hF18020C0 , 32'hDB38EE40 , 32'h0EA83B00 , 32'hF922E510 , 32'hF9489338 , 32'hF6711E30 , 32'hF3E10060 , 32'h07A50FB0 , 32'h027C6870 , 32'h02109664 , 32'hF27D9EA0 , 32'hEBBC2660 , 32'hFB055B10 , 32'hEFAD06A0 , 32'h0A1C2F70 , 32'hFC026890 , 32'h03C6819C , 32'hFC4BE580 , 32'hFA846E68 , 32'hF9A23FF8 , 32'hF921DC18 , 32'h02D2D248 , 32'hFF0925F1 , 32'hFFFD299B , 32'h1450D080 , 32'hFC0A71C8 , 32'hFE695860 , 32'h08BB3440 , 32'h0CEB1C70 , 32'h0375B8A8 , 32'h0BAFAF60 , 32'h03ACD0E4 , 32'hFBC029E8 , 32'h0BBED6D0 , 32'hF501FBF0 , 32'h0036BCFE , 32'hF9156C10 , 32'hFF4CDD8A , 32'h0A0DB820 , 32'h05DA2470 , 32'h000019D3 , 32'h13C7FB60 , 32'hFB915B70 , 32'h01B23B18 , 32'h0CDF3D70 , 32'h0BCB6270 , 32'hFFFEC303 , 32'hFBF79F10 , 32'h0590AC80 , 32'hF00AEBB0 , 32'h1EAC28C0 , 32'h0005044D , 32'hED0977C0 , 32'hFAE746C8 , 32'h01C59A44 , 32'h07FCD818 , 32'h0690EBC0} , 
{32'hFB075368 , 32'hF6B1FB90 , 32'h1686C6C0 , 32'h00000FC3 , 32'hFFFFD2ED , 32'h0287E500 , 32'h0006737A , 32'h12CF82A0 , 32'h0001B733 , 32'hE365B740 , 32'h1895DA20 , 32'hF0126360 , 32'h2E33C080 , 32'h051B8DC8 , 32'h0453E260 , 32'hFE7CD1D4 , 32'h12EE2900 , 32'h01A88364 , 32'hF20B97E0 , 32'hFFFC1863 , 32'h0E46C890 , 32'h05C5EF08 , 32'hEAC9A960 , 32'hFFFDC000 , 32'hEFBD9E20 , 32'hF884BE90 , 32'hEFC746C0 , 32'h0D584540 , 32'hF3D0CDD0 , 32'hF9326490 , 32'hF72330D0 , 32'h2373E540 , 32'hF8956B00 , 32'hE9918E40 , 32'hFFFDD775 , 32'hEAA4AEA0 , 32'h0CA1FE70 , 32'h0D36C8D0 , 32'h0D38AAC0 , 32'hED7BCF00 , 32'h0771D488 , 32'h010E1CF8 , 32'h006303C3 , 32'h058EF5E0 , 32'hF8227050 , 32'hF2D31AA0 , 32'h00DD0E08 , 32'h16EBE5A0 , 32'h01E72AC4 , 32'hF02F5C20 , 32'hF7A81DD0 , 32'h08A2BE70 , 32'hF7D17010 , 32'hFE6A6A58 , 32'hF9364750 , 32'h04ACA108 , 32'h132E2440 , 32'hF9E5E2F0 , 32'hF66D73D0 , 32'hF7E1DFC0 , 32'h0C119AC0 , 32'hFDC75268 , 32'h00B61611 , 32'hF78E2440 , 32'hEBAE3340 , 32'h0E9E3A70 , 32'hFFFD2A2B , 32'hFDEB4F00 , 32'h077112A0 , 32'h06D8E9D0 , 32'hFE58F5EC , 32'hF8BE0888 , 32'h04049838 , 32'h083D5E80 , 32'h12D67F60 , 32'hFB938568 , 32'h00976796 , 32'hF6294860 , 32'h01EFA370 , 32'hFD8FE79C , 32'hFB586270 , 32'hFB7C2720 , 32'h10442FE0 , 32'h0002B110 , 32'hED33CCA0 , 32'h02AA2010 , 32'h1B01A100 , 32'hFD157970 , 32'hE9BE6BA0 , 32'hFFFAF0A8 , 32'hFDE5AB74 , 32'hFF8A17EC , 32'h05C17FC0 , 32'hF48F8550 , 32'hFFFE8A9A , 32'h014693AC , 32'h05573200 , 32'hF4715260 , 32'h13B6F7E0 , 32'hFEC93CB8} , 
{32'hEC590C60 , 32'hF51AB140 , 32'h06D77030 , 32'h000478C1 , 32'h0001CE3D , 32'h0E955750 , 32'h0A5EDF50 , 32'hF7D13810 , 32'h0000BD5D , 32'h108239A0 , 32'hE6204B00 , 32'h091FACD0 , 32'hF5D81EA0 , 32'h188325C0 , 32'h06B1FF50 , 32'h0E450A20 , 32'hEB0009A0 , 32'h149E2A00 , 32'h0808A2B0 , 32'h0000D286 , 32'h0F31A270 , 32'h12643420 , 32'hF797FAA0 , 32'hFFFED9AB , 32'h048F3BF0 , 32'h025E97A8 , 32'hF485F5B0 , 32'hFF9FE31A , 32'hEE3B0AE0 , 32'hDAD4E600 , 32'hF172DD50 , 32'h19801680 , 32'h091A1680 , 32'hF07A4590 , 32'hFFFE5CAE , 32'h01DAA61C , 32'h073E2C18 , 32'hED4832E0 , 32'h024D7CA0 , 32'h18EBFB60 , 32'hFE3CDA74 , 32'hFEA4C3FC , 32'h02900D18 , 32'hF18935A0 , 32'hFF5B6DB2 , 32'h10C59E60 , 32'h043CD938 , 32'h0182B858 , 32'hF4886620 , 32'h06B99888 , 32'h0D1E9970 , 32'h026806E8 , 32'hECC0F2E0 , 32'h1A2EB240 , 32'hF15C8090 , 32'hFD083FF4 , 32'h0A5C1390 , 32'hF4F1C320 , 32'hF8205200 , 32'h00DE3C4E , 32'hDAEF2C00 , 32'hF74A0250 , 32'hFB00F970 , 32'hFE8EE6CC , 32'hEEF714C0 , 32'hFC4F11AC , 32'h00012ABF , 32'hF5A88280 , 32'hFDD0A894 , 32'h06649838 , 32'h05C38330 , 32'h01CB6D98 , 32'h003CCCA1 , 32'hFECF7124 , 32'hFF513A87 , 32'hF9B945F8 , 32'hF4932780 , 32'hED9B5060 , 32'h00B0E756 , 32'h0490F028 , 32'h01F7D1B0 , 32'hF06592D0 , 32'h0347ED34 , 32'h0005B22C , 32'hFFB09151 , 32'hECDD8EC0 , 32'hFFC21D70 , 32'h0B295880 , 32'hF54895D0 , 32'hFFFF29B7 , 32'hFCB9E774 , 32'hF81523F0 , 32'hE44E3560 , 32'hF7F175C0 , 32'h0003D427 , 32'hF1C9FAF0 , 32'h03E5F830 , 32'h11D88180 , 32'hFC510C74 , 32'hE87121E0} , 
{32'h03AFF9E8 , 32'h04B3A738 , 32'h17DD9D20 , 32'hFFFD28FB , 32'hFFFAE2CA , 32'h06D9BD58 , 32'h118434E0 , 32'hEF1ACAE0 , 32'h00002D6C , 32'h02447D84 , 32'h10E75360 , 32'h048B1F08 , 32'hF7A5D280 , 32'h09A1FDB0 , 32'h0DBF17C0 , 32'hED32BCA0 , 32'hFFC58F93 , 32'hFE3540C0 , 32'h07B47F08 , 32'h000005AC , 32'h029756DC , 32'hE6A2A160 , 32'hFF256E0D , 32'h00019FA3 , 32'hF1E3ED30 , 32'hF1C45850 , 32'hFE6055CC , 32'hFD719D4C , 32'h00E5708B , 32'hED545080 , 32'hF6CD9950 , 32'h101F0A40 , 32'h11ED22A0 , 32'h0C1D11F0 , 32'hFFFE7372 , 32'hF7355570 , 32'hF539ABE0 , 32'hF9631D40 , 32'hF779A720 , 32'hEC07FE80 , 32'h08ECF300 , 32'hFE8EE2D8 , 32'h0ACCCDE0 , 32'hEBD183E0 , 32'h00F3BF28 , 32'hFA8029F0 , 32'hF72958E0 , 32'hF379A810 , 32'hFE3A8548 , 32'h18E6CF40 , 32'h0B4BC650 , 32'h0082EE51 , 32'hF057EC60 , 32'hF48E0530 , 32'h1D0A26C0 , 32'hF8BC44B0 , 32'hFE47A3B4 , 32'h13040620 , 32'hF94465B8 , 32'hED3F7960 , 32'h04F1F8F8 , 32'hF8FBA3B0 , 32'hFFF757C7 , 32'h071D07E8 , 32'h1C332860 , 32'hFBCD2B90 , 32'h0004F024 , 32'hFC0953B8 , 32'hF69823E0 , 32'hF04D40E0 , 32'h0DB5C2C0 , 32'h02009A44 , 32'hF3650040 , 32'hDD974C40 , 32'h0E042760 , 32'h001A8728 , 32'hFF1407FE , 32'hE9207EC0 , 32'hF6F20540 , 32'h178D47C0 , 32'h1558FD20 , 32'hF3710390 , 32'h13ABDA40 , 32'hFFFF893F , 32'hF37E3C20 , 32'hFFD7DEB7 , 32'h19A03280 , 32'hEA6FBFA0 , 32'h1214F060 , 32'hFFFFCA9E , 32'h08C3EF40 , 32'h01798FD8 , 32'h10C65FC0 , 32'h097B9B70 , 32'hFFFF0C5E , 32'hF6F9E4E0 , 32'h04E34910 , 32'h02EEC374 , 32'hF57AE8D0 , 32'hFC9F9CF8} , 
{32'h0E085450 , 32'h0722E2D8 , 32'hF6770D40 , 32'hFFFED350 , 32'hFFFF126B , 32'h0583EEC0 , 32'h043F8F10 , 32'hFCA6601C , 32'h0002D584 , 32'h05BAE578 , 32'hF6B5CC60 , 32'h15A1C5E0 , 32'hFDA67380 , 32'hFAF13AA0 , 32'h1291FA60 , 32'h0BBC9C50 , 32'hF57C8FE0 , 32'h0735E890 , 32'hF772FFE0 , 32'hFFFC91EF , 32'h115F4D80 , 32'h1D6C4820 , 32'h0BE5F750 , 32'h00012E2A , 32'hE1DA98A0 , 32'hEBF62500 , 32'h07CAC580 , 32'h06FA0350 , 32'hE1103B80 , 32'hF23A8AF0 , 32'hEF1EDC00 , 32'hF9A21DA0 , 32'hF2A19840 , 32'hED6D9F20 , 32'hFFFE1184 , 32'hF4FE2210 , 32'hFF656B58 , 32'hF6D30F40 , 32'hF9CA5F60 , 32'h08E6B150 , 32'h1F50F120 , 32'hFDB24E54 , 32'hF1C2F920 , 32'h04E15370 , 32'hFB977E58 , 32'hF184A040 , 32'h0362F61C , 32'hEE6CE060 , 32'h16EE3BE0 , 32'h05D6C1D8 , 32'h0CE42F20 , 32'h09E1E690 , 32'hFEC21AA8 , 32'h09CB70A0 , 32'h132FD920 , 32'h0B6D7A50 , 32'h01F0FD70 , 32'h0D21C800 , 32'h00D2F898 , 32'hF75F0EF0 , 32'h12CA3AE0 , 32'hEDF50160 , 32'hE765F000 , 32'h0809E0E0 , 32'hFE2E91C8 , 32'h0A0B90F0 , 32'hFFFE6F2A , 32'h16FA7020 , 32'hFD2243A4 , 32'hF6C60430 , 32'hEE25E360 , 32'h03531668 , 32'hF4C2E570 , 32'hFB35B9B8 , 32'hFE00E1A8 , 32'hF78D3530 , 32'hEF389120 , 32'h09FD8200 , 32'hF689CA00 , 32'hFB6ADDA8 , 32'hE85B2100 , 32'h10ED9FC0 , 32'hF5064C60 , 32'hFFFE4676 , 32'h016E7650 , 32'h1826AC20 , 32'hF9C0ABC8 , 32'hFA3DA4C0 , 32'hFBA52F78 , 32'hFFFCB288 , 32'h1706CC40 , 32'h01911400 , 32'hFF67C182 , 32'hF2A4E890 , 32'hFFFF9500 , 32'h10BD24C0 , 32'hF83C8978 , 32'hFA087F78 , 32'hF4FAB880 , 32'h0DFF47C0} , 
{32'hF86B55A0 , 32'hFC8ED1B8 , 32'hFBCC3488 , 32'hFFFDCC0A , 32'h00041C8B , 32'h08AD2760 , 32'hF54FFA70 , 32'h00ED23C0 , 32'hFFFE64B7 , 32'hF3FDA8B0 , 32'h10018360 , 32'hFD0F7058 , 32'hF6F0A760 , 32'h1A1AEE40 , 32'h026229BC , 32'h0239658C , 32'hF8D29BB8 , 32'h01305F90 , 32'h02172D70 , 32'h00065028 , 32'h017B5DD4 , 32'hF2787350 , 32'h1E15CC40 , 32'h0001017C , 32'hEE74ABC0 , 32'h1D483920 , 32'hFB199448 , 32'h035E5A10 , 32'h128CABA0 , 32'hF0F174A0 , 32'h0E0B2E50 , 32'h07E4DCD8 , 32'h11822FC0 , 32'h09795480 , 32'hFFFD6074 , 32'h0A247040 , 32'h045A9B30 , 32'hF2F86340 , 32'hF38CF520 , 32'hE5744440 , 32'h2535D7C0 , 32'h00037366 , 32'hF8FB7798 , 32'h005FBE52 , 32'hF4B2B170 , 32'h02D9F150 , 32'h11DA0DA0 , 32'h10826260 , 32'hEA5B6C60 , 32'hF2CE2270 , 32'h1947F4E0 , 32'h045D4D70 , 32'h0E34BCB0 , 32'hE44E9040 , 32'hF1ACDFF0 , 32'hF312A4E0 , 32'h08383100 , 32'h00D668D3 , 32'hF30DFB40 , 32'hFA4FA0F8 , 32'hFDCC385C , 32'h02CAFDD0 , 32'hF3D39120 , 32'h01B27B98 , 32'h0DEACD70 , 32'h0573EC88 , 32'hFFFE814E , 32'hF9ED2F00 , 32'hFA0EB020 , 32'h00470DD0 , 32'hF1C72A00 , 32'h02B83AB8 , 32'hFCAA0498 , 32'h0DC60410 , 32'h105A7420 , 32'hEB82E400 , 32'hF241C5E0 , 32'h051CD050 , 32'h12609740 , 32'hE6B651A0 , 32'hFF59D0CC , 32'hFA8A8200 , 32'hF5927570 , 32'hFFFE02ED , 32'h0E69D2F0 , 32'h14D21C80 , 32'hECF50540 , 32'h00FEC27C , 32'hFD40D4EC , 32'h00006EFB , 32'h111C3340 , 32'hFACD9470 , 32'hFD4DA4DC , 32'hFA9381A8 , 32'hFFFCB838 , 32'hE7FD0320 , 32'hF1467B90 , 32'hFD1C274C , 32'h03EA7994 , 32'hF8CA8CA8} , 
{32'hFD069674 , 32'h0E7A8D80 , 32'h11781C00 , 32'hFFFEAE1E , 32'h00001918 , 32'h000280AF , 32'hFFA7077E , 32'h0AAFA560 , 32'h00028C99 , 32'hF5D4CCF0 , 32'hF81C6BA8 , 32'hF4C2FD00 , 32'h1213AB00 , 32'h10D33BC0 , 32'hFDDE5320 , 32'h05C462F0 , 32'h12860500 , 32'hF3956590 , 32'h035747F8 , 32'hFFFFE2D3 , 32'h13931260 , 32'hF37517E0 , 32'hFF7C39ED , 32'hFFFF9502 , 32'hEE162600 , 32'h071E8710 , 32'h0625DBF0 , 32'hFCE5C370 , 32'hEF3420E0 , 32'hF7B54840 , 32'h010B2838 , 32'hF160D9B0 , 32'h011A8394 , 32'h0B227F00 , 32'hFFFF1A0C , 32'h001B9B2D , 32'h07B09F70 , 32'h14E60EE0 , 32'hF0425970 , 32'h0892D7F0 , 32'hF2B51100 , 32'hFF0B559F , 32'hFE8B32D0 , 32'hF635AC40 , 32'hFF370E94 , 32'h04144188 , 32'h25E8EF00 , 32'hE5944C00 , 32'h06EB63E0 , 32'hFC7A9E40 , 32'h0FE55A20 , 32'hF2094200 , 32'hF363E460 , 32'h055DE040 , 32'h03402D90 , 32'hEFF0B460 , 32'h0C6FFEA0 , 32'h1C01F3A0 , 32'hF5FF6240 , 32'hFF660E52 , 32'hEC440C80 , 32'hEBF83560 , 32'h1614EEA0 , 32'hF8F455E0 , 32'hFA93C978 , 32'h023126D0 , 32'h00021EE2 , 32'hF439EFF0 , 32'hF820F6F0 , 32'hFD457CA4 , 32'h138BF8A0 , 32'hF318DAC0 , 32'h146D76E0 , 32'h0024F874 , 32'h0BED0570 , 32'h02EC2984 , 32'h04958BD0 , 32'h00524951 , 32'h050E2210 , 32'h018F32E8 , 32'h031BBDB4 , 32'hFDA150E8 , 32'hF33F9F20 , 32'h00019F93 , 32'h09CA4C90 , 32'h0E7DB3C0 , 32'hDAFB0B00 , 32'h06188848 , 32'hF2E998A0 , 32'h00018CE1 , 32'hFDF03FCC , 32'h074CCB48 , 32'h0EA8CA30 , 32'h1763A700 , 32'h0002ECF3 , 32'h299EA640 , 32'h01E216EC , 32'h05F10130 , 32'hFFD0D010 , 32'hFCF56BC8} , 
{32'hE545AF20 , 32'hF9EB1A08 , 32'h05F473F8 , 32'h00002FB2 , 32'hFFFC018A , 32'h0E1F5360 , 32'hF8EFCB50 , 32'h0BA98F90 , 32'h000682F2 , 32'hF7D0FC90 , 32'h017E7870 , 32'h03B213B4 , 32'h04549F50 , 32'hF4CA2E90 , 32'h0377A7C4 , 32'hE6E07680 , 32'h06AA5918 , 32'h0107452C , 32'hF7E072A0 , 32'hFFFEA936 , 32'h0C6550F0 , 32'hE71B56A0 , 32'h105AF6A0 , 32'h000027ED , 32'h0D0D2BE0 , 32'h02456628 , 32'hFCF64208 , 32'hEC31D560 , 32'hF3532DC0 , 32'hF9530E38 , 32'h01D91E0C , 32'hFDD4CEB8 , 32'hF94A5910 , 32'hED8DE620 , 32'h00032805 , 32'h01740FEC , 32'h008B57CE , 32'hE7B8A660 , 32'h242C9280 , 32'h05363298 , 32'hEB054F80 , 32'h0098C326 , 32'hF51DB130 , 32'hF64AE260 , 32'hF7B40540 , 32'hDABDF8C0 , 32'hF2604510 , 32'hF8DE1648 , 32'h0AEB4660 , 32'h048EF9D0 , 32'h0F4BDFB0 , 32'hFA40DD98 , 32'h094475B0 , 32'h0A0FE660 , 32'hF02DB1F0 , 32'hF2F00480 , 32'hFE072720 , 32'hF2B17300 , 32'h0785B0A8 , 32'h0B1F4740 , 32'h09F82540 , 32'hFD808F3C , 32'hFC1412AC , 32'hF7CF9800 , 32'h0D7D0050 , 32'h0DA3AC70 , 32'hFFFC320D , 32'hFDC18CE4 , 32'hF4FD2380 , 32'hF09E1DB0 , 32'h0BEAD2E0 , 32'h07D03888 , 32'h0537DD40 , 32'h026B8390 , 32'hF5EE1660 , 32'hF6D6A480 , 32'hF965DDA0 , 32'h023E703C , 32'h09AC0670 , 32'h2241C8C0 , 32'hEB648480 , 32'hEDD67BA0 , 32'hFF069DCB , 32'hFFFD7A16 , 32'h0FCCEDD0 , 32'h16ED1400 , 32'hEFA77D60 , 32'hEFD839C0 , 32'h0EB01060 , 32'hFFFDD242 , 32'hFAE17E28 , 32'h022E7398 , 32'hE9E2E660 , 32'h0C3A89D0 , 32'h00025546 , 32'hFBDA7610 , 32'hFC620DF4 , 32'hEA32B880 , 32'h0FCCE7C0 , 32'hFD4A87CC} , 
{32'h122A07C0 , 32'hFE5A02CC , 32'hFA4FEC68 , 32'h000648E7 , 32'hFFFF58B5 , 32'h14805D20 , 32'h023117D0 , 32'h05D5C4C8 , 32'h0004959D , 32'h09679EA0 , 32'hFE451B54 , 32'hE8BB5D20 , 32'h1022BDC0 , 32'h0EAF0EB0 , 32'hF850C4E8 , 32'hED185700 , 32'hE380A9C0 , 32'h13E969E0 , 32'h123E7740 , 32'h0002145F , 32'hF7125780 , 32'h1B04B580 , 32'hFBA3F3C0 , 32'hFFFB122B , 32'hF21926A0 , 32'hDA3D3DC0 , 32'hEEE8C620 , 32'hED5557E0 , 32'h163FF120 , 32'hFD431420 , 32'h01E4F000 , 32'h0700B5B8 , 32'hF4AB55E0 , 32'h07B626B8 , 32'h00008012 , 32'h03D6D8B8 , 32'h03283158 , 32'h00802561 , 32'h015ECA14 , 32'hF342E4F0 , 32'hFD294610 , 32'h01A9EB40 , 32'hFF461562 , 32'hEF4C6D40 , 32'h0A3F6D70 , 32'hEDCFCF40 , 32'h04B75058 , 32'h09AB66E0 , 32'h1492A800 , 32'hF8F89A10 , 32'h14A56560 , 32'h05F4A3B8 , 32'h13338A00 , 32'hFE2F75DC , 32'h01796534 , 32'h02ECE808 , 32'hEF26B200 , 32'hED4E87E0 , 32'hFCB3B19C , 32'hF4960150 , 32'hF43E2EF0 , 32'h197D9760 , 32'h0A2FC780 , 32'h053ECB00 , 32'hF805C1B8 , 32'h01EFB634 , 32'hFFFEF4CC , 32'hEA9A89C0 , 32'hFBDED678 , 32'h1AB61C80 , 32'h07133E30 , 32'h0CD20CD0 , 32'h02B7FA80 , 32'hF18B0B80 , 32'hF826AD60 , 32'hF361BAD0 , 32'h07295228 , 32'h047C3FC8 , 32'hEE02B980 , 32'hFC2A1140 , 32'hF4E70EE0 , 32'hFDEA7DD8 , 32'h0076E4E9 , 32'h000356BA , 32'h0693FF30 , 32'h0A09EF40 , 32'hEF9E4300 , 32'h089ED470 , 32'h15D8C3A0 , 32'hFFFF792A , 32'h09D05B90 , 32'h03720334 , 32'h13FE5A80 , 32'h05568978 , 32'h00081FDD , 32'h11C989A0 , 32'h091205A0 , 32'h063B6E30 , 32'h0CEC75D0 , 32'hF7A044B0} , 
{32'h011F3364 , 32'hFE837BD0 , 32'h132C6FE0 , 32'hFFF9DE61 , 32'hFFFCA23F , 32'h051D2648 , 32'h156D16E0 , 32'hD85F0040 , 32'hFFFF6E56 , 32'h07165380 , 32'h09F63D90 , 32'h0F0AFC70 , 32'h0103F458 , 32'h0679D708 , 32'hDEBF8B40 , 32'h0FBB9390 , 32'h06CF0C38 , 32'hE021FBE0 , 32'hF58CC770 , 32'h0001F327 , 32'h08852EB0 , 32'hF6DBBA60 , 32'h115B7580 , 32'hFFFDCC4B , 32'h0AA33990 , 32'hEF796920 , 32'hFF3DE4B5 , 32'hF4225230 , 32'h0FD6DB00 , 32'h032B65F0 , 32'hF3A09D20 , 32'h09E63D90 , 32'h03059204 , 32'hFD253388 , 32'hFFFB8CBB , 32'h00964704 , 32'h00B6A608 , 32'hFC2704E0 , 32'hEB81ED20 , 32'h1187BB40 , 32'hFFCE1F86 , 32'hFFFF7CD0 , 32'hF5C18E80 , 32'h04761678 , 32'h19774AE0 , 32'hF319CAE0 , 32'h016B417C , 32'h1C9F03A0 , 32'h019CE704 , 32'hFBC9E5B8 , 32'h0303E78C , 32'hFA1DD3B8 , 32'h0B931150 , 32'hED56A9A0 , 32'h006F2EA2 , 32'h0B9A7F70 , 32'hEDDF8780 , 32'h190CBA60 , 32'h034AD100 , 32'h15FD8100 , 32'hEC2DC060 , 32'hFDC0CBA0 , 32'hF5C56CB0 , 32'hF9499CF0 , 32'hE6F90DE0 , 32'h009B1BC7 , 32'h00000D73 , 32'hFA97BF30 , 32'hFF1D6CA3 , 32'hF9666A00 , 32'h0AB62A30 , 32'h07723E08 , 32'h025B9D10 , 32'h0EBC2210 , 32'h0420E6E8 , 32'h0022C7E6 , 32'hEA8B2FA0 , 32'hFC8462A0 , 32'hF5FACE80 , 32'hF8B42930 , 32'hECAEF600 , 32'h023EC224 , 32'h1723F620 , 32'hFFFEBC1F , 32'hF7D70510 , 32'h1B8F1720 , 32'h0B4AFE20 , 32'h0296B0EC , 32'h0314944C , 32'hFFFFC74E , 32'hF5CE6830 , 32'h06B9B5B8 , 32'hF0BF1000 , 32'h09B40BB0 , 32'h0000D26F , 32'h068EE800 , 32'h03E8C468 , 32'h03923B9C , 32'h0722DDA0 , 32'h09F35340} , 
{32'hFB239728 , 32'hED8C4800 , 32'hF8C99E28 , 32'h00037105 , 32'hFFFF9FF9 , 32'hFC80EDC8 , 32'hE6109260 , 32'hF701A670 , 32'hFFFEAA81 , 32'hFCD496B4 , 32'hF562EEC0 , 32'h075474F0 , 32'hFBD37818 , 32'hEBD396E0 , 32'hF316C670 , 32'h1D78CC00 , 32'h03D449F8 , 32'h13100C40 , 32'hF298B950 , 32'hFFFB1CAD , 32'h09FCCE40 , 32'hF16BCA20 , 32'hF0A1E910 , 32'h0003FFA4 , 32'hF344AF80 , 32'hF371E260 , 32'h0E4CF250 , 32'h13135980 , 32'h1F6E5020 , 32'h001DD4EB , 32'h04D54208 , 32'h14C50840 , 32'hF72CBC10 , 32'hF97A97B8 , 32'h000430D5 , 32'h1FB92960 , 32'hE32FDC20 , 32'h07B2DE80 , 32'h168BC720 , 32'h10A83A60 , 32'hFC7308D4 , 32'hFFAEE2CF , 32'hF9DF00D0 , 32'hF499BA90 , 32'hEC731A40 , 32'h119CB980 , 32'h0136C630 , 32'h0A9CBA30 , 32'h07A84468 , 32'hF56ECBA0 , 32'h1B76EA00 , 32'h0BFF2C80 , 32'hFDB50A1C , 32'hFF07755A , 32'hF2C7A7C0 , 32'h147A5F20 , 32'h08BA6FE0 , 32'h0EADBF30 , 32'h11C4FA00 , 32'hFBF43E08 , 32'h12739400 , 32'hF14532E0 , 32'hFF6965A9 , 32'h133CFFA0 , 32'h071383B8 , 32'hF5127E70 , 32'hFFFFEECE , 32'hED30CF00 , 32'hF982FB88 , 32'hFD7028A8 , 32'hFFF0DB9A , 32'hFD0405FC , 32'h02208F6C , 32'h0919B170 , 32'h127C5860 , 32'h0231B6B0 , 32'hF978FE28 , 32'hEE77D040 , 32'hF039FE10 , 32'h006DB2D4 , 32'hF977C2E0 , 32'hF33BB430 , 32'h0068FA36 , 32'hFFFB54A8 , 32'hFEEB0040 , 32'hF652A2B0 , 32'hF9332FD8 , 32'hFBF28CA8 , 32'h0ADF1FB0 , 32'h00042D76 , 32'h0933E6F0 , 32'h057B8620 , 32'h108DC600 , 32'h12BAF4E0 , 32'h0005A7E2 , 32'h07B258A8 , 32'h0A5B0370 , 32'hF5F88160 , 32'hFC3BD16C , 32'h01F527D4} , 
{32'hEDBA2F80 , 32'hF53A86E0 , 32'hF224DB10 , 32'h000291D5 , 32'hFFFD39F2 , 32'hF71BFD50 , 32'hFCDC0230 , 32'hE4DF2DC0 , 32'h000336EA , 32'h05E6A2D0 , 32'h03D2E2A0 , 32'h00F65271 , 32'hFEB666D4 , 32'hF8CE7770 , 32'h0A12C8F0 , 32'h026501FC , 32'h08E73760 , 32'hF97866F8 , 32'h05894208 , 32'h0003300A , 32'hF8174E38 , 32'h088A56E0 , 32'hF0C265A0 , 32'h0000B954 , 32'h00329C70 , 32'hFDC35AB4 , 32'h03C503B8 , 32'h078E53D8 , 32'hF96B32B8 , 32'hE3CE7600 , 32'h0CAF2050 , 32'h19BE3460 , 32'hF8E462D0 , 32'hE8650EA0 , 32'hFFFF79C6 , 32'h100D15C0 , 32'h09B8FFE0 , 32'hFD1D04C4 , 32'h0C4A4890 , 32'hE1F7C0A0 , 32'hE6C7A060 , 32'hFF98F220 , 32'hFDADB8A0 , 32'hFF0784C9 , 32'h07289438 , 32'h12828840 , 32'hF0C85D30 , 32'hE0B61680 , 32'h020D7274 , 32'hF9C6E2F0 , 32'h04BC4980 , 32'hFAB11FC0 , 32'hF987B7B8 , 32'hE07F9FE0 , 32'h0D21CC10 , 32'hF2504170 , 32'h00196772 , 32'h00FB6BDC , 32'h0EFC31E0 , 32'h1A43CFE0 , 32'h0D490B40 , 32'hFD1903BC , 32'h109806E0 , 32'hED22C5C0 , 32'hFF21EE0B , 32'hF52028B0 , 32'h0002D984 , 32'h074DEB00 , 32'hFF02165C , 32'h04E04310 , 32'hEA2146A0 , 32'h0F297880 , 32'h13126500 , 32'hEED30FE0 , 32'hFEC38158 , 32'hFCF97938 , 32'h04EDD330 , 32'h0A6774E0 , 32'h0299D824 , 32'hF34CCCF0 , 32'h026F8C6C , 32'h06192D90 , 32'h0EBBAA50 , 32'hFFFB01E4 , 32'h09D851E0 , 32'h24B6EB80 , 32'hFF4FD8A5 , 32'h1A0CB040 , 32'hFE51B3A8 , 32'hFFFEDAC3 , 32'h007B0EB5 , 32'h07D024F8 , 32'h038B5F24 , 32'hF75EB6D0 , 32'hFFFFD938 , 32'h01E47290 , 32'h06E78F40 , 32'h15681F60 , 32'hFD437DF4 , 32'hFA3FE0B0} , 
{32'h0356CCE8 , 32'h0744C898 , 32'hE401F9E0 , 32'h00010A34 , 32'h0008CEF3 , 32'hF644E610 , 32'h068C1628 , 32'hF5BE6A50 , 32'h0000C9F5 , 32'hE7E51080 , 32'hFFE725F8 , 32'hF57BEEF0 , 32'hFAA24DE8 , 32'hEB056240 , 32'h0077619E , 32'hF6A62CA0 , 32'h06020988 , 32'hF6847AA0 , 32'hFF773D46 , 32'h00043E96 , 32'h1B148B20 , 32'hFEDA175C , 32'h16E2CF00 , 32'hFFFCFE5B , 32'hF03BF450 , 32'hFB5B5778 , 32'hECCF5280 , 32'hF460A450 , 32'hF8B5F9D0 , 32'hF8CA9DD0 , 32'hFFDB9388 , 32'h030ABD74 , 32'h08D4B780 , 32'h016685EC , 32'hFFFF40DE , 32'h010F31C4 , 32'hFD295858 , 32'h025E0BAC , 32'h143BF820 , 32'h0AB333A0 , 32'h05CF0E10 , 32'hFFBAF549 , 32'hFDDE67A0 , 32'hFDC1DBD4 , 32'h0A096630 , 32'hE9373420 , 32'h0B4CDDC0 , 32'hF7170430 , 32'hF8C94088 , 32'h17BB9AC0 , 32'hF4A663D0 , 32'h069AA548 , 32'h00DD5375 , 32'hF2C935F0 , 32'h054BB9B0 , 32'h02169C6C , 32'hFDB5643C , 32'h1707F240 , 32'h10B1B660 , 32'hEE5A7940 , 32'h13DB5140 , 32'h1642EBC0 , 32'h00424C9C , 32'hFB3738E8 , 32'hF2F0DD70 , 32'hE1C67B40 , 32'hFFFD7D58 , 32'hF3097150 , 32'h07200A50 , 32'hF99C3BF0 , 32'hF951ECA8 , 32'h047DBE20 , 32'hF76B5FE0 , 32'h062454B0 , 32'hFDE2AC14 , 32'h00F3C6EE , 32'hFC9E6160 , 32'h0C1C18A0 , 32'hF66F4DA0 , 32'hF3B19510 , 32'h0939F260 , 32'hEB470260 , 32'h1278E640 , 32'h0001A0F5 , 32'h053B3F58 , 32'hD96D0D80 , 32'hF6461DE0 , 32'h16C63140 , 32'hF078D130 , 32'hFFFFCED9 , 32'h05769BB0 , 32'h020B4294 , 32'hF2A97760 , 32'h0324C338 , 32'h00002ADE , 32'h09BAE500 , 32'hED459640 , 32'h08279FD0 , 32'h1148A4A0 , 32'hDF5AF9C0} , 
{32'h00DCC4BD , 32'hF2FE4330 , 32'h0DDB84F0 , 32'hFFFEEAF4 , 32'hFFFE371D , 32'hE2CFFF20 , 32'h1CBB24C0 , 32'h04E2ACA8 , 32'h000495C2 , 32'h068A77A0 , 32'hF3FDEFE0 , 32'h0399E000 , 32'hF3272B30 , 32'hF3092A70 , 32'hF483F780 , 32'hFEFB8D00 , 32'h01204040 , 32'h03F38A30 , 32'h0549B2E8 , 32'hFFFE3777 , 32'hE3CF6FA0 , 32'hF95602B8 , 32'h0050FA39 , 32'h0001F18C , 32'h010005F4 , 32'h0B55C5E0 , 32'h112A2F20 , 32'hF9323910 , 32'h04BDFFF8 , 32'h08FB6B20 , 32'h18A4D940 , 32'h061AE9B8 , 32'hE35D4300 , 32'hF28F22F0 , 32'h00042F11 , 32'hEDB8FEE0 , 32'h07E31B00 , 32'hF407EF10 , 32'hF6702810 , 32'h06D179B8 , 32'hF99AA9A0 , 32'hFF3DC24A , 32'hEEA839E0 , 32'hFC38F8A4 , 32'h024B3FA8 , 32'hE1C89200 , 32'h044166A0 , 32'hF11EABB0 , 32'h00AC628F , 32'h0A3710B0 , 32'h136DEBC0 , 32'hF7C3DCA0 , 32'h023D8330 , 32'hFEA02850 , 32'h0232C8AC , 32'h043D40E0 , 32'h15138540 , 32'h09FF6FC0 , 32'h001705ED , 32'hF94811F8 , 32'h01D6BC04 , 32'h05546818 , 32'h120E1C80 , 32'h10C05D40 , 32'hE9C96000 , 32'h0CBC7CD0 , 32'hFFFE1C08 , 32'hF5BB73D0 , 32'h089EEBD0 , 32'hFFCAF799 , 32'h07950FE0 , 32'hFCBBD3BC , 32'hFE8B7374 , 32'h04C1F620 , 32'h1E6F2880 , 32'hFBE01720 , 32'h0DDDDA80 , 32'h08A89840 , 32'hF1BBF080 , 32'hFE4CA590 , 32'h11FCE400 , 32'hFB427750 , 32'hE98AECE0 , 32'hFFFE2ACC , 32'hE4B132C0 , 32'h06DC8840 , 32'hFD5B3288 , 32'h0BC907B0 , 32'hFFE47BCC , 32'h0000C144 , 32'h21D1DE80 , 32'h0129DAD4 , 32'hF3772CB0 , 32'hF1A11310 , 32'h00007EE0 , 32'hE68B7200 , 32'h0A81C130 , 32'hFECC9AFC , 32'h063547C0 , 32'hF5744770} , 
{32'h02BE1340 , 32'hF9BEBC58 , 32'h0CB84590 , 32'hFFFDB066 , 32'hFFFD00B4 , 32'hFBC049A0 , 32'h049EF150 , 32'hFFB7F845 , 32'h000189A4 , 32'h1390DFC0 , 32'hFD59EF64 , 32'hFA995668 , 32'hED4A31A0 , 32'hFE93928C , 32'h09AC51B0 , 32'hE1134EA0 , 32'h18607A40 , 32'hFE287BB8 , 32'h0493C608 , 32'h00002559 , 32'h095D60E0 , 32'hF47A2B40 , 32'hEFB19A00 , 32'h000170E1 , 32'hE4B61DE0 , 32'hF7EC03B0 , 32'h08EDDDE0 , 32'h10CE6720 , 32'hF1578560 , 32'hFF453840 , 32'hF00A6D80 , 32'hEE9C2B60 , 32'h015BE898 , 32'h09C4CE20 , 32'h00006AA0 , 32'h0D8D5C50 , 32'hF6080FF0 , 32'hF9FF68C0 , 32'h0C36F1F0 , 32'hFB22CC20 , 32'h0271FC7C , 32'h0171C948 , 32'h0B13BD80 , 32'h0A42A530 , 32'h0C1CFEF0 , 32'hF61CE370 , 32'hF9945D70 , 32'h0EAA21D0 , 32'h0F86D910 , 32'hEC3C4120 , 32'hFB6B2C70 , 32'hFD6A4148 , 32'hEF9ED340 , 32'hFF0B2EF0 , 32'hFE4AAD30 , 32'hF9CFA5C8 , 32'hFA6FED80 , 32'hF70CB910 , 32'hF269AB80 , 32'h097C3A40 , 32'h062B6AD8 , 32'hFA57B920 , 32'hED4FB8E0 , 32'hFA0FDA08 , 32'hFB3E6588 , 32'hFDCF2958 , 32'hFFFE021D , 32'hD827E8C0 , 32'hF6157350 , 32'h0D5D2260 , 32'h0C4FEAB0 , 32'hFC1D5550 , 32'h03108AE4 , 32'h0FA480E0 , 32'h0FA4DE90 , 32'h17B7D240 , 32'hFD1DAE68 , 32'h1EE45140 , 32'h09019420 , 32'hF068B0A0 , 32'hF3100B40 , 32'h0A1BBDE0 , 32'hEEF188E0 , 32'hFFFF05DF , 32'h15D9A500 , 32'hF99CAE20 , 32'h1A71F640 , 32'h07E93A38 , 32'h0B32B090 , 32'hFFFF2E4C , 32'h158DB320 , 32'h07CCFB38 , 32'hEEC501C0 , 32'h0916C2F0 , 32'hFFFA8385 , 32'hF6A0C620 , 32'h095520E0 , 32'h0FCC2F70 , 32'hF1146FE0 , 32'hF1B19C70} , 
{32'h01518EC8 , 32'hFE9A16EC , 32'hFFD124DC , 32'hFFFF8CCB , 32'hFFF7FF9D , 32'hEEC23460 , 32'hE4B72440 , 32'hFED88654 , 32'h00034B7D , 32'hF58FEF10 , 32'hE4B8C360 , 32'hC7E77880 , 32'h0B450600 , 32'h092F4AE0 , 32'h0B157820 , 32'hF00C60C0 , 32'hFE57EDC8 , 32'hFFE9FF7A , 32'hF365C1C0 , 32'h000007B8 , 32'h0D2BB520 , 32'hFC513668 , 32'hFBA7AA00 , 32'hFFFC4F0B , 32'hFD3E9A7C , 32'hEF6DBD20 , 32'hF9D01320 , 32'hF6B07440 , 32'h07AFF1B8 , 32'h1135F480 , 32'hF4D25EA0 , 32'hF90B48A0 , 32'hF5E1CBC0 , 32'h076CCDB8 , 32'hFFFBCC4D , 32'h0CA6F070 , 32'h099EA840 , 32'hE8189680 , 32'hE59D8C60 , 32'h0A823070 , 32'hEDE0F660 , 32'h00CF1F14 , 32'h021B8904 , 32'hFF0D7819 , 32'h06868C18 , 32'h053720A8 , 32'hF723B420 , 32'hFD7156C4 , 32'hFA64C960 , 32'h0BB59C40 , 32'h04281DD8 , 32'h0F9D8C30 , 32'hFB8B87B0 , 32'hEC0CDF00 , 32'h0003213F , 32'hF6F390F0 , 32'h09DDF330 , 32'h0A556BA0 , 32'hF1775E00 , 32'hFAB412F0 , 32'h009B61DE , 32'hED3DA680 , 32'hF68BACA0 , 32'h0F0D1880 , 32'hF5D276E0 , 32'hF90F49D0 , 32'hFFFC1E0C , 32'h15EE3080 , 32'h002D49AA , 32'h03DCA0BC , 32'hE80E8360 , 32'hF6BF3BC0 , 32'hF8F66C40 , 32'h0903DBA0 , 32'hF76EC280 , 32'h0088EA83 , 32'h03600888 , 32'h06E275A8 , 32'hE6E30BE0 , 32'h066173A8 , 32'hF83484A8 , 32'hEB3C4800 , 32'hFF85E09C , 32'hFFFE8163 , 32'hFD2EA95C , 32'h1458B840 , 32'h055F42B0 , 32'hF9097A60 , 32'hF4836220 , 32'h00018A6A , 32'hF568C2B0 , 32'hFD4D1F40 , 32'hF4F92EB0 , 32'h0DF87A00 , 32'hFFFEF58A , 32'hE1AE1E00 , 32'h07B44718 , 32'h05B03B18 , 32'hEE3E87E0 , 32'h00575298} , 
{32'h043D0650 , 32'h16AA4F60 , 32'hF1307990 , 32'h00000A3F , 32'hFFFC5B55 , 32'h10169100 , 32'h22B5BBC0 , 32'h04258B98 , 32'hFFFC862E , 32'hF1A3CB60 , 32'h034B3BFC , 32'h08602210 , 32'hFE4DFA28 , 32'hFCC0107C , 32'hF8851CF8 , 32'hFDDB2738 , 32'hF9FB8530 , 32'h06BA33D8 , 32'hE5D4FD80 , 32'h00089C95 , 32'h17B73AC0 , 32'h0E4755F0 , 32'h071D1950 , 32'h00072E9E , 32'h0D61EFF0 , 32'h09382480 , 32'h0C880CB0 , 32'hF3F53E50 , 32'h16FB9F60 , 32'h0D9B7FA0 , 32'hFB2B01A0 , 32'h0286038C , 32'h0B0DC850 , 32'h0086C2A3 , 32'hFFFF90D8 , 32'h0F1E8530 , 32'h032F74C8 , 32'hF71F2DB0 , 32'h133AEAE0 , 32'hED874EA0 , 32'hE4A53760 , 32'hFDD59D2C , 32'h0DF2C2B0 , 32'h0002C886 , 32'hE3F70740 , 32'h0066866B , 32'hFEBA82C0 , 32'hF67CAF70 , 32'hED19A920 , 32'h0B55D700 , 32'hF6B5B380 , 32'h0838C6E0 , 32'hE503E5E0 , 32'hFE75AF9C , 32'hF47896E0 , 32'h098282F0 , 32'hFCEE3EF8 , 32'h16D57280 , 32'hF73CD770 , 32'h07975C68 , 32'hF826C4B8 , 32'hF98B1AA0 , 32'hF18381E0 , 32'hF1E80950 , 32'hFF8B8DB7 , 32'h1708DF60 , 32'h0001EE6D , 32'hEDB45800 , 32'hF26A62B0 , 32'h1125D700 , 32'h06D72E50 , 32'hF53DEE10 , 32'hEC3DE7E0 , 32'hFD87F42C , 32'hF7FAE830 , 32'h0A1A7DC0 , 32'h0936AA60 , 32'h05F56F40 , 32'hEB2F2A00 , 32'hFFB1BF2F , 32'hF4A1C210 , 32'h04D3D360 , 32'hEF1A4980 , 32'h00010CFF , 32'hFDE11554 , 32'h0FC9D400 , 32'h00D98FBA , 32'hFE9AAFAC , 32'hF4C2D650 , 32'h0001D526 , 32'h0B2B8AE0 , 32'h06751A40 , 32'h191EA820 , 32'hE7F0A5E0 , 32'h0000AFAE , 32'hF7EA98F0 , 32'h012B0030 , 32'h0ECF3600 , 32'h065D3770 , 32'hFDEB4D00} , 
{32'hF9422398 , 32'h027C24D8 , 32'hFCF4AF90 , 32'hFFFA4B00 , 32'h0003AF24 , 32'hFFC92379 , 32'hF3EFCDC0 , 32'hF8FB0340 , 32'hFFFB250F , 32'hF1B0AAC0 , 32'hF7AD3180 , 32'hFC783F10 , 32'h070DD770 , 32'hFB4C3CE8 , 32'hE9155F40 , 32'h0DA78D00 , 32'h13D07160 , 32'h223D6EC0 , 32'h16C07160 , 32'h000307A7 , 32'h09925FA0 , 32'hFBE455A8 , 32'h08ACCE60 , 32'h0000574D , 32'hFA785640 , 32'hF827B5E8 , 32'h159F9800 , 32'hF0F31B50 , 32'h054E2838 , 32'h01958914 , 32'hFC17D354 , 32'hEC9AC260 , 32'h04A00838 , 32'hEB483820 , 32'hFFFE9DF2 , 32'hE9C9FCC0 , 32'h00F31458 , 32'hF7290580 , 32'hF7DF92E0 , 32'h00F16E52 , 32'h07FB7108 , 32'h01B600D4 , 32'hFFFEC469 , 32'hFD648228 , 32'hE7C72400 , 32'hF6DD9EF0 , 32'hEF21F7A0 , 32'hFC1C0118 , 32'h00CA7328 , 32'h15AD5D80 , 32'hEC7824C0 , 32'h00692EA7 , 32'h261B9280 , 32'hE7C5B740 , 32'h02E4C0A8 , 32'h0612B640 , 32'h04133660 , 32'hFB5DF880 , 32'hFF44ED52 , 32'h02F18820 , 32'hEA1FACE0 , 32'hF23C0410 , 32'h01014C90 , 32'hFCB8331C , 32'h087A3A60 , 32'h04F631B0 , 32'h00029831 , 32'hE5B72760 , 32'hF4F3C670 , 32'h0DDCDC80 , 32'hF0873DC0 , 32'hF4B7ADF0 , 32'h25EC7940 , 32'hF7E6D850 , 32'hECA220A0 , 32'h0212B060 , 32'hF3A66480 , 32'hF2607040 , 32'h0A737D60 , 32'h00F99636 , 32'h0BEBFBA0 , 32'h09CBA280 , 32'hFC553B14 , 32'hFFFE0ECF , 32'hFFF2282C , 32'hFE770434 , 32'h1C43BEE0 , 32'hFDB80264 , 32'hF51E2FC0 , 32'h0000C27F , 32'h0EF382B0 , 32'hFB919A68 , 32'hFF8FDFC3 , 32'h0096DAE4 , 32'hFFFFCB13 , 32'h0B390AF0 , 32'hFC00321C , 32'h033733EC , 32'hF3106420 , 32'hF0463540} , 
{32'hFFA164A0 , 32'hFB3C73E0 , 32'h12DE1E60 , 32'h0004316D , 32'hFFFB729B , 32'h05E78480 , 32'hEADED3A0 , 32'hF3DC7AB0 , 32'h00043AAA , 32'h06650A40 , 32'hF979DB60 , 32'hF037FFC0 , 32'hE8453D00 , 32'h0D8F3D80 , 32'hF725D9D0 , 32'hE2434240 , 32'h0319648C , 32'h19F07CE0 , 32'h0B69FA30 , 32'hFFFFC71A , 32'h06779C50 , 32'h1FC58E60 , 32'h1E35AF40 , 32'hFFFEBC02 , 32'h00048163 , 32'h214A5340 , 32'h000247C9 , 32'hF5CEBDE0 , 32'h0C7123D0 , 32'hFD94A1A4 , 32'h013279A4 , 32'hFD7D2218 , 32'h013BA038 , 32'h06FC70F0 , 32'hFFFCC668 , 32'h0B259D50 , 32'h0F3A1CF0 , 32'h063B89D0 , 32'h1004DF60 , 32'h15B8EB20 , 32'h01966558 , 32'h03518F6C , 32'h00B5216A , 32'hFA648ED8 , 32'hF34A5360 , 32'hFBA63F78 , 32'hF8DA1B68 , 32'hFC8EF81C , 32'h0D3B9280 , 32'hDFB3E8C0 , 32'hFA537F48 , 32'h02BA8418 , 32'hF89746F8 , 32'hFD9F9820 , 32'h0D855D40 , 32'h08306EF0 , 32'h097D1D80 , 32'h149ABFC0 , 32'h0BFE3D50 , 32'h021BB860 , 32'h0A9F5ED0 , 32'hF283B200 , 32'hF83993C8 , 32'hFF80F0CB , 32'h02ADEF30 , 32'h08440870 , 32'h0004006C , 32'h0F455C50 , 32'h02D8300C , 32'hF8C146C0 , 32'h16F30DA0 , 32'hF5B1AA70 , 32'h01D67A24 , 32'hE6FF31C0 , 32'hFFD01510 , 32'hF5BD92E0 , 32'h000C7966 , 32'h0BCF50D0 , 32'h072119F8 , 32'hF108C500 , 32'h03287A8C , 32'h0E5E8A50 , 32'h0BD4DFD0 , 32'h0000B2C9 , 32'hE2BD93E0 , 32'hFE2A10CC , 32'h11F11A60 , 32'h13656140 , 32'hFB4B5560 , 32'hFFFF0D24 , 32'hF12B5210 , 32'h0875F1C0 , 32'h035D2824 , 32'h0C5D1470 , 32'hFFFABE4E , 32'hFFDA128C , 32'h099A6D90 , 32'hF0E79DE0 , 32'h10135560 , 32'hFD490668} , 
{32'hF2660D90 , 32'hE4F78FE0 , 32'hFC25EAC4 , 32'h00087D81 , 32'hFFFE30C2 , 32'h05F26038 , 32'h10EA8DA0 , 32'h0AF90860 , 32'hFFFED9D8 , 32'hEECB6840 , 32'h14474300 , 32'h0BD37DF0 , 32'hEE1EE080 , 32'hE893AA20 , 32'hF31AAED0 , 32'hFD9117A8 , 32'hF7965610 , 32'h08D61E20 , 32'h07FE5B40 , 32'h00026F7E , 32'h0BA2E580 , 32'h1018A7C0 , 32'hF4C979B0 , 32'h00021495 , 32'hF1A7BC20 , 32'h018502D4 , 32'hFD9FEE40 , 32'hE7843060 , 32'hFA97BE80 , 32'h01AE4D8C , 32'hEE19E620 , 32'hFDB22B38 , 32'hF7808D50 , 32'h0A4BA4D0 , 32'h000072B4 , 32'hFBA3B118 , 32'hF408BAF0 , 32'h13919DA0 , 32'hEBDC3040 , 32'h065C76F0 , 32'hF2AF3D50 , 32'hFF6752C0 , 32'hE64383E0 , 32'hED2B5260 , 32'h0A7BF360 , 32'h06487C18 , 32'h065D4FA0 , 32'h160E96C0 , 32'hF0108C70 , 32'hF0853030 , 32'hFDF83440 , 32'h05D7EF78 , 32'h00B0D717 , 32'hFBE7C7C0 , 32'hF7039B90 , 32'h058B2240 , 32'hF5019350 , 32'hFDCE193C , 32'hFE5B94C4 , 32'hF136F030 , 32'h07C10828 , 32'h02EB1268 , 32'h0D7302E0 , 32'hF40C4980 , 32'h0D977660 , 32'h128F7520 , 32'h00002584 , 32'h080366D0 , 32'hFCA04754 , 32'hE175D6C0 , 32'hFE421A98 , 32'h028A3354 , 32'hFEF0EE24 , 32'hF5E859A0 , 32'hEECADA60 , 32'h021A5460 , 32'h0E84B050 , 32'h0DE0E560 , 32'h0ECDBF80 , 32'hFD99BF0C , 32'hFF03FC30 , 32'hE6B69860 , 32'hFF7A34F0 , 32'h000211F4 , 32'h0AE9A2E0 , 32'h09E624E0 , 32'h032B4D60 , 32'h07841328 , 32'hE4CF6380 , 32'hFFFA4894 , 32'h083B4000 , 32'h0321BDB4 , 32'h0231BF10 , 32'h0384113C , 32'h000214EE , 32'hF9B5A920 , 32'h1D30E3A0 , 32'h00010549 , 32'hD8DD3E00 , 32'hFB9E3180} , 
{32'h19172560 , 32'hDCEE3140 , 32'h0A5E5910 , 32'hFFFD2283 , 32'hFFFC80FF , 32'hEC81DCA0 , 32'h07328290 , 32'h0A7A8230 , 32'hFFFDCB26 , 32'hFCF44A1C , 32'h1A2DA7C0 , 32'hE6F87060 , 32'hF96F2DE0 , 32'hFF1F6CDD , 32'hE1CEAF80 , 32'h06BB1330 , 32'h027AA8B4 , 32'h1293C0A0 , 32'h138E1FE0 , 32'h0002D824 , 32'hFAA46AA0 , 32'hFE64A08C , 32'hF64B5040 , 32'h00032F75 , 32'h0044033D , 32'h08574010 , 32'hFB362320 , 32'hFFED8365 , 32'h008F5174 , 32'h026F2264 , 32'hEC7F3580 , 32'hF02D6120 , 32'h1B3D09C0 , 32'hFB408870 , 32'h0003A072 , 32'hFCEBDF00 , 32'hF7FEB270 , 32'h0205AD6C , 32'h05D4EE18 , 32'hFC1E0CC8 , 32'h01153BC4 , 32'h0065C8BE , 32'h01D21AD0 , 32'h0B17A570 , 32'h06DD3658 , 32'hFCEAB0D4 , 32'hFD27D2FC , 32'hE948AE20 , 32'hF75E1780 , 32'h00A6A4B7 , 32'h03DAC9E4 , 32'h04454E38 , 32'hF5275050 , 32'hFCFA81D4 , 32'hF1CD5090 , 32'hFDE52BC0 , 32'h043AF0B8 , 32'hFB110248 , 32'h00E7B278 , 32'h0CC400B0 , 32'hF00243B0 , 32'hEFEA8A60 , 32'hF0CB5420 , 32'hF9562A48 , 32'h011A73AC , 32'hE787DB40 , 32'hFFFF396D , 32'hFCC7805C , 32'h0A63C680 , 32'hE47C6D00 , 32'hF05E8340 , 32'h0630EA70 , 32'h016CF8F8 , 32'hF4A21CE0 , 32'h0E3CEAE0 , 32'hE6D90180 , 32'h05CB3100 , 32'h074E4048 , 32'hFA110DB0 , 32'h17278FA0 , 32'hD52791C0 , 32'h010B33F4 , 32'hFFCD0DD3 , 32'hFFFA7142 , 32'hF4C12B00 , 32'hF42C6000 , 32'hF247D770 , 32'hFFC2D69E , 32'h07CD6398 , 32'hFFFAB104 , 32'h037147A8 , 32'h0BF70A80 , 32'h0464CB68 , 32'hED0A9B20 , 32'h0004C7AF , 32'h0619ADA0 , 32'hF4850380 , 32'h113E1D40 , 32'h076EBB20 , 32'h0BBF80C0} , 
{32'h0191381C , 32'h0AF37180 , 32'h08B26880 , 32'hFFFC3E11 , 32'hFFFEBCFF , 32'h0936A0C0 , 32'h1003C2A0 , 32'h11D72780 , 32'h000065B8 , 32'hFC01320C , 32'hEEF567A0 , 32'hFBE28878 , 32'hFF86CE6A , 32'h0CAAC730 , 32'hE6EB5820 , 32'h0802C1B0 , 32'h01BEE614 , 32'h17891B80 , 32'h027F5754 , 32'h000014C0 , 32'h1348B580 , 32'hF4287990 , 32'h0179D9B8 , 32'h00004213 , 32'h05DDC8C8 , 32'hE4E858E0 , 32'h10A3FF80 , 32'h055A5130 , 32'hEB8EF240 , 32'hF8B224E0 , 32'hFF9E608F , 32'hFC22DAA8 , 32'hFC83951C , 32'h163BE5C0 , 32'hFFFE2F17 , 32'hFD0E721C , 32'h0746B540 , 32'h0B0D7600 , 32'h02BBE0BC , 32'h0F1D2260 , 32'hF6456450 , 32'hFF27427D , 32'h12575540 , 32'hF266D330 , 32'hF236AFE0 , 32'h09B459F0 , 32'h08D27E60 , 32'h0F9DE230 , 32'h0587A920 , 32'h09376460 , 32'h03D4153C , 32'h0C2887F0 , 32'hFAB48120 , 32'hF4105310 , 32'h014A3364 , 32'hFE5D37A0 , 32'hF60A5870 , 32'h0012353E , 32'hF203FE70 , 32'h1CD6A840 , 32'h1D4A65C0 , 32'h1C2DCF00 , 32'hF9254E50 , 32'hFA882208 , 32'h09971C00 , 32'hE23FC160 , 32'hFFFF1217 , 32'h16C1EDC0 , 32'h07373F60 , 32'hE90A6060 , 32'hFB7078E0 , 32'h0DBB66D0 , 32'h0FB41840 , 32'h0E9319B0 , 32'h05A608B8 , 32'hFA31C488 , 32'h008C877D , 32'h00DB438D , 32'h0C9CE590 , 32'hF3ACDEE0 , 32'h11D33200 , 32'h0787E220 , 32'hF1753840 , 32'h0001F406 , 32'hF0E68D50 , 32'h0FC1FDB0 , 32'hFD90F6FC , 32'hF7580EC0 , 32'h1185EFE0 , 32'hFFFD8AF3 , 32'hFC53804C , 32'h011E2DA4 , 32'hFF727F46 , 32'hE58B8220 , 32'h00010E0E , 32'hF6964AC0 , 32'h115C00A0 , 32'hFEEECA74 , 32'h103AD760 , 32'hEE42D020} , 
{32'h02189518 , 32'h09B46B90 , 32'hF9AEAD98 , 32'h0002DEB2 , 32'h000505AB , 32'hFEF2864C , 32'h0BEED4F0 , 32'hDF9FA180 , 32'hFFFB8A7A , 32'hFF744921 , 32'h08B94360 , 32'hFE93A59C , 32'hF8C799A0 , 32'h15C1E4A0 , 32'hEF333F80 , 32'hF2D84670 , 32'hFDE7BFD0 , 32'h0E7CEF70 , 32'hF6C068F0 , 32'hFFFC27A2 , 32'hFD26C0C8 , 32'hF28CDCE0 , 32'h04D03C60 , 32'h00031E35 , 32'h17A96820 , 32'hF1C44490 , 32'hF017A280 , 32'h0729AA98 , 32'hE06231A0 , 32'h06332BC8 , 32'h015C2570 , 32'hF1E132E0 , 32'hF0E2A290 , 32'hF3C1C8A0 , 32'hFFFC4605 , 32'hF878C070 , 32'hE4B81880 , 32'hFF96634E , 32'hFD4F3B50 , 32'hFDA81810 , 32'h04547738 , 32'h0128EF58 , 32'h02303B44 , 32'hF756A5F0 , 32'hF816C318 , 32'h09DE8AD0 , 32'hF79FE870 , 32'hFEC58EA0 , 32'hF69F4FE0 , 32'hEF9F4CA0 , 32'hEF8F3020 , 32'h19A3BE60 , 32'hFE65254C , 32'hF7E1BFA0 , 32'h01AF9760 , 32'hFC222F5C , 32'hFEE7F430 , 32'hE23DF480 , 32'h0921D180 , 32'hF171DDC0 , 32'h06A8E478 , 32'hEA7719A0 , 32'hFB2163D0 , 32'h147BEB40 , 32'hF2A3EF80 , 32'h0EBBA570 , 32'hFFF82FEA , 32'hE87312E0 , 32'h07428FC0 , 32'hF748E2A0 , 32'hF75F5E90 , 32'hFB7F2DB8 , 32'hF19DBC50 , 32'h006D107C , 32'h0EC94C10 , 32'h0539DB30 , 32'hEC329A60 , 32'h0EFAD0B0 , 32'h070EFBE0 , 32'h08427620 , 32'h1B271D40 , 32'hEB0B0420 , 32'hF0688250 , 32'hFFFBBC07 , 32'hF91AF178 , 32'h0EB30060 , 32'hECD79120 , 32'h16CD3D20 , 32'hFD6D3CBC , 32'hFFFF6D8B , 32'hE8C356C0 , 32'h07CEFEF0 , 32'h141A63C0 , 32'h00D16CF4 , 32'h00030860 , 32'h0A97C8B0 , 32'hFBD575F0 , 32'h010DE284 , 32'h07DA99D0 , 32'h03A30458} , 
{32'hEE9E1BC0 , 32'hF055D210 , 32'h012C3788 , 32'h000236A2 , 32'hFFFDB792 , 32'h003208A3 , 32'hFB1DB4B0 , 32'hE9255A40 , 32'hFFFD61E7 , 32'hFFA2CB62 , 32'h04DD5150 , 32'hE70A5E60 , 32'hFC865C0C , 32'h07517F70 , 32'hEF262540 , 32'h018B0410 , 32'h06C46CB0 , 32'hFFA14F36 , 32'hF28987B0 , 32'hFFFFB673 , 32'hEB44C120 , 32'hFFCB6EAE , 32'hF7E3C2C0 , 32'hFFFEB1BE , 32'hEB4A36E0 , 32'h008783C6 , 32'h004A0153 , 32'hEBB621C0 , 32'hF6060C40 , 32'hF7AC8D50 , 32'h095ACC40 , 32'hE7C0D840 , 32'hF15F24C0 , 32'h12B8B680 , 32'hFFFF9260 , 32'h01933988 , 32'hFE864888 , 32'hFD4FC3A0 , 32'h14029940 , 32'h06404570 , 32'h117E2780 , 32'hFE66FC88 , 32'h0FB3D690 , 32'h0E6E8040 , 32'h05E453B0 , 32'hFD830758 , 32'h1D58A7A0 , 32'hFD306F7C , 32'hE9729700 , 32'h0C3B92E0 , 32'hFF07326F , 32'hF4181BC0 , 32'hFE441848 , 32'h12E486A0 , 32'h0198A378 , 32'h0A049830 , 32'h03190E08 , 32'hF053F470 , 32'h06B76FB0 , 32'h087101B0 , 32'h0AB6BBB0 , 32'hFEBD4DF4 , 32'hF4D52160 , 32'hFDF88EAC , 32'h261BF480 , 32'h0B3909A0 , 32'hFFFFBA5F , 32'h0556FE08 , 32'h006097AF , 32'h1376A520 , 32'h09EE1960 , 32'h23011240 , 32'h01FA6C8C , 32'h055E5510 , 32'hFF6C0C45 , 32'h131D2FE0 , 32'hF1F55B70 , 32'hEC2D6340 , 32'hE32A9260 , 32'h0643C3D8 , 32'h040C5238 , 32'h0157B598 , 32'h0841B4E0 , 32'h000209C9 , 32'hFCDA294C , 32'h0B527B00 , 32'h01A5EA10 , 32'h0798E478 , 32'hDF7EC7C0 , 32'h00009974 , 32'h08414690 , 32'hFC7832C8 , 32'hFE286DA0 , 32'hF4CBB280 , 32'hFFFEC631 , 32'h041007D8 , 32'h11566EC0 , 32'h06DE56B8 , 32'h0B6773A0 , 32'h09E98990} , 
{32'hF854C0A8 , 32'hF2AA6830 , 32'hF51977F0 , 32'hFFFB1323 , 32'h000068DA , 32'h158CFC40 , 32'hEEDBCF80 , 32'h0E80B480 , 32'h00066A58 , 32'h0B53D5A0 , 32'h0938F120 , 32'hFD5A573C , 32'h0F22F410 , 32'hFD326168 , 32'h00E3E6C6 , 32'h084105C0 , 32'hFB453020 , 32'hEE315B00 , 32'h00CF880A , 32'h000455F5 , 32'hF8F4CAA8 , 32'h20AB4B00 , 32'h0C95AB90 , 32'h00005FF4 , 32'h0157DD98 , 32'hF1826670 , 32'h210158C0 , 32'hF2FF4A30 , 32'h03565FB0 , 32'hFDF4592C , 32'hF9CCD9D8 , 32'h07F764E8 , 32'hF0F27260 , 32'hFF192D45 , 32'h00016057 , 32'hF9DC1358 , 32'hF3956BD0 , 32'hEB6CE580 , 32'h059636C8 , 32'hF37849B0 , 32'h00B54FEF , 32'h013ECFB4 , 32'hFE6ED998 , 32'hF7C152E0 , 32'h08895EE0 , 32'hEC0E08A0 , 32'h015F604C , 32'h0A71D810 , 32'hE75FCBC0 , 32'h15E4E940 , 32'hF12B8DF0 , 32'hF675D180 , 32'hEC4467C0 , 32'hF95CF3B8 , 32'hE7C9FD40 , 32'hEF7D8E40 , 32'hF87A3DA8 , 32'h0018E9AB , 32'hF8774368 , 32'hFB5B0F58 , 32'h07CECD20 , 32'hE5E9EFA0 , 32'hFAE257C0 , 32'h10B790A0 , 32'h0C423900 , 32'hF02D6010 , 32'h0000599D , 32'h00D01FCA , 32'h16192240 , 32'hF4CF13A0 , 32'h1C987A40 , 32'hF91C2AB0 , 32'h14EF08A0 , 32'hFEF5E604 , 32'h19AD6B00 , 32'hFAAF1A90 , 32'h023981AC , 32'h04EBCD50 , 32'hF7C18EB0 , 32'hEE498C80 , 32'h0D3AF7E0 , 32'h063A58B8 , 32'hF46C2AF0 , 32'h000AFCDE , 32'h0142E810 , 32'hFDA8F984 , 32'h04C80E28 , 32'h0E3A1850 , 32'h0BA7EAB0 , 32'hFFFF9CA8 , 32'hE4C2DC40 , 32'h09F8DCA0 , 32'h015A1480 , 32'hFDA6D830 , 32'hFFFE313C , 32'h0851F1A0 , 32'hEC9103C0 , 32'hFE63209C , 32'hED7C5080 , 32'hFF96790D} , 
{32'hF5BF7020 , 32'h0D350FB0 , 32'h017D5360 , 32'h000673DA , 32'hFFFEA6DE , 32'hE7EBEFE0 , 32'hFA979C88 , 32'hFE2400A4 , 32'h000316B5 , 32'hFAD70DD8 , 32'h0AD3BE90 , 32'hF6BE6440 , 32'hFE03D5AC , 32'h0CCBD5E0 , 32'h018CACA8 , 32'h107945E0 , 32'hED803080 , 32'hFF8B2BC9 , 32'hE2FA11E0 , 32'h00026EFF , 32'hFE9FD308 , 32'h05D91470 , 32'hF8296E68 , 32'hFFFAC9BC , 32'h0572EE00 , 32'hE93B0AE0 , 32'h14776740 , 32'hF7C77040 , 32'hE7771500 , 32'h08A55190 , 32'hFE8142B8 , 32'hEDB0B960 , 32'hEE999A00 , 32'hFDBAD4D4 , 32'hFFFFDC03 , 32'h1BA9A660 , 32'h04154250 , 32'hFB1ECF78 , 32'h07AC74E8 , 32'h03B1134C , 32'h0398C708 , 32'hFF43FD4D , 32'h08162460 , 32'hEC597520 , 32'hF3F2C3A0 , 32'hFCD43EEC , 32'hFE1AB264 , 32'hF5855230 , 32'hF7D1F0E0 , 32'hEC5A5340 , 32'hFF46CDF1 , 32'hEA9B61C0 , 32'h00968834 , 32'hEA0E22E0 , 32'h0612D8A8 , 32'h0CAC1FC0 , 32'h0DE4FAC0 , 32'h0646DE30 , 32'hF94CD970 , 32'hF0CB8D10 , 32'hF5BB8C20 , 32'h222DCB00 , 32'h0D4941D0 , 32'hEDB16C00 , 32'hF87F54C0 , 32'hF840F690 , 32'h0006AD52 , 32'hF173F230 , 32'h08CC5F30 , 32'h025B056C , 32'h14BAACA0 , 32'h0C0E4980 , 32'hFCC7C5A8 , 32'hE352EF00 , 32'h05DEA898 , 32'hEB544560 , 32'hEC73C420 , 32'hFD07A8A0 , 32'h178998C0 , 32'hF9F77F20 , 32'hEF3536A0 , 32'hFA0077C8 , 32'hFD13BD9C , 32'hFFFFA3A9 , 32'h0291B174 , 32'hF0F0E320 , 32'h0A969390 , 32'hF1DFFCF0 , 32'hF7CAD840 , 32'h00088081 , 32'h01A05A40 , 32'h0CD4B3C0 , 32'hFA829DB0 , 32'h00FB6601 , 32'h0001F7F3 , 32'hEF2429E0 , 32'hEF5E5420 , 32'hFC891BA4 , 32'hF503E570 , 32'h18500860} , 
{32'h146D71C0 , 32'hF9F6D538 , 32'hED1A1960 , 32'hFFFE9C74 , 32'h0002C21E , 32'hD54262C0 , 32'h04482048 , 32'hFCD3E268 , 32'h0001C7CA , 32'h05375850 , 32'hF8D9A880 , 32'hFDA7C398 , 32'hF45C9A20 , 32'h02A47860 , 32'h0ABA9280 , 32'h0C574800 , 32'h12E09F40 , 32'hFB2C91D0 , 32'hFFC3D210 , 32'hFFFDA558 , 32'hF62D5150 , 32'h08CE8590 , 32'h023D0458 , 32'h00000E4E , 32'h05657B30 , 32'hE5E3DF00 , 32'h127E6780 , 32'hFE460EB4 , 32'hF3E25C30 , 32'hF796B780 , 32'h03D7FF80 , 32'hFC479F50 , 32'h1066AD80 , 32'h082AB990 , 32'h000906C2 , 32'h0CDD8AD0 , 32'h032AF2D0 , 32'hFD70AA28 , 32'h1C9B9E80 , 32'hFE6B9568 , 32'h0BE702B0 , 32'h001C52B3 , 32'hF6955D60 , 32'hF8AD1668 , 32'h0B55EEA0 , 32'h057CB520 , 32'hECB73B80 , 32'h131FC620 , 32'h05709FF0 , 32'hF8399A98 , 32'h0570B608 , 32'hFA30BB88 , 32'h1D756A20 , 32'hFFF51D37 , 32'hF839F358 , 32'hF9F94618 , 32'h0B5D6A70 , 32'h03532094 , 32'hDA768D40 , 32'hFFA7813F , 32'hEEC71FC0 , 32'hEC01A7C0 , 32'hFFB44536 , 32'hF8B93748 , 32'h07CAC498 , 32'h19034A40 , 32'hFFFC4674 , 32'h0EE12360 , 32'h0169EA58 , 32'hF05D4110 , 32'h12633980 , 32'hFAAC19A8 , 32'hEBE60EA0 , 32'h0396145C , 32'hFBC2AD88 , 32'h03305FA4 , 32'h13788960 , 32'hF8FD9418 , 32'hFD489950 , 32'hFE91A374 , 32'h05AECE90 , 32'hF8116D48 , 32'h0F4FEF60 , 32'hFFFD84B8 , 32'h07AB7488 , 32'h0774AFD0 , 32'hFB54BA10 , 32'hFAE40F28 , 32'hF7DC9E30 , 32'hFFFAB21F , 32'hF75DC960 , 32'h0297015C , 32'h119777C0 , 32'hF4DA9200 , 32'h00016F92 , 32'h09147930 , 32'hFF0A5427 , 32'hFA7AAB38 , 32'h1329A0E0 , 32'hD9A7EB40} , 
{32'h03176058 , 32'hF33B79A0 , 32'h0548BC50 , 32'h0001F4B3 , 32'hFFFF17EE , 32'hE9C2F020 , 32'h0A849120 , 32'hFB5806B0 , 32'h000560D7 , 32'hF9E1D620 , 32'h00D0C072 , 32'hFC25BF90 , 32'hFB33BBB8 , 32'h04661278 , 32'h085C5220 , 32'hFD230FD8 , 32'hE2ED2420 , 32'hFFA0154B , 32'hFDB4A134 , 32'hFFFADA3B , 32'h040CF400 , 32'h00FDB8B5 , 32'h0EFF3220 , 32'h0001299B , 32'h01107EB4 , 32'h130C8900 , 32'hE83FB660 , 32'h10C53320 , 32'hF13232F0 , 32'h0BD17F60 , 32'h0023AEAC , 32'h0DDE4F70 , 32'hFCD14160 , 32'h007A7914 , 32'h0001DABB , 32'hFC98C9E0 , 32'h09545C80 , 32'h00AB6414 , 32'h1019DF80 , 32'hF45C1A80 , 32'h0739ED70 , 32'hFFEB737C , 32'h02CD0408 , 32'hEA1183C0 , 32'hF8B8EDA8 , 32'hFDC91288 , 32'h05D68298 , 32'hFBC631A0 , 32'h1203F140 , 32'hFD6870C8 , 32'hEDEC63C0 , 32'h029DF7EC , 32'h11A6A4E0 , 32'h07DADA60 , 32'h00A8D3E6 , 32'hF8A542B0 , 32'hFCECE57C , 32'h01124578 , 32'hEFFA59E0 , 32'h103F1C40 , 32'h05290CF0 , 32'hF26D7960 , 32'h172138E0 , 32'h0B270050 , 32'h10183EA0 , 32'hEDB68800 , 32'h000B8A2A , 32'hE76F8A80 , 32'h02E6D5BC , 32'hF700A860 , 32'h1560B6E0 , 32'hF5E4A8A0 , 32'h16D9CA40 , 32'h1CAA0C00 , 32'hDD13A680 , 32'h0D56BE10 , 32'hF368D0F0 , 32'hFC7E03F8 , 32'hE7CE62A0 , 32'hE9B40D00 , 32'hFA56AC80 , 32'hF7242E60 , 32'h0EE140D0 , 32'hFFFAFBDA , 32'hEC73CC80 , 32'h05B774A8 , 32'hF5AD4EE0 , 32'hF1554C20 , 32'h05C93900 , 32'hFFFD7E9E , 32'h053D8850 , 32'h13AEDCC0 , 32'h02860058 , 32'hEEC5BCC0 , 32'hFFFF945F , 32'hFB251500 , 32'hFEEB3FC4 , 32'h03C8B52C , 32'hE2D5D7C0 , 32'h123131E0} , 
{32'h1801A7A0 , 32'h0D3EAFA0 , 32'hFE4673D0 , 32'h00050012 , 32'hFFFD7DC3 , 32'h0147309C , 32'hFB21E878 , 32'hFE6DF0AC , 32'h0007CA23 , 32'h0363AE8C , 32'hD55CE180 , 32'hFD635038 , 32'h0726DF70 , 32'h04FFD8F8 , 32'h03486564 , 32'hFB8A2FF8 , 32'h035EFDF8 , 32'hF4CEB8B0 , 32'hF80C94F0 , 32'h00043D2A , 32'hFE174868 , 32'hFD6A6224 , 32'h0381D4C0 , 32'h00012507 , 32'hEEAD60C0 , 32'h0200F6B4 , 32'hFB61F080 , 32'hF5447830 , 32'h0DACEE90 , 32'h09F2ED50 , 32'h0AA71BD0 , 32'h171CB960 , 32'hF8024A20 , 32'hFC3DA6D4 , 32'h0003C455 , 32'hEFC38180 , 32'hF6F4B9D0 , 32'hF8C70D68 , 32'hFCF1A770 , 32'hEF6458C0 , 32'h0239E0FC , 32'hFEBAC018 , 32'h105A4D40 , 32'h059B5990 , 32'h0E268590 , 32'hFC308F1C , 32'hEA75D940 , 32'h0C034500 , 32'hFC5827F4 , 32'hFD0F7380 , 32'hFB96F8C0 , 32'h0B171D00 , 32'hFF1F9941 , 32'h0E4D5EE0 , 32'hF23117A0 , 32'h096F25A0 , 32'h06510740 , 32'hFE95B634 , 32'h12DBE6A0 , 32'h0AD07360 , 32'hF3491E40 , 32'hFF40AB8A , 32'h1F3FAE00 , 32'h0744B560 , 32'h14830420 , 32'hEC19FCE0 , 32'hFFF8A1A0 , 32'h052215C8 , 32'hF8245760 , 32'hDCE85880 , 32'h0CA2FAB0 , 32'h0A3E0F80 , 32'hFBE62650 , 32'hEFB1B020 , 32'h030B711C , 32'h0EFA9D40 , 32'hE3EC0BA0 , 32'h05533628 , 32'h22B89040 , 32'h01F672FC , 32'hE7F05860 , 32'hFC3BB910 , 32'hEAA015E0 , 32'h000159B7 , 32'hFC839234 , 32'h0307F9F8 , 32'h04156DA8 , 32'h004C328C , 32'hE04CD840 , 32'h0004DEBF , 32'h0A5C9A40 , 32'h04EBE908 , 32'h0CD95F40 , 32'hFCD83CE8 , 32'h00042160 , 32'hFF04CD80 , 32'h01DF6BB0 , 32'h10F7B420 , 32'h0CA41960 , 32'hFB50A4A0} , 
{32'hF4CCEA30 , 32'h050C8A48 , 32'h039D6334 , 32'hFFFA944D , 32'hFFFDCB93 , 32'hEE2D28E0 , 32'h094876F0 , 32'h0EEBD270 , 32'hFFF96721 , 32'h0FFC4360 , 32'hE0CF1600 , 32'hF13E5CE0 , 32'h0E92D120 , 32'hE395F720 , 32'hE2FAF5E0 , 32'h0A2553D0 , 32'h0467A658 , 32'hF6329B20 , 32'h135C2260 , 32'h00067D2A , 32'h0A347790 , 32'hFFD7E920 , 32'h126935E0 , 32'hFFFF5DA9 , 32'hF7C9B150 , 32'hFE353298 , 32'hFA9623A0 , 32'hF3DB5840 , 32'hEA8EA140 , 32'h05D8E490 , 32'h010208DC , 32'hFC7ABC54 , 32'h0875C6A0 , 32'hF0C540E0 , 32'h000476E1 , 32'hFC025270 , 32'hF3A4F380 , 32'h0420C380 , 32'hF9C4C000 , 32'hE2303080 , 32'hF6252200 , 32'h0022AB39 , 32'hF30D9480 , 32'h01534C6C , 32'hFA170068 , 32'h01F6ECFC , 32'h12C5BBE0 , 32'h0B5A7480 , 32'hF22989F0 , 32'hE85A95A0 , 32'h20473700 , 32'h057B8B88 , 32'hFD0137A4 , 32'h15CE9720 , 32'h10F0E0E0 , 32'hF3229620 , 32'h07C22A18 , 32'hFE9E57F4 , 32'h04DF6520 , 32'h14F9DC40 , 32'h0447A3A8 , 32'h06CCF590 , 32'hF80D1768 , 32'hF9CA6A18 , 32'h0BA85B10 , 32'hFED2D578 , 32'h0005556C , 32'hF17E5E50 , 32'h100781E0 , 32'h06BB9F50 , 32'hFBEBC7B0 , 32'hF1DAADA0 , 32'hE363CA00 , 32'hEE39E620 , 32'hF2DD9450 , 32'h001A0DDB , 32'hED819720 , 32'hF782AA30 , 32'hF2C70610 , 32'hF8F557F8 , 32'h0637EF20 , 32'h095E2BF0 , 32'h07C93DF0 , 32'h00071B07 , 32'h07565638 , 32'hFF0C1BFF , 32'h111452E0 , 32'h098D6420 , 32'h0AD7EC40 , 32'h000160C8 , 32'hEDA060A0 , 32'hFB207998 , 32'h0C561560 , 32'h029E85E8 , 32'hFFF89070 , 32'hEF22DA20 , 32'hEEFF9EE0 , 32'hF519DE80 , 32'hF7A1E6F0 , 32'h016F6DD0} , 
{32'hF588D980 , 32'hE8DFB720 , 32'hF6DEB5F0 , 32'hFFF91AE5 , 32'hFFFC801A , 32'hFFF0B074 , 32'h16E95AE0 , 32'hF7973570 , 32'h000389E5 , 32'hE0EC4B80 , 32'hCFF4FA00 , 32'h04010E80 , 32'h07D26408 , 32'h08BBFAA0 , 32'hF13246D0 , 32'h05881CE8 , 32'hFE6B20A0 , 32'hE5378760 , 32'h0A071120 , 32'hFFFEEBA8 , 32'h0C47E2D0 , 32'h135D12A0 , 32'hEDC974E0 , 32'hFFF998B2 , 32'h0A3E1B60 , 32'h11524D40 , 32'hFA59EE70 , 32'h030546E8 , 32'h0C62C660 , 32'h02B8FDA8 , 32'hF0FBD990 , 32'hF6962540 , 32'hFABBD0E0 , 32'h064F2F70 , 32'h000364CA , 32'h13292DC0 , 32'hF702E670 , 32'hFC2BEE34 , 32'hFA46E0F0 , 32'h008B3E89 , 32'h0F571550 , 32'hFE55A9D4 , 32'h0479E810 , 32'hE72B0620 , 32'hFA7CA2A0 , 32'h01A59410 , 32'h072FD2F8 , 32'h07A855B0 , 32'h0E076230 , 32'h10A01980 , 32'hFA1BF1E0 , 32'hEDF3F160 , 32'h07821970 , 32'hF65F33E0 , 32'hFF1E6225 , 32'hDFCDD000 , 32'h12E18A60 , 32'hF3484ED0 , 32'hFCE8E5E4 , 32'hF75593B0 , 32'h0F235A40 , 32'h009E50EA , 32'h03E79EFC , 32'h054BF8E8 , 32'h0B018800 , 32'h0C9C2F00 , 32'h00107C3D , 32'h00FE8606 , 32'hECBE4180 , 32'h09691920 , 32'hF67EE3B0 , 32'h04E49EB0 , 32'hF456EBD0 , 32'hFC77A2B8 , 32'h10EE39C0 , 32'h059C9F58 , 32'h02C291B4 , 32'h160DB3A0 , 32'h128C9980 , 32'h0E1340F0 , 32'hF85E3A38 , 32'h04C07368 , 32'h0FF879C0 , 32'h00052629 , 32'hF3E376A0 , 32'hFA387930 , 32'h0EA07BB0 , 32'h039DEB2C , 32'h12884720 , 32'h0001B09A , 32'h01129C5C , 32'h05BC4D80 , 32'hFCE3ACCC , 32'hF4AE1DD0 , 32'h000319AB , 32'h106020E0 , 32'hFAA5BC10 , 32'hFE58E348 , 32'h0AA7DCC0 , 32'h10B183C0} , 
{32'hFCBB3ED8 , 32'hF9A92500 , 32'hD1EF5F80 , 32'hFFFCC9A4 , 32'hFFF6A087 , 32'hEFD1E340 , 32'h0647FBD0 , 32'hF67CC530 , 32'h0000492F , 32'h1585B940 , 32'hFB255880 , 32'h09AB1FA0 , 32'hF51A2870 , 32'h1E998360 , 32'h01B86478 , 32'h00BCF996 , 32'hFC654960 , 32'h05AD3590 , 32'h0F30F370 , 32'h00003ECA , 32'h08FB7C50 , 32'hEFC43DE0 , 32'hF13770F0 , 32'hFFF89744 , 32'hF9F18CA0 , 32'hFD7B6610 , 32'hF7941AF0 , 32'hF6185680 , 32'h05D9CB68 , 32'hF67D5780 , 32'h0A44B320 , 32'hF7C31290 , 32'h092653B0 , 32'hFC712FBC , 32'h00015E44 , 32'hEFEC4320 , 32'h09846850 , 32'h06125088 , 32'hFC059248 , 32'hF2FEE240 , 32'hF907BF80 , 32'hFC89A584 , 32'h0F886090 , 32'h0FC3D480 , 32'h04A5AF58 , 32'hFB352DF0 , 32'h031CB714 , 32'hF9B545C8 , 32'hFF5DBFC8 , 32'h00A8A680 , 32'h0D9533C0 , 32'h09C0FCA0 , 32'hF9E83FA0 , 32'h09A96470 , 32'hE1DC6440 , 32'h0D589670 , 32'h08933CA0 , 32'h19F7E6C0 , 32'hEB888BE0 , 32'hFFE31B33 , 32'h18F0F100 , 32'h16F5E620 , 32'hF9A95980 , 32'h06122898 , 32'hFA26EF80 , 32'h08283C70 , 32'hFFFEB56C , 32'h01373538 , 32'h00F3AEE6 , 32'h0366532C , 32'h0E6D3A60 , 32'hFB775C60 , 32'h1A8814E0 , 32'h09B4B1E0 , 32'hF84B4E68 , 32'hF9980B68 , 32'h01C3A7E0 , 32'h096FF7E0 , 32'h07E697C8 , 32'h146E8020 , 32'hF5C73030 , 32'hEC57BA00 , 32'h0059C828 , 32'hFFFDDFD3 , 32'hF2CFB430 , 32'h078D1EF0 , 32'h1D5664C0 , 32'h138FF660 , 32'hFFADCE98 , 32'h000567CB , 32'hF49BCB40 , 32'hF37B0C10 , 32'h09920D10 , 32'h06A2F4E0 , 32'h0003BC8F , 32'h0B6705E0 , 32'hF04ABD00 , 32'hE9410C00 , 32'hF2243340 , 32'h127F01C0} , 
{32'h1BC0B280 , 32'h0EAD8B90 , 32'h015AE070 , 32'hFFFD9208 , 32'h00057D39 , 32'h0620E190 , 32'hF87F3520 , 32'h02B552C4 , 32'hFFFE1C33 , 32'h002E7500 , 32'hF2457F70 , 32'h00EE7D41 , 32'hFF409ABC , 32'hFF4FE334 , 32'hFD91D384 , 32'h18026B80 , 32'h0CDE5E90 , 32'hF8DDA7A0 , 32'hFC2924E4 , 32'hFFFFA4A2 , 32'hF7EAD8D0 , 32'h10320C40 , 32'h01E20B50 , 32'h0004CB4D , 32'hFA84E578 , 32'h10C65CA0 , 32'hEB5B1560 , 32'h1A7BB6A0 , 32'h0B732940 , 32'h0900EFA0 , 32'hF4F60F00 , 32'hE80B1C60 , 32'h0D217650 , 32'hFC3884EC , 32'hFFFAC31B , 32'h05015BB8 , 32'h135CB780 , 32'hF55305B0 , 32'h14033260 , 32'h00271E61 , 32'hF85EB9D0 , 32'h01DCC184 , 32'h09FAF030 , 32'hE00166E0 , 32'h15E5A720 , 32'hF01197A0 , 32'hE8D5ACA0 , 32'h06613590 , 32'hF008E590 , 32'hF7A402F0 , 32'h078FA198 , 32'h044A82A0 , 32'hFC045038 , 32'h001685CC , 32'h0B80E810 , 32'hF0371F90 , 32'hEA8EF560 , 32'hF849C510 , 32'h00EBD2BE , 32'h07E0D3D0 , 32'h11200F60 , 32'h1789CF00 , 32'hF4013C90 , 32'hF55C1980 , 32'hF9156B80 , 32'h0D865690 , 32'hFFFFBE52 , 32'hF7B5DCF0 , 32'h0226BED4 , 32'hFB73EC30 , 32'hFCB074AC , 32'hF886DA18 , 32'h11887BE0 , 32'hFCE503B8 , 32'h1A795000 , 32'hF87E0278 , 32'hF5A0E480 , 32'hE86E1E40 , 32'hFA471880 , 32'h16AFB160 , 32'h0E07A0A0 , 32'hFFB63890 , 32'h023B4508 , 32'h00010382 , 32'hF7F38840 , 32'h08761770 , 32'hEF087DA0 , 32'h08A60EC0 , 32'hE8232040 , 32'hFFFBEF80 , 32'h0AA1C9A0 , 32'hFB2DBB48 , 32'hFE650ADC , 32'h01E70478 , 32'h0006FACD , 32'h02CB9A38 , 32'h0575CC78 , 32'hF41994D0 , 32'hDCCAF000 , 32'hFB143498} , 
{32'h05EA85C8 , 32'h04BCFF18 , 32'h10440480 , 32'hFFF7A5CB , 32'hFFF581F5 , 32'h06349D60 , 32'hF13F0B90 , 32'hF5D6C2F0 , 32'hFFFB9E68 , 32'hEFF966E0 , 32'h00671B22 , 32'h05D41088 , 32'h03560E8C , 32'h1AE5D400 , 32'hFDDAAF88 , 32'hFBA59E08 , 32'h0F186080 , 32'hFB9EBB48 , 32'h0C789210 , 32'hFFFF441E , 32'h077275D8 , 32'h14725380 , 32'hDC002540 , 32'h000273E0 , 32'h06252058 , 32'h0CC39EF0 , 32'h0E826E10 , 32'hF8FB97E8 , 32'h00E457C1 , 32'h0D4A7280 , 32'h090014E0 , 32'h02B521DC , 32'h02640BF4 , 32'hF37DA240 , 32'hFFFD3898 , 32'h078E4A28 , 32'hE230B620 , 32'h0161D834 , 32'h0B8C5D20 , 32'h0472B6B0 , 32'h0881DF00 , 32'hFF486B96 , 32'hF5ED9D70 , 32'h0F606DC0 , 32'h18E01E80 , 32'hFCA3C654 , 32'hFA9642E8 , 32'h01CAC164 , 32'hFB35BA30 , 32'hFF6B22FD , 32'h1636CF00 , 32'h087A51C0 , 32'h06E9D4F0 , 32'h0DCACEC0 , 32'h1018CCE0 , 32'hE9B3FEC0 , 32'hF223AD10 , 32'h21834A00 , 32'hFDB8FE2C , 32'hE7C9D9C0 , 32'h07B286C0 , 32'h04998178 , 32'hFEE62A84 , 32'hEE1F13C0 , 32'hFE06B390 , 32'h0CBE82A0 , 32'hFFF5F4B1 , 32'hFB598610 , 32'h0BED6890 , 32'hF9325258 , 32'hF6F602A0 , 32'h0568B1E8 , 32'h19980960 , 32'h011C9EE0 , 32'hDF5B4040 , 32'h09F613E0 , 32'hF136AD10 , 32'hFB28CFB0 , 32'hF965F388 , 32'hFC9F7E38 , 32'h09FF87A0 , 32'hF24AAB20 , 32'hE6572420 , 32'h000056B7 , 32'h00DC29BD , 32'hF7667C30 , 32'hFB7D60B8 , 32'hFB535FF0 , 32'h0F101F30 , 32'hFFFF9483 , 32'hF8EC0C28 , 32'h0F0D2260 , 32'h00A04AA2 , 32'hE8140BA0 , 32'h00097B65 , 32'hEA30DBC0 , 32'hFAEBFD48 , 32'h0569D6D8 , 32'h0F18C160 , 32'h04F0AC20} , 
{32'h250DE5C0 , 32'hECABDA80 , 32'h01DCFC48 , 32'h0004E08B , 32'h00063627 , 32'hFC35A1F8 , 32'h036A4260 , 32'hFFADAF08 , 32'h0005EFDA , 32'hFC2F1D90 , 32'hFB790550 , 32'h1240D300 , 32'h0D902B10 , 32'h022AC0DC , 32'h14B7C000 , 32'hF84BAD70 , 32'h0960DDA0 , 32'hFEC0A030 , 32'h017EC330 , 32'hFFFD05EA , 32'hFA3FD230 , 32'h076A02F8 , 32'h014336E8 , 32'hFFFF216A , 32'hFE66C3C0 , 32'h0959C5E0 , 32'h0194B0D4 , 32'hDEEDEC00 , 32'hF270ECB0 , 32'hE3BE61C0 , 32'hFF389170 , 32'hF5FCD7A0 , 32'h0809A900 , 32'h05B275B0 , 32'hFFFA30ED , 32'hFF39D8C3 , 32'hF8F26DF0 , 32'h05448CD0 , 32'hF25E5D60 , 32'h16BE4AC0 , 32'hE8E0E040 , 32'hFF16C839 , 32'h1683E800 , 32'h0BC932F0 , 32'hF40CC1B0 , 32'h008865C6 , 32'hEEC43B60 , 32'h0BB5A700 , 32'h0397381C , 32'hF2340010 , 32'hFB1EBD80 , 32'hFDAE84BC , 32'hF3A633F0 , 32'hEC53ABC0 , 32'hED3334A0 , 32'hFAB0DB38 , 32'h24910FC0 , 32'h007791DC , 32'h1F64A1A0 , 32'hEB720E60 , 32'hFB368110 , 32'h162B8160 , 32'h076CCB70 , 32'hFC6CA798 , 32'h0E674570 , 32'h04AFCC90 , 32'hFFF703A8 , 32'hEC0353C0 , 32'h0A76BB40 , 32'hFC44EE44 , 32'hF87E2B88 , 32'hFFAFE8E3 , 32'h004E5A04 , 32'h0F57B1C0 , 32'h028CD13C , 32'h03FA7CD0 , 32'hEEBE4600 , 32'hFB621858 , 32'hE638A900 , 32'hF6D9A320 , 32'h03DB4330 , 32'h113B7140 , 32'h0C7F2D80 , 32'hFFFB0AE6 , 32'h03D46A64 , 32'h10C75200 , 32'hF3A72FF0 , 32'hF10A5050 , 32'h0D65FA30 , 32'hFFF5975D , 32'hF72EAC10 , 32'hF580A7C0 , 32'h01E23E88 , 32'hF64E3D20 , 32'h0008AD99 , 32'hFD0C1DCC , 32'hFDC8F1C0 , 32'hF7DE2BB0 , 32'hF3577EC0 , 32'hFC398D54} , 
{32'hF12386F0 , 32'hFE9B5E54 , 32'hDC7E2D40 , 32'h00018A9F , 32'h00013AFB , 32'h022D1E5C , 32'hF06515C0 , 32'h04F0F968 , 32'hFFF99670 , 32'h033D8994 , 32'hFA3A5E88 , 32'hFEFC3174 , 32'hF501FFB0 , 32'hEA10FDE0 , 32'hF826B200 , 32'h0323DD0C , 32'hF63074D0 , 32'h03A71994 , 32'hF1E5BE20 , 32'hFFFEEF95 , 32'hFDAA7FE0 , 32'h0DFB61A0 , 32'h022F32F0 , 32'h0006E885 , 32'hF5CDAFC0 , 32'h09465250 , 32'hF199F880 , 32'h0B403EE0 , 32'hED6E5880 , 32'h140EE0E0 , 32'hF2311E60 , 32'h06355150 , 32'h0B07C2A0 , 32'h04310808 , 32'hFFFC75EA , 32'hFA15D190 , 32'hFC9A87E8 , 32'h11699980 , 32'hE9900B00 , 32'hF6EA83D0 , 32'hF03EFA30 , 32'hFF3F10F2 , 32'h156D14C0 , 32'hFFD74001 , 32'hFD6B5DE4 , 32'hEE758520 , 32'hF1C218D0 , 32'hFCF169F0 , 32'h0ABE39A0 , 32'hEAD39700 , 32'h009F4C11 , 32'hE3969FA0 , 32'hFA34D3C0 , 32'h023D9300 , 32'h08FBA720 , 32'h0755D738 , 32'hF5CE0130 , 32'h0BC46E50 , 32'hF32E6330 , 32'hEEA9DEE0 , 32'hEAFD26A0 , 32'hF9C43908 , 32'h05369688 , 32'hFD248F20 , 32'h15779A80 , 32'h0B1F56D0 , 32'hFFFBFF49 , 32'h03DC00A4 , 32'hF99173A0 , 32'hF72C8DA0 , 32'hF7E5DB90 , 32'h045B8AE0 , 32'h0C4192B0 , 32'h1BDEDDC0 , 32'h10EDEC20 , 32'hE321B300 , 32'hEB971FC0 , 32'hF83E0980 , 32'hF2F3AE60 , 32'h09C55C10 , 32'h14F884C0 , 32'hF74D6FE0 , 32'hF9CA6408 , 32'h00017907 , 32'h04439198 , 32'h062EE478 , 32'h10DE35E0 , 32'h02271660 , 32'h105AAF20 , 32'hFFFBF88A , 32'h00746B46 , 32'h07F106F0 , 32'hF837C3C0 , 32'h01CDD388 , 32'h00087326 , 32'hFE3C174C , 32'h0867A7A0 , 32'h185A5160 , 32'h238EBF80 , 32'hFF5861C5} , 
{32'hFE21F16C , 32'hFD9F764C , 32'hF346BC40 , 32'hFFFC9CF8 , 32'hFFFB04C2 , 32'hEEA9B660 , 32'hFBE26008 , 32'h151CDD80 , 32'hFFFD17B1 , 32'hFD2068C0 , 32'h09099E00 , 32'h02D3280C , 32'h005C7814 , 32'h133FEFC0 , 32'h085A1F10 , 32'h052562A8 , 32'hFD027BD4 , 32'h108DBCC0 , 32'hF2636C50 , 32'h00026C13 , 32'hFEF41B94 , 32'h01B160AC , 32'hF68484E0 , 32'hFFFACF10 , 32'h1E129280 , 32'hFF983A84 , 32'hE071BD80 , 32'hF620E5C0 , 32'hF8A09020 , 32'hFD6FBF18 , 32'h0707A808 , 32'hF26278C0 , 32'hF2325FA0 , 32'h0365CAD8 , 32'h0005F7B1 , 32'hFA81EA50 , 32'hFE72E450 , 32'hFD58B78C , 32'hEDC4F220 , 32'hE75FBB20 , 32'hFD7A5994 , 32'h052DDC10 , 32'hF55D6C90 , 32'hEEAEE2A0 , 32'hFAB835E8 , 32'h08F26830 , 32'h01DB8404 , 32'h08684A70 , 32'hF0000580 , 32'h00EF5E09 , 32'h0F1D50E0 , 32'hEB7A5080 , 32'h0676F050 , 32'h01DCB214 , 32'h0F42C500 , 32'h0D7B7EB0 , 32'hF457C760 , 32'h0C3FAD60 , 32'h1589C4C0 , 32'hF1DD8E80 , 32'h0A3294A0 , 32'hF8FCF388 , 32'hEE08D8E0 , 32'hFEBF2B88 , 32'h03708DD4 , 32'hFAC40008 , 32'h00017D07 , 32'h0102FC98 , 32'hEF63FC60 , 32'hF315AF80 , 32'h03A70F60 , 32'hF059E0B0 , 32'h10FB9FE0 , 32'hF854AB68 , 32'h0FE4DBE0 , 32'h2F913980 , 32'h005E8B13 , 32'hF1AC9070 , 32'hFB43DA20 , 32'hF9340AA0 , 32'hDD78E280 , 32'h16310A60 , 32'h00ABB7A6 , 32'hFFF934D7 , 32'hF7F75780 , 32'h0176B478 , 32'h02B49490 , 32'h08F8B590 , 32'h0BEEB4D0 , 32'h00071231 , 32'hFDE76840 , 32'h051B6308 , 32'hEBE30A00 , 32'h02131D44 , 32'h0003C7A7 , 32'h027988B8 , 32'hFE1563E8 , 32'h0109A2A4 , 32'h09FBAEA0 , 32'hE0198580} , 
{32'hF83F2590 , 32'hEF46DA80 , 32'hFD138AF4 , 32'h000CA1A7 , 32'hFFFD28AF , 32'hF46A6E60 , 32'h0094A293 , 32'hF9B36538 , 32'hFFFEEF55 , 32'hF0929590 , 32'hFE032D50 , 32'h08BD6230 , 32'hF7BD3460 , 32'hF08B3C90 , 32'h0B05F8B0 , 32'hF1848420 , 32'h0E7FE020 , 32'hFC0A5C58 , 32'h0E684A10 , 32'hFFFD1E46 , 32'h1264C7E0 , 32'h0CDA5C20 , 32'h13C96300 , 32'h00020603 , 32'h01DCE8E4 , 32'h015AC27C , 32'h09CA9220 , 32'h23754900 , 32'h05F975F0 , 32'h04416B80 , 32'hFA71C710 , 32'h014B54D4 , 32'h06A563B0 , 32'hF248F190 , 32'hFFFCB6E3 , 32'hF05D8D70 , 32'h11FB20A0 , 32'hEFF420E0 , 32'hF38E5100 , 32'h01B9D4E4 , 32'h0B043490 , 32'hFDD5D318 , 32'h1A935EE0 , 32'hF8437080 , 32'hFDFE864C , 32'hFDF8D318 , 32'h08DA7FA0 , 32'h001F94CD , 32'hF9886900 , 32'hFF8A46FC , 32'h0C2D8630 , 32'h0A45A5E0 , 32'h0F679330 , 32'hFC35026C , 32'hF12A1B20 , 32'h19B83840 , 32'h07EBE180 , 32'hF784ACF0 , 32'hF37D6B90 , 32'hF9BFEDA0 , 32'h00746237 , 32'h1279B980 , 32'h010C33EC , 32'hEB34F880 , 32'h037979B4 , 32'h048247C8 , 32'h00026CB7 , 32'hFD41593C , 32'h17E844A0 , 32'hFF0BD52D , 32'hFF5F0F2E , 32'h0C854510 , 32'hFF1D31BD , 32'hE14AF3A0 , 32'h08D473C0 , 32'h24949C00 , 32'h092695F0 , 32'hF415B960 , 32'hF14327C0 , 32'hF8D64D00 , 32'hFB1F7B88 , 32'hF50AB190 , 32'hE615A700 , 32'hFFFB0BBF , 32'h00DB7AC6 , 32'h05DE29E8 , 32'hF2A7FC40 , 32'hF97C3F40 , 32'h0D89C5D0 , 32'h0000FD0B , 32'hE09A5220 , 32'hFECDF080 , 32'hF7E38810 , 32'h11115260 , 32'hFFF746FA , 32'h07AA8908 , 32'h10487FE0 , 32'h140B6F80 , 32'h09332F50 , 32'h133E4120} , 
{32'hF48D3180 , 32'hFE3932C0 , 32'h1E225CE0 , 32'hFFFB1CFF , 32'h0004A793 , 32'h046E3600 , 32'hFDEFA3C4 , 32'h006B9DC3 , 32'h0002D4AF , 32'h0001CA70 , 32'hF8615DA0 , 32'h0B1CC7E0 , 32'hF6BAD0E0 , 32'hEFF6E400 , 32'h14189E80 , 32'h0F3BAC10 , 32'hFE6176B0 , 32'hFE2C2BE8 , 32'h041F4D18 , 32'hFFF88236 , 32'h03889538 , 32'h115C9D40 , 32'hFC0448EC , 32'h00064116 , 32'h01A719F4 , 32'hF89023F8 , 32'h02FE5B4C , 32'hF8327D40 , 32'hEE6CF760 , 32'h08905350 , 32'hFEA2352C , 32'h001DD6E8 , 32'h015C3320 , 32'hF7B1C6E0 , 32'hFFFC1E13 , 32'h0F2FD430 , 32'h1B979FC0 , 32'h0BC5B9E0 , 32'hEC25D9E0 , 32'hFED36864 , 32'h03F6EDA0 , 32'hFEE52748 , 32'h177B3880 , 32'h03EFA5BC , 32'h08628DA0 , 32'hF7E3C560 , 32'h0C2503A0 , 32'hEE6E8AA0 , 32'hF34F5110 , 32'hF2495CE0 , 32'hFBD95648 , 32'h01292A8C , 32'h1B210EC0 , 32'hED462FC0 , 32'hEB6D1660 , 32'hF3FBE7B0 , 32'hF3262170 , 32'hFE864978 , 32'h0FE15830 , 32'h03864BE8 , 32'h051C9218 , 32'hFD3DF418 , 32'hE5142F60 , 32'h1B4A5520 , 32'hF750B110 , 32'hF7020830 , 32'hFFFC47AF , 32'hFCFB5E24 , 32'hF4218A80 , 32'hF56AB8E0 , 32'h12626B20 , 32'hF7296330 , 32'h0EDC14B0 , 32'h007A6CCE , 32'hFF113683 , 32'h0FB3F270 , 32'hFF99E5E1 , 32'h07862F68 , 32'hFBBE1150 , 32'h128E19E0 , 32'hFD30E770 , 32'hF324F220 , 32'h0C939170 , 32'h0008BE84 , 32'h12456C00 , 32'hF48CF6A0 , 32'hFF57CC20 , 32'h08861BF0 , 32'h0120AB74 , 32'h00059BAB , 32'h0B83A450 , 32'hE8AB78E0 , 32'h2B81FC00 , 32'hF5FD1910 , 32'h00042313 , 32'hE7179640 , 32'h0486A5D8 , 32'hFB052D78 , 32'h18E9FEE0 , 32'h03A40544} , 
{32'h002ABBFE , 32'hF0BBC8D0 , 32'hFB8F3EB0 , 32'h00063B5D , 32'hFFFA87D2 , 32'hEEC29240 , 32'hEBBFFA80 , 32'hFC234960 , 32'h000B986C , 32'hFA7B63F8 , 32'h01EA5E84 , 32'hFF795BCB , 32'h025A6D24 , 32'hEA8DC820 , 32'h0E154F10 , 32'hF3F4AD10 , 32'hF700C1F0 , 32'hF08C6E20 , 32'h0A521B40 , 32'h00039E68 , 32'hFDBE4A00 , 32'h0518D918 , 32'hFEB135F8 , 32'hFFFDCDDB , 32'h079DAEF8 , 32'hF5CA2790 , 32'h1E26C900 , 32'h06EB9FD8 , 32'h05B35920 , 32'hF27AF580 , 32'h0481BE40 , 32'hF63A5300 , 32'h134AEE20 , 32'h029B4B20 , 32'h0000BEF0 , 32'hD8988980 , 32'hFB9D5BA8 , 32'hFD648AE4 , 32'h0261B484 , 32'hFE4CF344 , 32'hF993DC40 , 32'h00093038 , 32'hFECA22E8 , 32'hE3F38EA0 , 32'hFE4E0FB0 , 32'h116927A0 , 32'h187FC040 , 32'h165E1380 , 32'h17BC1860 , 32'hFA0EDFE0 , 32'h05407428 , 32'hFDCCFD88 , 32'hE2EDD500 , 32'hED7C6520 , 32'h119977A0 , 32'h0021EE45 , 32'hEDEE3840 , 32'hFECFB750 , 32'h0FAE5650 , 32'h017D9D78 , 32'hFEE0FF9C , 32'h0639B2A8 , 32'hF09E5AF0 , 32'h1007BEE0 , 32'hFB1D7768 , 32'h0C927A80 , 32'hFFF8070B , 32'hF5481560 , 32'hED80EC00 , 32'h0B8DEC90 , 32'h0B9CDE70 , 32'h089F2090 , 32'h04F7E280 , 32'h0D258C60 , 32'hEDF84920 , 32'hF9673748 , 32'hFBD2E900 , 32'hFE036D78 , 32'h0D454110 , 32'h12AC2A60 , 32'hF64D00E0 , 32'h01EB70AC , 32'hF7807580 , 32'hFFFD8E94 , 32'hE574DFC0 , 32'h014DB320 , 32'hF22A3E80 , 32'h00202B8E , 32'hE55D5B20 , 32'h000EFD92 , 32'hF912CB40 , 32'h016560BC , 32'h04DD24A8 , 32'hFC5CA1B0 , 32'h00050FC4 , 32'hECB2C700 , 32'hE9E98B00 , 32'h0EDFEC80 , 32'h0D39F5F0 , 32'hFED167D4} , 
{32'h01DBE170 , 32'h0C9B7050 , 32'h0C33DF80 , 32'h000414C1 , 32'hFFFE3BEA , 32'hFB56D0A8 , 32'hFED9E7F0 , 32'h0107F110 , 32'hFFF900CE , 32'hFAD8C6B8 , 32'hF38E6070 , 32'h1023A4C0 , 32'hFDF18390 , 32'hF12D2BA0 , 32'hF6BDF5A0 , 32'hECF02A60 , 32'hFBCF7930 , 32'h1338EFE0 , 32'h0262C620 , 32'h00083BA4 , 32'h0EE24910 , 32'hF8510210 , 32'h03CE40A8 , 32'hFFFE3A71 , 32'hFC944668 , 32'hEFA1BD80 , 32'h0E373690 , 32'h19BEDE60 , 32'h0AF2F2E0 , 32'hFC1FDF8C , 32'hF4CA6F70 , 32'hF63303E0 , 32'hFA5C3DB0 , 32'h0B271310 , 32'h00031D02 , 32'h03F13B54 , 32'hDBF7E1C0 , 32'h036E5950 , 32'h041B3660 , 32'hD613A500 , 32'hFE8C05D0 , 32'h01B41E44 , 32'h04BAAE10 , 32'h0B0C8D20 , 32'hFDCCA7EC , 32'h0A59F6D0 , 32'h03D10730 , 32'hF84CD330 , 32'hFAC00488 , 32'hFF07B6BE , 32'hF51CEEE0 , 32'hFE695E20 , 32'h055886C0 , 32'h06096D68 , 32'hEF0961C0 , 32'hF1033040 , 32'h099D2050 , 32'h01FC5754 , 32'h04939950 , 32'hF0BD9E50 , 32'hE5C75840 , 32'h14DA7B60 , 32'hFAD5B488 , 32'h0A58F480 , 32'hF6B6EB00 , 32'h0CEB5330 , 32'hFFF7952F , 32'h23E3DDC0 , 32'h127568A0 , 32'h053A3608 , 32'h130BCCC0 , 32'hF4A0B160 , 32'h17C46120 , 32'hF9E9C808 , 32'h00BD3D89 , 32'h012ABF94 , 32'hF0061FE0 , 32'h089A6BF0 , 32'hF5434720 , 32'h0425C730 , 32'hFE26BD50 , 32'h016C541C , 32'h25631780 , 32'h00072390 , 32'hF8608638 , 32'h07059A78 , 32'hEA5B6700 , 32'h0CCFC490 , 32'hF7594760 , 32'hFFFF97B3 , 32'h0D180770 , 32'h06A1C168 , 32'hE3ECA1E0 , 32'hFE1B6FD8 , 32'hFFFD0E10 , 32'hF95C35F8 , 32'h07484DD0 , 32'hFB37D7E8 , 32'h01431114 , 32'h027953F4} , 
{32'h0B5DDF80 , 32'h0DD39B30 , 32'h0B2FCCF0 , 32'hFFF9C39C , 32'hFFF162BF , 32'hFB08B130 , 32'h0F01AD20 , 32'hF86E6540 , 32'h000A17B0 , 32'hFFC6A4CE , 32'hDCDC4440 , 32'h147079C0 , 32'hF9B805A8 , 32'h04E01E20 , 32'hF84D5FB0 , 32'hF224F550 , 32'hF1D530A0 , 32'hF97D3E78 , 32'h02DCA940 , 32'h00063BD2 , 32'h0E23B230 , 32'hFF947B48 , 32'hFFDD82E9 , 32'hFFFF5FD1 , 32'hFF1C813E , 32'hF5F06C90 , 32'hFAE76D00 , 32'hFF5F375F , 32'hF410CAC0 , 32'h0E3DED90 , 32'h01218F94 , 32'h06EA3580 , 32'h0AB76260 , 32'h0A49D960 , 32'h0005BE06 , 32'h027A93D0 , 32'h06A035B0 , 32'hFDB03128 , 32'h04E2A5C8 , 32'hF5B674B0 , 32'hF83819F0 , 32'h036A060C , 32'hE3F07AA0 , 32'h0CA949F0 , 32'h11886C60 , 32'h010BFBF4 , 32'h02DD6114 , 32'h093A2F80 , 32'hF3F2FD80 , 32'hEF971DC0 , 32'hEABA5180 , 32'hFAFBE990 , 32'hF7F72D50 , 32'hF6866720 , 32'h04CBF240 , 32'h1BFC60C0 , 32'h0E3B90C0 , 32'hFB37BEA0 , 32'hFF396515 , 32'hF190EE50 , 32'h114E5AC0 , 32'hE57F95A0 , 32'hF9FCE580 , 32'h057F91D0 , 32'h17119460 , 32'hF9378168 , 32'hFFF82E8F , 32'hEB6BCFA0 , 32'h058F1948 , 32'h10539E80 , 32'hF27F5370 , 32'h11B96CA0 , 32'h2714C340 , 32'hF5B3B070 , 32'h084EE580 , 32'hEA298D60 , 32'h2987B440 , 32'hE8E8AC60 , 32'h013AB090 , 32'h01497530 , 32'hF8FB31A0 , 32'h02D8FD48 , 32'h0095B131 , 32'h00011E2E , 32'h0AA93C60 , 32'h00CE6174 , 32'hF1C505E0 , 32'hF79B4A40 , 32'hF6A40C00 , 32'hFFF932FC , 32'hFA202820 , 32'hFAB68078 , 32'hF586A2A0 , 32'h032AC16C , 32'hFFFC0A7B , 32'hF4596650 , 32'hF6F74EB0 , 32'hF4A58580 , 32'h0CF3C490 , 32'h0684F100} , 
{32'h01DBADB4 , 32'hEB1029C0 , 32'hFD2DBA90 , 32'hFFFFE2D6 , 32'h0000F8E4 , 32'h18D53AA0 , 32'hF100E150 , 32'hFCCD2D4C , 32'h0000A973 , 32'h0B06AE70 , 32'hF866C2A8 , 32'hF86B4098 , 32'h0A0ED270 , 32'hFF12E120 , 32'h02AC54C4 , 32'h17391920 , 32'h069264D0 , 32'h02A06CC0 , 32'hF69294D0 , 32'hFFF28A72 , 32'hFC0750A8 , 32'hF36C0090 , 32'h07593510 , 32'h00024612 , 32'hFBBB2500 , 32'h10C6B800 , 32'hEF8B2160 , 32'h1495D800 , 32'hE6863960 , 32'hEFED3240 , 32'h082F4CE0 , 32'hFD6FC764 , 32'hF8048CB0 , 32'h01262D98 , 32'hFFF18B63 , 32'hFB52C6A0 , 32'hE1C7E320 , 32'h036951E0 , 32'hFD1203D4 , 32'h0B4FBDA0 , 32'hF4FBA8A0 , 32'h0219210C , 32'h01849074 , 32'h0435AAB0 , 32'hFFD0DE5C , 32'hF21120A0 , 32'hF31D6D50 , 32'h0DE03260 , 32'hFA637C90 , 32'hFC546528 , 32'hF4B91480 , 32'h00F7C531 , 32'h05436B48 , 32'hEBB09C60 , 32'h087F85E0 , 32'hFA1A0038 , 32'hFBC8B5A0 , 32'h1C4DF500 , 32'hEF1A9220 , 32'h082D9C30 , 32'hF26DE7E0 , 32'h198EB540 , 32'hF531D1D0 , 32'h2231FE00 , 32'h0B474CB0 , 32'hFB241C20 , 32'h0004A414 , 32'hF46A2080 , 32'h02F2B090 , 32'h0B40DA30 , 32'h0938DE00 , 32'hEF661260 , 32'hF09F3210 , 32'hE1104B20 , 32'hEDE73C80 , 32'h06DC8DB8 , 32'h2B9F2A40 , 32'hFBFA0270 , 32'h03D06400 , 32'h00CAC707 , 32'hF7FCEA00 , 32'hF7BEB510 , 32'hF8CF37A8 , 32'hFFF5DAFC , 32'h029229A8 , 32'h0B373560 , 32'hFD56A12C , 32'h072A83A8 , 32'hF7B8AEA0 , 32'hFFFE4E32 , 32'h06D1F970 , 32'h06A23DB8 , 32'hF0295E70 , 32'hEB24C020 , 32'hFFF34552 , 32'h071C5998 , 32'h01F3498C , 32'h00BE9951 , 32'h0E0AB8B0 , 32'h0F6D9F50} , 
{32'hFE944CB4 , 32'h19319F20 , 32'hFC982290 , 32'h00024065 , 32'hFFFE8026 , 32'hF572EB20 , 32'h01A19768 , 32'h086EA050 , 32'hFFFEC010 , 32'h02CFC34C , 32'h0C809A30 , 32'h03E80DF4 , 32'hFBFD8E50 , 32'hE1BB24C0 , 32'h09639DC0 , 32'hF5B587B0 , 32'hFAC61F10 , 32'hFE0593E0 , 32'h022BCC98 , 32'h0005C8FC , 32'h02E1F67C , 32'hFC0938E0 , 32'h05277680 , 32'h0007346B , 32'hF946AAB8 , 32'h083D5410 , 32'hF5705420 , 32'hE8ACE680 , 32'h08201030 , 32'hED9B01E0 , 32'hFCB8F338 , 32'hFDFB3E10 , 32'hFF07D3E8 , 32'hFBFB17E8 , 32'hFFF90B5C , 32'h1897CC00 , 32'hEDEE15C0 , 32'hFAA2B520 , 32'hE7A4BE60 , 32'h0772DC18 , 32'h037CC754 , 32'hFFF675EE , 32'hFE191488 , 32'hF63068D0 , 32'hF7A01100 , 32'h01748F0C , 32'hEB3834A0 , 32'h00248CEF , 32'hF284D180 , 32'hF2E5AE50 , 32'h07922408 , 32'h0405F360 , 32'hFEFE0898 , 32'h0D641450 , 32'hF9246C40 , 32'hE1997060 , 32'h0F038450 , 32'hF3C84CF0 , 32'hE4BFCE40 , 32'h0B6385E0 , 32'h076D9E78 , 32'h0571AC90 , 32'hF0F8A3C0 , 32'h1518AC80 , 32'hE39BDA80 , 32'hFE706C2C , 32'h000055C1 , 32'hFAF808F0 , 32'hFA88F8F0 , 32'hF57F92E0 , 32'hFA71EB88 , 32'h2B99E000 , 32'h17A24EA0 , 32'h0159B7E8 , 32'hF8B8CE48 , 32'h0B4A3E10 , 32'h0D24ABC0 , 32'hEB974860 , 32'hFCC35A60 , 32'hF6B1C250 , 32'h05C85840 , 32'h0E942DC0 , 32'hF90D8AC0 , 32'h0008A0BC , 32'hEAAF2F00 , 32'hFC7BFD0C , 32'h0BB47E10 , 32'hF6C06450 , 32'hEFA36EA0 , 32'hFFF6FC10 , 32'h02912780 , 32'h19367DA0 , 32'h06B2E158 , 32'h09146C10 , 32'hFFF93EE9 , 32'h1171AD60 , 32'hF94512A8 , 32'h0590EB48 , 32'h11056040 , 32'h0B166940} , 
{32'hFC4F6D38 , 32'h1278F860 , 32'h01322230 , 32'h00059CF0 , 32'h0005734C , 32'hEEC05B40 , 32'h181CC740 , 32'h0E2ACB90 , 32'h000E815F , 32'hFAEFB1E8 , 32'h09ED6FA0 , 32'hFF4C7382 , 32'h030B9E88 , 32'h032848D8 , 32'hFEAB9B90 , 32'hF39E11C0 , 32'h08064520 , 32'hFEDFED38 , 32'h08DF1930 , 32'hFFFF24D9 , 32'h04705D58 , 32'h1356FA60 , 32'hEAB86440 , 32'h00042800 , 32'hFF84D793 , 32'h23E1DFC0 , 32'h07CC0D70 , 32'h10D7EC20 , 32'h03D5AA60 , 32'hF08E32B0 , 32'hF3CC8800 , 32'hF504AE10 , 32'hFA9027D8 , 32'hFF2388AE , 32'h000F6E50 , 32'h0BCD9A70 , 32'hEF02D160 , 32'h03830370 , 32'hFB7741F8 , 32'h0326E7E8 , 32'h05DCC6D0 , 32'hFD7EC620 , 32'hFB1931A8 , 32'h00C72236 , 32'h02A67C24 , 32'hF4B248B0 , 32'hFC20090C , 32'hFD515338 , 32'hF22B6AD0 , 32'h0818DFE0 , 32'hFD2A9260 , 32'h08A4C6A0 , 32'h09C4D7B0 , 32'hF15295E0 , 32'h116E1C80 , 32'h198C6CC0 , 32'h04D120A8 , 32'hFB087C90 , 32'h08D4C750 , 32'h13E86900 , 32'h0C9DABF0 , 32'h06538188 , 32'h0FB1E4B0 , 32'h2E7FE800 , 32'hFE31A138 , 32'hFF8B785C , 32'hFFFECD4A , 32'h0D35D6B0 , 32'h028AA1DC , 32'h10DE6A40 , 32'h1889DBE0 , 32'hFFBFE95E , 32'hFD0DA134 , 32'h0A209350 , 32'hFAB39538 , 32'hE4C3D2A0 , 32'hED640DC0 , 32'hED48F760 , 32'hFE3F03AC , 32'h04D53128 , 32'hEBE850E0 , 32'hF4C36A10 , 32'hF82875D0 , 32'hFFFC0524 , 32'h19429D20 , 32'h0B5680D0 , 32'h07E70FC0 , 32'hF7F060A0 , 32'h04F2FB18 , 32'hFFF72E12 , 32'hE53D2320 , 32'hF88437C8 , 32'h02974B78 , 32'h0297EA94 , 32'hFFFDA1F5 , 32'h05CC66F8 , 32'h03FFA808 , 32'h1038F7E0 , 32'hFD720770 , 32'hE49052C0} , 
{32'hFA182F10 , 32'h01C46EAC , 32'h0F64F6A0 , 32'h00036A36 , 32'hFFF8D7AF , 32'hFE9E2004 , 32'hF0200A80 , 32'hF0321CA0 , 32'hFFFE088A , 32'h041F5B38 , 32'hF38ACDE0 , 32'h0368B744 , 32'h036C9E44 , 32'hF4017CB0 , 32'hFF888275 , 32'hFD5FF300 , 32'h2128E440 , 32'hF7C21E40 , 32'h0815D150 , 32'hFFFFD7B7 , 32'hFAAFFDD8 , 32'h03E44604 , 32'hF9D0B330 , 32'hFFFAF710 , 32'h04BC9268 , 32'hFEFD9FFC , 32'hDC3F16C0 , 32'hF4652120 , 32'h06D0CEA8 , 32'hF7F692C0 , 32'hFD290044 , 32'hFD4C4DAC , 32'hF805E908 , 32'hFBC5F508 , 32'hFFF4D5D9 , 32'h074C1790 , 32'hFDF8F104 , 32'hF4536CB0 , 32'hF6341DB0 , 32'hF6004A30 , 32'h0993A7F0 , 32'hFC5E704C , 32'hF652B7D0 , 32'hE41784E0 , 32'h0201A9D4 , 32'h111B6180 , 32'h0375BF08 , 32'hF8713E90 , 32'hFD109B84 , 32'h0BE963F0 , 32'hF54594F0 , 32'hFFC26CAC , 32'hF8955218 , 32'h03C5B914 , 32'hF8D5E668 , 32'h23AFCE00 , 32'h1025A7E0 , 32'hF439FF00 , 32'h05F0F5C0 , 32'hF218E630 , 32'hFC562E60 , 32'h0E8D9820 , 32'hE2EEA5C0 , 32'hE7F85E40 , 32'h01A38FC0 , 32'hF126D0C0 , 32'h00042C97 , 32'h0A218370 , 32'h133D2360 , 32'hFC8B1FDC , 32'h1CBCDDC0 , 32'hEA9D33A0 , 32'hFB0A4980 , 32'h1CCBB9E0 , 32'hED8AC920 , 32'hE9342220 , 32'h0EC52900 , 32'hFED1D080 , 32'h0778EA28 , 32'h0434A708 , 32'h0C3E40E0 , 32'h005B3F84 , 32'hEE5CF3E0 , 32'h0007C6EF , 32'h05C5AD38 , 32'h11316E00 , 32'h04B8BEF0 , 32'hFD93CC98 , 32'h0BF9A5D0 , 32'hFFFCBEDD , 32'h17AEDA00 , 32'h19D3ACE0 , 32'h0E9CD9B0 , 32'hFB099C30 , 32'h0005010F , 32'h04E8E9A8 , 32'hF78F0070 , 32'h08D16B80 , 32'h033FAEC0 , 32'h04B88190} , 
{32'hF9EA7840 , 32'hDDA81C80 , 32'hFCD5920C , 32'h0009D199 , 32'hFFF77427 , 32'hFD63544C , 32'hFBCBF0A0 , 32'h0E50ED40 , 32'hFFFC8D85 , 32'h020F88B8 , 32'hEE4BAB40 , 32'h11EEA560 , 32'hFB6A9D10 , 32'h14E1B780 , 32'h155B2920 , 32'hFC9F956C , 32'h1288FE60 , 32'h0AB61F60 , 32'hFEE6B8C4 , 32'h000AF270 , 32'h052B7A98 , 32'hFEF4600C , 32'h08DC01D0 , 32'h000E0004 , 32'h05D01DB8 , 32'hF3FCFA30 , 32'hF79D9770 , 32'h1A57F380 , 32'h0D5748C0 , 32'h0DAD8520 , 32'hFC74E3C0 , 32'hFDD19BD4 , 32'hF2755A00 , 32'hF97DB990 , 32'h00002DEB , 32'hFF104DAC , 32'h0119A370 , 32'h03E41C94 , 32'hF358AAB0 , 32'h0030F924 , 32'hF6A7FC30 , 32'h0232073C , 32'hFFB372B8 , 32'h1E6F0180 , 32'hED02B7C0 , 32'h06BAFE68 , 32'h0C9B31C0 , 32'h095FD060 , 32'hE89F57E0 , 32'h0FB7A570 , 32'hEC011F80 , 32'hFE169884 , 32'h083511C0 , 32'h00E8B3DF , 32'h1BCCD820 , 32'hEAA19300 , 32'hFAF04730 , 32'hFFA3077F , 32'hFD1D3FA4 , 32'hFDE48FC0 , 32'h0354B7A0 , 32'h029768E8 , 32'h05F712B8 , 32'hF1AA36A0 , 32'hF32C2430 , 32'hFE0018F4 , 32'h00184616 , 32'hEC3788E0 , 32'hF97A3EE0 , 32'hE99D9AE0 , 32'h16D39980 , 32'h26A2A380 , 32'hF1866030 , 32'hFFC3E2C2 , 32'hF43DF000 , 32'hDDAA9B40 , 32'hFC68D0FC , 32'hFCDD3B64 , 32'hEBFF7220 , 32'h07EB1FA0 , 32'hFA748EF8 , 32'h1035BFE0 , 32'hFC3FFEBC , 32'h0003B0B9 , 32'h02AA8990 , 32'h0413FFE0 , 32'h013CB88C , 32'h0BC8FF50 , 32'hF7BA7400 , 32'h0009A43E , 32'h0474B150 , 32'h0D901980 , 32'h0D8B4D50 , 32'h0FA61810 , 32'h0007B3A1 , 32'hFC1B0438 , 32'hFF0DFACA , 32'hF338B560 , 32'hFEEA1580 , 32'hF4CFE540} , 
{32'h055F9E78 , 32'hFFFA832A , 32'h166D1F40 , 32'hFFF57EE3 , 32'h00096130 , 32'h0A27DE50 , 32'hF4E39300 , 32'hFFCFBA49 , 32'h00087A2A , 32'h02994DEC , 32'hF1B860E0 , 32'hFCF9EA8C , 32'h00533414 , 32'h192675C0 , 32'h0310E2C0 , 32'h051F4EE0 , 32'h0E406D80 , 32'h11FA9520 , 32'h0A8E0560 , 32'h00093373 , 32'hFF05A996 , 32'h02F6F120 , 32'h0E89E740 , 32'hFFFFD28F , 32'h00F2CAF9 , 32'hFD7C7F44 , 32'h1675AF40 , 32'h0B392470 , 32'hFEF715C8 , 32'hFB9C9AA8 , 32'hF9B739B8 , 32'h02C77B88 , 32'h07FF10F0 , 32'h0504CE50 , 32'hFFFF1869 , 32'h009E7138 , 32'h0DA4A110 , 32'hFF74AB87 , 32'hFE0A0480 , 32'hE99C91E0 , 32'hF5CCB350 , 32'hFE449658 , 32'hD3896AC0 , 32'hEE52B160 , 32'hF931CE28 , 32'hF70CB1F0 , 32'hF7151370 , 32'hE4AA1320 , 32'hF4C61440 , 32'hF77CD130 , 32'h00BBD41D , 32'hEFFA9A80 , 32'hF4EB91A0 , 32'hFFDAC28D , 32'hF7709090 , 32'h12B37000 , 32'hF27E92F0 , 32'h01BC4300 , 32'h01EE8998 , 32'hFCE61D2C , 32'hFA33DB10 , 32'h1D45EDC0 , 32'h09C8F910 , 32'h176C2DE0 , 32'h06C52570 , 32'h0AED67C0 , 32'h000805F4 , 32'hF9EB5DC0 , 32'hFFB9A47C , 32'hF0F72360 , 32'hEA826CE0 , 32'h1A9DBF80 , 32'hEBE4AE20 , 32'h271CC780 , 32'h0093415D , 32'h1A92DAE0 , 32'h0438FC08 , 32'h0B0886A0 , 32'hF687ED40 , 32'h040FCDC0 , 32'h00476B6C , 32'hFAE55878 , 32'h0BAE10F0 , 32'h000B2016 , 32'h0BC73B80 , 32'hF2D289C0 , 32'h12A8AA80 , 32'hFE31513C , 32'hF54BA900 , 32'hFFFBA5CA , 32'hEFEABE40 , 32'h0E5EC2A0 , 32'h01810964 , 32'hFA27EBA0 , 32'h0007982A , 32'h0E533820 , 32'hF9D2C398 , 32'hFFCAF7CA , 32'h00BCF316 , 32'h0BAC1690} , 
{32'h024478E0 , 32'h0EE789E0 , 32'h0663BE60 , 32'hFFF8A841 , 32'hFFEB6985 , 32'h01306654 , 32'h08C051E0 , 32'hF1079920 , 32'hFFFE1779 , 32'h07E130D0 , 32'h0CAA2DC0 , 32'hF00EF6A0 , 32'hFFA4FB9C , 32'hFD805388 , 32'hF76B5AC0 , 32'h05977908 , 32'h02EED204 , 32'h0481EE40 , 32'h088B0610 , 32'hFFF7AFD3 , 32'hF92BFF38 , 32'h06914918 , 32'h00ECA782 , 32'hFFFF840C , 32'hFE3587F0 , 32'hF6FB0080 , 32'h02861F78 , 32'h226A7880 , 32'h0B544E90 , 32'h0A01B0A0 , 32'h0BFCB7F0 , 32'hFD161FE4 , 32'hF6ED9DD0 , 32'hFE424A54 , 32'h0002507C , 32'h0D697010 , 32'h0017E4B8 , 32'hFEE9A958 , 32'hE1549C20 , 32'h014638B0 , 32'hF8B2D570 , 32'h03B74F3C , 32'h11AFE6A0 , 32'hEC695D80 , 32'hFB419CA0 , 32'h01634148 , 32'hFB1222F8 , 32'hFC191880 , 32'h006192F9 , 32'h0220474C , 32'h0E206FF0 , 32'hF983CCA8 , 32'hEB179BC0 , 32'h026EA254 , 32'hEF6DE4A0 , 32'hF0192340 , 32'hFAE4C450 , 32'hFBD1C2A8 , 32'h0D7F87C0 , 32'hF0E2BF40 , 32'h14BF79E0 , 32'hEAE0C660 , 32'h08CA68D0 , 32'hF846A6E0 , 32'h0ABFAD80 , 32'h0B986A20 , 32'hFFE5ED0A , 32'hEC2B4D20 , 32'h19D2A5E0 , 32'hEE4C6140 , 32'h0C1C12E0 , 32'h04AA95D8 , 32'hFAA23ED8 , 32'h01F74374 , 32'hDCF5FC00 , 32'hF71AB040 , 32'h085CDBE0 , 32'h03613470 , 32'h016B5018 , 32'hF583A680 , 32'hF2E5AA40 , 32'hFEF2FF44 , 32'h0675BD68 , 32'h000A8100 , 32'h040261D0 , 32'h04B18F70 , 32'h0D0C2420 , 32'hF3BCAC80 , 32'hF2DF2670 , 32'hFFFC05C2 , 32'h0B875FE0 , 32'hD1CFB300 , 32'hE2CC9760 , 32'hF31FB410 , 32'hFFFFBF49 , 32'h14437B60 , 32'hF0A79820 , 32'hF6098F90 , 32'h1400E1A0 , 32'hF382FBE0} , 
{32'h07A25650 , 32'h08F710E0 , 32'hFDA07398 , 32'hFFFB6426 , 32'hFFFCC426 , 32'hFD303848 , 32'hE2E94C80 , 32'hF1300F50 , 32'hFFFFFA00 , 32'h0D88C7C0 , 32'hF57F5F60 , 32'h01D825B4 , 32'hF7683500 , 32'hFDBA36E4 , 32'hFE0E66F4 , 32'hFBBACA30 , 32'hF4714820 , 32'h0BF3BF20 , 32'hFE0DA57C , 32'h0014FF62 , 32'h01345E98 , 32'hF724CD30 , 32'hEC2A0D00 , 32'h00000669 , 32'h00BB7D43 , 32'h1E0651C0 , 32'h24DA7440 , 32'hDCD98000 , 32'h0085DB34 , 32'h09BDC990 , 32'hFE641B98 , 32'h060A1308 , 32'hFA6A6860 , 32'hF0030430 , 32'hFFF99A14 , 32'hF20FFC60 , 32'h03D94CC0 , 32'h091A7270 , 32'hFCC75E58 , 32'hEFAA3B80 , 32'h1188C980 , 32'hFF47F0E0 , 32'h04BB9630 , 32'hEDADE960 , 32'hFC43E9C0 , 32'h0517F148 , 32'h0A071BD0 , 32'h093798C0 , 32'hFF9D2035 , 32'h09A348B0 , 32'hE1A20A20 , 32'h078DBDC0 , 32'hF5D66590 , 32'h09D3B270 , 32'h106BC280 , 32'hF71B7B70 , 32'hFFF85AA3 , 32'hFA9269E8 , 32'hE5861BE0 , 32'h006DF1B0 , 32'h11293A80 , 32'h0F251EB0 , 32'hFEF4FA34 , 32'hF8052C38 , 32'hEC69CBA0 , 32'hFB43F718 , 32'hFFFA182F , 32'hEC1F74A0 , 32'h02F27110 , 32'hE7B4E0C0 , 32'hFB42D9B0 , 32'hF01BBCB0 , 32'hF0F8D530 , 32'h0226AC04 , 32'h0B329550 , 32'hFA0F7008 , 32'h05DB1490 , 32'hEF8BFDC0 , 32'hF5C98410 , 32'hFD2E7BCC , 32'hEC29D080 , 32'hFCBB9118 , 32'h17A14180 , 32'h000C6390 , 32'h18122640 , 32'h0E2C74E0 , 32'hF4ACDB20 , 32'h03DC99B0 , 32'h07ED2E20 , 32'h00023E46 , 32'h014F70FC , 32'hEEB5D3A0 , 32'hF4212080 , 32'h02EB305C , 32'h0003AE5B , 32'h0A9B71B0 , 32'h13886D80 , 32'h058724B0 , 32'h0FB49720 , 32'h069DC938} , 
{32'hF701FDD0 , 32'h0BCBAF50 , 32'h04FD6278 , 32'h0009AC58 , 32'hFFFA7B1D , 32'h19A7C540 , 32'hFD1B24E8 , 32'hFF19A39B , 32'hFFF9C6CB , 32'hFBECF208 , 32'hF81BF8D8 , 32'h03F7D014 , 32'h079AFA90 , 32'hF7C72730 , 32'hFD440AE8 , 32'h047D68E8 , 32'hF71072F0 , 32'hEFD472A0 , 32'h027BF894 , 32'hFFF36F75 , 32'h03C7C618 , 32'hF6840660 , 32'hEBFCC780 , 32'h00008146 , 32'h08A4D720 , 32'h08549C00 , 32'h06F01268 , 32'hF757B9B0 , 32'h023D1768 , 32'hFBB20A88 , 32'h0AD53580 , 32'hF5CBC050 , 32'hFF2718E9 , 32'hF51B53F0 , 32'hFFEFB8C7 , 32'h04AB6AE8 , 32'h10244160 , 32'h0883D200 , 32'h07CC44C8 , 32'hF44C9960 , 32'h02F5A604 , 32'hFF08A07F , 32'h320E4D40 , 32'h05C33E20 , 32'hFBAAC930 , 32'hF9CA21D0 , 32'h08469140 , 32'hFF64F993 , 32'h07454BE8 , 32'hF8F30CA8 , 32'h0D37F0B0 , 32'h026FA608 , 32'h0C885B20 , 32'hFD1BBE5C , 32'h1605FCC0 , 32'h158C7E80 , 32'h00DB2B5E , 32'hFEAFFCF0 , 32'hFD1DDA8C , 32'hF6752220 , 32'hECC7EA80 , 32'hF1ACF780 , 32'hF667B710 , 32'h15D56E00 , 32'h0611F348 , 32'h0DE5FD50 , 32'hFFFD2A9C , 32'hF953F0C8 , 32'h28ADBF00 , 32'hEACFC7C0 , 32'hF0F99FF0 , 32'h1922B560 , 32'hF659C5A0 , 32'h0D98D6F0 , 32'hFAC6A0A0 , 32'hFFB0BD09 , 32'h1721AF60 , 32'h08166F00 , 32'h07B65FC0 , 32'hFE9D8454 , 32'hF0FEC640 , 32'hFD57DBAC , 32'h0B6B5310 , 32'h0006967A , 32'hF1353F70 , 32'hFE03FFEC , 32'hFDE8BE80 , 32'h0D2236D0 , 32'h03016314 , 32'hFFFFDD50 , 32'h0048EC9D , 32'h1E8EB000 , 32'hFA9919B8 , 32'h05B8E908 , 32'h0004D9C8 , 32'hFD912FAC , 32'hF9E7D870 , 32'hF5DB9570 , 32'hE3C03200 , 32'hE115B760} , 
{32'hF704CA60 , 32'hFB089370 , 32'h16EF1600 , 32'h00153661 , 32'hFFFB5EA6 , 32'hF86D68A0 , 32'h1A704C20 , 32'hF829F040 , 32'h00000480 , 32'h0602CD60 , 32'h03CD2B64 , 32'hFDB177AC , 32'hF6D6A1F0 , 32'h026AA2FC , 32'h0B8361C0 , 32'h01FE5C84 , 32'hFB7D3D30 , 32'hFFD6F5DD , 32'hF8376618 , 32'h00061BC0 , 32'hF7AF9310 , 32'h042C83A8 , 32'h0A3C50E0 , 32'h00038CCB , 32'hF363DD30 , 32'hF0688EE0 , 32'h0D227100 , 32'hFF398E0C , 32'h05FA5580 , 32'hEE6C67A0 , 32'h04A89EC0 , 32'h046D4348 , 32'hFDD56DE4 , 32'hF8B25880 , 32'hFFFD82C3 , 32'h0D2907D0 , 32'hF0BEA790 , 32'hF2F26760 , 32'hFACE6CE0 , 32'hFDC5D494 , 32'hFCD8F90C , 32'h01CCFDB4 , 32'h196C71A0 , 32'h00BFC54D , 32'hFDBC540C , 32'hFE0A6240 , 32'hFAFFF9E8 , 32'h01A92CD8 , 32'hF93CCA18 , 32'h0AB73810 , 32'h005679E4 , 32'hF863E9F0 , 32'h134B77A0 , 32'h19FBFB20 , 32'h13A2E900 , 32'hF77897E0 , 32'hF7A2E270 , 32'hFA6FAD50 , 32'h09C31690 , 32'hFA58D3F0 , 32'h038552B4 , 32'h165F70E0 , 32'hFFF7B974 , 32'hF7BAB790 , 32'h169DE7E0 , 32'h01B96364 , 32'h00025A4C , 32'hFAA4F6B8 , 32'hF34E0200 , 32'hFAA547F0 , 32'hE19E6CE0 , 32'hCD5E8EC0 , 32'h0DB6B920 , 32'h19137600 , 32'h04D897D0 , 32'hE6EC4F60 , 32'h14969D00 , 32'h0801C120 , 32'hFE3145B0 , 32'hF5E06FE0 , 32'hEB3B7C00 , 32'hFF27D3D1 , 32'hF3E44360 , 32'hFFFD1417 , 32'hF58879D0 , 32'hF6C42230 , 32'h00477E53 , 32'h04A0A260 , 32'hE4CCFD00 , 32'h000A52DB , 32'hE132E760 , 32'h0B101D60 , 32'h06FB0410 , 32'h12081800 , 32'h0005C642 , 32'h0261BB2C , 32'h074F7F10 , 32'hFD413928 , 32'h0BEE7B40 , 32'h0726AA88} , 
{32'h08104830 , 32'h0FE292C0 , 32'hED6ED6C0 , 32'hFFFA1711 , 32'h000D1161 , 32'h1E502D80 , 32'hFBF188F0 , 32'hF75D8BB0 , 32'h0006AE35 , 32'h06387F60 , 32'hFF86F754 , 32'hF2345420 , 32'h03B61190 , 32'hF498ECA0 , 32'h02902500 , 32'hFE872918 , 32'hE3F4B8A0 , 32'h06D54D28 , 32'hFCCE1CDC , 32'hFFEC09A5 , 32'hF9376B80 , 32'hF5004200 , 32'h021C4F54 , 32'hFFF93669 , 32'hF2B92000 , 32'h0CA43170 , 32'h146830E0 , 32'h1D3767A0 , 32'hF57C0B10 , 32'hFCEF71C0 , 32'hFDCB8CA0 , 32'hEE42B220 , 32'hFD248474 , 32'hF657B1D0 , 32'hFFF9805A , 32'h02DEC314 , 32'hFC495540 , 32'h034B9B84 , 32'hE2BA4DE0 , 32'h086747C0 , 32'h06BA3990 , 32'h0567A7E0 , 32'hE4D42500 , 32'h01F9D180 , 32'h08D83510 , 32'hF67ABFB0 , 32'hFA8DB548 , 32'hFE5DA7EC , 32'h016A1C9C , 32'h09332080 , 32'h01C3ADE4 , 32'h100F8EA0 , 32'h0ABA7B20 , 32'h017003D0 , 32'hFFC2EF15 , 32'hF7F21FF0 , 32'h1A150C20 , 32'hFF25EF3D , 32'h12145900 , 32'h005798C3 , 32'hFEDB2CC4 , 32'hFF1B5AFF , 32'h01BC5F08 , 32'hD086C640 , 32'h061CC988 , 32'hF8E33A38 , 32'h0012A9BD , 32'hFACDCC10 , 32'hFB8251B8 , 32'h0B308C90 , 32'h17E33100 , 32'h07921808 , 32'h024FBBF4 , 32'h1478EB60 , 32'h0C1F8220 , 32'h0DDC6A90 , 32'h117427A0 , 32'hF9DA4888 , 32'h062847B0 , 32'h0C78F4C0 , 32'hEE40D6E0 , 32'hF67BA600 , 32'h111ADAA0 , 32'h000442B7 , 32'hF0476110 , 32'h02192A24 , 32'h058F93B8 , 32'h07D00EA0 , 32'h04FF0D18 , 32'h000824DB , 32'hEB3EE380 , 32'h116EE0C0 , 32'h174EEBC0 , 32'hF2D91EA0 , 32'h00053056 , 32'hEB9CD540 , 32'h0453CDA8 , 32'hFD262E1C , 32'h000ABEBF , 32'hF0529C60} , 
{32'h054E22C8 , 32'hF79D8C70 , 32'h0CDBA2A0 , 32'h00081D63 , 32'h000D2B59 , 32'hFF1CC377 , 32'hF1419790 , 32'h13328440 , 32'hFFFD22CA , 32'h09A753A0 , 32'hF401BCC0 , 32'h0E50C1E0 , 32'hF4245B60 , 32'h0A0B4670 , 32'h06BBCD98 , 32'hFB82E138 , 32'hF10C6CC0 , 32'h03B36724 , 32'h0AE20830 , 32'hFFF1C462 , 32'hF4616490 , 32'h004DEF10 , 32'h0EDCEDB0 , 32'hFFFBCFBD , 32'h0C5013E0 , 32'hFF95E2E7 , 32'hFCD00538 , 32'hFA0BE458 , 32'hFF420287 , 32'h00C15FC3 , 32'hEFB77C20 , 32'h0D0C0220 , 32'hFCA54E28 , 32'h092202F0 , 32'h0009D40C , 32'hFB146F48 , 32'hD27B3CC0 , 32'h07840E80 , 32'hF885AAF0 , 32'h063EACC8 , 32'h041766D0 , 32'h05990920 , 32'h217C1700 , 32'hF5020F50 , 32'h0B2904B0 , 32'hEE5AFC60 , 32'h0D318360 , 32'hEED2ADE0 , 32'hF8C25FE8 , 32'h004F98EA , 32'h0BE91180 , 32'hFAD68558 , 32'hFE464F04 , 32'hE3401180 , 32'hF525E6A0 , 32'h126AF2C0 , 32'hF92F91F0 , 32'hFD26E6B4 , 32'hF216E9A0 , 32'h14886BC0 , 32'h19A4BCE0 , 32'hEBB88620 , 32'h1874FE80 , 32'hE1CFA3A0 , 32'hEDDE3CC0 , 32'h066F4A40 , 32'h00035944 , 32'h050637D0 , 32'h0AD099E0 , 32'h17F19460 , 32'hEF152BC0 , 32'hF5786B10 , 32'hF4E32AF0 , 32'h08EC1FB0 , 32'hFA7E1580 , 32'h0C3AEB30 , 32'hFD823F94 , 32'hF2501D60 , 32'h03F0B65C , 32'h0DF16140 , 32'hFFE94454 , 32'h052A1588 , 32'h086BA8A0 , 32'h0001C4FF , 32'h0C7F6AB0 , 32'hFE7D2D60 , 32'h04236F98 , 32'hFEF30890 , 32'hEB6C9860 , 32'h000F7F2E , 32'h082DF830 , 32'h1826E620 , 32'h02F66734 , 32'hFE031E6C , 32'hFFEEC5A0 , 32'hFF5CD685 , 32'hF57C8630 , 32'hEEF6D980 , 32'h08DA1820 , 32'hF9EF6328} , 
{32'hF6B8EFC0 , 32'h070C6818 , 32'h049DB9F8 , 32'hFFF6D1B5 , 32'hFFFEE8FD , 32'h031C2028 , 32'hF6FC2910 , 32'hEB4EF320 , 32'h0006EC03 , 32'hF3D9BC00 , 32'hFF17067C , 32'h02956CB8 , 32'hFCC19CA4 , 32'h058846E8 , 32'h173F4640 , 32'h08313C80 , 32'hFB238210 , 32'hFEEA0EB0 , 32'hEDD99A60 , 32'hFFF6DD59 , 32'h0545B968 , 32'h0CA01520 , 32'h0362E494 , 32'h000133EB , 32'h02BE4A74 , 32'h0478CF28 , 32'hEE28ECA0 , 32'hF9DBB138 , 32'h06E40FF8 , 32'hF71C92A0 , 32'h00FD5A80 , 32'hF1FC2290 , 32'h0A1A1060 , 32'h04C43CE8 , 32'hFFF7C626 , 32'hFE65D5D8 , 32'hDF8F7380 , 32'hFAE5F280 , 32'hFEA21728 , 32'hFF3E099A , 32'hFB87B6F0 , 32'h0042A3C8 , 32'hE3E9BF00 , 32'h03091104 , 32'hF3186B90 , 32'hFFA490BE , 32'h105BB680 , 32'h01CC4958 , 32'h1A2263E0 , 32'h003F1F90 , 32'hF23A2E20 , 32'hEB4B96E0 , 32'h02D285F8 , 32'h0606FB28 , 32'hFD1B169C , 32'hFE79E614 , 32'hF770A6E0 , 32'hFCE47598 , 32'hF083F8E0 , 32'h1DCC9880 , 32'hFB74E9B8 , 32'h094AF7E0 , 32'h0A7AB810 , 32'hFBE47E98 , 32'h02AEBFAC , 32'h00E2A2FF , 32'hFFFD1692 , 32'hFA360B20 , 32'h392BFF00 , 32'hF9C88F70 , 32'hF2C398E0 , 32'h028CF4E0 , 32'h0D6AC910 , 32'hF7B69E70 , 32'h1360AA20 , 32'h02F7C880 , 32'h0100C39C , 32'h1099EE80 , 32'hF5BD5650 , 32'h0ED81510 , 32'hF3C447A0 , 32'hFC462058 , 32'hF3D08480 , 32'h000FE7C7 , 32'hF170D170 , 32'hFF546DFA , 32'h0D112140 , 32'hF793B090 , 32'h005BAF68 , 32'hFFF5C3A7 , 32'h08940180 , 32'hDCAF2E40 , 32'h1A94F480 , 32'h0C524000 , 32'hFFE38BCE , 32'hF44353A0 , 32'h02F0C658 , 32'h039C1390 , 32'h0153C6FC , 32'hE97C9420} , 
{32'hFB6E3718 , 32'h1898E020 , 32'h07F4D030 , 32'h000D8BBC , 32'h0011EB80 , 32'h02D553AC , 32'hF0D6A280 , 32'hF2633BA0 , 32'hFFF960FD , 32'hFA284270 , 32'h055B2970 , 32'hFA7BD460 , 32'h0F2E1D90 , 32'h0269C208 , 32'hFA9D5000 , 32'h06AF1DC0 , 32'h09CD31E0 , 32'hF3F3E600 , 32'h0586AA00 , 32'h000F806F , 32'hF893C780 , 32'h0B5D2160 , 32'h115E9FE0 , 32'hFFE914B3 , 32'h030B3748 , 32'h056D4760 , 32'hFDA25418 , 32'h0AB42680 , 32'hF9B5B9B0 , 32'h000A146E , 32'h04E87758 , 32'hF57A5B20 , 32'hF81EA318 , 32'hF95A1C18 , 32'h000C02D4 , 32'hF7D836A0 , 32'hE7877F60 , 32'hEFC81660 , 32'hFD5D0CA8 , 32'h0099DAD4 , 32'hFC99E49C , 32'hFDBF3758 , 32'h0DDC49D0 , 32'h096FCE60 , 32'h0F25E0A0 , 32'h0F848FC0 , 32'h189B54A0 , 32'hF9836BB8 , 32'h0BF0CA50 , 32'hF4757CA0 , 32'hF7AC51B0 , 32'hFC80022C , 32'hFBF1BD50 , 32'h07242DC0 , 32'hE6EAE420 , 32'h18B88D20 , 32'h079409B0 , 32'hF6E1FA40 , 32'hF4385DD0 , 32'h068646D8 , 32'h08B2B0E0 , 32'h0C8AB520 , 32'h0AAEE100 , 32'h004306FA , 32'hFA2847C0 , 32'h0E5B1E00 , 32'h0005741A , 32'hFCAB1AF0 , 32'hC0D76140 , 32'hE2017820 , 32'hF7754150 , 32'h053CDAF8 , 32'h06EED6C8 , 32'hEB0B3B60 , 32'h028D4EB8 , 32'hEE7C8140 , 32'h0E70ED10 , 32'h06178C90 , 32'hE2D56740 , 32'hF7C9E950 , 32'hFF15606F , 32'hF7B00EB0 , 32'h07A24310 , 32'hFFF0A6B4 , 32'hFD1730D4 , 32'hF789FE70 , 32'h078BCA30 , 32'hFD07AD34 , 32'h1152DA80 , 32'hFFF609E0 , 32'hFFC1E231 , 32'h05F3B740 , 32'hFC826318 , 32'hF1493840 , 32'hFFEDE484 , 32'hF66F8300 , 32'hFA726A40 , 32'hF940E058 , 32'hF21D8770 , 32'hE7DF1260} , 
{32'h00E8FC5C , 32'h0CCCFBC0 , 32'hF9B51880 , 32'hFFEF998E , 32'hFFF42D2F , 32'hF819B100 , 32'h07106C30 , 32'hF359C980 , 32'hFFF31D95 , 32'h05562D08 , 32'h03A987D0 , 32'hFBD6E7A0 , 32'hFA774FF0 , 32'h005ACDA4 , 32'h0B685F00 , 32'h0C9FFD80 , 32'hFCD797EC , 32'h017F276C , 32'hFE532338 , 32'hFFFF1711 , 32'h00D8FF6B , 32'hFD764CAC , 32'hFA3885B0 , 32'h0004E473 , 32'hFACA50A8 , 32'h04C70830 , 32'h06676BC0 , 32'h08452520 , 32'h07540D90 , 32'hFD2901B0 , 32'h043B3788 , 32'hFD26254C , 32'hFD410100 , 32'h0D1DF820 , 32'hFFFAE08A , 32'hEF3ABF80 , 32'h21EF0940 , 32'h00B709A1 , 32'hF3A0D330 , 32'h0AAFE440 , 32'hFDD76B5C , 32'hFFB1FD85 , 32'hF3ED8EC0 , 32'h0AAEF270 , 32'hFF88075E , 32'h07D445B0 , 32'h0AF33800 , 32'h0DDC7540 , 32'h02B725C4 , 32'h035D6DD8 , 32'hF90896F8 , 32'hF50A1CD0 , 32'hF3FF6050 , 32'h039C9EC4 , 32'hE21BE800 , 32'hED47FDC0 , 32'hF7F4B1C0 , 32'hF7B942A0 , 32'h0D8DAB50 , 32'h0440B7D0 , 32'h0F9A7520 , 32'h026FB460 , 32'hFD9885A0 , 32'h0DA89B30 , 32'h063D09D0 , 32'h09158130 , 32'hFFFA41B1 , 32'hF7775990 , 32'h17203B80 , 32'h07476710 , 32'hEE8B0780 , 32'hE95200E0 , 32'h00E2D4E4 , 32'hE111DA20 , 32'hF783A9F0 , 32'hF7B2CE60 , 32'hEC029E00 , 32'hFCFB3F04 , 32'hFA25D970 , 32'h0A72EE60 , 32'hFCA6BD50 , 32'hF6977040 , 32'h02F144C8 , 32'h000BB987 , 32'h10C50760 , 32'hFF2653CA , 32'h08B92F30 , 32'hF221E3E0 , 32'h04BA8408 , 32'hFFF985D4 , 32'h08512F60 , 32'h4A4CB080 , 32'hFE28A000 , 32'h0101C878 , 32'h0001EB9F , 32'h02821B38 , 32'h0B34A450 , 32'hF6A7DE40 , 32'h112D68A0 , 32'hEEA82C80} , 
{32'hFF5AD539 , 32'h00BA4344 , 32'hFE596C00 , 32'h0010217F , 32'hFFE682BA , 32'hFF19035B , 32'h02EC93BC , 32'hFDFBCEA8 , 32'h00047540 , 32'hFDF12564 , 32'hFEA2B730 , 32'h016D3D44 , 32'h011C92E0 , 32'hFEE897F8 , 32'h00A0FD75 , 32'h003C7D66 , 32'h032F2EDC , 32'hFD14525C , 32'h0015705A , 32'h00105474 , 32'hFFB2B93A , 32'h01470458 , 32'hFD3D9548 , 32'h0015D89A , 32'hFF2C79E0 , 32'h01697A4C , 32'h012B14BC , 32'hFD9F4FB8 , 32'hFF4E596B , 32'hFD5CAD3C , 32'h0082964E , 32'h00CB6D56 , 32'h00CD9518 , 32'h005F446B , 32'h007B95EE , 32'hFFAF1B93 , 32'h02D5A07C , 32'h001CED97 , 32'h0197CDCC , 32'h002045F7 , 32'h00B4EE7D , 32'h7EF9CF80 , 32'h00CD6CCD , 32'h001E63AA , 32'hFE360E70 , 32'h01CA9E14 , 32'h020EBFD4 , 32'hFE4C6A1C , 32'h00949E41 , 32'h024B4920 , 32'h01516FC4 , 32'h0107A844 , 32'hFF1E9610 , 32'h02127138 , 32'hFE011220 , 32'h0386FFA4 , 32'h008076DA , 32'h00FAC693 , 32'hFDE8B418 , 32'h01035598 , 32'hFE4EADB4 , 32'h03235258 , 32'hFECC3644 , 32'h0311AAB0 , 32'hFFC7E000 , 32'h00D09B18 , 32'hFFC8B7DD , 32'h019CB974 , 32'hFEED7C84 , 32'hFCD735B0 , 32'hFFCD3FD8 , 32'h01A289DC , 32'hFE9B2F48 , 32'h0062CB19 , 32'hFF87B867 , 32'hFE283D18 , 32'hFD093294 , 32'h014F93B0 , 32'hFF5823EE , 32'hFFB17BF8 , 32'h02272004 , 32'hFC7FBD38 , 32'hFE8492BC , 32'hFFEC4FC6 , 32'h019C1A14 , 32'h0028C5FD , 32'h00B95CEE , 32'hFEC8E3F8 , 32'h025509B8 , 32'hFFB2E815 , 32'h015F5974 , 32'hFFA39F99 , 32'h01C8AB38 , 32'hFFD49AB1 , 32'h00127099 , 32'h005042B2 , 32'h003F3347 , 32'h032719C0 , 32'hFE478988 , 32'h045BED90} , 
{32'hFFFA5434 , 32'hFFF25219 , 32'hFFFA9CED , 32'h04B1F888 , 32'h0B359900 , 32'h00003650 , 32'hFFFE1CF5 , 32'h00058D3F , 32'h1818C720 , 32'h0000DC3E , 32'hFFF9CABB , 32'h0000AB8B , 32'hFFFDED7F , 32'h0008AB6A , 32'hFFFD5B44 , 32'h0001C0A7 , 32'hFFFBA096 , 32'h0003081D , 32'h0002D4B1 , 32'hE39526C0 , 32'h00009BDF , 32'hFFFB6740 , 32'h00021074 , 32'h07A9D2F0 , 32'h0004544F , 32'hFFFA6853 , 32'h00039205 , 32'h00031DC8 , 32'h0005A72F , 32'h00071C67 , 32'h00000116 , 32'hFFFFEC60 , 32'hFFFD72B4 , 32'hFFFDA62D , 32'hFDEFF3B4 , 32'hFFFFD8A7 , 32'h0006D6E1 , 32'h00000C1E , 32'hFFFDCB1B , 32'hFFFB7565 , 32'h000007A0 , 32'hFFC2BFE4 , 32'h0001A097 , 32'hFFFE4A00 , 32'hFFFA0D2C , 32'h00061C22 , 32'h0000B89E , 32'hFFFED5FA , 32'hFFF7E551 , 32'h00088B35 , 32'h00009877 , 32'hFFFBD65E , 32'h00084AD1 , 32'h0001D5B8 , 32'h0010FE95 , 32'hFFFB9D5A , 32'h000018B6 , 32'h0005618B , 32'h0004706E , 32'hFFFC8D79 , 32'hFFFEBCD1 , 32'h00049B8E , 32'h00000C82 , 32'hFFF11491 , 32'hFFFD5028 , 32'hFFF90D6C , 32'hACF29880 , 32'hFFFB3AAE , 32'hFFE87C83 , 32'h0002F921 , 32'h0007CAAE , 32'hFFFF5D48 , 32'hFFF99EF2 , 32'h00054336 , 32'h0002E9DE , 32'hFFFF51E2 , 32'hFFFE8534 , 32'hFFFC453F , 32'h00023A8C , 32'h0003A063 , 32'hFFFA71FB , 32'h00052EC0 , 32'h00028DC9 , 32'h13AC80E0 , 32'hFFFD4DD5 , 32'hFFFACC16 , 32'hFFFF9480 , 32'h000B90A4 , 32'hFFFFDEF7 , 32'hBADF7880 , 32'hFFFBAFAB , 32'h0012C7A2 , 32'h00062F76 , 32'h0001319D , 32'hCBD47C00 , 32'hFFFE018D , 32'hFFFFDC69 , 32'hFFFC39A7 , 32'hFFF94D9B , 32'h00091ADA} , 
{32'hFFF8A17F , 32'hFFF8F3EB , 32'h00040BEC , 32'hCE734A40 , 32'h46AC0700 , 32'hFFFE2AE4 , 32'h0001C4A9 , 32'hFFFD92D2 , 32'hDDCACD40 , 32'hFFFCD73A , 32'hFFFD079F , 32'hFFFDAB40 , 32'h0000C0E3 , 32'h0002635A , 32'h0004E74F , 32'hFFFAC4F4 , 32'hFFFC6B28 , 32'hFFFAEBF4 , 32'h0002DDED , 32'h2A6E7000 , 32'hFFFE7F05 , 32'h00023EBB , 32'h00020DA5 , 32'h39112680 , 32'hFFFF8070 , 32'h00000359 , 32'hFFF8828E , 32'h00059F6C , 32'hFFFC40E4 , 32'hFFFCE36B , 32'h0003FBAC , 32'h000035D6 , 32'hFFF7A5D7 , 32'h00020B5C , 32'hFF857FFA , 32'h00030121 , 32'hFFFAEBC2 , 32'hFFFB1BC3 , 32'h00002EBF , 32'h0005212E , 32'hFFFCF03E , 32'hFFFD85B8 , 32'h000515A5 , 32'hFFFF0481 , 32'h0000C671 , 32'h00019E0A , 32'h0002ACAE , 32'h000271C7 , 32'h0007DBFB , 32'hFFFFC5CA , 32'h00022644 , 32'h0001AF28 , 32'h0001B233 , 32'hFFFE479F , 32'h0003EF21 , 32'h000A122A , 32'h0006BA8D , 32'h00004D98 , 32'hFFFCE5E5 , 32'h00010A22 , 32'h0002E856 , 32'hFFFF76CF , 32'h00037FCF , 32'hFFFAFFBE , 32'h000492B1 , 32'hFFFF4645 , 32'hD8FF4B40 , 32'h0003621E , 32'h00016A91 , 32'h0005113B , 32'h0006BF63 , 32'h000158E7 , 32'h00022361 , 32'hFFFA12CF , 32'hFFFC31C0 , 32'hFFFE7283 , 32'h000C5D08 , 32'h00022F0B , 32'h00016E11 , 32'hFFFFF7E4 , 32'hFFF450E7 , 32'hFFFE9AF7 , 32'hFFFF60D8 , 32'h0DD78A90 , 32'hFFF4FB9E , 32'h00043395 , 32'h0004FEB7 , 32'hFFFD160B , 32'h000115EC , 32'h0EE57960 , 32'hFFFD0951 , 32'h0000CE9D , 32'hFFFF8E4B , 32'h0003F541 , 32'h1BC95BE0 , 32'h0000091D , 32'hFFFBF04F , 32'h000003DB , 32'hFFF9E9A5 , 32'h00016E26} , 
{32'hFFF853FD , 32'h0002B944 , 32'h0002C820 , 32'hC28A8380 , 32'hC2218E80 , 32'h00098769 , 32'hFFF25DBC , 32'h00033C42 , 32'h283C19C0 , 32'hFFFFD868 , 32'h0002B51D , 32'h00018240 , 32'hFFFF6C38 , 32'hFFFC2013 , 32'h0003350C , 32'h00031877 , 32'hFFF97FD2 , 32'h00013D7A , 32'hFFFCE141 , 32'h09BBFB50 , 32'hFFFC9F2F , 32'hFFFF94A8 , 32'h000EE389 , 32'h13026E20 , 32'h00002B47 , 32'h0001B95F , 32'hFFFB11A7 , 32'h0003DCC9 , 32'hFFFBCA62 , 32'hFFFB9707 , 32'hFFFDAC6D , 32'hFFFFDD66 , 32'hFFFE5B83 , 32'hFFFC98E0 , 32'h2974B140 , 32'h00001869 , 32'hFFEF3754 , 32'h000043AE , 32'hFFF9ECD2 , 32'h000482EF , 32'h0004AED1 , 32'hFFA86E6C , 32'h000E9363 , 32'h000093F6 , 32'hFFFE9356 , 32'hFFFE90E5 , 32'h0007AD26 , 32'hFFFD0C14 , 32'hFFFE6EA2 , 32'hFFFCB2E9 , 32'hFFFADFE1 , 32'h0000C26B , 32'h0008288F , 32'hFFFC620A , 32'h0001CC8B , 32'h0004CF33 , 32'h00016301 , 32'hFFF74E74 , 32'hFFFA7503 , 32'h0006F669 , 32'hFFFB7169 , 32'h000858BA , 32'h0003E2E2 , 32'hFFF38F01 , 32'hFFFA35BF , 32'hFFFFC962 , 32'hEE0DF940 , 32'h00027001 , 32'hFFFE008D , 32'h00073B5B , 32'hFFFDCF36 , 32'hFFFC4FFD , 32'hFFF7AFA6 , 32'hFFFD7B9C , 32'h00047502 , 32'h0006E518 , 32'h00081361 , 32'h00038767 , 32'hFFFCFFD3 , 32'hFFFD5CF7 , 32'h0003AA81 , 32'h0001DC4C , 32'h0004B4FA , 32'hDEDA16C0 , 32'hFFF87166 , 32'hFFF9540F , 32'h00004A53 , 32'h000736FE , 32'hFFF9882E , 32'hE1E6CDA0 , 32'hFFFEE246 , 32'h00075B69 , 32'h000522C3 , 32'h00068935 , 32'h338FBE40 , 32'hFFFD1777 , 32'h0000E8E8 , 32'hFFFC2E3F , 32'hFFF93788 , 32'hFFF982BA} , 
{32'hFFFBD049 , 32'hFFFFA642 , 32'hFFFFA662 , 32'h127C52C0 , 32'hE2E05E00 , 32'hFFFDED0D , 32'h0001DAEC , 32'h00075808 , 32'hE3C10D00 , 32'hFFFBAF7C , 32'hFFFCD474 , 32'h00050B34 , 32'hFFFF0A0A , 32'h0001AA85 , 32'h00016F33 , 32'h0002B24A , 32'h000217B6 , 32'hFFFDC528 , 32'h0002699B , 32'hF83C4800 , 32'h0000EB63 , 32'h00054BBC , 32'h000B59A9 , 32'hD6C900C0 , 32'hFFFF276A , 32'h00097B3F , 32'hFFFE7A09 , 32'h00060F79 , 32'hFFFB8447 , 32'hFFFDE0E0 , 32'hFFF846E1 , 32'h000208F2 , 32'h000452D5 , 32'h0004B72E , 32'hCD10A700 , 32'h00041B29 , 32'hFFF91767 , 32'hFFFEF303 , 32'h00038F07 , 32'hFFFFBDAF , 32'h0000A5E0 , 32'h001CBE12 , 32'hFFEE90F5 , 32'h00019153 , 32'hFFFC57D0 , 32'hFFFA626F , 32'h000547FD , 32'hFFFA2B87 , 32'hFFFCB27B , 32'h000578A1 , 32'hFFF92B1C , 32'hFFFC4BF4 , 32'h0005A010 , 32'hFFFF527E , 32'h0000C144 , 32'h00009269 , 32'h0004AB53 , 32'hFFF8F23D , 32'hFFF66AEF , 32'h0010AF2E , 32'h00021963 , 32'h0000CD84 , 32'h0009FB04 , 32'h0002A885 , 32'hFFFDA8C2 , 32'hFFFB4F25 , 32'hB31B5A80 , 32'h00018FDC , 32'hFFF8CDBE , 32'h000385D5 , 32'h0004713E , 32'h00068920 , 32'hFFFAE59F , 32'hFFFB367E , 32'h000813E8 , 32'h0001427C , 32'h000216E1 , 32'h0000AFDE , 32'hFFFA1F90 , 32'hFFFE8583 , 32'h00012238 , 32'h00050DBC , 32'h0002B289 , 32'hED9491C0 , 32'h00013B99 , 32'hFFFCA271 , 32'h0009AFFD , 32'hFFFD6C12 , 32'h00048588 , 32'h249B3A80 , 32'hFFFE1342 , 32'h0001BBB6 , 32'h000A6082 , 32'h000046CE , 32'h31820680 , 32'hFFFF0B33 , 32'h0002DD22 , 32'h00004ACB , 32'hFFF84B4B , 32'hFFFF304D} , 
{32'hFFF95E40 , 32'h00068104 , 32'h000103F0 , 32'hEE1D1940 , 32'h36C26F80 , 32'hFFFB07BF , 32'h000522B5 , 32'hFFFB44B7 , 32'h4EA1CC80 , 32'hFFFCF94E , 32'h00016476 , 32'h0002A04B , 32'hFFFC5903 , 32'hFFFF12CD , 32'hFFF9D5FB , 32'h0000D2A9 , 32'h0008E93E , 32'h0003B269 , 32'h000197B1 , 32'hC902D940 , 32'h0005B6EC , 32'hFFFFC0B9 , 32'h00003AAD , 32'hF10CB170 , 32'hFFFD0ED9 , 32'h00016AAE , 32'hFFFD3594 , 32'hFFF8D248 , 32'h00079243 , 32'h00048FA2 , 32'hFFFCEFE6 , 32'h00017682 , 32'hFFFEC1D6 , 32'h00007579 , 32'h07D25DA8 , 32'hFFFF89C2 , 32'h000549E8 , 32'hFFFDA1EE , 32'h0000A934 , 32'hFFF5FD1B , 32'hFFFCA14F , 32'h0023B981 , 32'h00036362 , 32'h00059605 , 32'hFFFD5D0C , 32'h000C7B55 , 32'h0001C9D3 , 32'h00068AC1 , 32'hFFF8D96F , 32'hFFFE449C , 32'hFFFC37FD , 32'hFFFCE783 , 32'hFFF8D5D8 , 32'h000C16A3 , 32'hFFFFE071 , 32'hFFF81ADA , 32'hFFFD98F8 , 32'hFFFD8191 , 32'hFFF99DD3 , 32'hFFFAC626 , 32'hFFFDED12 , 32'h0003614C , 32'hFFF72431 , 32'h0000D032 , 32'h00001073 , 32'h00045A2B , 32'hF6C709F0 , 32'hFFFFE91B , 32'h000795F4 , 32'hFFF454E8 , 32'hFFF862F7 , 32'h00031CE3 , 32'h0001AC00 , 32'hFFF6BDE7 , 32'hFFF95D55 , 32'hFFF41DE7 , 32'h0000A47E , 32'hFFFF42CB , 32'hFFF506BC , 32'hFFFBB07D , 32'h0002A2C8 , 32'h000267C6 , 32'hFFFD52BC , 32'hEB9563C0 , 32'h0003F5D1 , 32'h0001D41A , 32'h000474B0 , 32'hFFFF1AD3 , 32'h0004AA6D , 32'h36CD8BC0 , 32'h00080848 , 32'h00067F22 , 32'hFFF98968 , 32'h000340D1 , 32'h0849F5F0 , 32'h0006A808 , 32'h0004CB87 , 32'h0002AD9B , 32'h0000766F , 32'h0003674E} , 
{32'hFFFC624E , 32'h0000EDF9 , 32'hFFFF8E1F , 32'h0BB2BD60 , 32'h26564780 , 32'hFFF68B1E , 32'h0002326C , 32'h00022BF6 , 32'h1EC42940 , 32'h0004A558 , 32'hFFFEA2DF , 32'h00001C22 , 32'hFFFB52AC , 32'h00012CB5 , 32'hFFFFA5B6 , 32'hFFFEF908 , 32'hFFFE9DA3 , 32'hFFFB84D9 , 32'h00000EA2 , 32'h0C08CBC0 , 32'h0002A95F , 32'hFFFE17B3 , 32'hFFFE7559 , 32'hF6DEA280 , 32'h00033AA4 , 32'hFFF9E654 , 32'h0006570D , 32'h0001E452 , 32'h00058ED5 , 32'h00070335 , 32'h000584B4 , 32'h0002498E , 32'hFFFEAE93 , 32'h00027396 , 32'hBA6ED080 , 32'hFFFCB87F , 32'hFFF67E55 , 32'h0001758A , 32'hFFFE8A0A , 32'hFFFA3350 , 32'h00006F1E , 32'h00237AFD , 32'h0004310B , 32'h0000C99B , 32'h000041F7 , 32'h00024EC6 , 32'h00092DB8 , 32'hFFFE1757 , 32'hFFFCBEC0 , 32'h000059F3 , 32'h0005D21E , 32'h00005D6C , 32'hFFFDE1A6 , 32'h0001AD94 , 32'hFFFB6A8B , 32'h0000D8F0 , 32'hFFF9E3A8 , 32'hFFFFA08D , 32'hFFFDE62A , 32'h000518C1 , 32'h0008B445 , 32'hFFF489C5 , 32'h00016A20 , 32'hFFFE3A83 , 32'h00004CA3 , 32'h00028F57 , 32'h1FD09CC0 , 32'h0002F1BB , 32'h0005B305 , 32'h0006C99F , 32'h00019329 , 32'hFFFA1014 , 32'h0000BEEF , 32'hFFF6C09B , 32'hFFFAF08B , 32'h000213BD , 32'hFFFC1D50 , 32'h0001B135 , 32'h00028DFF , 32'h0002F759 , 32'hFFFCAD1F , 32'h0002C9A0 , 32'hFFFD9FB3 , 32'hECB90840 , 32'h000068C8 , 32'hFFFB692F , 32'h0003E1BF , 32'hFFFBD1E4 , 32'hFFFBDCBC , 32'hBB42BC80 , 32'h000530D4 , 32'hFFF8D572 , 32'hFFF91B46 , 32'h00046990 , 32'h3384BA40 , 32'hFFFC99CD , 32'hFFFCE700 , 32'hFFFC6578 , 32'h0008EB90 , 32'hFFFE4A32} , 
{32'hFFFF358F , 32'hFFF6443C , 32'h00003955 , 32'hBF52DE00 , 32'h02CA66B8 , 32'hFFF4DB40 , 32'h0003A10F , 32'h000400B5 , 32'hEFCB60C0 , 32'hFFFEE52D , 32'h00066460 , 32'h0004695E , 32'hFFFD90D9 , 32'hFFFB5369 , 32'h00058927 , 32'hFFF9DA11 , 32'h0002ABB1 , 32'h0001FD17 , 32'hFFFD1FD9 , 32'hE77D3180 , 32'hFFFFD7C1 , 32'hFFFD7F44 , 32'h00055A20 , 32'hBE2F9F80 , 32'h00004593 , 32'h00000155 , 32'hFFFEFD9F , 32'h00023B88 , 32'h00028D27 , 32'hFFFADA04 , 32'h00016501 , 32'h0003EE84 , 32'hFFFE43B8 , 32'hFFFBC53E , 32'hFE492290 , 32'h000194FD , 32'hFFF99CEE , 32'hFFFD69D4 , 32'h000562A1 , 32'h00024CA6 , 32'hFFFC4592 , 32'h002047D3 , 32'h000E8ACF , 32'h00070B51 , 32'hFFFE54E1 , 32'h0002D68B , 32'hFFFA2E3C , 32'h000185E7 , 32'hFFFC2B9B , 32'hFFFCB660 , 32'h000111D0 , 32'h0004F70A , 32'h000256FD , 32'hFFFC8921 , 32'h000B3D2C , 32'h000CDE2C , 32'hFFFEDE79 , 32'h00002FF0 , 32'hFFFD7FCF , 32'h0002272E , 32'hFFFE6E90 , 32'h0001EE0D , 32'h00041BF2 , 32'h0003EA24 , 32'h00025562 , 32'h000288A9 , 32'h0DC164D0 , 32'hFFFFC943 , 32'hFFEECD7C , 32'hFFFD9C1F , 32'hFFFFC1B0 , 32'hFFFEF276 , 32'hFFFFF694 , 32'hFFFB2495 , 32'hFFFE4AAF , 32'hFFF904F6 , 32'hFFFE6B02 , 32'h0001BC70 , 32'hFFFD4B11 , 32'hFFFB567D , 32'hFFFEA1D6 , 32'hFFFF317F , 32'hFFF4985C , 32'h4F8A7F80 , 32'hFFFDF164 , 32'h0000E49A , 32'hFFF17B9D , 32'h0000D68E , 32'hFFF9E774 , 32'hF2671690 , 32'hFFFB4091 , 32'hFFFDCDD1 , 32'hFFFE34CF , 32'h0002FF6F , 32'h1128C880 , 32'hFFFF4785 , 32'h00035B30 , 32'h00066CB6 , 32'hFFFC9A8C , 32'h000487A9} , 
{32'hFFFD2AB4 , 32'hFFFA5DB0 , 32'hFFFD4E35 , 32'h2080E580 , 32'h07C39BB0 , 32'h000C3514 , 32'h0002B30D , 32'hFFFD8DDA , 32'h34E839C0 , 32'h00040CB1 , 32'h000730A6 , 32'hFFFC98D8 , 32'hFFFE5125 , 32'hFFFD7F16 , 32'h0003134E , 32'h000B0BE6 , 32'hFFFF9914 , 32'hFFFFD75E , 32'hFFFF4051 , 32'h5A1D0B00 , 32'h00009D1D , 32'hFFF799D8 , 32'hFFFDDFE5 , 32'hD4F3A4C0 , 32'h000092EA , 32'h0004BB4C , 32'hFFF4C579 , 32'h000D0308 , 32'hFFF9E505 , 32'h000366B3 , 32'hFFFE15B2 , 32'hFFFA4458 , 32'hFFFFD8A7 , 32'h00001FCB , 32'h1C52FFE0 , 32'h00029291 , 32'h0001903B , 32'h0003E0F5 , 32'hFFFC3E2F , 32'h000B84D2 , 32'h00004D20 , 32'hFFDFC2EE , 32'h0003168E , 32'h000743C7 , 32'hFFFC054B , 32'hFFFCE432 , 32'hFFF72E26 , 32'h00014AEE , 32'h0004D124 , 32'hFFFE6AA6 , 32'h0006728C , 32'h00014F0C , 32'h0009743F , 32'hFFFA2D3F , 32'h0002C6D1 , 32'hFFFAFDA4 , 32'hFFFEDBC0 , 32'h0005FB5D , 32'h0000D5C2 , 32'hFFFFC2A1 , 32'hFFFFAF1E , 32'hFFF559B3 , 32'hFFFCFEB0 , 32'hFFFD3983 , 32'h0002CE6A , 32'h000030C4 , 32'hEBD5DC60 , 32'hFFFE9F57 , 32'h0011A484 , 32'h00057E4F , 32'hFFFE2C7D , 32'hFFFB502F , 32'hFFFE1093 , 32'hFFFF4DE2 , 32'hFFFE1945 , 32'h000B551C , 32'h0002FDC8 , 32'hFFFCBC95 , 32'h0002511F , 32'h0007A1B4 , 32'h0005EADE , 32'h0001F99F , 32'hFFFDD61E , 32'h22208A00 , 32'hFFFAD2E9 , 32'h00019C3B , 32'h00013450 , 32'hFFFE7464 , 32'h0003306E , 32'h0A512E80 , 32'h00060DE0 , 32'h00089749 , 32'h0004D010 , 32'hFFFA792C , 32'h03CD83C0 , 32'hFFFEDEA6 , 32'h000330F5 , 32'hFFFBE8B8 , 32'h0000DC93 , 32'h0000CF1A} , 
{32'hFFFE99FA , 32'hFFF99477 , 32'h00053AD4 , 32'hDE0FCF00 , 32'h20164F80 , 32'h0005BABF , 32'hFFFFA3E1 , 32'h00016526 , 32'hDEF387C0 , 32'h0003644A , 32'hFFF96D53 , 32'h00022E7F , 32'hFFF8DAC0 , 32'hFFFC33D2 , 32'h00066568 , 32'hFFFD081C , 32'hFFFA1749 , 32'h0000477F , 32'hFFFD94D9 , 32'h16B6DC40 , 32'h00064092 , 32'h00047DF8 , 32'hFFF7F42C , 32'hBD903280 , 32'hFFFD7F3F , 32'hFFFC680B , 32'h00058F2F , 32'hFFFFE316 , 32'h0005927C , 32'hFFFFE778 , 32'hFFFE9132 , 32'h0003BF7C , 32'hFFFE0E35 , 32'hFFFF03CE , 32'h163EA740 , 32'h0004D693 , 32'h000ADDB5 , 32'h00061643 , 32'hFFFA2AE3 , 32'hFFFEE09D , 32'hFFFC03E2 , 32'hFFEC44A9 , 32'h0003B415 , 32'hFFF96660 , 32'hFFFA03C7 , 32'hFFFC4B25 , 32'hFFFAD1FC , 32'h00027550 , 32'hFFF9F0A6 , 32'h00053F69 , 32'hFFFF3420 , 32'hFFFF0B8A , 32'hFFFF9763 , 32'h0006977D , 32'h00081091 , 32'hFFF3F1A1 , 32'hFFFB8036 , 32'hFFFF54A8 , 32'h00067E7F , 32'hFFF8EE98 , 32'hFFFDC8E2 , 32'hFFFE4D51 , 32'hFFFC64CA , 32'h0001D63D , 32'h0001B98E , 32'hFFFEF136 , 32'hFD7A6230 , 32'hFFF9704C , 32'h00174E92 , 32'hFFFE1B6F , 32'h0006C8AB , 32'h0005CA0B , 32'hFFFF01FD , 32'h000AE99C , 32'hFFFCAFEC , 32'hFFFBCEB6 , 32'hFFFFB554 , 32'hFFFD8644 , 32'h0005946A , 32'h000528F5 , 32'hFFFC5B2A , 32'h00010593 , 32'hFFFA8991 , 32'hB2066500 , 32'hFFFEDBF5 , 32'h0003C841 , 32'hFFFF83D0 , 32'h000341D9 , 32'hFFF6BB33 , 32'hEDACF9C0 , 32'h000144C0 , 32'h0004466A , 32'h00092331 , 32'h0005E1AB , 32'hDC744E40 , 32'h00001070 , 32'h000364EB , 32'hFFFFF8EB , 32'h00079B21 , 32'h0003621E} , 
{32'hFFFE64CA , 32'h0001E50F , 32'h00037F7D , 32'h36382F80 , 32'h1FF75B60 , 32'h000631AD , 32'hFFF5DF35 , 32'hFFF9D2D8 , 32'hE174CE20 , 32'h00039024 , 32'hFFFCD4DD , 32'hFFFDCDD8 , 32'hFFFD8E80 , 32'h00020C3E , 32'hFFFFEE01 , 32'hFFFF6E9E , 32'hFFFFEB4B , 32'h00008E09 , 32'hFFFAA21B , 32'hDD23FF40 , 32'h0005CC97 , 32'hFFFAD53A , 32'h00058215 , 32'hF5D6FEF0 , 32'hFFFEFB54 , 32'h00028A7B , 32'h0000476A , 32'hFFFD99D0 , 32'h0000C5CA , 32'h0000CC21 , 32'h000213F6 , 32'h00007C97 , 32'h0004E7DD , 32'h00020297 , 32'h4C962B00 , 32'hFFFFEEF7 , 32'h0002D42F , 32'hFFFB7477 , 32'hFFF8250B , 32'hFFFB8925 , 32'hFFFE8638 , 32'hFFA27454 , 32'hFFF6A824 , 32'hFFFF9966 , 32'hFFFF9ECB , 32'hFFFE307F , 32'h00036808 , 32'h0005A246 , 32'h000002E6 , 32'h0002FFF8 , 32'hFFF7C199 , 32'hFFFB5EAE , 32'hFFFB66DE , 32'hFFFCFA97 , 32'h00079B06 , 32'hFFF56A04 , 32'hFFFE0DF3 , 32'h00035F6D , 32'hFFFAEB51 , 32'h0005BEFB , 32'h0003D566 , 32'hFFFED325 , 32'hFFF89191 , 32'h00004969 , 32'hFFFD05F4 , 32'hFFFE252D , 32'hFA6F3BE8 , 32'hFFF9815E , 32'h0010A802 , 32'h00034E66 , 32'hFFFE3766 , 32'hFFFEDE55 , 32'h00050970 , 32'hFFF7E314 , 32'h00000AE7 , 32'h0005EF42 , 32'h00075C9F , 32'h0003284A , 32'h0001E4F2 , 32'hFFFFE524 , 32'hFFFB6339 , 32'h0004F339 , 32'hFFFDF451 , 32'h02B102BC , 32'hFFFC81B2 , 32'h0002E8E2 , 32'h0006A538 , 32'hFFFDFBB8 , 32'hFFFE18DF , 32'hE4097FA0 , 32'h00033A59 , 32'hFFFDC142 , 32'hFFFF5263 , 32'h0000498A , 32'h3B094480 , 32'hFFFD056F , 32'hFFFEC50E , 32'hFFFD4519 , 32'h00050DAA , 32'h0004001F}
};

logic signed [31:0] VT_3 [10][10] ='{
{32'hC3322280 , 32'hCBF809C0 , 32'h0FD8FC60 , 32'h2AAF9C00 , 32'h05207198 , 32'hFBE72948 , 32'hB8CF5C80 , 32'h2533BEC0 , 32'hFF0B2E64 , 32'h258E18C0} , 
{32'h28D97640 , 32'hBB452D00 , 32'h08DE5A00 , 32'h2A998180 , 32'hDC3B8D40 , 32'h1259CCE0 , 32'h07420990 , 32'hCE6C4E00 , 32'h3E3C8E00 , 32'hF6179A60} , 
{32'hC91ECB80 , 32'h1F27BFE0 , 32'h01FCA088 , 32'h332A5500 , 32'hD64C5F00 , 32'h19B580E0 , 32'h16BE6B60 , 32'h19A839A0 , 32'h08E6F560 , 32'hB1BCF480} , 
{32'h3D6545C0 , 32'h046B4568 , 32'h0481A2D0 , 32'h25499C40 , 32'h05B1BEA0 , 32'hACD64080 , 32'hEBE318C0 , 32'h3214E780 , 32'h02AD29BC , 32'hDBB92C00} , 
{32'h20F4D840 , 32'hDFF43400 , 32'hC855A0C0 , 32'h0AF42B10 , 32'hD2E241C0 , 32'h23D98A40 , 32'h21628780 , 32'h3DFC3100 , 32'hD54FDC00 , 32'h1EDD6480} , 
{32'h0B162860 , 32'hDF136B00 , 32'h63D03D80 , 32'hD8D1AF40 , 32'hDF1DAA40 , 32'h07F9C800 , 32'h0BB80300 , 32'h13F86DE0 , 32'hD74E6700 , 32'hED80EEA0} , 
{32'h15EC3740 , 32'h1F362B80 , 32'h0795CD40 , 32'h38464040 , 32'hE7B308A0 , 32'h062E0810 , 32'hDE787200 , 32'hC30E19C0 , 32'hB1B4ED80 , 32'h0A6252D0} , 
{32'h049B8B68 , 32'h34793DC0 , 32'h0635C500 , 32'hE51FCD20 , 32'hA84F6F80 , 32'hF30DE430 , 32'hDAA04480 , 32'h0927D2C0 , 32'h2BDA15C0 , 32'h27D89F00} , 
{32'h27AB5980 , 32'h040C41B0 , 32'hF076D420 , 32'hE2D6E140 , 32'h1138A400 , 32'h43365B80 , 32'hB1ABAF00 , 32'h100A2300 , 32'h04AE0928 , 32'hCE43F340} , 
{32'h1EDC9940 , 32'h2DE93A00 , 32'h334B5C40 , 32'h306B1800 , 32'h282B3F40 , 32'h30CC7880 , 32'h14CF8CC0 , 32'h20DA5DC0 , 32'h1D804600 , 32'h2C648340}
};

logic signed [31:0] US_0 [784][37] ='{
{32'hFFF92C07 , 32'h0000EB1A , 32'hFFFD5D02 , 32'hFFF09627 , 32'hFFFD1ED7 , 32'h000137F3 , 32'hFFFF0105 , 32'hFFFFAC32 , 32'h0002A16B , 32'h0000B006 , 32'h0001687E , 32'h0002324F , 32'hFFFEF4DD , 32'hFFFC66D8 , 32'hFFFCF97F , 32'h00031C7D , 32'hFFFDF35C , 32'hFFFB8C79 , 32'h000D898A , 32'hFFF70456 , 32'h00041BA1 , 32'hFFF780F4 , 32'hFFFCF3C8 , 32'hFFFC32C2 , 32'h0000D003 , 32'hFFFDE045 , 32'hFFF972BC , 32'h000C2CA0 , 32'hFFFC52DC , 32'hFFFEF738 , 32'hFFFE0916 , 32'hFFFA231C , 32'hFFFFEA46 , 32'h00011683 , 32'h0002E45A , 32'h0002F83E , 32'hFFF5B3ED} , 
{32'h0001D23B , 32'h0003D490 , 32'hFFF8F4A3 , 32'h000EF5FC , 32'h000596AB , 32'hFFFC116C , 32'h0002EED5 , 32'hFFFD2B87 , 32'h0005D47B , 32'h00007936 , 32'h000555C3 , 32'h00045662 , 32'hFFFE7DAB , 32'h0004C286 , 32'hFFFC855B , 32'hFFF58246 , 32'hFFF9C4FC , 32'hFFFC5859 , 32'h0001F4B4 , 32'h00034042 , 32'hFFFF9A6F , 32'h0001F38E , 32'h0003BD72 , 32'hFFF8E959 , 32'h00082B58 , 32'h00008ECE , 32'h000748C1 , 32'h00010EEE , 32'hFFFFF703 , 32'hFFFDEE48 , 32'hFFFCE1FD , 32'h00019807 , 32'h0004B340 , 32'hFFF93DBF , 32'hFFFF674C , 32'hFFFB2591 , 32'hFFF72B85} , 
{32'hFFF87A29 , 32'hFFFD6EAF , 32'hFFFD719C , 32'h000975B2 , 32'hFFFE42D9 , 32'h0008E51B , 32'hFFF702FF , 32'hFFFDB5C7 , 32'hFFFE1E75 , 32'hFFFC1BE7 , 32'hFFFFE398 , 32'hFFFAF7A6 , 32'h00028A8A , 32'h00000815 , 32'h000AD994 , 32'hFFFE0040 , 32'h0000249B , 32'h000660E2 , 32'h0000542B , 32'hFFFD5EDC , 32'h00014929 , 32'hFFFE34A9 , 32'hFFF42699 , 32'hFFFBD23A , 32'hFFFD0D68 , 32'hFFFC0269 , 32'h00045490 , 32'h0001A92A , 32'hFFFDD25E , 32'h0004462A , 32'h00085A3C , 32'hFFFCB090 , 32'hFFFA56C5 , 32'hFFFE9CC4 , 32'hFFF7EE3B , 32'hFFFBA668 , 32'h0008AF46} , 
{32'hFFFAF134 , 32'h00070E00 , 32'hFFF4D7AB , 32'hFFFCAD04 , 32'h0001AC8D , 32'h00006F54 , 32'hFFF79915 , 32'hFFFE0A3F , 32'h0008757B , 32'hFFFC725C , 32'hFFFF5858 , 32'h0000A6C8 , 32'h00009263 , 32'hFFFF8017 , 32'hFFF78467 , 32'h00118363 , 32'h0000778A , 32'h0003426F , 32'hFFFDB5B6 , 32'hFFF7077D , 32'h00010CF2 , 32'h000899E2 , 32'h0008105F , 32'hFFFE6748 , 32'hFFFDF3BA , 32'hFFFE01E2 , 32'h000355E1 , 32'h000521DE , 32'hFFFB8AD8 , 32'h00024FF1 , 32'hFFFF58F1 , 32'h00007886 , 32'h0003FC22 , 32'hFFFC491A , 32'h00006298 , 32'hFFFF783C , 32'h0002C7EB} , 
{32'hFFFF6588 , 32'h000190AE , 32'hFFFCE5D8 , 32'hFFFDE233 , 32'hFFFF76E7 , 32'h0009832B , 32'h00072142 , 32'h0000AC62 , 32'h0003029D , 32'hFFFA4AD2 , 32'hFFFBDC66 , 32'h00021CE0 , 32'h0007A836 , 32'hFFF48410 , 32'hFFFE8F3D , 32'hFFFA3865 , 32'hFFFA109C , 32'h00014F26 , 32'h00072952 , 32'hFFFD53B2 , 32'hFFFCE1E4 , 32'h0009B840 , 32'h000323FA , 32'h000232BB , 32'hFFF8F525 , 32'h0003829B , 32'h00036634 , 32'hFFFCEDCA , 32'hFFFACC09 , 32'hFFF7AE4C , 32'h00061C79 , 32'hFFFB074A , 32'h00077CEA , 32'h0001D36F , 32'hFFFD4651 , 32'hFFFDF8E2 , 32'hFFFA7F62} , 
{32'h000914CE , 32'h000C7058 , 32'hFFFBE0F9 , 32'h0003822F , 32'h000807B4 , 32'hFFFB338C , 32'hFFFA4590 , 32'h00029BFB , 32'hFFFF2088 , 32'h0000E9D2 , 32'h00076171 , 32'h00022962 , 32'h00035893 , 32'hFFF7C364 , 32'h000505A8 , 32'h0006F175 , 32'hFFFFF298 , 32'h0000EE18 , 32'hFFFB4CEF , 32'h000A8FD7 , 32'hFFFC3382 , 32'h00008862 , 32'h0001F09B , 32'h00044BDC , 32'hFFFBE79D , 32'h00037DDB , 32'h00005DBC , 32'h0001CEB9 , 32'hFFFD68E7 , 32'hFFF64300 , 32'h00020DBF , 32'h0000773F , 32'h0008492C , 32'h00015727 , 32'h00031857 , 32'h000437C1 , 32'hFFF49659} , 
{32'h000186A9 , 32'h000233E1 , 32'hFFFEA02B , 32'hFFFAF67E , 32'hFFFABD9C , 32'hFFF5E2B0 , 32'hFFFABBD6 , 32'h00022EF9 , 32'h00060C2F , 32'hFFFFD50D , 32'h00023469 , 32'hFFFE3FB5 , 32'h00059780 , 32'h0004550B , 32'hFFF8925B , 32'hFFF4802C , 32'h00019D5B , 32'h00005243 , 32'hFFF44F80 , 32'h0003FD1D , 32'h00027E60 , 32'h000B836D , 32'h0001AA44 , 32'hFFF79874 , 32'hFFFB5F81 , 32'hFFF4A442 , 32'hFFFDC27C , 32'hFFF763B6 , 32'hFFFE3D14 , 32'hFFFC48FB , 32'h00014B1E , 32'hFFFF23E2 , 32'h00098B1D , 32'hFFFD3A45 , 32'h00001F9E , 32'h00052D97 , 32'hFFFEDD51} , 
{32'h00021606 , 32'hFFF6FA2D , 32'hFFF97EE6 , 32'hFFF62294 , 32'hFFFF0A7E , 32'hFFFD243A , 32'h0005F8BE , 32'hFFFADE21 , 32'h000194BA , 32'h000481A9 , 32'hFFF48880 , 32'hFFFE52AB , 32'h0004216B , 32'hFFF9E9CF , 32'hFFFC6F77 , 32'h0002D822 , 32'h00080065 , 32'h0000EFD4 , 32'hFFFAAD70 , 32'hFFFA5686 , 32'hFFFD83FC , 32'hFFFE196E , 32'hFFFE5E31 , 32'h0003A59A , 32'hFFFA4530 , 32'h0000C597 , 32'h0006A528 , 32'hFFFABAF6 , 32'hFFFFCE31 , 32'hFFFADBB9 , 32'h000975D9 , 32'h000594EF , 32'hFFF8D98A , 32'hFFFFFC40 , 32'hFFF34DF8 , 32'hFFFEE909 , 32'hFFFD0733} , 
{32'hFFF92845 , 32'hFFF813BA , 32'hFFFCC331 , 32'hFFFF86C4 , 32'hFFFD7075 , 32'h0002BE6A , 32'hFFFD5584 , 32'hFFF92BF5 , 32'h0007D4AC , 32'hFFFC36FF , 32'h00016B52 , 32'hFFFCC66E , 32'h0001617F , 32'h000353F5 , 32'hFFF7D298 , 32'hFFFDEC7A , 32'hFFF9FEC5 , 32'hFFFEB103 , 32'hFFFE2811 , 32'h0001C3C7 , 32'h00047E72 , 32'h00006769 , 32'hFFFFA6A2 , 32'h00016907 , 32'h0004A583 , 32'h00050304 , 32'hFFF9444F , 32'hFFF71905 , 32'h0002385E , 32'h00026D0F , 32'h0000B754 , 32'hFFFB6225 , 32'hFFF85CB0 , 32'h0000B628 , 32'h0007D9DB , 32'h0009741F , 32'hFFFC0615} , 
{32'h0006F0D0 , 32'hFFFA0456 , 32'h0000B475 , 32'hFFFE6CDD , 32'h000520B0 , 32'h000485E9 , 32'h0007056D , 32'hFFFCDC48 , 32'h0006104A , 32'h0004077C , 32'h000134AB , 32'hFFFF6F4E , 32'hFFFD24A9 , 32'hFFF838C3 , 32'h00049FB4 , 32'h0005250B , 32'h00058A82 , 32'hFFFD7940 , 32'h0000D821 , 32'h00031A8C , 32'hFFFD0238 , 32'h00085E48 , 32'hFFFBD952 , 32'h00050E18 , 32'hFFFFE97D , 32'h00085AF0 , 32'hFFFCBCF5 , 32'hFFFED0C0 , 32'h0003D43D , 32'hFFFFEC68 , 32'h0007473C , 32'h00034F1F , 32'h00003353 , 32'h0005DB08 , 32'h000469DD , 32'h00076FD2 , 32'h0006F241} , 
{32'hFFFE5B1C , 32'hFFF8719D , 32'h00005398 , 32'h00043206 , 32'hFFFFC794 , 32'hFFF9F530 , 32'h0003BC9C , 32'h00080F58 , 32'hFFFCFAD8 , 32'hFFFFCEAB , 32'hFFFF965C , 32'hFFFAB806 , 32'hFFFDCCF8 , 32'hFFFCE9ED , 32'h00053016 , 32'h00030095 , 32'hFFFD9966 , 32'hFFF927A1 , 32'h0002CB34 , 32'hFFFBDA97 , 32'h000183CE , 32'hFFFE7F61 , 32'h00040B7F , 32'hFFFF03C9 , 32'hFFFD9980 , 32'hFFF9352B , 32'h0005444C , 32'h00007295 , 32'hFFF35683 , 32'hFFFE995D , 32'hFFFED542 , 32'hFFFF23C2 , 32'h00030B95 , 32'hFFFF5BDF , 32'h0005901F , 32'hFFFFEA19 , 32'h00062984} , 
{32'hFFFCB286 , 32'h0005CAC4 , 32'h0002DD85 , 32'hFFFF14A7 , 32'h000280D5 , 32'hFFFFB16A , 32'hFFF902E1 , 32'h00014E4C , 32'hFFFF7586 , 32'hFFFD973E , 32'h0007AA3A , 32'hFFFA9E92 , 32'hFFF72092 , 32'hFFFAB093 , 32'h0001207F , 32'hFFFB5EF2 , 32'hFFFCC416 , 32'h00069164 , 32'h0003DD2A , 32'h000774EF , 32'h00081EF6 , 32'hFFFF5346 , 32'h0008FFDF , 32'h00015ED2 , 32'hFFFF761E , 32'h0003D20C , 32'hFFFFEEE2 , 32'h00031417 , 32'hFFFB0EB5 , 32'h00055F32 , 32'h000457F5 , 32'h0001F2E8 , 32'h0000B330 , 32'h000415CF , 32'hFFFD338A , 32'hFFFD57D4 , 32'hFFFFBA20} , 
{32'h0003945C , 32'h0002B920 , 32'h0008F446 , 32'hFFFCCCE2 , 32'hFFF9E2FF , 32'h0009AF2A , 32'h0002F54C , 32'hFFFB2016 , 32'hFFFCA79F , 32'h0004C197 , 32'h00033A8E , 32'hFFFF777A , 32'hFFF7FC37 , 32'hFFFB7920 , 32'h00020FBD , 32'h00014D6D , 32'h0000284F , 32'h000403C4 , 32'hFFFE6A26 , 32'h000A03C4 , 32'hFFFCEB6F , 32'h000061E9 , 32'hFFFFAF6D , 32'hFFFC4363 , 32'h0004CB7B , 32'hFFF6E93F , 32'hFFFC6120 , 32'hFFFBC7E8 , 32'h0001A2D2 , 32'h0005E3E3 , 32'h00082978 , 32'h000227B9 , 32'h0006A66E , 32'h0003AD5A , 32'hFFFB4564 , 32'hFFFDE88C , 32'hFFFB851D} , 
{32'hFFFCE6A3 , 32'hFFFAD1C0 , 32'h00008B38 , 32'hFFFD3E31 , 32'hFFFE447F , 32'h000A64DB , 32'hFFFDDADD , 32'hFFF3E612 , 32'hFFFA6E16 , 32'hFFF9EC23 , 32'hFFFB6370 , 32'hFFFDF535 , 32'hFFFDB9AB , 32'hFFFE2DD4 , 32'hFFFAB959 , 32'h00030563 , 32'h00045FA4 , 32'hFFFEEE0B , 32'h0006E99B , 32'h000378C2 , 32'hFFFEE1A3 , 32'hFFFF6A41 , 32'hFFF70648 , 32'h0002E16F , 32'h0001179C , 32'h0006B461 , 32'hFFFB7EAC , 32'h0000309C , 32'h0008CECC , 32'h00044EDB , 32'hFFFEFA5A , 32'hFFFD6C90 , 32'hFFF2F4B6 , 32'hFFFFFDCE , 32'h00020671 , 32'hFFF97A12 , 32'hFFFEAD8E} , 
{32'h0003A11A , 32'hFFFE4898 , 32'h00080835 , 32'h000131E1 , 32'h000080A4 , 32'h00014B15 , 32'h00006EB4 , 32'hFFF9AE3D , 32'h00066DA8 , 32'h0006E54E , 32'hFFFE621A , 32'hFFFE4B4D , 32'hFFFB12A5 , 32'hFFFF6E8D , 32'hFFFAF66F , 32'h0000DA0B , 32'hFFFFC834 , 32'h0000358B , 32'hFFF88DBD , 32'h00085B95 , 32'hFFFCFA1F , 32'h0004BEE6 , 32'h000305EF , 32'h0000F602 , 32'hFFF94E38 , 32'hFFFFAB29 , 32'h0002B080 , 32'hFFFBEB72 , 32'hFFFBBBEA , 32'hFFF6E497 , 32'h000C6807 , 32'h0002BEC5 , 32'hFFFC6B30 , 32'hFFFEEB49 , 32'h00022187 , 32'hFFFC83E6 , 32'hFFFB7BA4} , 
{32'h0002FD85 , 32'h0004CA70 , 32'h0000735E , 32'h000027CE , 32'hFFFE8B4F , 32'h0004B3AF , 32'hFFFC4FD0 , 32'hFFF88BFD , 32'h000FD0F3 , 32'h00042B05 , 32'hFFFB7C38 , 32'h0006E72C , 32'hFFFCACF5 , 32'hFFFF42A9 , 32'h00038211 , 32'hFFFEAC65 , 32'h00018E73 , 32'hFFFBE1E1 , 32'h0002BF03 , 32'h000891EE , 32'h00083EA2 , 32'hFFFFE680 , 32'h0007AE9C , 32'h00002E18 , 32'hFFFF00F3 , 32'hFFFCEF8E , 32'h000586B7 , 32'hFFFE468A , 32'h0004F5CA , 32'hFFFD1FED , 32'hFFFF42FE , 32'hFFFFD84A , 32'h00046BC0 , 32'hFFFBFD0A , 32'hFFF73D59 , 32'hFFFAB181 , 32'h00074C98} , 
{32'h00063113 , 32'h0008E052 , 32'h0009CE70 , 32'hFFFFD4F3 , 32'h00079788 , 32'hFFFC7630 , 32'h000A9B9E , 32'h0008E7AB , 32'hFFFF273B , 32'h0007CAA9 , 32'hFFFF9C63 , 32'hFFF3D094 , 32'hFFFF8DC3 , 32'hFFFEC355 , 32'hFFFB14A2 , 32'h00004D90 , 32'h000712A1 , 32'hFFFEF595 , 32'h000493A3 , 32'h000B5B81 , 32'h00061E2D , 32'h0008CFDA , 32'hFFF97D4F , 32'h000038D5 , 32'h0000BAA9 , 32'hFFF6C5EC , 32'hFFFD6B47 , 32'h00048E1F , 32'hFFFEA175 , 32'h00021FA3 , 32'hFFF89CE5 , 32'h00026F12 , 32'h0005C2F1 , 32'h0000DF90 , 32'h00024B56 , 32'hFFFA00D7 , 32'hFFFE5DB1} , 
{32'hFFFC1EA5 , 32'hFFFFED88 , 32'hFFFF90AC , 32'h000321F0 , 32'h00018A9C , 32'h0003B1B2 , 32'hFFF31239 , 32'hFFF8F724 , 32'hFFF962F3 , 32'hFFFD46CB , 32'h0000C2C7 , 32'h0000984A , 32'hFFFA6962 , 32'hFFFFEBF9 , 32'h000043A1 , 32'h00004096 , 32'h0007BE79 , 32'hFFFC95DA , 32'h000533D0 , 32'h000823C9 , 32'h000200DC , 32'h000259BC , 32'hFFFE66E7 , 32'hFFFB7448 , 32'h0003DEBD , 32'hFFFCEE37 , 32'h0005845C , 32'h0000C812 , 32'h000209FC , 32'hFFFE06F4 , 32'h000489D7 , 32'hFFFAECF8 , 32'h000376C7 , 32'hFFFE917C , 32'hFFFCB1E0 , 32'hFFFDDB13 , 32'h0001965F} , 
{32'hFFFA5F25 , 32'h00073CBF , 32'h0000839A , 32'hFFFCC17A , 32'h00032892 , 32'hFFFA75EF , 32'hFFF7AD66 , 32'h0004E48E , 32'h000865F2 , 32'hFFFE05AB , 32'hFFFD124B , 32'h0000F733 , 32'h0005E660 , 32'h00027B03 , 32'hFFFC65DD , 32'hFFFA949E , 32'hFFF858FD , 32'hFFF898E0 , 32'hFFFEE54D , 32'h00048B1F , 32'hFFFEE46C , 32'hFFF68E69 , 32'h0002BC01 , 32'hFFFAAD4C , 32'h0004F80B , 32'h00046103 , 32'h0000AE47 , 32'h000225DD , 32'h00059240 , 32'h000035A0 , 32'hFFFCFD6D , 32'h00014F38 , 32'hFFFC5112 , 32'h0004DD02 , 32'h00035EA0 , 32'h00034623 , 32'hFFFCB0AB} , 
{32'hFFFDDC66 , 32'h000ACA8C , 32'hFFFC01B2 , 32'h0002871D , 32'h0001F7E0 , 32'h000832C4 , 32'h00049988 , 32'h000105BF , 32'hFFF29ADF , 32'hFFFC66BE , 32'hFFFD980D , 32'h00017053 , 32'h00034F6E , 32'hFFF9283D , 32'h000EDA47 , 32'hFFFE79A8 , 32'hFFFE9484 , 32'hFFFB2D31 , 32'h00042F1D , 32'h0004469A , 32'h00033C7B , 32'h000119F1 , 32'hFFFEFEF3 , 32'hFFF6F233 , 32'hFFFCD2F5 , 32'h0001C474 , 32'h0003A518 , 32'h0005306A , 32'hFFFEB0A2 , 32'hFFFD30FC , 32'h000035EE , 32'hFFFC4153 , 32'h00060FAE , 32'hFFF5728E , 32'h000343DD , 32'h000711A1 , 32'hFFFCEE3B} , 
{32'hFFFF747D , 32'hFFF9407F , 32'h000325ED , 32'h0000FA15 , 32'hFFFD5AEC , 32'hFFFDA5FE , 32'h000142B9 , 32'h00026E9E , 32'h00018BEA , 32'h0007563C , 32'h0004B46B , 32'h0005D2E2 , 32'h0005A3E8 , 32'h00012E53 , 32'h00019207 , 32'h000C7098 , 32'hFFF9B86E , 32'h00015DF4 , 32'hFFFC6944 , 32'h00022BCB , 32'h00022245 , 32'h0000E18E , 32'h0008EECD , 32'h00005BFF , 32'hFFFEEFDB , 32'h0001DF0A , 32'hFFFBB062 , 32'hFFFD4273 , 32'hFFF7C684 , 32'hFFFABD5B , 32'hFFFF4DCC , 32'hFFFBE7EC , 32'h0006ABA5 , 32'hFFFE6A82 , 32'h000619E5 , 32'hFFFC7B53 , 32'hFFFFD14B} , 
{32'h0000B6FA , 32'hFFFEB38D , 32'hFFFFBA6C , 32'h00039A45 , 32'hFFFC77D7 , 32'hFFF40F2B , 32'hFFF8C9C5 , 32'h00043FC7 , 32'h0004B84F , 32'hFFF1E798 , 32'hFFFAE591 , 32'h000400AE , 32'hFFFE593A , 32'h00033A6E , 32'hFFFF8841 , 32'h00010E7C , 32'hFFF95B77 , 32'h00005275 , 32'hFFF73969 , 32'h0000C684 , 32'h00026229 , 32'h0008353C , 32'hFFF85F3D , 32'h0004D4A3 , 32'h0001B4EA , 32'h00050612 , 32'hFFFF6E47 , 32'h000BF647 , 32'hFFFCE762 , 32'h0002B6C9 , 32'h0002D288 , 32'hFFF54277 , 32'hFFFD3EDC , 32'hFFFA721A , 32'hFFF7D54D , 32'hFFF80C79 , 32'hFFFC35CF} , 
{32'h000B1EB3 , 32'hFFF9B1E2 , 32'hFFFA5F11 , 32'hFFFF91B3 , 32'h0001C3AB , 32'h0001BF32 , 32'hFFFF61DD , 32'hFFF97F44 , 32'hFFF7E853 , 32'h00059D05 , 32'hFFFECC19 , 32'hFFFF7BF6 , 32'hFFF715C5 , 32'h000559CE , 32'hFFF60BCA , 32'hFFF660BD , 32'h0000B44F , 32'h0001FE47 , 32'h00080E6E , 32'hFFF9DC01 , 32'h0003EFB9 , 32'h000214F8 , 32'h000228F7 , 32'hFFFF1B0A , 32'h0008254B , 32'h0006AA73 , 32'hFFFBF5A0 , 32'h000B48F3 , 32'h0004551F , 32'hFFFFA74C , 32'h00003B5D , 32'h0000C52B , 32'h00023EB7 , 32'hFFFB0DD1 , 32'hFFF7BC42 , 32'hFFFF4F68 , 32'h00033E6F} , 
{32'hFFFCD686 , 32'hFFFBD672 , 32'hFFFDB474 , 32'hFFF5CA7A , 32'h00016B89 , 32'h000010FE , 32'hFFFEE560 , 32'h000C4B2A , 32'hFFFF991A , 32'h00041746 , 32'hFFF9DAC0 , 32'hFFFD5568 , 32'hFFFA729D , 32'hFFFDF41C , 32'hFFF9EE41 , 32'h00021155 , 32'h00015A47 , 32'h000093F8 , 32'h0005EE7C , 32'hFFFE6AF7 , 32'h0001BCA4 , 32'hFFFF1652 , 32'hFFFF79AC , 32'hFFFF08D6 , 32'h0001FDEB , 32'h00085970 , 32'hFFFFF2B9 , 32'h000054FD , 32'h0004DA63 , 32'hFFFF3E73 , 32'h0003600A , 32'h0001270A , 32'hFFFBD4BF , 32'h00086829 , 32'h0004B6F9 , 32'hFFFEE1F2 , 32'h00005725} , 
{32'hFFFAE293 , 32'h0008B4CC , 32'hFFFA5746 , 32'h0000530A , 32'hFFF8C091 , 32'h000A2A3A , 32'hFFFF3BAF , 32'hFFF99914 , 32'hFFFDC7F0 , 32'hFFF75BA0 , 32'h0000FE95 , 32'hFFFA853B , 32'hFFFD475A , 32'hFFFD73F8 , 32'hFFFFBA19 , 32'h0004F113 , 32'h00031F72 , 32'h0009A28C , 32'hFFFE5758 , 32'hFFFCD9BB , 32'h00054B1F , 32'h0003C112 , 32'h0006C5DD , 32'h00002450 , 32'hFFFA11C7 , 32'hFFFDEAE3 , 32'h0009DE0C , 32'h00046DFE , 32'hFFF94268 , 32'h00088360 , 32'hFFFDE7F5 , 32'h0006D516 , 32'hFFF9759B , 32'h000014F6 , 32'hFFF7ECA4 , 32'hFFFBF108 , 32'h000199EF} , 
{32'hFFFDCF15 , 32'h0007F5B7 , 32'hFFF8F076 , 32'h0002351D , 32'h0002237F , 32'hFFFC7E23 , 32'hFFFFF7AF , 32'hFFFA9578 , 32'h0001710F , 32'hFFFD877A , 32'hFFFE0FA1 , 32'h00032848 , 32'hFFFE37DA , 32'h0002CCAE , 32'h0005B9F6 , 32'hFFF58EE3 , 32'h00016BEB , 32'hFFFE5E4D , 32'hFFFD4C6F , 32'h0003EE05 , 32'h00047B48 , 32'h00099150 , 32'h000058B4 , 32'h0001FE53 , 32'hFFFE2094 , 32'hFFFCF6E8 , 32'hFFFB05B8 , 32'hFFFA7C5D , 32'hFFF9B54C , 32'hFFFE3859 , 32'h0005F964 , 32'hFFFB3153 , 32'h00014871 , 32'h0001B384 , 32'h00013C3C , 32'h0001050A , 32'hFFF608D9} , 
{32'hFFFC63F8 , 32'hFFFF6323 , 32'hFFF8B840 , 32'h00027867 , 32'h0000D84C , 32'hFFF9E12F , 32'h000354EC , 32'hFFFD3E20 , 32'h0000B695 , 32'hFFFCEF77 , 32'hFFFD6509 , 32'hFFF9F754 , 32'h00045078 , 32'h000742F5 , 32'h00017F1A , 32'h00064838 , 32'hFFFFA7E9 , 32'h0007B17D , 32'hFFFE1B53 , 32'hFFF813C3 , 32'h00063448 , 32'h00079F2B , 32'h0001BAF7 , 32'hFFFC4C0A , 32'h0004E21A , 32'h00066041 , 32'hFFF98C18 , 32'hFFFB454B , 32'hFFF8B996 , 32'h0003671C , 32'h0001531A , 32'h00029CA3 , 32'h00065BAF , 32'h00028935 , 32'h0000B2D4 , 32'h00041AEB , 32'hFFF46A62} , 
{32'hFFF4813E , 32'h00040217 , 32'hFFFDB838 , 32'hFFF931BB , 32'h00040EF9 , 32'h0001B482 , 32'hFFFEE3A3 , 32'h0006D8B3 , 32'hFFFD3D15 , 32'hFFF74449 , 32'h0007AC6D , 32'hFFFB9D8F , 32'hFFF46169 , 32'hFFFABD6C , 32'h000C99D6 , 32'h0001D101 , 32'h0008B253 , 32'h0000CCED , 32'h0001D422 , 32'hFFF941EE , 32'h0005C605 , 32'hFFFBAE1A , 32'h0000EE9A , 32'h000072BC , 32'hFFFF679A , 32'hFFF6E412 , 32'hFFF98E85 , 32'h00025102 , 32'hFFFCA044 , 32'h00024AD4 , 32'hFFFF8344 , 32'h00045C1C , 32'h0003CE22 , 32'hFFFC4654 , 32'hFFFD2A51 , 32'h0001CF68 , 32'hFFF7DB8A} , 
{32'h0002E5AC , 32'hFFF61557 , 32'hFFFB154A , 32'hFFFF57CC , 32'hFFFDD10A , 32'h00020269 , 32'hFFFCD824 , 32'hFFFF44B4 , 32'hFFF9162F , 32'h00066142 , 32'h0008B6DF , 32'h00013977 , 32'hFFFCC9AC , 32'h000260DE , 32'hFFF50D4C , 32'hFFFE0474 , 32'h00022C1E , 32'hFFFC131F , 32'h000195E6 , 32'hFFF58F5E , 32'hFFF0A2A4 , 32'h000425CC , 32'hFFFEF6AF , 32'hFFFBC87C , 32'hFFFAA9E1 , 32'h00009855 , 32'hFFFAA7C9 , 32'h00051CAC , 32'h0004855D , 32'hFFFB4677 , 32'hFFFB15E3 , 32'hFFF34ED6 , 32'h0003E6D1 , 32'h0000F821 , 32'hFFFE5C2E , 32'h0001DCC1 , 32'h0007B09F} , 
{32'h0003AB51 , 32'hFFF3AAD5 , 32'hFFFDC42D , 32'h00038F6D , 32'h00050C8E , 32'h00056419 , 32'hFFFE5C19 , 32'hFFF69881 , 32'hFFFF2587 , 32'h000381A5 , 32'hFFFFFF9B , 32'h000702DB , 32'hFFFB1625 , 32'h0003147C , 32'h00091736 , 32'h00020038 , 32'h0002E17D , 32'h00005E21 , 32'h00024DD8 , 32'hFFFA0C73 , 32'h0006B1D5 , 32'hFFFE92DF , 32'hFFFE94DA , 32'hFFFD1461 , 32'hFFFF6850 , 32'hFFFD084F , 32'h0004433C , 32'h00045364 , 32'h0007FC27 , 32'hFFFEE233 , 32'h00031471 , 32'h0003FD21 , 32'hFFFD2DE4 , 32'hFFFA7176 , 32'h0001255D , 32'hFFFD9DE1 , 32'hFFFE69AF} , 
{32'hFFFDD734 , 32'h0000DE60 , 32'hFFFF43EF , 32'hFFFD9926 , 32'hFFFA69D2 , 32'h0004A7BC , 32'h0004819C , 32'hFFF669D6 , 32'h0003E62F , 32'h00034AC7 , 32'h0003B7B6 , 32'h0003A3C4 , 32'hFFFB0D61 , 32'hFFFF66F6 , 32'hFFFDAD7B , 32'h0006C898 , 32'hFFFDD93A , 32'h0001431E , 32'hFFFFAC05 , 32'h0002BA76 , 32'hFFFD2166 , 32'hFFFF835E , 32'hFFF1D41B , 32'h0002936C , 32'hFFFEE9A1 , 32'h00030208 , 32'hFFF4A50E , 32'h0009F8E0 , 32'hFFFD0078 , 32'h0003FE44 , 32'hFFFD08B2 , 32'hFFFF160A , 32'h00016E8A , 32'h0007843C , 32'hFFFF828C , 32'h000285BF , 32'h00001F24} , 
{32'hFFFC1753 , 32'hFFFC7297 , 32'hFFF870AD , 32'h00064A35 , 32'h000D1453 , 32'hFFF6FD0A , 32'hFFFD5AAE , 32'h0001F67E , 32'h000936C1 , 32'h0003FB15 , 32'h0004E81C , 32'hFFFE9939 , 32'h0002FB06 , 32'h0002537B , 32'h0000E8AC , 32'h0003CDED , 32'h0006C499 , 32'h00000023 , 32'hFFFC875A , 32'h0003B12D , 32'hFFF6E85C , 32'h00005C8E , 32'h0002C2DC , 32'h00035FCA , 32'hFFFE0448 , 32'hFFF7CB9F , 32'hFFFAB2A3 , 32'h00028B2D , 32'hFFF882C2 , 32'h0007B2CA , 32'hFFFAEFCD , 32'h0000B89D , 32'h000B7A7F , 32'h0006FAF2 , 32'h0001F06A , 32'hFFF90AA5 , 32'h0003B93A} , 
{32'h00004645 , 32'hFFFFE466 , 32'hFFFEC509 , 32'hFFFD59F1 , 32'hFFFF1DB6 , 32'hFFFD1817 , 32'h00050F28 , 32'h00052AFC , 32'hFFFAB42F , 32'h0002E077 , 32'h000073E7 , 32'hFFF2DAC0 , 32'hFFFFDA9F , 32'hFFFDC816 , 32'h000A4F6F , 32'hFFFE0182 , 32'h0000455C , 32'h00076E6C , 32'hFFFCA254 , 32'h00088F37 , 32'h00035C6B , 32'hFFFE67FA , 32'hFFFDE424 , 32'h0000E471 , 32'h0002FD91 , 32'hFFFC6BA9 , 32'h0001AA27 , 32'hFFFD97E9 , 32'h0001ACF8 , 32'h00027F03 , 32'h0006E783 , 32'h00090376 , 32'h00038957 , 32'h00070038 , 32'hFFFAB4C0 , 32'h0003C789 , 32'hFFFEB650} , 
{32'h000127C9 , 32'h00009239 , 32'hFFFB1C1F , 32'h00031DF0 , 32'hFFF4B355 , 32'hFFF8516A , 32'hFFFEF191 , 32'h0003A69D , 32'hFFFEB4FA , 32'hFFFBF74D , 32'h00008D17 , 32'hFFFDD2FD , 32'h00038DEC , 32'hFFFD7895 , 32'hFFFF9364 , 32'h00044A0F , 32'hFFFDA130 , 32'h0008EF52 , 32'h0003AAA3 , 32'h0002DAE2 , 32'hFFFFA7C2 , 32'hFFFBCE38 , 32'h00011211 , 32'h0005EBEE , 32'h000D5A5C , 32'h00032A5F , 32'h00044AA6 , 32'h0000B851 , 32'h0002CBB7 , 32'h00054389 , 32'h000182EB , 32'hFFFD9F84 , 32'h0000B708 , 32'h000148DB , 32'hFFFFD2D9 , 32'h0001BE4C , 32'hFFFF35D3} , 
{32'h0008E447 , 32'h0002193F , 32'hFFFC4BA6 , 32'h0000D3A0 , 32'hFFF9478B , 32'hFFFB88AE , 32'hFFFADE2D , 32'hFFF9EB12 , 32'hFFFFB053 , 32'h0003C5FB , 32'hFFFDB4B7 , 32'h0003EDAE , 32'hFFF81AD1 , 32'hFFF5A09B , 32'h000ECA26 , 32'h00022117 , 32'h00069AA2 , 32'h000B4FDE , 32'hFFF91000 , 32'h00042510 , 32'h00018A53 , 32'hFFFF19D4 , 32'h000283A3 , 32'hFFF8A780 , 32'h000E5745 , 32'hFFF4414A , 32'hFFFBF504 , 32'hFFFC173C , 32'hFFFF9818 , 32'hFFFBE902 , 32'hFFFD6339 , 32'h0006346F , 32'h00048FE0 , 32'hFFFBF537 , 32'h00012115 , 32'hFFFDB060 , 32'hFFFA267C} , 
{32'hFFFA3767 , 32'h00074E2C , 32'h000329F8 , 32'hFFFBCBBB , 32'h000225BD , 32'hFFF6BF30 , 32'hFFF94BDD , 32'h000624C1 , 32'hFFFE3B39 , 32'h0006D64A , 32'hFFF6561E , 32'hFFFDB1DA , 32'hFFFF7573 , 32'hFFFAEE6F , 32'h0000796C , 32'h0008A6AA , 32'hFFFDF00A , 32'hFFFC8D17 , 32'h000438EC , 32'hFFF30FF8 , 32'hFFFE2CAD , 32'h00090374 , 32'hFFF71B6C , 32'hFFFE5775 , 32'hFFFCF9C5 , 32'h0007454C , 32'h00000F87 , 32'h000708DE , 32'h0003B52C , 32'hFFFE57AC , 32'h00011ADF , 32'hFFFE4EBB , 32'hFFFFFDBA , 32'hFFFB7548 , 32'h0001DF1F , 32'hFFF60531 , 32'h00023E41} , 
{32'h0001A3E6 , 32'h0000425F , 32'hFFFE054E , 32'h00013A21 , 32'h00026C87 , 32'h0000F0BD , 32'hFFFF9005 , 32'hFFFBDF7F , 32'h00013EC1 , 32'h00024E45 , 32'hFFFB9D1C , 32'h0004DA1D , 32'hFFFAC55A , 32'h0002E946 , 32'hFFFFDD90 , 32'hFFFA7190 , 32'hFFFE418F , 32'h0006528D , 32'hFFFE5DD9 , 32'h0007001A , 32'h0004C565 , 32'hFFFFEE41 , 32'hFFF33B4D , 32'hFFFE67BF , 32'hFFFC40ED , 32'h00090187 , 32'hFFFA5202 , 32'h00017120 , 32'hFFF799E8 , 32'hFFF973C3 , 32'h00036CC9 , 32'h00031D74 , 32'hFFFEF7BD , 32'hFFFBA382 , 32'h0002AF88 , 32'h0000E35A , 32'h0001C655} , 
{32'h00019D5B , 32'hFFFF32D2 , 32'h00008E2B , 32'h0008EED1 , 32'h000487F5 , 32'hFFFD5C57 , 32'h00007D0A , 32'h0006626C , 32'hFFFBE170 , 32'h0003DF6D , 32'hFFFF39BE , 32'h00045E89 , 32'hFFFAA92E , 32'h00002591 , 32'h00089CA5 , 32'h00091035 , 32'hFFFC4BE2 , 32'hFFFEF6AA , 32'h000508DD , 32'hFFFB7B6F , 32'h0003493F , 32'hFFFE14EE , 32'h0002D48B , 32'h00046F57 , 32'h00032B6B , 32'h000296D8 , 32'h0000BA03 , 32'h000067B5 , 32'hFFF99B19 , 32'h00096CDE , 32'h00046298 , 32'h0001F97B , 32'hFFFB8E22 , 32'hFFFF5E54 , 32'h0000DCF6 , 32'h0006B169 , 32'h000B8AC2} , 
{32'hFFFF1D2E , 32'h000A0F1B , 32'h00026469 , 32'h00025F18 , 32'h0000A8C8 , 32'h000684CD , 32'h00015FBA , 32'hFFF8834A , 32'h000319F2 , 32'h0002CAE9 , 32'hFFF62B19 , 32'h0002A26E , 32'hFFFF4236 , 32'h000652C5 , 32'h00053B00 , 32'hFFF50E24 , 32'hFFFA0180 , 32'h00000390 , 32'h0005529A , 32'h00075A44 , 32'h0003EBFB , 32'hFFF9F0C0 , 32'h0004A93D , 32'hFFFCEFD7 , 32'h00095B7E , 32'h000044D0 , 32'hFFFC2C1A , 32'h000364A2 , 32'hFFFF0533 , 32'h00005D4B , 32'h00003B54 , 32'h00060DEB , 32'hFFFF856E , 32'hFFFAEB79 , 32'hFFFE7AD9 , 32'h0001E4E7 , 32'h0002C4B6} , 
{32'hFFFC0C82 , 32'h0001BB1C , 32'hFFFF5887 , 32'h0006D5EA , 32'hFFFF8D3A , 32'hFFF4CD43 , 32'h0001F556 , 32'h0006F424 , 32'hFFFE8E1D , 32'hFFFFCE93 , 32'hFFF92DDF , 32'hFFF891A5 , 32'h00043E70 , 32'h00053C88 , 32'hFFFDAC8B , 32'hFFFE1D60 , 32'h0003F0B9 , 32'h00016267 , 32'h000003EA , 32'hFFFEF67A , 32'h00040E24 , 32'hFFFD770D , 32'hFFFD840E , 32'h0000CE99 , 32'hFFFB6493 , 32'hFFFC7344 , 32'h00010F20 , 32'h000232E5 , 32'hFFFB563A , 32'h00012DAA , 32'h0009E7CF , 32'hFFFF40A6 , 32'h00060908 , 32'h0006B66B , 32'h00071D38 , 32'hFFFC8CC3 , 32'hFFFF1C69} , 
{32'hFFF95731 , 32'h0005C4F9 , 32'hFFFBFB3D , 32'h0006E43A , 32'h0004006D , 32'h00064731 , 32'hFFFC9C49 , 32'h00028A06 , 32'h00031500 , 32'h000171CF , 32'h00068744 , 32'hFFFCBB2B , 32'hFFFB7A91 , 32'h0002D2E8 , 32'h00000005 , 32'h00043F2E , 32'hFFFF5AC6 , 32'hFFFED904 , 32'hFFFF8095 , 32'hFFFFC2A2 , 32'hFFFB8453 , 32'hFFFBF76D , 32'hFFFAF4C1 , 32'hFFFE2E2E , 32'h0002D3F0 , 32'h0003227A , 32'hFFFE4F80 , 32'hFFFE9ED2 , 32'h0002F024 , 32'hFFFD28A7 , 32'h0006CF70 , 32'hFFF7566E , 32'h00013C7D , 32'h000E7874 , 32'hFFFE2074 , 32'h0000621D , 32'hFFFE66F1} , 
{32'hFFFDA5B6 , 32'h0002F356 , 32'h000734B4 , 32'h0006CDB6 , 32'h000241EB , 32'h0000641A , 32'hFFF4DF91 , 32'h00039278 , 32'hFFFF3A6F , 32'h0004FB82 , 32'hFFF7B486 , 32'hFFFF3C5A , 32'hFFFEC9F8 , 32'h00027334 , 32'hFFFD3DCB , 32'h0005E976 , 32'h00041D0F , 32'hFFFD6B09 , 32'hFFFAD0C3 , 32'h0000931F , 32'hFFFA74EF , 32'hFFFBB1F2 , 32'hFFFC3220 , 32'h00042200 , 32'hFFF94F9F , 32'h00030534 , 32'hFFF9B7C0 , 32'hFFFFB02B , 32'hFFF9E5D7 , 32'h000784E7 , 32'h0007B520 , 32'h00060D63 , 32'hFFFEE913 , 32'hFFFD60F3 , 32'hFFF719C6 , 32'h00011457 , 32'h0003D40A} , 
{32'h00029C21 , 32'hFFFE39C4 , 32'h000835EB , 32'h0005C251 , 32'h0001B1F0 , 32'hFFFBD64F , 32'h0003B3CE , 32'h0001A06C , 32'hFFFC99EB , 32'h0009B62F , 32'hFFFEF180 , 32'hFFFD73E6 , 32'h0001C83F , 32'h0004AEA2 , 32'hFFFC2285 , 32'h00005B6B , 32'h0000E50B , 32'h0001619F , 32'hFFF72026 , 32'hFFFBC56A , 32'hFFFE1EE5 , 32'hFFFBAAFE , 32'h00073F6D , 32'h0003C4BD , 32'hFFFE607E , 32'hFFFBF8C0 , 32'hFFFBB18E , 32'h0000C7A2 , 32'hFFF92C35 , 32'hFFFBF384 , 32'h00076344 , 32'h000659D4 , 32'hFFFFC57B , 32'hFFFB1105 , 32'h00066796 , 32'hFFF601CF , 32'h0003032F} , 
{32'hFFFA868E , 32'hFFFE037C , 32'h0006EC18 , 32'h0003B86C , 32'hFFFCDAAB , 32'hFFF92616 , 32'hFFFC5C86 , 32'hFFFFF2F8 , 32'h00054C3B , 32'hFFFDADE7 , 32'hFFFEAF6E , 32'hFFFD469E , 32'h0005FDA6 , 32'h0001D4C6 , 32'hFFFA3B65 , 32'hFFFC535E , 32'h0007FB5C , 32'hFFFDD88F , 32'hFFFD1E54 , 32'hFFFAED0F , 32'hFFFAB810 , 32'h0004BDDC , 32'h0002DAE3 , 32'hFFFBE693 , 32'h00057DBD , 32'hFFFE9509 , 32'h00022C71 , 32'h00091EC8 , 32'hFFF660F9 , 32'h0001D8EB , 32'hFFFF02FF , 32'hFFF7E388 , 32'hFFFC8E22 , 32'hFFF74E45 , 32'hFFFBC6CB , 32'hFFFBB6DE , 32'hFFF4599C} , 
{32'hFFF2DDC6 , 32'hFFFDEBA5 , 32'hFFFEE89D , 32'h00047934 , 32'hFFFAC46A , 32'hFFF35F61 , 32'h00007911 , 32'h00000C9B , 32'h0006B322 , 32'h0007FB5F , 32'hFFFB00F7 , 32'h000125D6 , 32'hFFFF18A0 , 32'h00083986 , 32'h000D6B86 , 32'h00077051 , 32'hFFFDF856 , 32'hFFFC2E2B , 32'hFFFD9510 , 32'hFFFC18DB , 32'h000608F8 , 32'h00036D4C , 32'hFFFE53E3 , 32'hFFFCCED5 , 32'hFFFCEFF1 , 32'hFFFD5B88 , 32'h00060715 , 32'hFFF5072A , 32'h00074CAC , 32'hFFFEEC26 , 32'hFFFA39D2 , 32'h000B6A38 , 32'h000078F0 , 32'h0002AE7F , 32'hFFFDBEAD , 32'hFFFFC2C7 , 32'hFFFB37AA} , 
{32'h0005CE82 , 32'h00026E81 , 32'h000113C8 , 32'hFFFCA232 , 32'h0006C2A9 , 32'hFFFF715A , 32'hFFF6F112 , 32'h000912F3 , 32'h000211B2 , 32'h0001C76A , 32'hFFFFFA04 , 32'hFFFFE339 , 32'h0003A6D5 , 32'hFFFF8293 , 32'hFFFFA967 , 32'h00046414 , 32'h00020E46 , 32'hFFFDA6AC , 32'hFFFE7C1C , 32'h000294FA , 32'h0000EC6F , 32'hFFFE8ACA , 32'hFFF3999B , 32'h00013C37 , 32'hFFF9D96C , 32'h0000733E , 32'h0001ED46 , 32'h00050828 , 32'h00028B23 , 32'h0002F32C , 32'h000060ED , 32'h00060657 , 32'hFFF388FE , 32'h0004ABA9 , 32'hFFFE2AB0 , 32'h00012C7A , 32'h0003B9D7} , 
{32'hFFF8B8F5 , 32'h00037FCF , 32'hFFFE3A52 , 32'h00002880 , 32'h00026DFC , 32'hFFF74DB9 , 32'h000BEDAE , 32'h000287C7 , 32'h000C164E , 32'hFFFFB239 , 32'h00060AB7 , 32'h0001138D , 32'hFFFAB011 , 32'h00006C55 , 32'hFFFAA7E7 , 32'hFFFA3B6E , 32'h000370B5 , 32'h0001DF37 , 32'hFFFCED79 , 32'hFFFDCF8B , 32'h0004BF50 , 32'h000598D3 , 32'h0000362B , 32'h0002C626 , 32'hFFF9C30E , 32'hFFFB6892 , 32'h000117EE , 32'hFFFD4F5D , 32'h00015F7F , 32'h0001639F , 32'hFFFE62B1 , 32'h0002DE5C , 32'h0004BFCA , 32'h000234FD , 32'hFFFA2CD0 , 32'h0002175E , 32'hFFFACB2E} , 
{32'h00035D2B , 32'h0001B1D7 , 32'hFFFF2371 , 32'hFFF3ED8F , 32'hFFFE7515 , 32'h00019602 , 32'hFFFCC6B6 , 32'hFFFB759C , 32'hFFFBC50E , 32'h0000B783 , 32'h00078F0C , 32'hFFFDCDB3 , 32'h000D04EE , 32'hFFFE93CB , 32'h00055B3D , 32'hFFFFE6CD , 32'hFFF6B80A , 32'h00049EF7 , 32'h00027B6E , 32'h00017AAF , 32'hFFFA91E7 , 32'h0005A08B , 32'h0000F85B , 32'hFFFDE7DF , 32'h00084618 , 32'h0008025F , 32'hFFF982EF , 32'hFFFC683F , 32'hFFFFEECA , 32'hFFFEEB3C , 32'h00014323 , 32'h00039BC4 , 32'hFFFA6032 , 32'h00063018 , 32'h00068B85 , 32'hFFFBC608 , 32'hFFF4DE19} , 
{32'h0009EF1B , 32'h0004F062 , 32'h00027F6A , 32'h001185F4 , 32'hFFF82739 , 32'h00055CD0 , 32'hFFFFA40E , 32'h00032533 , 32'h000479C0 , 32'hFFFDBBCD , 32'h000DBAC5 , 32'h000BCF01 , 32'h00034157 , 32'h000AF32F , 32'hFFFEBB79 , 32'hFFF6A7A7 , 32'hFFFBF3B7 , 32'h00053E0B , 32'hFFF95C10 , 32'h000635A2 , 32'hFFF902A5 , 32'hFFFE1F76 , 32'hFFFC7D79 , 32'hFFFEC991 , 32'hFFF54F8E , 32'h00011B9D , 32'h0006DDD8 , 32'h00014072 , 32'hFFF9CCE2 , 32'hFFFCA68B , 32'hFFFC42EC , 32'hFFFA89A2 , 32'h00014D66 , 32'h00075E44 , 32'h000125FD , 32'hFFFB51E3 , 32'h00044A4F} , 
{32'hFFFAE082 , 32'h00007C74 , 32'h000225A0 , 32'h00075EDE , 32'hFFFD7284 , 32'h0007E06A , 32'hFFFFDA66 , 32'h0002AA61 , 32'h00049631 , 32'h00017730 , 32'h000AB8C4 , 32'h000153EA , 32'h0000A3FD , 32'hFFFF13E2 , 32'hFFFD1A68 , 32'hFFF9E4C6 , 32'h0004A443 , 32'hFFFEB76A , 32'hFFFB40C6 , 32'hFFF8055E , 32'hFFFCF569 , 32'hFFFCBCB2 , 32'hFFFDCE5F , 32'hFFFA833F , 32'h00027D16 , 32'h000025AC , 32'h0001EF85 , 32'hFFFF295B , 32'h0000BC86 , 32'hFFFB2B5E , 32'h000B43DF , 32'hFFF901BF , 32'hFFF4413B , 32'h00004FCA , 32'hFFFCD646 , 32'h000162E2 , 32'h00023C50} , 
{32'hFFFFC5FA , 32'h0002DCA4 , 32'h00009A4E , 32'hFFFEFE30 , 32'hFFFD53E0 , 32'hFFFE2E19 , 32'hFFFF9CB2 , 32'hFFFA68DC , 32'hFFF718BB , 32'hFFFFA0F1 , 32'h0000F79C , 32'hFFFE1C40 , 32'hFFF88FF4 , 32'hFFFBEE9D , 32'h00057576 , 32'hFFF536AC , 32'hFFFD2B24 , 32'hFFFEA7EE , 32'h0001FB4B , 32'hFFFA4286 , 32'hFFF602FF , 32'hFFF8A8A2 , 32'h000445E0 , 32'hFFF57545 , 32'hFFFC89F2 , 32'h000A9574 , 32'h00066B49 , 32'hFFFC80E6 , 32'hFFFEBE30 , 32'hFFF9FE84 , 32'hFFFB9BFB , 32'hFFFE44BF , 32'h00033B2B , 32'h00071E46 , 32'hFFFED1F4 , 32'h00024E3F , 32'hFFFD6E81} , 
{32'h0009730F , 32'hFFF6B190 , 32'hFFFABA6C , 32'hFFF9229E , 32'h00063114 , 32'h00017EAD , 32'hFFFD9E09 , 32'hFFFA2579 , 32'hFFFE61D4 , 32'h0003E303 , 32'h000009B7 , 32'hFFFFF1A0 , 32'hFFFDD91A , 32'h000261EB , 32'h0001653F , 32'hFFFA0E75 , 32'h000260C7 , 32'hFFFDD33D , 32'h0006086D , 32'h00053400 , 32'hFFFB243B , 32'hFFF60EDA , 32'hFFFF39E0 , 32'hFFFAEB59 , 32'h00003A3B , 32'h00000F47 , 32'hFFFFDCFF , 32'h00014103 , 32'hFFF4B8F4 , 32'h0003C028 , 32'h000A61B8 , 32'h00034D19 , 32'hFFFF6D8C , 32'hFFFFCFE6 , 32'hFFFFDD01 , 32'h00047140 , 32'hFFFA26E6} , 
{32'hFFFAD697 , 32'hFFFFC3CB , 32'hFFFAE58C , 32'h00062B88 , 32'hFFF829B7 , 32'hFFFCE18C , 32'hFFF8D927 , 32'hFFFC2916 , 32'hFFF47570 , 32'h0000B03D , 32'h0003912B , 32'hFFFCF58E , 32'h001132CE , 32'hFFF71160 , 32'hFFFB52A7 , 32'hFFFCE69E , 32'hFFFCB1E8 , 32'hFFFD4615 , 32'h0000E76D , 32'h00071A93 , 32'hFFFDFD5C , 32'h0008F9DC , 32'h0002919E , 32'hFFFCF0F2 , 32'h000AFF23 , 32'hFFFE06E7 , 32'hFFFEAFD7 , 32'hFFFB3D6C , 32'h0003DF5D , 32'h0005DDA3 , 32'hFFFD5E8C , 32'hFFF99E29 , 32'hFFFF0B28 , 32'h00105D01 , 32'hFFFA48D0 , 32'h00009AF1 , 32'h000041BD} , 
{32'h00056E90 , 32'hFFFB76F6 , 32'hFFF777E8 , 32'hFFFF47CF , 32'h000633F0 , 32'hFFFE25C7 , 32'hFFF55189 , 32'h000088B5 , 32'hFFFB00D8 , 32'h00032044 , 32'hFFFCE69A , 32'hFFFC8A00 , 32'h00050301 , 32'h000082CB , 32'hFFFE94EB , 32'h00079317 , 32'hFFFB0CA4 , 32'hFFFBFCEF , 32'h0000A714 , 32'hFFFEBF04 , 32'h0009F0E5 , 32'hFFFAE7AF , 32'hFFFF01E6 , 32'hFFFBF23A , 32'hFFFD5D2D , 32'h00002D90 , 32'h000A3CFA , 32'h00028F4D , 32'h0000DE83 , 32'hFFF89909 , 32'h0004204A , 32'h0002AED3 , 32'hFFFF1841 , 32'hFFF7DCED , 32'h0002ADB1 , 32'h00068283 , 32'h00015DBB} , 
{32'h00015163 , 32'h0003683A , 32'h00022A98 , 32'hFFFF5852 , 32'h0001E150 , 32'h000509F5 , 32'h00043600 , 32'hFFFE246C , 32'hFFFC81DC , 32'hFFFBD479 , 32'h000104D8 , 32'h000301E7 , 32'h000348A5 , 32'hFFFCFDB4 , 32'h0004371B , 32'h00016AFA , 32'hFFFD2DEF , 32'hFFF9CF01 , 32'hFFF5FA4C , 32'h0001B725 , 32'hFFFFA0FE , 32'hFFFDC904 , 32'hFFFD7C8B , 32'hFFFE4136 , 32'h0002BA7B , 32'h000160C9 , 32'hFFFED27F , 32'hFFFB3D21 , 32'hFFFDBC99 , 32'hFFFF7334 , 32'hFFFA6BC6 , 32'h00053CA3 , 32'h000522C5 , 32'hFFFE2B6B , 32'hFFFBCA7E , 32'h000488AD , 32'hFFFCB154} , 
{32'h0006E321 , 32'hFFFC05ED , 32'h000123FC , 32'hFFF6775C , 32'hFFFDC000 , 32'h000A320B , 32'h00099457 , 32'h000497BC , 32'h0001BE04 , 32'hFFFBF285 , 32'h0005E0E6 , 32'hFFFC422E , 32'hFFF3F06B , 32'h00017695 , 32'hFFF8336A , 32'hFFF864E8 , 32'h0006DF05 , 32'h000153A7 , 32'h00023730 , 32'hFFFDCE86 , 32'h0001FC51 , 32'h00024C44 , 32'hFFFA2031 , 32'h00029263 , 32'hFFFA7722 , 32'hFFFC43FB , 32'h00096193 , 32'hFFFE4027 , 32'h0000F258 , 32'h0005A4D4 , 32'h0000D60D , 32'h0001C3E9 , 32'h0000454F , 32'h00065B53 , 32'hFFFEFAB6 , 32'hFFFDD5D6 , 32'hFFFD6C0C} , 
{32'hFFF91BF2 , 32'h0005919A , 32'h0006A0D8 , 32'hFFF4936D , 32'hFFFD0231 , 32'h0006DBF5 , 32'hFFFAAF4B , 32'hFFFB0189 , 32'hFFFD8B81 , 32'hFFF5A875 , 32'hFFFC2676 , 32'hFFFB14BC , 32'h0001871D , 32'hFFFE3AA1 , 32'h000072F0 , 32'h000288E1 , 32'h000123CE , 32'hFFFAC725 , 32'hFFFF36A6 , 32'h00028444 , 32'h00069A58 , 32'hFFF8B30C , 32'hFFFBF6D7 , 32'hFFFF9B1A , 32'h0001E9FD , 32'hFFFF950E , 32'h0003475B , 32'hFFF591EE , 32'hFFFF810F , 32'h0007A5B3 , 32'hFFF9515B , 32'h0003EE2F , 32'h00034418 , 32'h00000086 , 32'hFFFBDBDB , 32'h00020776 , 32'h00033D90} , 
{32'hFFFEEF04 , 32'hFFFC81A2 , 32'h0001C452 , 32'h0003BAD8 , 32'hFFFE5B35 , 32'hFFFFA789 , 32'hFFFB126E , 32'h0001D65F , 32'h00017861 , 32'h00045FA3 , 32'h00047737 , 32'hFFFEC790 , 32'h00019A07 , 32'h000165BE , 32'hFFF83425 , 32'hFFFF36F9 , 32'h00001C2D , 32'h000DD8DD , 32'h00027BD3 , 32'h000C932B , 32'hFFF912C3 , 32'h00027799 , 32'hFFFECE97 , 32'h0005A699 , 32'h0002ED68 , 32'h0000B3F3 , 32'h0000170A , 32'hFFFF989A , 32'hFFFA851D , 32'h00009005 , 32'hFFF978C9 , 32'hFFFE215D , 32'h000AC865 , 32'hFFFCBA79 , 32'hFFFE1D97 , 32'hFFF0C83B , 32'hFFF537E5} , 
{32'h00020DE9 , 32'h000C7D21 , 32'hFFFEA25F , 32'hFFFC3F37 , 32'hFFFD7444 , 32'hFFFC3E0B , 32'hFFFDFC96 , 32'hFFFE1A7A , 32'h00029775 , 32'hFFFA8B90 , 32'hFFF9A714 , 32'h00070FAA , 32'hFFFDD684 , 32'hFFF9155A , 32'h00012D42 , 32'h0002824C , 32'h00005374 , 32'hFFFD5C51 , 32'hFFFED401 , 32'h00047CEB , 32'h000468DD , 32'h00004604 , 32'h0005558A , 32'hFFFBCE73 , 32'hFFFBBE12 , 32'h0003356E , 32'hFFFE1403 , 32'h000011F1 , 32'hFFFF1EB1 , 32'hFFFBD28E , 32'hFFFEA6B5 , 32'h0004F26A , 32'hFFFD902A , 32'h00064718 , 32'hFFFA1142 , 32'hFFFC306F , 32'h000233DF} , 
{32'h000290EA , 32'h0000184F , 32'h00019248 , 32'h000102D7 , 32'h0005D62A , 32'h00005D43 , 32'hFFF9EDF2 , 32'h00027721 , 32'h00034BFF , 32'hFFFF5CB5 , 32'hFFFA7E68 , 32'h0006B8CF , 32'h000304BB , 32'h0005F295 , 32'hFFFE1C52 , 32'h00006061 , 32'hFFFE21F7 , 32'h0003B358 , 32'hFFF87F11 , 32'hFFFE1AA7 , 32'h0000F60A , 32'hFFFE64C9 , 32'h0000D69E , 32'h00053D7A , 32'h0001EC5F , 32'hFFFD17AA , 32'h000076A4 , 32'h00094F4D , 32'hFFFF5586 , 32'h000362BD , 32'h0002EDF9 , 32'h0005E611 , 32'hFFFCA3A1 , 32'h00031AA1 , 32'hFFF93DAC , 32'h000095AC , 32'hFFF9A2A6} , 
{32'hFFFA9867 , 32'hFFFB5EFE , 32'hFFFD3A4B , 32'hFFFED453 , 32'hFFFF9569 , 32'h00017A60 , 32'h00054284 , 32'h00007FF9 , 32'hFFFBCA15 , 32'h0002809C , 32'h0001C84B , 32'hFFFA26D6 , 32'hFFFC415F , 32'hFFFD4F63 , 32'hFFFD9E15 , 32'h000AF4EE , 32'h00002F2F , 32'hFFFE5417 , 32'h000BDD74 , 32'h000068A4 , 32'hFFF30CBA , 32'h000CBF76 , 32'h000ABFD6 , 32'hFFF6913D , 32'hFFFB2D25 , 32'hFFFE9DD7 , 32'h0001CEE0 , 32'hFFFFB242 , 32'hFFF91283 , 32'h0002CA12 , 32'hFFFAE6B7 , 32'hFFFF0188 , 32'h000B091F , 32'h0001EFE6 , 32'hFFFE39E1 , 32'h00017D5B , 32'hFFFC2762} , 
{32'hFFF733BA , 32'h00088E3D , 32'hFFFA35C8 , 32'h000173FC , 32'h000165AA , 32'hFFFCB8CE , 32'h00011F4C , 32'h0007F6DC , 32'hFFFADDE2 , 32'h0004BB5B , 32'hFFFF5675 , 32'h0000F40C , 32'h0004B6A5 , 32'h000A8B52 , 32'h000304BA , 32'h00006062 , 32'h00031815 , 32'hFFF81D20 , 32'h0007ACB2 , 32'h00016E31 , 32'hFFFCC989 , 32'h000453A5 , 32'h00069724 , 32'hFFFF4BAF , 32'hFFF9930B , 32'hFFF67DDB , 32'h0004E44C , 32'h00087C65 , 32'hFFFF36B1 , 32'h00040DCE , 32'h00065F83 , 32'h000476FB , 32'hFFFE48F5 , 32'h0007FAB3 , 32'h00011CA4 , 32'hFFFFE070 , 32'h0001A4AA} , 
{32'h00030A65 , 32'h00027D4E , 32'hFFFEDA26 , 32'hFFFA9454 , 32'h0005BD0B , 32'hFFFC9BA9 , 32'h00004AB2 , 32'hFFFE5784 , 32'hFFFECCB7 , 32'hFFF77054 , 32'hFFFFF78E , 32'h00014165 , 32'hFFFF055A , 32'hFFFD7353 , 32'h0000C8FA , 32'h0004DEE7 , 32'hFFFDC268 , 32'hFFF8795F , 32'h0007D9AA , 32'h00033C86 , 32'h00068AC8 , 32'h0001C84D , 32'h00059299 , 32'hFFFEEB50 , 32'hFFF9C2F4 , 32'h00037AF1 , 32'hFFFE3A11 , 32'h0007148D , 32'hFFFE1541 , 32'hFFFE7A1F , 32'hFFFB1056 , 32'hFFF5059D , 32'h00002CBE , 32'h00042034 , 32'hFFFAC39E , 32'h00070960 , 32'hFFFC9A66} , 
{32'hFFFDDCB6 , 32'hFFFDEA42 , 32'h00054D1F , 32'h00088ABB , 32'h000B015A , 32'h0003D3F4 , 32'h00067D13 , 32'h0006717C , 32'h00002822 , 32'h0001F7A2 , 32'h000895D9 , 32'hFFFC3C36 , 32'h00032F8B , 32'hFFF4E71D , 32'hFFFDD9A0 , 32'h00010358 , 32'h00001503 , 32'h00052DE9 , 32'h0001E3FA , 32'hFFF80811 , 32'h000152A8 , 32'hFFFFCDAF , 32'h00095805 , 32'h0000D4AC , 32'h00016BA9 , 32'h0000B4A6 , 32'h00029AE1 , 32'hFFFED31C , 32'h000259F5 , 32'h0003F9D3 , 32'hFFF7804A , 32'h000452D0 , 32'h0003C61E , 32'h00028D9C , 32'h0000FB45 , 32'h00044B2D , 32'hFFFABEF2} , 
{32'h000021E6 , 32'hFFFC3883 , 32'hFFFE3C77 , 32'hFFFE6F18 , 32'hFFFAFFD4 , 32'h0003C1AE , 32'h0004FB87 , 32'hFFFD043B , 32'hFFFC7796 , 32'hFFFFC1B9 , 32'hFFFC0455 , 32'h000012E8 , 32'hFFF64B9F , 32'hFFFAC0A3 , 32'h000254DB , 32'hFFF16FC1 , 32'h0006645B , 32'h00017582 , 32'hFFF7D7C7 , 32'hFFF78AD5 , 32'h0001D532 , 32'h00025B15 , 32'hFFFB2A09 , 32'hFFFF37AF , 32'hFFFF7C55 , 32'hFFFEF4DA , 32'h0004FDDB , 32'h0001E61E , 32'h0007291C , 32'h00066C2F , 32'hFFFADF8D , 32'h00007943 , 32'hFFFF9DA5 , 32'hFFFB6F29 , 32'hFFFEAB9F , 32'hFFFA32F5 , 32'h00015C36} , 
{32'hFFFF110F , 32'hFFFB4270 , 32'hFFFE0279 , 32'hFFFF9AB4 , 32'hFFFE161F , 32'h0002E2DF , 32'h00010626 , 32'h0001660F , 32'h000AEAAA , 32'hFFFCE432 , 32'h0008EA1D , 32'hFFFA8FF6 , 32'h0005426E , 32'hFFF40883 , 32'hFFF7072D , 32'h0007BEE6 , 32'hFFFA80AF , 32'hFFFDB4EF , 32'hFFFE5885 , 32'hFFFFE7E0 , 32'hFFFB3171 , 32'h0006E46C , 32'hFFFC4726 , 32'hFFFD7B7B , 32'h0001D11A , 32'h0002372B , 32'h00021E10 , 32'h0005E928 , 32'h00020C91 , 32'h0000B482 , 32'hFFFC12C8 , 32'hFFF8BB67 , 32'h00024805 , 32'h000B43F1 , 32'h0000E8E0 , 32'hFFFE0D9E , 32'h0005F742} , 
{32'hFFFFFDA9 , 32'h000413B1 , 32'h00042366 , 32'hFFFDEA7E , 32'h000347ED , 32'hFFFD92E8 , 32'hFFFEA165 , 32'h00065ADD , 32'h0003EADF , 32'h0001E808 , 32'hFFFE42F5 , 32'h00029352 , 32'h0000804A , 32'h0002768F , 32'hFFFF19E3 , 32'h00058D0B , 32'h0002350C , 32'hFFFFB728 , 32'h000281D3 , 32'h0001A638 , 32'h00071A74 , 32'hFFFD0102 , 32'h0002CFD3 , 32'hFFFFD0E6 , 32'h00050FD7 , 32'h0003C10D , 32'hFFFB2540 , 32'h0000349D , 32'h000243E1 , 32'hFFFDD8E0 , 32'h00001152 , 32'hFFFF9FB4 , 32'hFFFB4932 , 32'h00049899 , 32'hFFF818F4 , 32'h00007B48 , 32'hFFFA1F82} , 
{32'h0005563A , 32'h00014195 , 32'h0000CC53 , 32'hFFFF64EC , 32'hFFF51603 , 32'hFFFD9F13 , 32'hFFFE04C7 , 32'h00001742 , 32'h00066DD2 , 32'h0006D227 , 32'hFFFFBCE0 , 32'h0002025F , 32'hFFFAE1E3 , 32'h00013389 , 32'hFFFF3C1A , 32'h00054067 , 32'h00017204 , 32'hFFFA365D , 32'h00072E05 , 32'h00016B91 , 32'hFFFBC0B7 , 32'hFFFCA428 , 32'h0001FB42 , 32'h00093F2D , 32'h000415BC , 32'h000595B4 , 32'h000389DC , 32'hFFFEDD1A , 32'h00012DC6 , 32'hFFFEA050 , 32'h000226AE , 32'h0000A77E , 32'hFFFC7C9F , 32'h0004D523 , 32'h000444A5 , 32'h0000019B , 32'h0004CAFD} , 
{32'hFFFC4238 , 32'h0002C76F , 32'hFFFB8A07 , 32'hFFFD0B4F , 32'h0002DCFE , 32'hFFFD2912 , 32'h00020C23 , 32'h0001339D , 32'hFFFE9282 , 32'h00005E5C , 32'h0002079C , 32'h00026DBF , 32'h00066F66 , 32'h0004B947 , 32'h00002C0A , 32'h00073A17 , 32'hFFFFBE0A , 32'h0002AA01 , 32'hFFF94E5A , 32'h000294BE , 32'h0002791F , 32'hFFFF1091 , 32'hFFFB4346 , 32'h0000D5EE , 32'h00004CEA , 32'h0000A333 , 32'h00060A83 , 32'h0000FF45 , 32'hFFFE44E8 , 32'hFFFE75ED , 32'h00078177 , 32'h00065F3F , 32'h00004D9B , 32'hFFFB7345 , 32'hFFFCF3AA , 32'h0003DB15 , 32'hFFFBA9CE} , 
{32'hFD58A920 , 32'hFFE7A65F , 32'hFE387634 , 32'h05BA6E48 , 32'h00642313 , 32'h0066ECAE , 32'hFF2A288D , 32'h06077310 , 32'hFE96DE50 , 32'h002AB3AE , 32'h0094D2E9 , 32'h02996994 , 32'h01A3FB28 , 32'hFFF64098 , 32'hFE99402C , 32'hFF6ECFB7 , 32'h00D2CFAA , 32'h01710410 , 32'hFBED8B10 , 32'h0118A210 , 32'hFF1D6511 , 32'h0214C6B0 , 32'hFCD858A4 , 32'h004C7E7C , 32'h00AF24B5 , 32'hFE7DF85C , 32'hFE1A16AC , 32'h00AA5090 , 32'h0008696A , 32'hFF46537C , 32'hFECEDD98 , 32'h0121D3AC , 32'hFE060974 , 32'hFC9C3C6C , 32'h03AD8588 , 32'hFB70EC18 , 32'hFDF8BD44} , 
{32'hFFFBB7D2 , 32'h0005E316 , 32'hFFFE9D1D , 32'hFFFEB186 , 32'h00016F5D , 32'h0005A5D5 , 32'h0001B031 , 32'hFFFE72A5 , 32'hFFFEFDE2 , 32'hFFFBB00D , 32'hFFF7C93E , 32'hFFFEEE1A , 32'h000066ED , 32'hFFFF2A1B , 32'hFFFDBF42 , 32'hFFFFB381 , 32'hFFFF0158 , 32'hFFFC55B1 , 32'h000400A9 , 32'hFFFB3448 , 32'h00034F50 , 32'h0001FD2F , 32'h00001E2F , 32'h0001ECBC , 32'h000098B8 , 32'h00036FBA , 32'hFFFFC352 , 32'hFFF988BA , 32'h00040EDC , 32'hFFFBEBF8 , 32'h00019D31 , 32'h0006D32D , 32'hFFFC581C , 32'hFFFB0354 , 32'hFFFDFD38 , 32'h00048238 , 32'hFFFF6337} , 
{32'hFFFFD83B , 32'hFFF7247F , 32'h00023393 , 32'h00005451 , 32'h00079A74 , 32'h0003D2B8 , 32'h000764D0 , 32'hFFFE95B8 , 32'hFFFAAB90 , 32'hFFFF84E6 , 32'hFFFEB711 , 32'h00045836 , 32'h00061E71 , 32'h000117AD , 32'h0002A8E2 , 32'h00018EA9 , 32'hFFFE5A07 , 32'hFFFF031E , 32'hFFFE821A , 32'hFFFF1683 , 32'h00036ADF , 32'hFFFE54FD , 32'hFFFB6D9F , 32'hFFFB1442 , 32'h00036B47 , 32'h00033A13 , 32'h0004F470 , 32'h00076E07 , 32'hFFFEE174 , 32'hFFFF5510 , 32'hFFF93738 , 32'h0002CE3F , 32'hFFFBBEC0 , 32'hFFF8EEC8 , 32'hFFFC1C0B , 32'h000B5DC7 , 32'hFFFD79D1} , 
{32'hFFFFE41A , 32'h00020F67 , 32'h0000E542 , 32'h000145A1 , 32'h00026CDE , 32'hFFFE98BF , 32'h00007774 , 32'h0000A33A , 32'hFFFE3EB7 , 32'hFFFDBFD7 , 32'hFFFE979C , 32'hFFFD9B84 , 32'hFFFED03A , 32'hFFFC59A6 , 32'h0003274F , 32'h00070687 , 32'hFFFC393C , 32'h00040EF6 , 32'h0004A506 , 32'hFFFB997C , 32'hFFFF24D1 , 32'h00082B9C , 32'h0006BD4F , 32'h00097352 , 32'hFFFA0B7F , 32'h0006C086 , 32'h00074EE2 , 32'hFFFEFC75 , 32'hFFFC1C11 , 32'h000037BB , 32'h00055DEE , 32'h00002706 , 32'h0004B862 , 32'h00028941 , 32'hFFFFB244 , 32'hFFFEAE6E , 32'h0004BCEA} , 
{32'h0004DF9A , 32'h00020BCF , 32'h0001406A , 32'hFFFE8535 , 32'h00014850 , 32'hFFFC5D63 , 32'h0002AE8E , 32'hFFFCEBA2 , 32'h00011AE0 , 32'hFFFA57B9 , 32'h000119C3 , 32'h00029E6B , 32'hFFFF6ECD , 32'h00013C65 , 32'hFFFAA173 , 32'hFFFDEA82 , 32'h0000D7E4 , 32'hFFFF6860 , 32'h00063AD4 , 32'hFFFB3426 , 32'hFFF93B94 , 32'hFFFF9DBE , 32'h0003AADD , 32'h000186ED , 32'hFFF7C825 , 32'hFFFD0206 , 32'h00049523 , 32'h00069115 , 32'hFFFFC204 , 32'h000694AF , 32'h000079DB , 32'h0002E569 , 32'h0002397C , 32'hFFFCAF15 , 32'hFFFBC954 , 32'hFFFB5742 , 32'h0002D623} , 
{32'h00026E26 , 32'h000260D6 , 32'hFFFED2FA , 32'hFFF7798F , 32'hFFFCFD97 , 32'h0004EB65 , 32'hFFFB5157 , 32'hFFFA07AA , 32'hFFFE2CCC , 32'hFFFEEBFB , 32'hFFFD1D0B , 32'h00029DBB , 32'h0000DF56 , 32'hFFFF9CCB , 32'h00053A85 , 32'h00065D25 , 32'hFFFB3BB4 , 32'hFFF95BE1 , 32'hFFFE1B41 , 32'h000120EE , 32'hFFFD876B , 32'hFFFE9B0D , 32'hFFFC0ECC , 32'h0000CA94 , 32'h0002B966 , 32'h00013419 , 32'h00023F87 , 32'h0002A63E , 32'h000021DA , 32'h0000A20A , 32'h0006B234 , 32'hFFFD1FDD , 32'hFFFE4DAC , 32'hFFFAD2C3 , 32'hFFFDF1FA , 32'h0002CFED , 32'h00069951} , 
{32'h0002388F , 32'hFFFBA332 , 32'h00051A18 , 32'hFFFC83FE , 32'hFFFA3F27 , 32'hFFFEFB7A , 32'hFFF799BD , 32'hFFFCA666 , 32'h00001096 , 32'hFFFFCA6E , 32'h000123E7 , 32'hFFF8F7E8 , 32'h00021ABA , 32'hFFFB34BA , 32'h0001B493 , 32'h0005B2CD , 32'h0002633F , 32'hFFFFC9FB , 32'hFFFD3B18 , 32'h0002A673 , 32'hFFF98335 , 32'hFFF6270F , 32'hFFF81F87 , 32'h000273CC , 32'hFFF5341D , 32'hFFFCF37C , 32'h00014C2B , 32'h0001F2D2 , 32'hFFF93D40 , 32'hFFFB15AC , 32'hFFFD0DF2 , 32'h00005713 , 32'h000745B6 , 32'h0001E18E , 32'hFFFD2372 , 32'hFFFC70E3 , 32'h000146CE} , 
{32'hFFFA8E84 , 32'h0008DA5A , 32'h000344C5 , 32'h00042F6D , 32'h0001A3A1 , 32'hFFFB524E , 32'h00015113 , 32'hFFFE3517 , 32'hFFF93F35 , 32'hFFF9FB78 , 32'h0003A938 , 32'h0000D854 , 32'h00049995 , 32'h0004886A , 32'h0005E761 , 32'h00036689 , 32'hFFF9B256 , 32'h000298C6 , 32'h00021EB9 , 32'h000802F0 , 32'hFFFEBE5F , 32'hFFFDCBA9 , 32'h000787CB , 32'hFFF6B9A0 , 32'hFFF9F147 , 32'hFFFC96DF , 32'hFFF345F0 , 32'h00000141 , 32'hFFFF7A03 , 32'h000508D5 , 32'h0000F37D , 32'hFFF9BC6F , 32'hFFFAB0E1 , 32'hFFFF8379 , 32'hFFFA0246 , 32'h00064D0F , 32'hFFFC35A1} , 
{32'hFFFF06B1 , 32'h0003D070 , 32'h00010B7E , 32'h00030615 , 32'hFFFFA18E , 32'hFFFE04F5 , 32'h0007332E , 32'hFFF74458 , 32'h00018130 , 32'hFFFDB342 , 32'h000150B0 , 32'hFFFC9F64 , 32'h000205F2 , 32'h0001A73F , 32'h0009CF2E , 32'h0000C6AD , 32'hFFF96663 , 32'h000796AF , 32'hFFFEDC67 , 32'hFFFC9BD6 , 32'h000781E7 , 32'hFFF76172 , 32'hFFFD3A4E , 32'h0004D5E8 , 32'h00073542 , 32'h0004890C , 32'h0005B66A , 32'h0003C7DE , 32'h00047273 , 32'hFFFAC71B , 32'h00047419 , 32'hFFFEA669 , 32'h000200E1 , 32'h000162C8 , 32'hFFFDA8E4 , 32'h00008EBD , 32'hFFFE8F7D} , 
{32'h0001DAC2 , 32'hFFF7819A , 32'hFFFDEC34 , 32'h000158D5 , 32'hFFFFA57F , 32'h0001E17C , 32'h0008B975 , 32'hFFFC9395 , 32'hFFFF876D , 32'h000400F1 , 32'hFFFFB433 , 32'hFFFA5128 , 32'h0007ACA7 , 32'hFFF901B7 , 32'h00007D81 , 32'hFFFFF42A , 32'hFFFBD60B , 32'hFFFB068C , 32'h00021242 , 32'h000461BC , 32'hFFFEDCCF , 32'hFFFD790D , 32'hFFFE9257 , 32'h0005507F , 32'hFFFD13B1 , 32'h00049956 , 32'hFFFCCBCE , 32'h000063DE , 32'h0001D337 , 32'hFFFE23FE , 32'h00043A28 , 32'h00056A67 , 32'hFFFD7E1A , 32'hFFFB3D51 , 32'h00019FD7 , 32'h000320BB , 32'hFFF8B0BD} , 
{32'hFFFFEF08 , 32'hFFF0040C , 32'h000CF270 , 32'hFFFC023C , 32'hFFF7F3D1 , 32'hFFFA9E7F , 32'h000A4FC7 , 32'h000553F8 , 32'hFFFE2C52 , 32'hFFFD3342 , 32'hFFFFE5FA , 32'h00054D52 , 32'h000806DF , 32'h0005B075 , 32'hFFF710FA , 32'h00009E9F , 32'hFFFA3F55 , 32'h0009150D , 32'h000314EF , 32'h00032733 , 32'hFFFE6877 , 32'hFFFA2026 , 32'h0002358E , 32'hFFFC37ED , 32'h0005625E , 32'h000AD4C6 , 32'hFFFEAA82 , 32'hFFFCBCB7 , 32'h0002F6F6 , 32'hFFF93E67 , 32'hFFF53503 , 32'hFFFE2313 , 32'h000B908B , 32'hFFFC2A53 , 32'hFFF01A5F , 32'h00041B58 , 32'h00006B7F} , 
{32'h00030230 , 32'hFFF99551 , 32'hFFFFA7A1 , 32'hFFFE7DDB , 32'h0007318B , 32'h0004C676 , 32'hFFFBAA22 , 32'h00017FF3 , 32'hFFFED30E , 32'hFFFAC141 , 32'h000A926C , 32'hFFFF5ACE , 32'h00049486 , 32'hFFF9F4A0 , 32'h0002E44C , 32'hFFF74E4B , 32'h0008F924 , 32'h0005E923 , 32'hFFFEE456 , 32'hFFF900B2 , 32'h000246DB , 32'hFFFB1A11 , 32'h00087A91 , 32'hFFF0BF99 , 32'h00010CAD , 32'hFFFD462A , 32'h0000B41B , 32'h0009FFA0 , 32'hFFF6D66D , 32'h0004CCD6 , 32'h0004EBDC , 32'h00000DB2 , 32'h00029DCC , 32'h000553DC , 32'hFFF9F493 , 32'hFFF186D5 , 32'hFFFC79B8} , 
{32'h00032427 , 32'h0001F134 , 32'h0009B3CC , 32'h0002717B , 32'h0001F7FC , 32'h0006BF26 , 32'h00030C47 , 32'hFFFE16AC , 32'hFFFF0725 , 32'hFFFF5BA4 , 32'hFFFF5B11 , 32'h0005966A , 32'hFFFB2F6E , 32'hFFFEC701 , 32'hFFF811DF , 32'h00000688 , 32'h00009AF3 , 32'h0002E391 , 32'h0007B8A1 , 32'hFFFC251F , 32'h0002D7C5 , 32'h000113A3 , 32'hFFFFAA30 , 32'hFFFC2594 , 32'h00033C6F , 32'hFFFF75C5 , 32'hFFF4B39A , 32'hFFFD33D7 , 32'h00072A02 , 32'h00080811 , 32'h00009D06 , 32'hFFFCFED8 , 32'hFFFF3D14 , 32'h000049B5 , 32'hFFFAE67E , 32'hFFF5F9D6 , 32'hFFFF308D} , 
{32'h0002C288 , 32'hFFFF32C6 , 32'h00019821 , 32'h0000F055 , 32'hFFFAD155 , 32'h000748AE , 32'h00019F29 , 32'hFFF9A603 , 32'h0001ED00 , 32'hFFFE6BFD , 32'h0002961E , 32'h00008E4E , 32'h00001FE5 , 32'hFFFDF7E9 , 32'hFFFFFE56 , 32'h00006B43 , 32'h00006759 , 32'hFFF98D66 , 32'h00061DDC , 32'h0000733A , 32'hFFFCAA63 , 32'hFFFE814C , 32'h00014367 , 32'h00018030 , 32'hFFFF5C9D , 32'hFFF9D312 , 32'h0000D061 , 32'hFFFF9108 , 32'h00013562 , 32'hFFFFF90F , 32'hFFFCCE9C , 32'h000240E6 , 32'hFFF5809F , 32'h00048C40 , 32'hFFFE670D , 32'hFFFF870C , 32'h0001029C} , 
{32'h0001BA98 , 32'h0002243E , 32'h000686DD , 32'h0003594B , 32'h0000FD4D , 32'hFFFB82C4 , 32'hFFF7A37A , 32'h00011375 , 32'h000680F9 , 32'hFFFED404 , 32'h00043226 , 32'h0003A37C , 32'h00019A18 , 32'hFFFBCC18 , 32'hFFFDA412 , 32'hFFFF7B65 , 32'h000926DB , 32'h0001D105 , 32'hFFFC73AA , 32'h0000A315 , 32'hFFFE662E , 32'h0001F3E1 , 32'h00013E8B , 32'h0007DCE5 , 32'hFFFC291E , 32'h000552E3 , 32'h0004C495 , 32'h00034634 , 32'hFFFF49FC , 32'hFFFDEA5D , 32'hFFFE2EF4 , 32'h0004DFED , 32'hFFFB4A85 , 32'hFFFEF8E7 , 32'h0001DCBB , 32'h00022971 , 32'h00001EA2} , 
{32'h000445D8 , 32'hFFFD32A7 , 32'hFFF934C0 , 32'hFFFEAC92 , 32'hFFFDE887 , 32'h0000BA86 , 32'h0000CABB , 32'hFFFE1F45 , 32'h0006FFC8 , 32'hFFFB8CF1 , 32'h0006BCA4 , 32'hFFFCD832 , 32'h0002E81B , 32'hFFFCCB6E , 32'h00022F41 , 32'h0007AAC6 , 32'hFFFC9873 , 32'hFFF9CDE1 , 32'hFFFF781F , 32'h000562FB , 32'h00018066 , 32'h00061F09 , 32'hFFFE3F56 , 32'hFFFF4CF1 , 32'hFFFF9198 , 32'hFFFBC4EE , 32'h0007E6D3 , 32'h00036111 , 32'h0002A8E1 , 32'hFFF8FE19 , 32'hFFFF8E15 , 32'h00058CE4 , 32'h0000E419 , 32'h0000C92B , 32'h000061BE , 32'h000310E1 , 32'h00044D2B} , 
{32'h0002F144 , 32'h0005387D , 32'h0007E5A8 , 32'hFFFF04F6 , 32'hFFFCB6A8 , 32'h000A9EB1 , 32'hFFFB49CB , 32'h0006AA19 , 32'hFFFDFBCC , 32'hFFFFE85D , 32'hFFFB444C , 32'h00092022 , 32'h0007F7E1 , 32'h0003E9A4 , 32'hFFF4E451 , 32'hFFFD63E2 , 32'h0006D767 , 32'hFFF73D86 , 32'hFFFDBBFD , 32'h000252FF , 32'hFFF91DA1 , 32'h00021EE5 , 32'hFFFF6690 , 32'h00018CBD , 32'h000042F3 , 32'hFFFBEF71 , 32'hFFF90525 , 32'h00050B44 , 32'h00026454 , 32'h000999B7 , 32'hFFF7B5D8 , 32'hFFFE945B , 32'hFFFF7370 , 32'h000135DA , 32'hFFFCBA7F , 32'h000786C3 , 32'hFFF80379} , 
{32'h00048FD0 , 32'hFFF740ED , 32'h0002B2BA , 32'hFFFEFAA5 , 32'hFFF5F835 , 32'h00041FF2 , 32'h0003A05B , 32'hFFFB9AE9 , 32'h000593DD , 32'hFFFC282F , 32'h000414AE , 32'hFFFF17E4 , 32'h00033FC4 , 32'h0000180F , 32'hFFF68502 , 32'h00014664 , 32'hFFFC83F8 , 32'hFFF60C49 , 32'h000BC1CA , 32'h00007711 , 32'h0000831C , 32'hFFFCB4F1 , 32'h0006E848 , 32'hFFFE63CF , 32'h0004EE94 , 32'hFFFE8D9A , 32'h00050431 , 32'h0001834F , 32'hFFFD14A1 , 32'h00002E9E , 32'h0002CD33 , 32'h00015D3C , 32'h0002179F , 32'h0003876A , 32'h000177A3 , 32'h00041324 , 32'h000436B1} , 
{32'hFFFFA64C , 32'h0005347D , 32'h00050FE3 , 32'h000B7AE0 , 32'hFFFEDB52 , 32'h00033FF9 , 32'h0002C418 , 32'h00015528 , 32'hFFF75F29 , 32'hFFF67683 , 32'h0000C5D6 , 32'hFFFB9853 , 32'h00007EC6 , 32'hFFF7F374 , 32'hFFFF75DB , 32'h00031F8A , 32'h000037F7 , 32'h00048506 , 32'hFFFFC611 , 32'hFFF75969 , 32'hFFFD1B3F , 32'h00039930 , 32'h0000820C , 32'h000219DE , 32'h000700BE , 32'hFFFAAED1 , 32'hFFFE9356 , 32'hFFFEC017 , 32'hFFFCC398 , 32'h00003D81 , 32'h0007D9FD , 32'h00015A27 , 32'hFFFDD892 , 32'hFFF92AD8 , 32'h0004DEC6 , 32'h00082FA8 , 32'h00064B94} , 
{32'hFFFEDBE9 , 32'h0001FAED , 32'h00072FB5 , 32'hFFFFEA4D , 32'hFFFE18DC , 32'hFFFDEFEE , 32'hFFFA2B3A , 32'h00038912 , 32'hFFFD1EDE , 32'h00067D93 , 32'h0000BF98 , 32'hFFFAA5A6 , 32'h000350F7 , 32'hFFFD9F94 , 32'h0001AE42 , 32'hFFFB3095 , 32'hFFFD4F13 , 32'h0001EB62 , 32'hFFFACD12 , 32'hFFFC35D2 , 32'hFFFD9331 , 32'hFFFEF22E , 32'h0001F175 , 32'h00037567 , 32'hFFFC2F48 , 32'h00025390 , 32'hFFF8FA00 , 32'hFFFD7E93 , 32'h0003500B , 32'h000A34EC , 32'h00003DAC , 32'h00075483 , 32'h0008909B , 32'hFFFEDE18 , 32'hFFF94871 , 32'h00051743 , 32'h0002D597} , 
{32'h000799DA , 32'h0001314A , 32'hFFFFEA6E , 32'h0003EB00 , 32'hFFFBC6FF , 32'hFFFE2B40 , 32'h0002C3C1 , 32'h000035DD , 32'hFFF6D2EE , 32'h0003094A , 32'hFFF9FC3E , 32'hFFFCDE3D , 32'hFFFD42A6 , 32'hFFF8BCB5 , 32'h000636C8 , 32'hFFFC13B6 , 32'h000135DE , 32'hFFF7DEAF , 32'h00025CEC , 32'hFFF9F4F9 , 32'h00006B4D , 32'h00045019 , 32'hFFF8A05A , 32'h000184CC , 32'h00056131 , 32'hFFFD885C , 32'h0000694E , 32'h0004149B , 32'hFFFB7111 , 32'h0001AD9D , 32'h000066BF , 32'hFFFDEA25 , 32'hFFFDB51C , 32'h0009395A , 32'hFFFBF268 , 32'hFFF875F9 , 32'hFFFCBC50} , 
{32'h000350E9 , 32'h00012ED1 , 32'h0003E110 , 32'hFFFECC9D , 32'hFFFFB705 , 32'hFFFEE0FD , 32'hFFFF64E9 , 32'h0007794E , 32'hFFFAE64E , 32'hFFFD4262 , 32'hFFFCFF3D , 32'h000389E2 , 32'h00030C8B , 32'hFFFE19CA , 32'hFFF6A622 , 32'h000467CC , 32'h0000D4D1 , 32'h000004C4 , 32'hFFFDAD0B , 32'h0005721A , 32'h0001C607 , 32'h00034089 , 32'h00023F06 , 32'hFFFF27C9 , 32'h00043A0D , 32'hFFFE73C1 , 32'h00020C60 , 32'hFFF9EB66 , 32'h0003A7AF , 32'hFFFE1A64 , 32'h0002D1D5 , 32'hFFFFEAAC , 32'hFFFC4F5C , 32'h0002484D , 32'hFFFD619C , 32'hFFFE356E , 32'hFFFEF963} , 
{32'hFFFF4600 , 32'h0002256A , 32'hFFF4635B , 32'hFFF84EEB , 32'hFFFB0B28 , 32'h0005F26D , 32'hFFF9D809 , 32'h0004790E , 32'hFFFF363D , 32'h0008A859 , 32'hFFF9FABF , 32'h000083BB , 32'hFFFAACA1 , 32'h000414A4 , 32'h00021EAC , 32'hFFFFE918 , 32'h00094BDE , 32'h00058870 , 32'h000178AA , 32'h0004AEBF , 32'hFFFD60B8 , 32'h00039641 , 32'hFFFFE1FD , 32'h00075994 , 32'h00016AC0 , 32'hFFFB0CCD , 32'h00059A99 , 32'hFFF958B8 , 32'hFFFBB4D6 , 32'h0005FE5C , 32'h000871FE , 32'h0008800F , 32'h0009CD5B , 32'hFFFBB6BF , 32'h00003F8C , 32'h0001764B , 32'h00038EF5} , 
{32'hFD4B1550 , 32'hF7DB5920 , 32'hFB3F7630 , 32'h08895E10 , 32'hFE0A6668 , 32'hFF1DA6EA , 32'hFD7B9654 , 32'h04AF2DF0 , 32'h0A572D30 , 32'hFD9B2C30 , 32'h015F887C , 32'h084A5370 , 32'hFDF75F18 , 32'hFD6914A8 , 32'h01CD749C , 32'hF78405A0 , 32'h03006294 , 32'h01E7DD64 , 32'hF88BB2F0 , 32'hF5C5FE10 , 32'h08564D50 , 32'h009B59BB , 32'hFE7047F4 , 32'h0C729F30 , 32'hFFD25BD0 , 32'h06482060 , 32'h0C2604F0 , 32'h032DB4E0 , 32'h02B56D84 , 32'h014DD6A8 , 32'h00C372FF , 32'hFB053EC8 , 32'hF8657B98 , 32'h04C62F08 , 32'hF9D0ECA0 , 32'h04241C88 , 32'hFC0E246C} , 
{32'h00017EE3 , 32'h00023F7F , 32'hFFFB9E0C , 32'h00026D89 , 32'hFFFBF7F5 , 32'h0003A726 , 32'hFFFFF090 , 32'hFFFCE76D , 32'h00054410 , 32'hFFFF6CDB , 32'h0000086B , 32'hFFFC762B , 32'hFFF8CEC7 , 32'h0005D40E , 32'h0002834A , 32'hFFFD5E60 , 32'h00013F56 , 32'hFFFFD29A , 32'h00021C6E , 32'h0000CA9B , 32'h0002CB55 , 32'h00019049 , 32'hFFFE0C58 , 32'hFFFC9902 , 32'h00025D12 , 32'h0004FFCF , 32'h0002C7C0 , 32'hFFFFAAC4 , 32'h0001DE27 , 32'hFFFE44BC , 32'hFFFEA907 , 32'h0001D8ED , 32'h0002A4CD , 32'h0002A404 , 32'h0007AFC6 , 32'hFFFEA99B , 32'h0000B5C4} , 
{32'hFCECD8CC , 32'hF6C63300 , 32'hFA9EFE20 , 32'h09AE3850 , 32'hFDC603DC , 32'hFF00C340 , 32'hFD2C73B8 , 32'h05459EE8 , 32'h0BB9F890 , 32'hFD4CB9A0 , 32'h018E2DF8 , 32'h095F39D0 , 32'hFDB72F34 , 32'hFD10FCF0 , 32'h020E3430 , 32'hF6600A90 , 32'h036C28F0 , 32'h022A7EA0 , 32'hF7847EF0 , 32'hF4677F70 , 32'h096678E0 , 32'h00B3F851 , 32'hFE398D28 , 32'h0E20E860 , 32'hFFCB7279 , 32'h071C6828 , 32'h0DCA9710 , 32'h03A11F78 , 32'h030F8404 , 32'h017AB830 , 32'h00DADFA1 , 32'hFA5CD208 , 32'hF75AB970 , 32'h056DFAD8 , 32'hF9015198 , 32'h04B6BB60 , 32'hFB84CC50} , 
{32'hEA798F80 , 32'h102A46E0 , 32'h084C6030 , 32'hF9084508 , 32'h06B07B98 , 32'hEB5EF360 , 32'h0A36DE10 , 32'hFAC06920 , 32'h165B9BA0 , 32'hFD748974 , 32'hE84EAE40 , 32'h06FDE2F8 , 32'h0FA23E80 , 32'h05C26818 , 32'h06953710 , 32'h0379FC70 , 32'h09D72E60 , 32'h013E21A0 , 32'h00E64564 , 32'hFC5C012C , 32'hFD2A7004 , 32'hFD582A18 , 32'hF9C068C8 , 32'hFFC72E88 , 32'hFBB66850 , 32'hFAEF7410 , 32'h10A52DA0 , 32'hF0FE1630 , 32'h00A0E866 , 32'h0A5378F0 , 32'hF3D23630 , 32'hF9D79C30 , 32'h09B82AE0 , 32'hFA6964C8 , 32'h03479EAC , 32'h03D4C2E4 , 32'hFE106190} , 
{32'h0B179920 , 32'hEB5E9760 , 32'hFEA5FC14 , 32'h0405F400 , 32'hFB1290E0 , 32'hFB3F7BD0 , 32'hF898BB48 , 32'h0D171BA0 , 32'h17446E60 , 32'h005F6017 , 32'hFE92C140 , 32'h103E8F40 , 32'h0008C9C6 , 32'h0B848210 , 32'h062EFF80 , 32'hECFFCFC0 , 32'h067FB9F8 , 32'hFDF3B3FC , 32'hEAE00FA0 , 32'hEFE2ACA0 , 32'h0318E300 , 32'h06BD2C58 , 32'hFBD535F0 , 32'h09F4BA40 , 32'h087203E0 , 32'hFD597C0C , 32'h0D236050 , 32'hFB4520B8 , 32'h02B97B98 , 32'hFCA12C34 , 32'h02186958 , 32'hF5453210 , 32'hFE0B0D50 , 32'h16697EC0 , 32'hF6A14350 , 32'h041354C0 , 32'hFAD0DF58} , 
{32'h211B1FC0 , 32'hF05E1B30 , 32'hF8636D60 , 32'h04084118 , 32'h0031C363 , 32'hFEAF5524 , 32'h0C427B00 , 32'hF8BA6D40 , 32'h07E9F500 , 32'h07AB58C8 , 32'hFB531DD0 , 32'hFD89DE60 , 32'h036AEF48 , 32'h27F2CE40 , 32'hFB739618 , 32'hF7510260 , 32'h0C4DB3A0 , 32'h0B5F98C0 , 32'hEC295E40 , 32'hFDAF6824 , 32'h004A449F , 32'h09630540 , 32'h13571D20 , 32'h05BE8D50 , 32'h080E4D50 , 32'hFA8D9328 , 32'hF922C748 , 32'hE45B69A0 , 32'h05A474B0 , 32'hF8EA3040 , 32'hE91EC580 , 32'hFB844738 , 32'h120CC540 , 32'h0DE30F90 , 32'hF940F690 , 32'h025EB5D8 , 32'h01D6249C} , 
{32'hFCA247E8 , 32'hF23644C0 , 32'hF84689F8 , 32'h0E785760 , 32'hFCBAC2B4 , 32'hFB2B3358 , 32'hF934D768 , 32'h10E75CA0 , 32'h0E55F1E0 , 32'h00BE75E3 , 32'h023E3850 , 32'h0EA45490 , 32'hFBF17198 , 32'hF9CE84C0 , 32'h07054F30 , 32'hEED05500 , 32'h094B0100 , 32'h04E5BD98 , 32'hF4CFC7B0 , 32'hEA949F80 , 32'h0BB124B0 , 32'h0625CEE0 , 32'hFEEDA730 , 32'h19084760 , 32'hFF5C3763 , 32'h08DCE6D0 , 32'h1D625D60 , 32'h04BC1D60 , 32'h0B572B60 , 32'h07C51BA8 , 32'h08A98A80 , 32'hF7287F60 , 32'hEE4520E0 , 32'h0AFA29A0 , 32'hF33979A0 , 32'h05D57818 , 32'hFF8B2FC3} , 
{32'h08419010 , 32'hF88604F0 , 32'h00CA62CA , 32'h006DBFAB , 32'hFA60ACB8 , 32'hFC695DC0 , 32'hFE3D0FB0 , 32'hFD0B2928 , 32'hDBDC3980 , 32'hF81616B8 , 32'h03564244 , 32'hF1805910 , 32'hE8B0E660 , 32'hF7BCFEE0 , 32'hF377C120 , 32'hE2EC4A00 , 32'h1274C0E0 , 32'hFC0BC4A4 , 32'h11AA6E40 , 32'h0983AFC0 , 32'h00D3EE85 , 32'h0F8026D0 , 32'h113DC880 , 32'h0A10A990 , 32'h0C612490 , 32'hF25AEBB0 , 32'hF5AC7E00 , 32'h01DBA868 , 32'h046A4210 , 32'hFA464F48 , 32'h0ED4F680 , 32'hFF61367E , 32'hF33BCE60 , 32'h07D6E7A8 , 32'hE9B97760 , 32'hFCB25D8C , 32'h02E327B0} , 
{32'hFD5C7684 , 32'h015F5614 , 32'hFEF40014 , 32'h01D757B0 , 32'hFE533C08 , 32'h00562353 , 32'hFF28E0AB , 32'h0082E79F , 32'hFED24E1C , 32'h03A80D98 , 32'hFDE8250C , 32'hFEBE6830 , 32'hFD6F3EE4 , 32'hFF96CA88 , 32'h012F15C0 , 32'hFFBE96ED , 32'h00E8E1A5 , 32'hFD709AE8 , 32'hFB37F738 , 32'hFF9C0359 , 32'hFC2794D4 , 32'h04ED8810 , 32'hFF1063F3 , 32'hFE7E1990 , 32'hFEA7F80C , 32'hFE6A3A50 , 32'hFE3F97D4 , 32'hFF7074C8 , 32'hFEF7EF2C , 32'hFEBD4F78 , 32'hFDCDB130 , 32'hFCF1256C , 32'h0092FFE6 , 32'hFF8CA0E4 , 32'h01C9EAD8 , 32'h013B823C , 32'h004EFB94} , 
{32'hFF206A5E , 32'h02F95D6C , 32'h08143180 , 32'h012529DC , 32'hFE573F48 , 32'hDADFB840 , 32'h08FAA020 , 32'h0DF930E0 , 32'hDB17FEC0 , 32'hF65A49D0 , 32'hFBEBBF50 , 32'hF9CAF010 , 32'hFF4B6B01 , 32'hFF9F63D1 , 32'h02529C2C , 32'hE7BE8180 , 32'h12F97F60 , 32'h065595F0 , 32'h106785C0 , 32'hFE05BD48 , 32'hF5CC42F0 , 32'h1E4599C0 , 32'h056EC3F0 , 32'h0B859F70 , 32'h0BFBA9D0 , 32'hFCC70F24 , 32'h026BEBC0 , 32'h11717FC0 , 32'hFE8245B4 , 32'hF9DD5410 , 32'h031C629C , 32'h027430B4 , 32'h044A5AA0 , 32'h0596B518 , 32'hEAFE2E20 , 32'hF46B6670 , 32'hF9A71BA0} , 
{32'h0ADC24A0 , 32'hFB36FF60 , 32'h0A7AEC30 , 32'hE47656C0 , 32'h04BBB470 , 32'hFBCF99A8 , 32'hFAAE7DE0 , 32'hE5658EE0 , 32'h0A82F330 , 32'h294AE840 , 32'h0EEC2D00 , 32'hFF4E87CF , 32'hEA1C8060 , 32'hF501AE20 , 32'hF6C50380 , 32'hE974B6A0 , 32'h0CC3E830 , 32'h07D7A428 , 32'hF0F51080 , 32'h091B7EA0 , 32'hF7DA6880 , 32'hFAEA4CD8 , 32'hE01951C0 , 32'h09328810 , 32'hF40ACE90 , 32'hE7F10800 , 32'h0713C5B0 , 32'h2095F000 , 32'h122C3C60 , 32'hF92A65A8 , 32'h01450C5C , 32'hFFEC5CFA , 32'hF677D790 , 32'hEF98F660 , 32'h103DB9C0 , 32'h08E30050 , 32'hFFD3EC27} , 
{32'hE9941760 , 32'h0AE9F9E0 , 32'hF6580D60 , 32'h0F97CBA0 , 32'h01095088 , 32'h0A68D1D0 , 32'hFE073BBC , 32'h0A2DCD90 , 32'hF1BCD3D0 , 32'hF982C1F8 , 32'h0195FF70 , 32'h02B1FDE0 , 32'hFF6666B8 , 32'hEC2CDF40 , 32'hF6CDFC50 , 32'h051A5110 , 32'hFB6AC718 , 32'h025E5048 , 32'h0341B5A4 , 32'hFFE5ED9A , 32'h05ECD8F8 , 32'hF8D81F28 , 32'hF7176C10 , 32'hFF0B80C9 , 32'hFC133FFC , 32'h0108554C , 32'hFFECAB57 , 32'h12B9E480 , 32'hFD6FB874 , 32'h000EFC94 , 32'hFD04F71C , 32'h0478AF80 , 32'hF5014870 , 32'hEF9BA4E0 , 32'h0B2C6510 , 32'hF67F7E40 , 32'hFA2FDE30} , 
{32'hF691B4B0 , 32'h061E5AE8 , 32'hFCA5BC14 , 32'h025AE240 , 32'h00204F34 , 32'h053B4708 , 32'hFFC08445 , 32'hFF0C2833 , 32'hF9AD1E50 , 32'hFC0A1D24 , 32'h004C99EF , 32'hFEAC80A0 , 32'hFDE13F48 , 32'hF5176A40 , 32'hFC59CAC0 , 32'h03678960 , 32'hFC88F6C0 , 32'hFFB7CDBE , 32'h06407E18 , 32'hFEBE5C60 , 32'h0454DE20 , 32'hF9AFEA50 , 32'hFE9BB034 , 32'hFF1848E4 , 32'hFD08C6EC , 32'h023B1674 , 32'h020D5130 , 32'h099F4470 , 32'hFE913284 , 32'h00CDAE9E , 32'hFFB23EFF , 32'h012D5B54 , 32'hFC1228B8 , 32'hFAA14C20 , 32'h022CDF0C , 32'hFFCB543E , 32'hFF0D90EA} , 
{32'hECD885E0 , 32'h0C6B72B0 , 32'hF92425F8 , 32'h04C0E4E8 , 32'h0042A15D , 32'h0A998B10 , 32'hFF833764 , 32'hFE08B5B0 , 32'hF32B2410 , 32'hF800C310 , 32'h00973B59 , 32'hFD411848 , 32'hFBB8DC08 , 32'hE9E10FA0 , 32'hF8A01EC0 , 32'h06E65B38 , 32'hF8FBDAD8 , 32'hFF72B414 , 32'h0CB518B0 , 32'hFD6E5488 , 32'h08C5B650 , 32'hF335D6C0 , 32'hFD3034FC , 32'hFE287F58 , 32'hF9F5F0C0 , 32'h047F1818 , 32'h04291760 , 32'h137E8FA0 , 32'hFD230154 , 32'h01A64B18 , 32'hFF60B53E , 32'h0260047C , 32'hF80A28C8 , 32'hF5142280 , 32'h046B18C8 , 32'hFF8FF07E , 32'hFE13A664} , 
{32'h00037A23 , 32'h00001965 , 32'h0001B9F3 , 32'h0002ACA0 , 32'h0009FF9B , 32'h00020A83 , 32'hFFFF9327 , 32'h000152B9 , 32'h0003DCF7 , 32'h00011A2B , 32'h00012B11 , 32'h00013ACA , 32'hFFFDCE7C , 32'hFFFF1219 , 32'hFFFCF111 , 32'h00010284 , 32'hFFFFF44C , 32'hFFFB05AF , 32'hFFFB7A14 , 32'h00052FC8 , 32'hFFFF682A , 32'hFFFE7852 , 32'h0004837F , 32'hFFFE1A1F , 32'h000417E4 , 32'hFFFFCB30 , 32'h0000CC57 , 32'hFFFFE6C9 , 32'hFFFF33D4 , 32'hFFFF795D , 32'hFFFEFD17 , 32'hFFFBF4BD , 32'h000157D0 , 32'h00004290 , 32'hFFFDD427 , 32'hFFFFD13E , 32'hFFF9BE9A} , 
{32'h0000CC7B , 32'h0005B28F , 32'hFFFFD3EE , 32'h0003006E , 32'h0000A106 , 32'hFFFFE15B , 32'hFFF818D4 , 32'h0007F90C , 32'h0003846B , 32'hFFFE366F , 32'hFFFA9D26 , 32'hFFFEF996 , 32'h000AD5BA , 32'h0005DB08 , 32'h0004D41F , 32'hFFFDD345 , 32'hFFFBE053 , 32'hFFFE727A , 32'h0003B0E8 , 32'hFFFAB53C , 32'hFFFA31EF , 32'hFFFEF23A , 32'h00054887 , 32'h00011CE7 , 32'h0000134E , 32'hFFFB44BC , 32'h0000EC13 , 32'hFFFF086D , 32'hFFFF068E , 32'hFFFCA078 , 32'hFFFA075F , 32'hFFFFE2F3 , 32'hFFFED2E4 , 32'hFFFA8770 , 32'hFFFD3183 , 32'hFFFD2852 , 32'hFFFE4FF9} , 
{32'h0001672B , 32'hFFFBA3F2 , 32'h0001910C , 32'h00054818 , 32'h00044810 , 32'hFFF9DDE7 , 32'hFFFFD04C , 32'h00055AF8 , 32'h000339A9 , 32'hFFFD299C , 32'hFFFD27D2 , 32'h0003C65C , 32'hFFF93186 , 32'h00043DE1 , 32'hFFFF9AB8 , 32'h0004722D , 32'hFFFF47AC , 32'h0002C7D6 , 32'hFFFFF324 , 32'hFFFD839B , 32'h000239F9 , 32'h00059A0F , 32'h0004CA27 , 32'h0007C736 , 32'h00012FA5 , 32'hFFFBBFD6 , 32'h000562FF , 32'h00041AF0 , 32'h00035602 , 32'hFFFD9295 , 32'h00046E63 , 32'h00022632 , 32'h00048F2D , 32'hFFFCD892 , 32'h0002F4A6 , 32'hFFF8AB9B , 32'hFFFAE50C} , 
{32'hFFFE5BF8 , 32'hFFFDE9F5 , 32'h0002BE67 , 32'h00051F55 , 32'hFFFE33AD , 32'h0000C50D , 32'h000820DD , 32'h00036DCF , 32'hFFFCB86D , 32'hFFFECBA5 , 32'hFFFE1697 , 32'h00011448 , 32'hFFF8C7A3 , 32'hFFF5BBE8 , 32'h0002DDD7 , 32'h00039995 , 32'h0004790A , 32'hFFF8F4CA , 32'hFFFED8A6 , 32'h000A80E1 , 32'h000330D5 , 32'hFFFD1AC6 , 32'h0008BD4C , 32'hFFFB8368 , 32'h00027260 , 32'hFFFF3EA4 , 32'h00013875 , 32'h0003FD76 , 32'h0002D596 , 32'h000312BF , 32'hFFFED15F , 32'h0002CC97 , 32'h0001E8F5 , 32'h0006AA24 , 32'h0003575F , 32'h000060A3 , 32'hFFFCFE29} , 
{32'h0000B731 , 32'hFFFC1406 , 32'h00052E4B , 32'hFFFE5518 , 32'hFFFF374A , 32'h00030795 , 32'hFFFD623D , 32'h0003F797 , 32'h0006E5E3 , 32'h0003E445 , 32'h0002488D , 32'h00037588 , 32'hFFF8ADCE , 32'h000113CC , 32'hFFF84623 , 32'h00011FBB , 32'hFFF8429A , 32'hFFFFA055 , 32'hFFFF7947 , 32'h0003654F , 32'h00024DB7 , 32'h000006AE , 32'h00004BD4 , 32'hFFF885F4 , 32'hFFFB6592 , 32'h00019584 , 32'hFFFDBE68 , 32'h000045BB , 32'h0008C8D5 , 32'hFFF8287E , 32'h000667DD , 32'hFFFE1A33 , 32'hFFFE84B9 , 32'h00062ECA , 32'hFFF91AAB , 32'hFFF7817D , 32'hFFFD2F22} , 
{32'h00010DD2 , 32'hFFFA0883 , 32'h0003CE35 , 32'h00066C61 , 32'h000101B7 , 32'hFFFBA33E , 32'h000390A0 , 32'hFFFCE674 , 32'hFFFBC9C6 , 32'h0004F3A0 , 32'h0007FD64 , 32'h00013C31 , 32'hFFFE0611 , 32'hFFFCAF0E , 32'hFFFC8EDE , 32'hFFFFC389 , 32'hFFFA5D2A , 32'h00030F9D , 32'h000500FF , 32'h0007DD5C , 32'hFFF638B6 , 32'hFFFD42E1 , 32'h0007E09B , 32'h00042932 , 32'h0004B4F8 , 32'h000371D5 , 32'h0002FDBE , 32'h0005704A , 32'h00015252 , 32'h0001371A , 32'hFFFB34B1 , 32'hFFFF0358 , 32'h0004CBE8 , 32'h0004B71A , 32'h0003E15D , 32'h0005CCCF , 32'hFFFDF573} , 
{32'h000509CF , 32'hFFFEBC2B , 32'hFFF8691E , 32'hFFF697E4 , 32'hFFFA4557 , 32'h00031E76 , 32'h0000497D , 32'h00093C30 , 32'hFFF7F3EC , 32'hFFFDF341 , 32'h0006655A , 32'hFFFB0B3E , 32'hFFFFE345 , 32'h0001E891 , 32'h00006AC1 , 32'hFFFE2A22 , 32'hFFFC5FDF , 32'h000A7BA3 , 32'h000AC2A9 , 32'h0000F892 , 32'h0000F8FB , 32'hFFFC7323 , 32'h00013F9F , 32'h0000A1D5 , 32'hFFFFB527 , 32'hFFF8BCEC , 32'h0003974A , 32'h00057671 , 32'h000154B4 , 32'h0007BB0D , 32'h00064153 , 32'h000A6127 , 32'h0008F682 , 32'hFFFC4E86 , 32'h00086CAD , 32'h0004130B , 32'hFFF66C19} , 
{32'h000471DB , 32'h00005ED4 , 32'hFFFFFB40 , 32'h0000475D , 32'hFFFF5FAE , 32'h0000E4E7 , 32'h0004E0A0 , 32'hFFF89BAD , 32'hFFFF6952 , 32'hFFFC47E1 , 32'hFFFF4959 , 32'h000309A5 , 32'hFFFE62B8 , 32'h000364BC , 32'hFFFC6DCB , 32'hFFFA0029 , 32'h0002A4CC , 32'hFFFFCDAF , 32'h00056688 , 32'hFFFECB1C , 32'h0004A4B8 , 32'hFFFD7F70 , 32'hFFF9E6F8 , 32'h0002C54D , 32'hFFFCF0C8 , 32'hFFFECAC0 , 32'h0000C76D , 32'hFFF680C7 , 32'h0001A9EE , 32'h000E6F19 , 32'h00006C4B , 32'h0000477A , 32'h00012D13 , 32'h00058FDF , 32'h00039960 , 32'hFFFFB9C6 , 32'h00027C9A} , 
{32'hFFFF8C1D , 32'h00036EA9 , 32'h00006740 , 32'hFFFE2268 , 32'hFFFBF431 , 32'hFFFFE22B , 32'h000210C8 , 32'h0003B6C3 , 32'hFFF72ACD , 32'hFFF97F07 , 32'h00009DDD , 32'h0003CFD9 , 32'hFFFCFDBE , 32'h0005DC6F , 32'hFFF7DAE5 , 32'hFFFFAE7F , 32'hFFFA79E2 , 32'hFFFFF952 , 32'h0007B83B , 32'h000AA772 , 32'h0006706E , 32'h00023B76 , 32'h0006DDFE , 32'hFFFEFB9A , 32'h00017874 , 32'h0008659E , 32'hFFFF040E , 32'hFFFCD2E2 , 32'hFFFFC453 , 32'hFFFDE96F , 32'h000103F3 , 32'hFFFBBC0D , 32'hFFFAA50D , 32'hFFFD91A3 , 32'hFFFF0D16 , 32'h00068304 , 32'h00046A04} , 
{32'hFFFC42B1 , 32'h00026D3C , 32'hFFFEF906 , 32'hFFFE410B , 32'hFFFE3933 , 32'hFFF69A86 , 32'hFFFB426A , 32'h00017CF1 , 32'hFFFBCC03 , 32'h00036A1C , 32'h0001C756 , 32'h00049357 , 32'h00090325 , 32'h0002E679 , 32'hFFF43B49 , 32'hFFFD60BE , 32'hFFFE6F51 , 32'h0001B58F , 32'hFFFE6D97 , 32'hFFFC40FB , 32'h000172D8 , 32'hFFFDBCFC , 32'hFFF9EEF9 , 32'hFFFEDD83 , 32'hFFFEDA90 , 32'h0000CD83 , 32'h0002A84E , 32'hFFFE34B3 , 32'hFFFF5869 , 32'h0007AF7A , 32'h00039013 , 32'hFFFD593B , 32'hFFFF3C84 , 32'h00043938 , 32'h0002152B , 32'h00030B62 , 32'h0000E155} , 
{32'hFFFF76EC , 32'hFFFF033A , 32'h000190A5 , 32'hFFF20FB3 , 32'hFFFDDDBB , 32'h0001AB8A , 32'h000694BF , 32'hFFFBB6BA , 32'h0007541B , 32'hFFFD9C16 , 32'h0002BE92 , 32'hFFF7FD62 , 32'h00068DB8 , 32'h0002FC87 , 32'h0000D60D , 32'hFFFBB6A4 , 32'hFFFBBDDF , 32'h0009E336 , 32'h00003C66 , 32'hFFFA1792 , 32'h000038B1 , 32'hFFFC5EBA , 32'h0004B948 , 32'hFFFBA735 , 32'h00023898 , 32'h0001A0BA , 32'hFFFDC6BB , 32'hFFFEE373 , 32'hFFFA4167 , 32'h00010986 , 32'h0006D4DA , 32'h0004F371 , 32'h00033E43 , 32'h0004233E , 32'hFFFEED48 , 32'hFFFA93C5 , 32'h00032260} , 
{32'hFFFD15EF , 32'hFFFE4A76 , 32'h0004FBB7 , 32'h00059D5F , 32'h0004EEBC , 32'h0002BA1B , 32'hFFFF03D1 , 32'hFFFDEE1B , 32'h0000A937 , 32'h00063D6C , 32'hFFFD17F9 , 32'h0000332E , 32'h0004738A , 32'h0001CB5E , 32'hFFFE27B8 , 32'h00006688 , 32'hFFFEEF4E , 32'h00007394 , 32'h00008A20 , 32'h0000CEEB , 32'hFFFA3D3A , 32'hFFFEF7BB , 32'h00033812 , 32'hFFF7CEA9 , 32'h00044DC4 , 32'h0000C002 , 32'h00062B57 , 32'h000225CB , 32'hFFFC7E2C , 32'hFFFAD173 , 32'h00036357 , 32'hFFFB934E , 32'hFFFAC534 , 32'hFFFCA482 , 32'hFFFFD615 , 32'hFFFCC55C , 32'hFFFFBADA} , 
{32'h00375827 , 32'hFFEF6E6A , 32'h0001591E , 32'hFFF48EB3 , 32'hFFE12966 , 32'hFFF91A5A , 32'h00045CA1 , 32'hFFDB80D1 , 32'h00148D2C , 32'h000CD101 , 32'hFFD35830 , 32'hFFF59BDF , 32'hFFBC5EA9 , 32'h001DE14A , 32'hFFF5FDB8 , 32'h000E4480 , 32'h002884D1 , 32'hFFF98C7D , 32'hFFD50334 , 32'h00152E65 , 32'hFFDADBB8 , 32'h00089FEE , 32'h0015F930 , 32'h001F333A , 32'h000AB358 , 32'h000C45AE , 32'hFFFF9333 , 32'hFFD856E2 , 32'h000B389C , 32'h000317DC , 32'hFFEFD719 , 32'hFFF1BB19 , 32'h001464C5 , 32'h001FB6FF , 32'hFFD7626D , 32'h0007350C , 32'hFFF7CC48} , 
{32'hF79F2EB0 , 32'h0675B868 , 32'h043C8D88 , 32'hFFCA7DB7 , 32'h04F68210 , 32'hF58A3F10 , 32'h05D4A2E0 , 32'hFD9A5470 , 32'h0C4EF4E0 , 32'hFE8A27CC , 32'hF68B0820 , 32'h0247E1E0 , 32'h07CBC788 , 32'h01F50960 , 32'h059833B0 , 32'h0896C1F0 , 32'h0343AD08 , 32'h01A99F94 , 32'h005D75F3 , 32'hF762CD80 , 32'hFDDE01E4 , 32'hFE197478 , 32'hF720C0F0 , 32'h00E9C0F6 , 32'h00906D49 , 32'h000E4118 , 32'h0A62EFE0 , 32'hFEC9DBF8 , 32'hFEF7A908 , 32'h020608F0 , 32'hFA331610 , 32'h02D36DA4 , 32'h0C116EE0 , 32'hFCF8D3AC , 32'h0602A118 , 32'hFF4815CF , 32'hFD62443C} , 
{32'h02CE8068 , 32'h07FF8960 , 32'h05745D48 , 32'h07A83018 , 32'h046F2008 , 32'h01710344 , 32'hF48F3EC0 , 32'h022127A0 , 32'h024CB820 , 32'hFE22BEE0 , 32'h03370FC4 , 32'h077CF930 , 32'hFBE482D0 , 32'h0E96B150 , 32'hFA49F638 , 32'h02340120 , 32'h0A4180D0 , 32'hF0ED12C0 , 32'h085C3990 , 32'h0729CD48 , 32'hF9B85BE8 , 32'hF9EEC7D0 , 32'h014121F0 , 32'h0262403C , 32'hFD57DA58 , 32'h060577C0 , 32'h08978390 , 32'h06E96EF8 , 32'h04389C98 , 32'hF4CF4630 , 32'hFD646A08 , 32'hFE4DB5C8 , 32'h04957528 , 32'h003CF44A , 32'hFCBADB14 , 32'h03515AD8 , 32'hFEC126E0} , 
{32'hFBAF7968 , 32'hF3E59B80 , 32'hF8EC68C0 , 32'h0B9810A0 , 32'hFC4F61D4 , 32'hFE4BF3C0 , 32'hFD2D28EC , 32'h0701B160 , 32'h0F0FE520 , 32'hFC37A6E4 , 32'h022AEDA8 , 32'h0BAB64E0 , 32'hFD1DE8B4 , 32'hFCC0BC18 , 32'h029426EC , 32'hF3C57F80 , 32'h04398120 , 32'h02FF9F38 , 32'hF5988170 , 32'hF1669DC0 , 32'h0BE37480 , 32'h016F7150 , 32'hFDF565D0 , 32'h11CF3A80 , 32'hFF93B9F4 , 32'h08D1BC40 , 32'h11E27240 , 32'h05731FF8 , 32'h024AFE7C , 32'h02050B40 , 32'h01E961E8 , 32'hF88BDF98 , 32'hF4F03300 , 32'h06431568 , 32'hF6AF2BF0 , 32'h064CA5F0 , 32'hFAABCFE0} , 
{32'hE8241660 , 32'h03D24F44 , 32'hEC0A0360 , 32'hFFB2CD40 , 32'hFAAA3368 , 32'h4CA6F180 , 32'h0DE1FE40 , 32'h016E81B0 , 32'h59BFFF00 , 32'hAF32B580 , 32'hD9809DC0 , 32'h15723200 , 32'h13297D40 , 32'h33A7FD80 , 32'hE32A43A0 , 32'hDB0DB000 , 32'h05EAF400 , 32'h2309C080 , 32'hD0370300 , 32'h118BA780 , 32'h0EB68DB0 , 32'h00966BD4 , 32'h24749D40 , 32'h2D817780 , 32'hF5F3EEF0 , 32'hF311E330 , 32'hE3D15A20 , 32'hFAAEF730 , 32'h0359C0E8 , 32'h1C79ED20 , 32'hD5555C40 , 32'hEE87C980 , 32'hFA903228 , 32'h01589034 , 32'h1F185200 , 32'h1AD66EC0 , 32'h15DB44A0} , 
{32'h006213FD , 32'hF621D470 , 32'h0E2DD2A0 , 32'h08EF0500 , 32'h010EE4CC , 32'hE5572CC0 , 32'h03F1CD58 , 32'h0D8412C0 , 32'h0BEA6640 , 32'hE94A4040 , 32'hF84E3188 , 32'h0EB25C20 , 32'h092ED950 , 32'h0F4883F0 , 32'h02FEFC98 , 32'hF17850E0 , 32'h150BDF60 , 32'hFFC4920B , 32'hE991EA00 , 32'hFB7D8D18 , 32'hFD0BC650 , 32'hF7BB9C90 , 32'h0647FD58 , 32'h0A433880 , 32'hFC9FC5FC , 32'hF3EBD5B0 , 32'hEFAD9600 , 32'hF69C4790 , 32'hFDF6BDD0 , 32'h0BC46B30 , 32'hF9D36320 , 32'hFF4CDD52 , 32'h0D766B40 , 32'h0317575C , 32'h0EBCE940 , 32'h0815B5C0 , 32'h09D72A00} , 
{32'h0D7754A0 , 32'hF666A1F0 , 32'hFDBB167C , 32'hF3BDB4E0 , 32'hF5199300 , 32'hFD086B0C , 32'h0213B754 , 32'hFFC4B2A9 , 32'h18E01F60 , 32'h14F43380 , 32'hE6A8F080 , 32'h0E200500 , 32'hF29F5DB0 , 32'h30DB1C40 , 32'hF5AE4140 , 32'h04142850 , 32'h129D7480 , 32'h18E86D80 , 32'hDF195F00 , 32'h0E12D580 , 32'hF1DBAE20 , 32'hF055CC70 , 32'h2AFE6700 , 32'h1122A380 , 32'hFC6E7CE8 , 32'h081BE9E0 , 32'hEB836580 , 32'hE9179A20 , 32'h00248547 , 32'hF532D070 , 32'hE8400360 , 32'hFF55AE19 , 32'h0AD08060 , 32'h13029280 , 32'hE1C757E0 , 32'h0785C1D0 , 32'h0453AAF8} , 
{32'h160A07A0 , 32'h0B45F330 , 32'hEA284480 , 32'hF27D3FA0 , 32'h038CDBE8 , 32'hD95418C0 , 32'h08C62AD0 , 32'h1AF6BD40 , 32'hF198EA80 , 32'h28B11400 , 32'hFC84EE80 , 32'h0A77B1F0 , 32'hE1BFCBE0 , 32'h216E8000 , 32'hEF8DB000 , 32'hFE8E0B7C , 32'h224F4400 , 32'h08EA0EC0 , 32'hE518CE20 , 32'h188DA640 , 32'hEF2C2F80 , 32'hD4B7F6C0 , 32'h1DC624A0 , 32'hFD3D0638 , 32'hFE80B97C , 32'h0CB48430 , 32'h02B63B54 , 32'hEBEDCCE0 , 32'hE189E400 , 32'hF4D62A70 , 32'hFC8B9304 , 32'hF6FF56A0 , 32'h204A6D40 , 32'h1BDCA380 , 32'hF5AB6B30 , 32'h05465F28 , 32'h0623C1B0} , 
{32'h05FB9F00 , 32'h0C2247E0 , 32'h03DF5A8C , 32'h009FB6C3 , 32'h0CD556B0 , 32'hDA2086C0 , 32'h18CD8CC0 , 32'hE5F93380 , 32'hEBF9C780 , 32'h2903F680 , 32'h05679F00 , 32'hFE974EAC , 32'hE662A420 , 32'h00D6A183 , 32'hF743FD40 , 32'hFAB46928 , 32'h04F8F630 , 32'h036D034C , 32'hEE0C3E40 , 32'hEDDBFAA0 , 32'hE3F17780 , 32'h0542D680 , 32'h1809B800 , 32'h0756C518 , 32'h089DBFE0 , 32'h0E8246A0 , 32'h1EEF2C60 , 32'h024C02C0 , 32'hD77C4C40 , 32'h0D73F610 , 32'hF04A85B0 , 32'hF0B89AD0 , 32'hE4A15A60 , 32'h09926FD0 , 32'hF20332C0 , 32'hEDD90F00 , 32'hFE621964} , 
{32'h018B9FB0 , 32'h1D20F2C0 , 32'hE21FCFE0 , 32'h16D5F4A0 , 32'h066E0E48 , 32'hD9A75740 , 32'h09E7A310 , 32'hE7C46340 , 32'hEC023DC0 , 32'h00B01531 , 32'h043E7EC8 , 32'hD0BB2E80 , 32'hFCDDCFC0 , 32'h06B9C0C0 , 32'hF91C4338 , 32'hE38873A0 , 32'h06BBEB58 , 32'h209211C0 , 32'h0A9FF7F0 , 32'hFC5A383C , 32'h05B4E9A0 , 32'h12DFC4A0 , 32'h0BC1B000 , 32'h2785E2C0 , 32'h1B80A2C0 , 32'hDAC25BC0 , 32'h05AFB790 , 32'h146F72E0 , 32'hEDBB4860 , 32'h04A7DA88 , 32'hEFD3FFA0 , 32'hFF5EBEB5 , 32'h11AAFCE0 , 32'h19363600 , 32'hDA5C2300 , 32'hFD6C5414 , 32'h00922051} , 
{32'hEBA90640 , 32'h2B6EA9C0 , 32'h037DB8C4 , 32'h066CDF60 , 32'h1979E440 , 32'hEBC28460 , 32'h1DC26400 , 32'hE94163E0 , 32'hE4AD28E0 , 32'h16B5C720 , 32'hEC5D1AC0 , 32'hF1C55AD0 , 32'hE2991060 , 32'h11F97D00 , 32'hEFD5F160 , 32'hDB2D8040 , 32'hF707C990 , 32'h0A7CBC80 , 32'h1F261120 , 32'hEDBE5540 , 32'h0236E334 , 32'h192F26E0 , 32'h0419D3B0 , 32'h27E4AD00 , 32'h23DB9540 , 32'hDCD79D80 , 32'h0512E868 , 32'h0AA022D0 , 32'h1121C2C0 , 32'hF82C4C98 , 32'hF15A3A10 , 32'h0073FC5E , 32'h08F27810 , 32'h0B0A41B0 , 32'hD5597940 , 32'hF754AE10 , 32'hF68FB6A0} , 
{32'hE3561E60 , 32'h21F18300 , 32'hE7EF7320 , 32'h07616188 , 32'h035A9190 , 32'h2B2C9180 , 32'h17A996C0 , 32'hF48FA360 , 32'h15AD55A0 , 32'hFBCF7B30 , 32'hF9720490 , 32'hE7827E80 , 32'h118B2520 , 32'h1D02EDE0 , 32'hF2A63650 , 32'hE49E8080 , 32'hDCC0BE40 , 32'h1CB5B9C0 , 32'hFC0881FC , 32'h06D73120 , 32'hFBB31A10 , 32'h28077E00 , 32'hEFD10800 , 32'h2A9CD740 , 32'hF8BBDDF0 , 32'hFA5E3358 , 32'hFBC13928 , 32'h1E075200 , 32'h12B99E00 , 32'h06C33DF0 , 32'hFF6CBE89 , 32'hFDF4318C , 32'h19EF57C0 , 32'h0B8EFD20 , 32'hFBF9AD90 , 32'hE6D58EC0 , 32'hED2CE140} , 
{32'hF8ADCAD0 , 32'h043D0288 , 32'hFA069088 , 32'hF2BDAAF0 , 32'h0377792C , 32'h20E16980 , 32'h08272480 , 32'hEADC4400 , 32'h207DA880 , 32'h075846C8 , 32'hF4206C20 , 32'hE9DA3E80 , 32'hF71D30F0 , 32'h025525D0 , 32'h019A6878 , 32'hE880D3A0 , 32'h0244415C , 32'h02EB7CC0 , 32'h1339E000 , 32'h0A06B7C0 , 32'h07EDFC58 , 32'h118BB2C0 , 32'hF11BF470 , 32'h173418E0 , 32'h0E3219B0 , 32'hFA84EDD0 , 32'hF5657450 , 32'h09CCB750 , 32'h060804A8 , 32'h10B562A0 , 32'hFF6B3A11 , 32'h03408BF8 , 32'h0FBAB400 , 32'hFF11C8F2 , 32'h0665CCC0 , 32'hFD4343A8 , 32'hFC4CF42C} , 
{32'hEBC74540 , 32'hFF499649 , 32'h01F2F1F8 , 32'hF3591CC0 , 32'h032962A0 , 32'h0706FE48 , 32'hF5310570 , 32'h05727BB0 , 32'h02C32ECC , 32'hFAEEE110 , 32'hFE14A45C , 32'h05FB5178 , 32'hF939EF18 , 32'hF80EB7C8 , 32'hFA1510D8 , 32'h0370BC98 , 32'hFC3AAF2C , 32'h086A54D0 , 32'h01EBBBBC , 32'hF9845EC0 , 32'hFB987A78 , 32'hFCECB358 , 32'h0BB5E460 , 32'h090861E0 , 32'h00270F4A , 32'hFFAA60A2 , 32'hF86C9D90 , 32'h07325828 , 32'hFB99E710 , 32'hF556B620 , 32'hFB7E0F40 , 32'h09EAA8B0 , 32'hF73A1C80 , 32'hFE51AC98 , 32'hFCE67868 , 32'h0168FF6C , 32'h02B4FC98} , 
{32'hFEB4E9F8 , 32'hFFE9C78B , 32'hFE1F012C , 32'hFFB56C2A , 32'h001D1E74 , 32'hFE737AC4 , 32'hFF28BCF0 , 32'h02FBED0C , 32'h0066325F , 32'h0138D460 , 32'h02F18C3C , 32'h0082A77A , 32'hFDB9F2A8 , 32'h00CCD42E , 32'hFEE7984C , 32'h00942017 , 32'hFFDCEE81 , 32'hFDA40A84 , 32'h00B1084B , 32'hFF554EE5 , 32'h0210DB30 , 32'hFFD72797 , 32'hFF11CD20 , 32'hFDB91AB4 , 32'h00F654BF , 32'hFF3EE9BA , 32'h02E66258 , 32'hFD83985C , 32'hFFF9A929 , 32'hFEF35140 , 32'h02563608 , 32'h0017A15E , 32'hFC4A74D0 , 32'hFD93BA4C , 32'h0238DE08 , 32'hFF66CB7E , 32'hFD8CB95C} , 
{32'hED01BBC0 , 32'h109DBA20 , 32'hF1B75FF0 , 32'h058D1C58 , 32'h01BCFD18 , 32'h265ACB80 , 32'hFCE22F6C , 32'hF414FA80 , 32'h16C1BE60 , 32'h0C74DC80 , 32'h0386E568 , 32'h0284E5F8 , 32'h00806DC6 , 32'h02BDE56C , 32'hFCB14574 , 32'h11296380 , 32'hE757A620 , 32'hFF9A43A4 , 32'hE9449FA0 , 32'hFBB82750 , 32'hF954AD80 , 32'hEC583620 , 32'hFB0C62B8 , 32'hF95D1508 , 32'hEE450520 , 32'hFDD26164 , 32'hFE9AB7D0 , 32'hF40FFE00 , 32'h09DE8E30 , 32'h04118C18 , 32'hFBC97F08 , 32'hFBD64248 , 32'hFC852D30 , 32'h0383E764 , 32'h11460060 , 32'h046A9738 , 32'hFC8145F8} , 
{32'h04ACEB10 , 32'h0BA42B50 , 32'h09417A20 , 32'h03D04A08 , 32'hF0CA29E0 , 32'hFE3B8434 , 32'hFA0063D8 , 32'hFF067482 , 32'h00E22B88 , 32'hFD407BBC , 32'hFE57A860 , 32'hF9A33718 , 32'h04219AB8 , 32'hFC062A0C , 32'hFD393470 , 32'hFC540E5C , 32'hFFD8CA28 , 32'h06691D90 , 32'h000BD345 , 32'hFB60CC88 , 32'hFFA79882 , 32'hFFD63D0B , 32'h003F4DBB , 32'hFEA4B854 , 32'hFFFBE33C , 32'h0289D6C0 , 32'hFF4DB069 , 32'hFD6A7074 , 32'h058F19F0 , 32'hF7876930 , 32'h00F5DB4D , 32'h0102D868 , 32'hFF3A5267 , 32'h006D582A , 32'h05583000 , 32'h06F87C78 , 32'h012CC9F0} , 
{32'h000A6DC2 , 32'hFFF75217 , 32'h0003AA70 , 32'hFFEE8E2F , 32'hFFEBB832 , 32'hFFFACB16 , 32'h0019ECC1 , 32'hFFFBBFA5 , 32'h0006F60E , 32'h0001520F , 32'hFFF35944 , 32'hFFFCC6D2 , 32'hFFF56EA5 , 32'hFFFB91F0 , 32'h0000121D , 32'h0000F3B5 , 32'h0003CFBA , 32'h000775BA , 32'hFFE3E206 , 32'hFFFFA453 , 32'h00024B5D , 32'h000B7D26 , 32'h0001A457 , 32'hFFFFC3A6 , 32'h000E8C5B , 32'hFFF9C3A9 , 32'hFFF828C4 , 32'hFFEDC1CE , 32'h0001D828 , 32'h0002A03A , 32'hFFFFC57A , 32'hFFFFDE82 , 32'hFFFBC4E5 , 32'h00034FE0 , 32'hFFFC7ECC , 32'hFFFA8DDF , 32'h000091D1} , 
{32'h001AE627 , 32'h0014A687 , 32'h0052E52E , 32'h002EAC78 , 32'h0032990E , 32'h00299B15 , 32'hFFE396EE , 32'h000B5E90 , 32'h00262A18 , 32'hFFE53822 , 32'h0003A1F7 , 32'h001AF5B7 , 32'hFFEF4DA0 , 32'h0060730E , 32'hFFED384A , 32'hFFC77CD9 , 32'h003963B3 , 32'hFFA14874 , 32'h0043BF0B , 32'h002DD7FD , 32'hFFDAD5C4 , 32'hFFB086C6 , 32'h001EEF5D , 32'h0013B300 , 32'hFFEE8771 , 32'h0003C4A3 , 32'h002516F7 , 32'hFFDE9FAD , 32'h00154E5D , 32'hFFCBC48C , 32'h00161175 , 32'h000FA414 , 32'h002CF3EF , 32'h003A40AE , 32'hFFE97E50 , 32'h000BB930 , 32'hFFCD4644} , 
{32'h00029E49 , 32'h0007454D , 32'hFFF75122 , 32'h0005982C , 32'h00043593 , 32'hFFFEEA83 , 32'hFFFF80A9 , 32'hFFFD8424 , 32'hFFF81A5E , 32'h0006C4DF , 32'hFFFB45A9 , 32'h000532EA , 32'hFFFE554F , 32'h00009940 , 32'h00012517 , 32'hFFFF91A4 , 32'h00000D53 , 32'hFFFEBD7E , 32'hFFFDE096 , 32'hFFF9B9D3 , 32'hFFFC3886 , 32'hFFFF98D6 , 32'h00020D86 , 32'hFFFE7099 , 32'h00023B66 , 32'hFFFA4CF2 , 32'hFFFA8958 , 32'hFFFCB474 , 32'h0002A5EE , 32'hFFFF7469 , 32'h000499F5 , 32'h000279AC , 32'h00045604 , 32'h00076100 , 32'h0002B2A9 , 32'hFFF932C7 , 32'hFFFCF3DA} , 
{32'h000111D2 , 32'hFFFA3CF8 , 32'h0004E613 , 32'hFFF7D155 , 32'h0002B8D4 , 32'h00034661 , 32'hFFFA2C10 , 32'hFFFEB5F6 , 32'hFFFBE8D0 , 32'hFFFAD816 , 32'hFFFABF4C , 32'h0002CB39 , 32'h0000E9E3 , 32'hFFF5BA98 , 32'h00064B20 , 32'hFFFA9447 , 32'hFFFBE195 , 32'hFFFBA142 , 32'h00057705 , 32'hFFF4E831 , 32'hFFFCD6AF , 32'hFFFAD45E , 32'h0002400E , 32'h0003D423 , 32'h00058941 , 32'hFFFBD8EA , 32'h00057C81 , 32'hFFFE7FFB , 32'hFFFD3290 , 32'h00018189 , 32'h000710C2 , 32'h0007DC64 , 32'hFFFF4AA4 , 32'hFFFF34D7 , 32'hFFFFB8D5 , 32'hFFFB49C9 , 32'hFFFEEAEC} , 
{32'h0005A3E9 , 32'hFFFD5CCB , 32'hFFFF1B5F , 32'h0001180F , 32'h0001A67A , 32'h0000E200 , 32'hFFFA1852 , 32'h0004B8E0 , 32'h00015B85 , 32'h00094EED , 32'h00049592 , 32'hFFFBC004 , 32'hFFFC5ED0 , 32'hFFFF79E3 , 32'hFFF81F32 , 32'h000D9A33 , 32'h0007D286 , 32'h0004EDA5 , 32'hFFFECB52 , 32'h00052019 , 32'hFFFC9C5E , 32'hFFFD0887 , 32'hFFFF1DBC , 32'hFFF49992 , 32'h00029677 , 32'hFFFF78E9 , 32'h0000DBF4 , 32'h00000209 , 32'h0002DB50 , 32'h0003513D , 32'h0001CC6D , 32'hFFFB7AFE , 32'h0001CB96 , 32'hFFFBEB4F , 32'h0003B0BB , 32'hFFF88A37 , 32'hFFFBD64D} , 
{32'h000B0F18 , 32'h0007CEC5 , 32'hFFFDC2C3 , 32'hFFF93155 , 32'h00009A8E , 32'h0002EE47 , 32'hFFFC3703 , 32'h00023AB2 , 32'hFFF71875 , 32'h00022AD0 , 32'hFFF77F5C , 32'h00046727 , 32'hFFFF3412 , 32'h0005BB02 , 32'hFFFC9880 , 32'hFFF7DBEE , 32'h000DA686 , 32'h000A0B54 , 32'h00020ECD , 32'h000174BC , 32'hFFFFD5CB , 32'h00052848 , 32'hFFFF26F0 , 32'h000070D5 , 32'hFFFEE087 , 32'h00000242 , 32'h0001A9CF , 32'hFFFE82BF , 32'hFFFD8ABA , 32'h000122E5 , 32'hFFFAD1F6 , 32'hFFFDFF16 , 32'hFFF7F568 , 32'h000263D5 , 32'h00004DBD , 32'hFFFA5048 , 32'hFFF8D3AA} , 
{32'hFFFA7C04 , 32'h0009934E , 32'h0004ABD8 , 32'h00011E8E , 32'hFFFEEDF5 , 32'hFFFBE541 , 32'h00037370 , 32'h00047BD2 , 32'hFFFEF5F7 , 32'h00006297 , 32'h00009F94 , 32'hFFFFF4C9 , 32'h0007F13E , 32'h0002F17D , 32'hFFFEB8F9 , 32'hFFFEF82D , 32'hFFFDEAD9 , 32'h0000E634 , 32'h0001D224 , 32'hFFFEE62D , 32'h000C438E , 32'hFFFBCB6D , 32'h00007FA9 , 32'h0005C979 , 32'hFFFF5B46 , 32'h00023192 , 32'h0002C7C5 , 32'hFFF7995C , 32'hFFFF49A9 , 32'h0002E02C , 32'hFFF703EC , 32'hFFFC6EA6 , 32'h0003F0C3 , 32'hFFFC6FB0 , 32'h0006A47C , 32'hFFFCD154 , 32'h000097B9} , 
{32'h00078475 , 32'hFFFFC103 , 32'hFFFA72F7 , 32'hFFFD2399 , 32'hFFFDAA52 , 32'hFFFCB580 , 32'hFFFFB303 , 32'h00073610 , 32'hFFF4FFBB , 32'hFFFCA115 , 32'hFFFB8624 , 32'h000006C8 , 32'hFFFD2502 , 32'hFFFDBBB8 , 32'hFFFEC828 , 32'hFFFF0550 , 32'h00025152 , 32'h00059D6B , 32'hFFFAAFA1 , 32'hFFF62A0B , 32'h00086B21 , 32'h0008364B , 32'h00087B7C , 32'h00015027 , 32'h0007464F , 32'hFFFE9831 , 32'hFFFD9CBB , 32'hFFFE7794 , 32'h0004809B , 32'h00001A31 , 32'h0000B08E , 32'h0000A0C2 , 32'h0004DF18 , 32'h00043C57 , 32'h00050201 , 32'h00071BBC , 32'h000235E4} , 
{32'h000814C3 , 32'h0000CEF3 , 32'h0000D957 , 32'h00049F90 , 32'h00019313 , 32'h00080A3B , 32'h0002BC1B , 32'hFFF577ED , 32'h00038573 , 32'hFFFC8C04 , 32'h000A421E , 32'hFFFBCE70 , 32'hFFFEE5D6 , 32'hFFFE5C25 , 32'h00046860 , 32'hFFF54DF3 , 32'h0004C903 , 32'hFFFE6580 , 32'hFFFEC928 , 32'hFFF51B41 , 32'h00039D53 , 32'hFFFD63EF , 32'hFFFDFC42 , 32'h0002F498 , 32'hFFFCFEDF , 32'h00015CA7 , 32'hFFF8A61E , 32'h00016A90 , 32'h00050E7F , 32'h0003BAA0 , 32'h0003D9FD , 32'h000770C7 , 32'hFFFCA568 , 32'h000030D5 , 32'h00005406 , 32'h0001D692 , 32'h00049F38} , 
{32'hFF8E778E , 32'h005F0134 , 32'hFFB45430 , 32'h003DC92E , 32'h00080090 , 32'h003A55E7 , 32'hFFFA9F37 , 32'h0001AFCF , 32'h000160AB , 32'h002BC717 , 32'hFFD3BA2E , 32'hFFD921A5 , 32'hFFF5BD65 , 32'hFFDC5D3E , 32'hFFE23ABB , 32'hFFFBE8C4 , 32'hFFD6A4A4 , 32'hFFF62D0D , 32'hFFD85408 , 32'hFFFE88F4 , 32'hFFCD2B83 , 32'h001AED45 , 32'hFFEDB6FE , 32'h00001797 , 32'hFFFA35B2 , 32'hFFD4B467 , 32'hFFF24F83 , 32'hFFF360FB , 32'h00414CD3 , 32'hFFEA7F02 , 32'hFFF649C9 , 32'hFFE3C238 , 32'h001131FD , 32'h002ACF23 , 32'h00015160 , 32'h0020E45E , 32'hFFE8C204} , 
{32'hF28C2140 , 32'h0A7FF3F0 , 32'h03F4B7C8 , 32'h01C5949C , 32'h073D5360 , 32'hF0C11950 , 32'h09A07D10 , 32'hFDB88CF0 , 32'h136BACA0 , 32'hFD58DDBC , 32'hF0D6CF40 , 32'h027CC1A8 , 32'h09C2D570 , 32'h0350F8E8 , 32'h0A19C390 , 32'h0D6CB510 , 32'h00DE8B80 , 32'h056173E8 , 32'h0136864C , 32'hF0F4AB80 , 32'hFADFDE90 , 32'hFA84DC98 , 32'hF2E6AC20 , 32'h00F4EBA2 , 32'hFDBD3D04 , 32'hFEDABED0 , 32'h0DF35B90 , 32'hFDC93E4C , 32'hFEC95A54 , 32'h051504B0 , 32'hF7DCCE90 , 32'h05DCAA38 , 32'h1250E1C0 , 32'hFC034590 , 32'h0847C080 , 32'hFC385678 , 32'hFD5828D4} , 
{32'hFFA42A98 , 32'h00E4D13D , 32'hFDE5736C , 32'h0204D268 , 32'hFFB6BD69 , 32'h000001FF , 32'h012314F8 , 32'h00DE31D3 , 32'h0170983C , 32'hFF795375 , 32'hFE231B28 , 32'hFE941038 , 32'hFD79D5AC , 32'h00B7902A , 32'h01B47680 , 32'h00D5039A , 32'hFD2C3364 , 32'h0239A1C4 , 32'h00B04DCF , 32'hFE1410D0 , 32'hFDAAAE10 , 32'hFE080A88 , 32'h005060C9 , 32'h0036FF34 , 32'hFD847984 , 32'hFEDE3FC4 , 32'hFEAB3B94 , 32'hFEE58BE0 , 32'h00413A54 , 32'h01D6C9C4 , 32'hFFECE6F1 , 32'h018CFCF8 , 32'h00DBC040 , 32'h00D1FAEE , 32'hFEDDD900 , 32'hFE12FD00 , 32'h01071328} , 
{32'hF0A3FA70 , 32'h083EC1F0 , 32'h045A4A28 , 32'h0FB93960 , 32'h006E5843 , 32'hEE55FC80 , 32'h0FBB6FE0 , 32'h01CADB74 , 32'h0398DE98 , 32'hE61DA820 , 32'hE6800820 , 32'h0D9FDC90 , 32'h19688B40 , 32'h08D5EA90 , 32'h10293E40 , 32'h13897680 , 32'hFFE51B91 , 32'h03E57368 , 32'hF740FFD0 , 32'hF3132D00 , 32'hF669D1E0 , 32'hF9ED4158 , 32'h0181F85C , 32'h0C349890 , 32'h0086DDA1 , 32'h0CF8E9F0 , 32'h11A2A0E0 , 32'hF95F88A8 , 32'hF8527228 , 32'hF8B48BA0 , 32'hFD49BD60 , 32'h0D033640 , 32'h0BFC18B0 , 32'hF01ED190 , 32'h0256B8EC , 32'hFB3F0100 , 32'hF6403B20} , 
{32'hE9EF4680 , 32'h0F9E3690 , 32'h04C9B130 , 32'hF7C296B0 , 32'h00ED1758 , 32'hEC8195C0 , 32'h084F66D0 , 32'h012372FC , 32'h1671D660 , 32'h00409F5A , 32'hDDCF7280 , 32'h04F6E9E0 , 32'h098B7CA0 , 32'h04377950 , 32'hFE752BD8 , 32'hF5F81D10 , 32'h0B906B50 , 32'hFEBBFE00 , 32'h0301EA5C , 32'h0D7DD750 , 32'hFC48A328 , 32'hFDC8E488 , 32'h0587CE28 , 32'hFF3A818B , 32'hF69CD720 , 32'hF5E7FEE0 , 32'h0AC54030 , 32'hE4F51BA0 , 32'h05191C60 , 32'h0EDF9110 , 32'hF56BAE70 , 32'hEEBE0CA0 , 32'hFA2DB0F8 , 32'hFA062A28 , 32'hFB894C98 , 32'h09859820 , 32'h02FF974C} , 
{32'h02BB97AC , 32'hFF2337E3 , 32'hFB4EC028 , 32'hFB6F0D68 , 32'hFE8C3C40 , 32'h18AEFF00 , 32'hFF7417F9 , 32'hFAEAB948 , 32'h1991F3A0 , 32'hFAED75A0 , 32'h0049E154 , 32'h033FA79C , 32'h056DA978 , 32'h070C6CF0 , 32'hFAF64F40 , 32'h0727B058 , 32'hF5210920 , 32'hFBC4E850 , 32'hF4543110 , 32'h09966630 , 32'h028943D8 , 32'hF9D17B68 , 32'hFEC68484 , 32'hF7C595C0 , 32'hF85EE748 , 32'hF9073D68 , 32'h019A9908 , 32'hFB4CCD38 , 32'hFCFBB614 , 32'h070F86D0 , 32'hF615FBB0 , 32'hF74A6B30 , 32'hFD43B464 , 32'h040E0530 , 32'h13C42280 , 32'h094DCBF0 , 32'hFFE0B316} , 
{32'hF295B590 , 32'h0A478260 , 32'hF506D840 , 32'h01E18D14 , 32'hFE0640B0 , 32'h1DD564E0 , 32'hF7D4CBC0 , 32'h00F7C4D0 , 32'h0EB73910 , 32'h05337B58 , 32'hFDDAC37C , 32'h07396470 , 32'hFF45366D , 32'h00199E79 , 32'hFC229E50 , 32'h04467528 , 32'hED595800 , 32'hF9353E10 , 32'hEC302D20 , 32'hF4646F00 , 32'hFA4E1138 , 32'hF0B300E0 , 32'hF6572400 , 32'hF3F64120 , 32'hFA663980 , 32'hF3F24D10 , 32'h013E12AC , 32'hFF6FD1A2 , 32'h04859618 , 32'hFD3D1A80 , 32'hFE75EA44 , 32'hF8B09388 , 32'h00B21934 , 32'h1004CEE0 , 32'h0B642A90 , 32'h00E0F629 , 32'hFA82C490} , 
{32'hE99D1BE0 , 32'h1E3859C0 , 32'hF686A1E0 , 32'hEF0384A0 , 32'h060E81B8 , 32'hEDB1BB20 , 32'hF7B77330 , 32'h0FC4BB50 , 32'h19F40540 , 32'hF5265D50 , 32'hE6989260 , 32'hF8D34758 , 32'h0B1DDDD0 , 32'h07DDE898 , 32'h1BF3E960 , 32'h0B1A4710 , 32'h0E08BA70 , 32'h02828A7C , 32'hFB207FC8 , 32'hF8BFD3A0 , 32'hFC0FC880 , 32'h025598E0 , 32'h1D4047E0 , 32'hFCB7ED3C , 32'hF61E0810 , 32'h03789164 , 32'hED875060 , 32'hF1860A00 , 32'hEF455020 , 32'h09CE97F0 , 32'hF1F30D70 , 32'hFAC839B8 , 32'h00644A7D , 32'h0167B598 , 32'hE907AFA0 , 32'h14A3E5E0 , 32'hFF18788D} , 
{32'hF4F58700 , 32'h104E3CC0 , 32'h04620C38 , 32'hF4773C50 , 32'hF83B1758 , 32'hD0C23840 , 32'h174AB9A0 , 32'h0ADE3F20 , 32'h1CE85C40 , 32'h281B03C0 , 32'hE5C34D40 , 32'h11A61980 , 32'h2150FEC0 , 32'h31B3DA40 , 32'h1016E020 , 32'h11FC18E0 , 32'h2C5AC7C0 , 32'h0E48B190 , 32'hF9D15810 , 32'hF7680310 , 32'hFB8764C0 , 32'h06AD4800 , 32'h19E245A0 , 32'hCB9AA780 , 32'h0A9A2640 , 32'hD2EA2480 , 32'h21133480 , 32'hCA1B1780 , 32'h0D364810 , 32'hF6E337F0 , 32'h13EE9F60 , 32'hF8A113E8 , 32'hE710A3E0 , 32'h070DE230 , 32'hF9221E50 , 32'h13D536E0 , 32'h05021AC0} , 
{32'hF17C7630 , 32'h1F7E7AC0 , 32'h1E6EC980 , 32'h0E53F790 , 32'hFF63A360 , 32'hCD784E40 , 32'h26F26700 , 32'h0CBC2440 , 32'h07F1EBE0 , 32'h0DA8D690 , 32'hDF738C00 , 32'hFEF4E494 , 32'h21933340 , 32'h31F6F180 , 32'h04D9F738 , 32'h014DCB24 , 32'h10B1A4C0 , 32'h1472F640 , 32'hFA3873F8 , 32'hD861B040 , 32'hE8026E00 , 32'h0BB8AB70 , 32'h0F89AAF0 , 32'hF0AB4290 , 32'h21D08400 , 32'hDD9B1640 , 32'h24140240 , 32'h16399720 , 32'hFB103A58 , 32'h189799A0 , 32'h2B6A0800 , 32'hFAC16A00 , 32'hE9AA71E0 , 32'hFE58776C , 32'hD6C27900 , 32'hEF9B1000 , 32'h09FF9E30} , 
{32'hE41626E0 , 32'h0D25ECA0 , 32'h05B2A768 , 32'h02850358 , 32'h02166034 , 32'hE4ECD4C0 , 32'h0F955F40 , 32'hFB458418 , 32'hE7405860 , 32'hFFB12A82 , 32'hFF23302B , 32'h009648A1 , 32'hFF614B17 , 32'h1AF583C0 , 32'h0A2980E0 , 32'hE7AB2B20 , 32'h0E62F030 , 32'h0BE90130 , 32'hFA757E08 , 32'hEF177680 , 32'hF73C6EA0 , 32'h007A8C34 , 32'h13B5EB20 , 32'hE2FD1320 , 32'h327BAF00 , 32'hF1A3A130 , 32'h0604A5C8 , 32'h1D382DE0 , 32'hF6C77400 , 32'hFD45B7D0 , 32'h0F81CED0 , 32'hE5B879E0 , 32'h076D9D88 , 32'h0368B928 , 32'hD720CE40 , 32'h0832D6D0 , 32'hFB2E3F60} , 
{32'hED74E2C0 , 32'h00F7ABE5 , 32'h0824AC20 , 32'h12F62D80 , 32'hF872DFA0 , 32'hC78C1F80 , 32'h12C02A60 , 32'h17543F00 , 32'hE24142E0 , 32'hE8D21660 , 32'hF1AC0F50 , 32'h05F16FB0 , 32'hF2C8FF10 , 32'h2AB394C0 , 32'hFE421298 , 32'hEBCA6D20 , 32'h13848820 , 32'h134F6420 , 32'h0A73C6D0 , 32'hE0BD5DA0 , 32'hFBCBF1F0 , 32'h02546EE4 , 32'h121D6C40 , 32'hF31505F0 , 32'h324CF7C0 , 32'hE8440A40 , 32'hF1095B30 , 32'h3249F780 , 32'hFCCEC760 , 32'h0618E2D0 , 32'h202AE200 , 32'hE8804740 , 32'h076410F8 , 32'hF79106E0 , 32'hE1E121C0 , 32'h14888000 , 32'h046BE2E8} , 
{32'hC9ED26C0 , 32'h1CD4ECE0 , 32'hF11CE390 , 32'hF1F5C040 , 32'hF2E3E070 , 32'hF3693660 , 32'h093D1FF0 , 32'h1335B800 , 32'h069745A8 , 32'h2098E740 , 32'hFC58770C , 32'hFA5CF1F0 , 32'hE8A298A0 , 32'h3A560000 , 32'hFCF9F3E4 , 32'hFD5DD938 , 32'hE56EDC40 , 32'h13EFB780 , 32'hF6137B00 , 32'hE57CBF80 , 32'hF5CA9F20 , 32'h09A5D110 , 32'h03AFB998 , 32'hFCEDD51C , 32'h19ECD520 , 32'hEFAAFE20 , 32'hDBE41240 , 32'h149B6440 , 32'hFC515348 , 32'hDF075E80 , 32'h07BE3EC8 , 32'hFBCC5558 , 32'h0222A33C , 32'hF8B84168 , 32'hF7532A30 , 32'h247D5C80 , 32'h0E330710} , 
{32'hC632D080 , 32'h275096C0 , 32'hE6D39FE0 , 32'h027ADD04 , 32'h00D73BC4 , 32'h160A1DA0 , 32'h25CC1A00 , 32'hF44E1E40 , 32'h35445580 , 32'h00E27057 , 32'hE16D57A0 , 32'hF1091120 , 32'h1EC3BC40 , 32'h29400940 , 32'hFB2C4568 , 32'hEA0CB5A0 , 32'hE8BE1AC0 , 32'h1D3A01E0 , 32'hF3C2BD60 , 32'hF8D7B418 , 32'h093E99D0 , 32'h21E50440 , 32'hF315B1E0 , 32'hF87302E8 , 32'h1ABCCE40 , 32'hFB682D20 , 32'hF9F006C0 , 32'h0EF479C0 , 32'h18109E60 , 32'h0C92C2C0 , 32'h2B9D75C0 , 32'h132D8860 , 32'h0E70DCD0 , 32'hEAD82E80 , 32'h0E8773D0 , 32'hF1F50DA0 , 32'h024FC1DC} , 
{32'hE794E4E0 , 32'h121AD6C0 , 32'hD8A0A280 , 32'hE94A6140 , 32'hF3583520 , 32'h1F4E0A80 , 32'hF9AFED38 , 32'hEBCC0100 , 32'h162A4320 , 32'h3E3CB700 , 32'hE50279C0 , 32'hC8B7E740 , 32'hE54892C0 , 32'h12D2E0C0 , 32'hF03EB660 , 32'h15FBD500 , 32'hDA380A40 , 32'h12EFD1E0 , 32'h3A48DE40 , 32'hFDBCC220 , 32'hFA6B1A78 , 32'h48B3F880 , 32'hDA6950C0 , 32'h14ED6280 , 32'h1365A080 , 32'h2B3A53C0 , 32'h1B764A60 , 32'h144D26A0 , 32'h1A76BF60 , 32'hDF66BD00 , 32'h04DA4DD8 , 32'h0816DD40 , 32'hE9D83D60 , 32'hFF18C50A , 32'hF669F460 , 32'hF8F1F030 , 32'h14CCF8A0} , 
{32'hD327B640 , 32'hFC3E9538 , 32'hC82345C0 , 32'hF774DDA0 , 32'hDF285A80 , 32'hF1DE2B30 , 32'h10AC0060 , 32'h01EF5750 , 32'h004E3EA7 , 32'h0F698480 , 32'h0E8060B0 , 32'h0946A2B0 , 32'h0352AAD4 , 32'h162A6860 , 32'h04039B68 , 32'hF0EB88A0 , 32'h12485320 , 32'hEDB64400 , 32'h16CF1540 , 32'h0DDD4D30 , 32'h04510CF0 , 32'h12744D60 , 32'hFB22F6A8 , 32'hFCA719C4 , 32'h038DA01C , 32'h0A1BCE60 , 32'hFCF6C898 , 32'hE73EF120 , 32'h1A667A60 , 32'hEC937DA0 , 32'h17C55420 , 32'h2E5CE740 , 32'hDF4E2EC0 , 32'h0AA4AB80 , 32'h0095B6E3 , 32'hFED7DA84 , 32'hF89FA4A0} , 
{32'hF4AE7F20 , 32'h067A8FF0 , 32'h05787B48 , 32'hF874FD90 , 32'h16911840 , 32'hFCC211A4 , 32'hEFB5FFE0 , 32'h02FC15D4 , 32'h07579410 , 32'h27C97CC0 , 32'h09F7BF80 , 32'hF246C5B0 , 32'hF5503D00 , 32'hFDE5FBD0 , 32'hF6523C50 , 32'hF8769BB8 , 32'h08E32D40 , 32'h07AA1080 , 32'h08F85BD0 , 32'hFC9C4278 , 32'hF5DF42A0 , 32'h070EF978 , 32'hD616C540 , 32'h0305D76C , 32'hFCBB36DC , 32'h0CC3A510 , 32'hF4C0C360 , 32'hF6B59590 , 32'hF57045B0 , 32'h171DF640 , 32'h0DE32490 , 32'h0A58CDA0 , 32'hEF17AAC0 , 32'h0303A834 , 32'h0036D0D5 , 32'h084011B0 , 32'h0DBFDBB0} , 
{32'hF48BA580 , 32'h0AAC90A0 , 32'hF9C38CE8 , 32'hEF65B260 , 32'h0048E6B5 , 32'hFC60908C , 32'hFA1215A0 , 32'h064CBF38 , 32'h05A3AB40 , 32'h1C456DA0 , 32'h0F42DB90 , 32'hF4DDC630 , 32'hDD1BCBC0 , 32'hFDEC0A2C , 32'h01B3A898 , 32'h03D722DC , 32'hEF817320 , 32'h01F9F6D0 , 32'h19DDD520 , 32'hF1BED450 , 32'h14386FA0 , 32'hFB93A978 , 32'hE8CE6C60 , 32'hFBEFB758 , 32'h00C43851 , 32'hFB9A9CE8 , 32'hFAC13FF8 , 32'h09F73A60 , 32'hFB3B7478 , 32'h001E329E , 32'hF8A15780 , 32'hF81D4538 , 32'hF2A86B50 , 32'hFD197098 , 32'h0C9917E0 , 32'h168A5E20 , 32'hFDCDC1A4} , 
{32'h000C26C2 , 32'h00768C81 , 32'hFFE2DA59 , 32'h0019B750 , 32'h0027169C , 32'h000EFFD0 , 32'hFFB6E190 , 32'h000ED820 , 32'h00175118 , 32'hFFFAC5B4 , 32'h0002FBEF , 32'h00881684 , 32'hFF5C464D , 32'h00A483C7 , 32'hFFC341A2 , 32'h0004F480 , 32'h00E3A184 , 32'hFF2433EA , 32'h003E769E , 32'h009329EE , 32'hFFD174F9 , 32'hFFF98466 , 32'h00272D96 , 32'h0048CC77 , 32'h00647B59 , 32'h00AD3CBE , 32'h004D64C7 , 32'hFF8F1193 , 32'h00461E1E , 32'hFF69C612 , 32'h003F6740 , 32'h005CC7A6 , 32'h00470F75 , 32'h000EEEC1 , 32'hFFD30519 , 32'h00667955 , 32'hFF859CB7} , 
{32'hEF80E580 , 32'h0E823330 , 32'hFCA69178 , 32'h0766CC28 , 32'hFCEDE608 , 32'h06AE9418 , 32'hFB3469C8 , 32'hFBAFC9D0 , 32'hF9C08BF8 , 32'hF799D280 , 32'h076A0B60 , 32'hFBE63380 , 32'hF9883B28 , 32'hEE599800 , 32'hF79351E0 , 32'h04EF0050 , 32'hF9E2C860 , 32'h00BF1039 , 32'h09F18770 , 32'hFDD0856C , 32'h074FC358 , 32'hF4FAD2C0 , 32'hFE885AE4 , 32'hFE006604 , 32'h008D8AAF , 32'h05BE0AA8 , 32'h005B7653 , 32'h0E1E2370 , 32'hF914DAC0 , 32'h0389D02C , 32'h0186ADBC , 32'h07EC8030 , 32'hFAB1DE88 , 32'hF927C098 , 32'h019F027C , 32'h03B8BCD4 , 32'hFBB1CEC8} , 
{32'h002B7E6F , 32'hFFE0B93C , 32'h00600613 , 32'h00707663 , 32'h003C3CFE , 32'h003D19B3 , 32'hFFD37B2E , 32'hFFEE4F37 , 32'h000A431A , 32'hFFF46D22 , 32'h00194827 , 32'hFFA91B97 , 32'hFFFDF6F3 , 32'h008A0206 , 32'hFFDE4A87 , 32'h0006A089 , 32'h00A8FECA , 32'h0009BDDC , 32'h000BD087 , 32'h0060919E , 32'hFF722EE5 , 32'hFF9BB8D5 , 32'hFF642C08 , 32'h0024B6CF , 32'h00108A8E , 32'h00197950 , 32'hFFC75DBA , 32'hFF9948FF , 32'h0005BD4A , 32'hFF528BC7 , 32'hFFCF787C , 32'hFFC4E48B , 32'hFFEEC7C0 , 32'h001FF4BF , 32'hFFAB6D9C , 32'h0056B10F , 32'h003C14AC} , 
{32'h0010D851 , 32'hFFFA1D1A , 32'h0005643B , 32'hFFFD7E54 , 32'h000575EF , 32'h000B5993 , 32'h000AED7F , 32'hFFDF3724 , 32'h000DBA45 , 32'hFFFF48FF , 32'hFFEB66F9 , 32'hFFE978C9 , 32'hFFE70ACD , 32'h0002C5AC , 32'hFFE98AB9 , 32'hFFFDC029 , 32'h0013D5A8 , 32'h000003BB , 32'h00029684 , 32'hFFFE0318 , 32'hFFF8EC3D , 32'h000696CA , 32'h000DE92F , 32'h000A1DC4 , 32'h0001551D , 32'hFFEEA3BA , 32'h0005F53B , 32'hFFEA7CC4 , 32'h000397AF , 32'h00003679 , 32'hFFF63617 , 32'hFFFA92AB , 32'h00051FF4 , 32'h000D1C67 , 32'hFFFCD84C , 32'hFFFA0860 , 32'h0004AFD7} , 
{32'hFFFEC378 , 32'hFFF88961 , 32'hFFFEA1FB , 32'hFFFF2DE5 , 32'h00087A23 , 32'hFFFEA8F0 , 32'h00006D08 , 32'hFFFD6F72 , 32'h00011BB1 , 32'hFFFA55FC , 32'hFFF97EA3 , 32'hFFFDE0B5 , 32'hFFFC7FC0 , 32'hFFFB37E1 , 32'h0001FBBA , 32'h00059ECB , 32'hFFFE94A9 , 32'hFFFB13F6 , 32'h00084FC1 , 32'hFFFDB2CD , 32'h00040C8D , 32'h0008EFF3 , 32'h00071E4D , 32'hFFF7A470 , 32'h00030001 , 32'hFFFF9BDC , 32'h000CAADB , 32'hFFFC41AC , 32'hFFFE9C5C , 32'hFFFA6B05 , 32'hFFF74506 , 32'h0002BF4A , 32'h00025B4F , 32'hFFFE8E1D , 32'h000298E8 , 32'hFFFC1EF5 , 32'h00043D17} , 
{32'hFFFB822C , 32'hFFFCF643 , 32'hFFFFEF99 , 32'h00002921 , 32'hFFFA7107 , 32'h000461F3 , 32'h0004EE4C , 32'hFFFD24D8 , 32'hFFF773F4 , 32'hFFFB949C , 32'h00003A78 , 32'h00025295 , 32'hFFFC1BB8 , 32'h00036644 , 32'h0003990E , 32'hFFFC2B82 , 32'hFFF87EB6 , 32'hFFFE0BD3 , 32'hFFF91357 , 32'hFFFF5BB5 , 32'h00039707 , 32'hFFF6F17D , 32'h00054830 , 32'hFFFB17D3 , 32'h000A9F9B , 32'hFFFEBAA4 , 32'hFFFA2EE6 , 32'hFFFFB3CC , 32'hFFFAE5CB , 32'hFFFCA104 , 32'h0001C254 , 32'h000107ED , 32'hFFFD9E60 , 32'hFFF6D8B9 , 32'hFFF76679 , 32'h0004BB6C , 32'hFFFA9112} , 
{32'h00038CA9 , 32'h000407E7 , 32'h0003DE88 , 32'hFFFF3B50 , 32'hFFF95A66 , 32'hFFFC7906 , 32'hFFFC3545 , 32'hFFFD5380 , 32'hFFFB692A , 32'h00010D8C , 32'hFFFE1129 , 32'hFFFF8203 , 32'h0007A6EE , 32'hFFFDD948 , 32'h000A2FD8 , 32'hFFFFC1F5 , 32'h000069C8 , 32'h000B2542 , 32'h0006A4F8 , 32'hFFFB7DAD , 32'hFFF781FB , 32'hFFFCA976 , 32'hFFFFD992 , 32'h000188B2 , 32'hFFFF8D96 , 32'h00023CB0 , 32'h0000F9B8 , 32'h0004263D , 32'hFFFD18BB , 32'hFFFE25B1 , 32'hFFFE33B5 , 32'hFFFBC769 , 32'hFFFD275B , 32'h0004B01E , 32'hFFFE3A61 , 32'h00070710 , 32'h00001ED0} , 
{32'hFFFF7BCE , 32'hFFF53DB2 , 32'hFFF9D093 , 32'h00045EB3 , 32'h0000C84F , 32'hFFFD79B8 , 32'hFFF581CD , 32'hFFFD63DF , 32'h0005DD37 , 32'h0000513A , 32'h00042395 , 32'h0005A405 , 32'hFFFD1032 , 32'h0006BDF5 , 32'hFFF99DDC , 32'hFFFE7DAF , 32'h0002B3D2 , 32'h0005197A , 32'h0003EF81 , 32'hFFF95F54 , 32'h0006163F , 32'hFFFC6076 , 32'h00044DCE , 32'h00016C84 , 32'h0001B807 , 32'hFFFBAA70 , 32'h00042FDF , 32'hFFFF05F7 , 32'hFFF8EE3C , 32'h000E966E , 32'h000007F1 , 32'h00020F80 , 32'hFFFB5239 , 32'hFFFCCB7B , 32'hFFFF1EB8 , 32'hFFFC3B30 , 32'h000553F8} , 
{32'hFFFD5005 , 32'h00009517 , 32'hFFFBD393 , 32'hFFFF8615 , 32'hFFF8C6B3 , 32'hFFFAE5AF , 32'hFFFAEDDD , 32'hFFFE1687 , 32'hFFFFC058 , 32'hFFFA6558 , 32'hFFF855C6 , 32'h000137C0 , 32'h0005EDC9 , 32'hFFF7381D , 32'hFFFCD9AC , 32'hFFFCE7FA , 32'hFFFEA958 , 32'hFFFAC840 , 32'h0002B191 , 32'h00012A12 , 32'hFFFFED08 , 32'h0004032F , 32'h00047A73 , 32'hFFF1FAC3 , 32'h000410FF , 32'h000108AE , 32'hFFFB182F , 32'hFFFEC918 , 32'h0000D588 , 32'h0000DAE2 , 32'h00022BCC , 32'h0000A606 , 32'hFFF661BB , 32'hFFFDB505 , 32'hFFFFC1E5 , 32'hFFF6EB2F , 32'h0001D678} , 
{32'h0004A857 , 32'hFFFACAC9 , 32'hFFF83706 , 32'h00010AF3 , 32'hFFF912B1 , 32'h000324AA , 32'hFFFAA8D2 , 32'h000100D5 , 32'h00029409 , 32'hFFFCBABF , 32'h0007D9C9 , 32'hFFFBA564 , 32'hFFFBD494 , 32'hFFFDD850 , 32'hFFF9C0DC , 32'hFFFA2692 , 32'h00036E02 , 32'h0002E613 , 32'hFFFF35B6 , 32'hFFFD45A9 , 32'h0002FBBB , 32'h0000101A , 32'hFFFFBA84 , 32'hFFFE85BD , 32'hFFF9E662 , 32'hFFF96692 , 32'hFFFB0FDA , 32'hFFFE3D9C , 32'h0002A8C0 , 32'hFFF89F0E , 32'hFFFE73E3 , 32'hFFFD4E2E , 32'hFFFE36D9 , 32'h00021527 , 32'h00003BDF , 32'h00078D91 , 32'h000820CE} , 
{32'hFFF76434 , 32'h001B26DD , 32'h00053040 , 32'h00072C26 , 32'h000123F1 , 32'h0013CEA1 , 32'hFFFA0E6F , 32'h000057C4 , 32'hFFFD1CD5 , 32'h000014F4 , 32'h0009DCC6 , 32'h000B7579 , 32'hFFFC94FF , 32'hFFFC888C , 32'hFFF8AAC0 , 32'h00041EA2 , 32'h000417B5 , 32'hFFFF8873 , 32'hFFF1134E , 32'hFFF8751E , 32'h00012217 , 32'h0007F4A8 , 32'hFFFE59AE , 32'hFFFA372D , 32'hFFF507F5 , 32'hFFFD6D8B , 32'hFFFBDF25 , 32'h00026CBE , 32'h0002DCD2 , 32'hFFF6BEBB , 32'hFFF9B603 , 32'h00019EBC , 32'h00065865 , 32'h000AF0A5 , 32'hFFFA7BA3 , 32'hFFF181E7 , 32'hFFF6CB68} , 
{32'hF328F1D0 , 32'h09D415C0 , 32'h0453F370 , 32'h016462B4 , 32'h06F694C8 , 32'hF11A7A50 , 32'h09268490 , 32'hFE10CCD0 , 32'h126A58E0 , 32'hFD9CACE4 , 32'hF1694C00 , 32'h029B4A00 , 32'h09924A10 , 32'h031C3B14 , 32'h0994D910 , 32'h0C73E6B0 , 32'h01C0C908 , 32'h04A10A08 , 32'h01234504 , 32'hF20947C0 , 32'hFBA19090 , 32'hFB42DCD0 , 32'hF2F46FD0 , 32'h00E8D147 , 32'hFE590C78 , 32'hFEC401F4 , 32'h0D94A060 , 32'hFE1691D0 , 32'hFED36EEC , 32'h0468ABF8 , 32'hF8153D00 , 32'h058A4660 , 32'h11A5A620 , 32'hFBCBAAE8 , 32'h0849C600 , 32'hFCA0D2EC , 32'hFCFBF6F0} , 
{32'hF13C1F80 , 32'h06877DE8 , 32'h07409068 , 32'h025027C0 , 32'h09E977C0 , 32'hF8C5A058 , 32'h030B4EA0 , 32'hFFE3AABE , 32'h109BD240 , 32'hFFBB55BE , 32'hEDED4440 , 32'hF91BCFE0 , 32'h06B040F8 , 32'h0423EED0 , 32'h0BD5E500 , 32'h0D01A2F0 , 32'h07868490 , 32'hFF6899AA , 32'h02AC8F84 , 32'hF1D52870 , 32'h09C42B50 , 32'hFC2398B0 , 32'hF8326E28 , 32'h029F2C48 , 32'h032261C0 , 32'hFDC638DC , 32'h02BCF4CC , 32'h00035BA3 , 32'hFCC34AE0 , 32'hFF0C3EFD , 32'hFDD417C4 , 32'h09DB0290 , 32'h0F369900 , 32'h08517370 , 32'h0894F710 , 32'hFD34B69C , 32'h06153440} , 
{32'hEDB43FE0 , 32'h04715E40 , 32'hF37A2430 , 32'hFECA3D94 , 32'h120357A0 , 32'h24C53800 , 32'h1095F580 , 32'hEE93E680 , 32'h4734CF00 , 32'hFB153D18 , 32'hEE27D6C0 , 32'h05D50BF0 , 32'h11F55160 , 32'h1A2F7FC0 , 32'h035E863C , 32'h1C8243C0 , 32'hE7E10A00 , 32'h08B31BF0 , 32'hF0E2B8F0 , 32'hF3FA47C0 , 32'h01EC4754 , 32'hF0D90EB0 , 32'hEABE18C0 , 32'hFDF86C9C , 32'hFDE03F98 , 32'h0AA68A80 , 32'h0AD99150 , 32'h058430A0 , 32'hFEFFB134 , 32'h13CB8BC0 , 32'h010A41CC , 32'h00EAC22E , 32'h12AC3820 , 32'hF4B78770 , 32'h10C9CB80 , 32'hFA0A1EE0 , 32'hF5977A20} , 
{32'hFF16A49C , 32'h0C04EFC0 , 32'hF0AF7A10 , 32'hF76661A0 , 32'hFC4D3E68 , 32'h46E15700 , 32'h0E4D1A60 , 32'hE2C979E0 , 32'h3E014C40 , 32'hE9B10B80 , 32'hF04AF670 , 32'h0033D25C , 32'h03D7A934 , 32'h0AAA2070 , 32'hFF529258 , 32'hFC4FF1E0 , 32'hE248ECA0 , 32'hFDFD1058 , 32'hFA82FBA0 , 32'h0ACF3790 , 32'h0ACBC6B0 , 32'hF5010B80 , 32'hF61378F0 , 32'h04A29F40 , 32'hF92B2630 , 32'h17C013E0 , 32'hFC4E2DD4 , 32'h04A10378 , 32'h044BF588 , 32'h0F63EDE0 , 32'h07B0C808 , 32'h006264DF , 32'h04959930 , 32'h09A7C990 , 32'h0F7E07B0 , 32'h0BC5A400 , 32'h0BDE8230} , 
{32'hFE9C99A0 , 32'h1FB34420 , 32'hF5682350 , 32'hF58DA9D0 , 32'hEBCE9E60 , 32'h3BF63E80 , 32'h23EED100 , 32'hF9459FF8 , 32'h5BF05980 , 32'hDB298780 , 32'h02A2932C , 32'h0E4FF640 , 32'h147186A0 , 32'h0F0202D0 , 32'h139FCD20 , 32'h24D4DE80 , 32'h01F2B294 , 32'h153B2480 , 32'hFD82074C , 32'h22768E00 , 32'h03C2CA58 , 32'h18B876C0 , 32'hEEC0C0E0 , 32'h15053D20 , 32'hEEF90240 , 32'h0246E5CC , 32'h0B1A2190 , 32'h013C59AC , 32'h0325B8AC , 32'hFD8E6C48 , 32'h0FBAD820 , 32'hE6391AE0 , 32'h1D58C960 , 32'hF71D3730 , 32'h136762C0 , 32'h0434FBC0 , 32'hF4915BB0} , 
{32'hD6FEFA80 , 32'h3DEEBB40 , 32'hFD902CA0 , 32'hD2EECFC0 , 32'hEC42A4C0 , 32'h03A25C28 , 32'h0A836050 , 32'h0480EC28 , 32'hFA20C720 , 32'h1515AD40 , 32'hD96FD2C0 , 32'h058BE208 , 32'h2B352400 , 32'h11763FE0 , 32'h04AB1088 , 32'h17A5CD40 , 32'h03AD70A0 , 32'hE4B76200 , 32'hE94CD7E0 , 32'h161AD380 , 32'h0811AEB0 , 32'hF27A4BA0 , 32'hEA2D14C0 , 32'h0E96E490 , 32'h11385F00 , 32'hCC76FE00 , 32'h16960F60 , 32'hD03A9B80 , 32'h0B828B60 , 32'h2E01D580 , 32'hFF280F88 , 32'hE59888A0 , 32'hDCB94680 , 32'hED64E600 , 32'hD338CA00 , 32'h167ECE40 , 32'h10247840} , 
{32'hFF2A1441 , 32'h1B031980 , 32'h087D79F0 , 32'hE7C15260 , 32'hFA9E0A10 , 32'hFB0F9FE0 , 32'h008FA031 , 32'h0A9DA9B0 , 32'h0932EC70 , 32'hFB9AC678 , 32'hDB003DC0 , 32'h027AABF0 , 32'h0E810F50 , 32'h0DA22390 , 32'h11C498C0 , 32'h1F1F9D60 , 32'h00422567 , 32'hDDCD4340 , 32'hEA011FE0 , 32'h1566CF20 , 32'hFBFDB700 , 32'hEA1BE820 , 32'hEB9380C0 , 32'h059830D8 , 32'hF7CAF8E0 , 32'hFFBA28E2 , 32'h122F1540 , 32'hE92D3560 , 32'hF9F1B470 , 32'h1CDAA920 , 32'hFE76EF18 , 32'hE9FFF200 , 32'hDFBDA980 , 32'hECA63A60 , 32'hDAC1E380 , 32'h17C22460 , 32'h1112D880} , 
{32'hECEF8A60 , 32'h2F1EF500 , 32'h092F1E00 , 32'hE0934080 , 32'h0C4DC910 , 32'hD9E40F00 , 32'hFEAEB6E0 , 32'h0F0D1950 , 32'hEB1B7C40 , 32'h0C069CA0 , 32'hE7C795A0 , 32'h1794CF60 , 32'h0792CBB8 , 32'hF580AC20 , 32'hF50B1680 , 32'hE2939980 , 32'h0194E5D4 , 32'hF17D0CC0 , 32'h09674740 , 32'h11F82EE0 , 32'h053EDD48 , 32'h03003BDC , 32'h0DA51690 , 32'hEC078200 , 32'hEBD35660 , 32'hF3528610 , 32'h27AD5500 , 32'hE4AF5EC0 , 32'hFE3ED0F0 , 32'h0A80A7B0 , 32'hD4F1FA80 , 32'hE5DBB6C0 , 32'hDDA9C800 , 32'hF9CDBAF0 , 32'hF9B6EBF8 , 32'h090F4370 , 32'h08608590} , 
{32'hED6B5CC0 , 32'h24775940 , 32'h19EDB4C0 , 32'hF7AEA670 , 32'hEEBC3EA0 , 32'hCAB35300 , 32'hFFD32B42 , 32'h168B0D40 , 32'hEBDE7400 , 32'hF7C5BBE0 , 32'hE8798A40 , 32'hFC15C77C , 32'h0BCC5520 , 32'hF4F3C490 , 32'hF7756090 , 32'hDE7925C0 , 32'h18ABD200 , 32'h08EB1640 , 32'h15A1FFA0 , 32'h08D45F50 , 32'hF72E8450 , 32'h0EC6EF50 , 32'h01F9449C , 32'hF567A4C0 , 32'h013AADCC , 32'hFB435CB0 , 32'h09E16CD0 , 32'hFE764EE0 , 32'h107B69C0 , 32'h009D38F9 , 32'h0832C530 , 32'hE78C1320 , 32'hEDBC0720 , 32'h0E62F400 , 32'hE6016780 , 32'h00F34BC9 , 32'h0E3A4AB0} , 
{32'hDF036780 , 32'h2CCD1640 , 32'hF79EE430 , 32'hEFD1C3C0 , 32'hF0391EE0 , 32'hC710C500 , 32'h10623FC0 , 32'h2757D000 , 32'hC76CED40 , 32'h03D4F92C , 32'hE4ACF120 , 32'h057A36D8 , 32'h04AE9AF8 , 32'h09B37460 , 32'hF29BD910 , 32'hD00FB6C0 , 32'h13538F00 , 32'hFB161E00 , 32'h15E2F200 , 32'h1B07D6A0 , 32'h08A6D2C0 , 32'h30874DC0 , 32'h1988A880 , 32'h109FFEA0 , 32'hF8A03FE8 , 32'h0891CC90 , 32'h0E3C2670 , 32'hFADE2690 , 32'hF0B55860 , 32'h0655CA80 , 32'h0F605340 , 32'hF743C2B0 , 32'h06133C70 , 32'h110FA440 , 32'hEF17DB20 , 32'h002F323D , 32'hF7DD0A50} , 
{32'hC116B6C0 , 32'h3ACDC180 , 32'hF6057E60 , 32'hF6D269B0 , 32'hFB3AD1D0 , 32'hDBBF71C0 , 32'h11EC7500 , 32'hFB2D81B8 , 32'hC193E3C0 , 32'h1000AC20 , 32'hD8AD3C40 , 32'hEB0D93A0 , 32'h1CFE4E20 , 32'h22E84D80 , 32'hEFC63CC0 , 32'hE3F4D300 , 32'h1BAD3FE0 , 32'h0BF6B330 , 32'h1C11FDE0 , 32'h2C08D080 , 32'hF19BDA10 , 32'h2D624600 , 32'h31F66540 , 32'h04F77498 , 32'hDCF2D4C0 , 32'h047A0A78 , 32'hFBA0F7D8 , 32'hD46B6800 , 32'h13CE1020 , 32'h0B0EE2E0 , 32'h024E2EBC , 32'hFB487360 , 32'hF0A810D0 , 32'hECC45B80 , 32'hFA451578 , 32'hEE163820 , 32'h1D9DD080} , 
{32'hDA142600 , 32'h10581AA0 , 32'h040EE118 , 32'hFA93F000 , 32'h04E00B28 , 32'h150FD7A0 , 32'h1743C6A0 , 32'hDF5A3000 , 32'h1C5E6860 , 32'hEC0C45A0 , 32'hD6C74540 , 32'hEBF45B40 , 32'h1563C820 , 32'h1B70FC40 , 32'hEC4A76E0 , 32'hD7C827C0 , 32'h1161F020 , 32'h0CC23BB0 , 32'h134A5C80 , 32'h36F39A80 , 32'h0F019B50 , 32'h1B6D2780 , 32'h076A0398 , 32'h0670EF88 , 32'h07D9FDF8 , 32'h0E6EA710 , 32'hF6333DA0 , 32'hFCB9DB10 , 32'h0E62C850 , 32'h14892640 , 32'h148B3D80 , 32'hF7FB5DF0 , 32'hED8482A0 , 32'hE851BE20 , 32'hEBEFCF60 , 32'h0C766330 , 32'h0382DB10} , 
{32'hE34447E0 , 32'h23780000 , 32'h053249D0 , 32'hEF658B60 , 32'hF61C18A0 , 32'h188AF160 , 32'h07048680 , 32'hF2D24740 , 32'hFD5CEFCC , 32'h0022FADB , 32'hF1522EF0 , 32'hED0E2680 , 32'h1B2576C0 , 32'h0D6A0930 , 32'hF4400AE0 , 32'hEC2C1D00 , 32'hF97BE618 , 32'h1AFBC4C0 , 32'h14097660 , 32'h32E50940 , 32'h01C8405C , 32'h10D9B9E0 , 32'hFE46B05C , 32'h0F0A39B0 , 32'hF90296B8 , 32'h0C80F140 , 32'hEC2F8580 , 32'h1425E7A0 , 32'hF65326C0 , 32'hF6A29F70 , 32'hFB0260E0 , 32'h114DCB60 , 32'h0E956670 , 32'hFD93AAEC , 32'hF7CE0D90 , 32'h0A636610 , 32'hFEE5DEC0} , 
{32'hBE2E8080 , 32'h4AC4F800 , 32'hE71417A0 , 32'hF526DE00 , 32'h050D9AC0 , 32'h28049640 , 32'h0E329120 , 32'hE5DC9800 , 32'hD9B3BBC0 , 32'h1F9CE040 , 32'hF2B2B4F0 , 32'hE5BC2280 , 32'hEF27C520 , 32'hF1B0D860 , 32'hD5DCF800 , 32'hFFFBA696 , 32'hE36979E0 , 32'h07F8FC78 , 32'h1961A760 , 32'h1A9A4200 , 32'hF61247D0 , 32'hEB7EFB60 , 32'h01E601A8 , 32'hFDA6BB4C , 32'hE0F58C00 , 32'hE9C00720 , 32'h084A0170 , 32'h12698140 , 32'hF38E7AC0 , 32'hFD90CE20 , 32'hE8CCAB80 , 32'h043B1060 , 32'h1BAD30C0 , 32'h0FAAF080 , 32'h1AD88680 , 32'hFC429C44 , 32'hF9ADFC98} , 
{32'hF5E74B30 , 32'h2031B580 , 32'hFA658178 , 32'hE1497880 , 32'h08F2C580 , 32'h118923A0 , 32'h0294B5C4 , 32'hF2DFC8F0 , 32'hF91C50B8 , 32'h30550380 , 32'h0C7DF840 , 32'hDC0E0A40 , 32'hFDCCF42C , 32'hFCF9C590 , 32'hFA9F6D68 , 32'h0C718DA0 , 32'hE6416280 , 32'h02671A7C , 32'h2DA1A680 , 32'h13F39720 , 32'hED0E4B20 , 32'h2451DF80 , 32'hF982BB50 , 32'hEFDA62C0 , 32'h09262B10 , 32'h056C0CC8 , 32'h11108F40 , 32'h098ACD30 , 32'hFDE0203C , 32'hED1CBC00 , 32'h08D0FD20 , 32'h211CC380 , 32'hF5359A20 , 32'h0087410B , 32'h06F4A808 , 32'hFDBFA628 , 32'hEE8D3A00} , 
{32'hE6FD0CC0 , 32'h247BA580 , 32'hEE5F3860 , 32'hDE226000 , 32'h0A67F470 , 32'h234BF700 , 32'hFBCEEDA0 , 32'hF4FF92D0 , 32'h120BA880 , 32'h415F2600 , 32'h179DCD20 , 32'hE690D720 , 32'hEC73DDC0 , 32'hDB636080 , 32'hFDB1A848 , 32'h13E2C300 , 32'hE45969C0 , 32'h0B3B7570 , 32'h2E1511C0 , 32'h0EA46240 , 32'h16503480 , 32'hFEB1EE0C , 32'hF0272150 , 32'hEC51E840 , 32'hE90E9D80 , 32'h25EEF180 , 32'h125E0440 , 32'h1C3BFB80 , 32'hEA369E20 , 32'h0BEF0270 , 32'hE8AEECC0 , 32'hF82827B8 , 32'hEF400F40 , 32'hF59B5760 , 32'h0CF86D40 , 32'h090DA860 , 32'hF7A233B0} , 
{32'h09173360 , 32'h0F6D0770 , 32'hFA5E8C28 , 32'hDBBAB180 , 32'hFB2DFD20 , 32'hFBBE1BB8 , 32'h09D54A00 , 32'hFA194568 , 32'hFD74ADA8 , 32'hFE73543C , 32'hF88D1F28 , 32'hFA0DF5C8 , 32'hF8BBE260 , 32'hFDD5EF18 , 32'h01B183A4 , 32'hFF0A3C11 , 32'hF3A7E0E0 , 32'hF5124BD0 , 32'h136F9080 , 32'hF88F7EC0 , 32'h00B481C9 , 32'hF4FD93A0 , 32'h1A951DC0 , 32'hFF404094 , 32'hF4ECBFC0 , 32'h12EE37A0 , 32'h113F7FE0 , 32'h019A734C , 32'hF586F910 , 32'h049C2BE8 , 32'h0B3C8030 , 32'hF710CB30 , 32'h16FDED80 , 32'h0B0B6480 , 32'hF09C0B80 , 32'h19A963C0 , 32'h01725EDC} , 
{32'h051C3700 , 32'h02D6C7F0 , 32'h0D6A2360 , 32'hF53B1C10 , 32'hFB849408 , 32'hD92669C0 , 32'hF783B1D0 , 32'h136D86A0 , 32'hED18C680 , 32'h1A2E4AC0 , 32'h1BBEDE40 , 32'hFDE431B4 , 32'hEED74C80 , 32'h15CE8E20 , 32'h14A6CFA0 , 32'h148C6860 , 32'hE1784F00 , 32'hFA9A05F0 , 32'h0A6DE830 , 32'hECC3B960 , 32'hFA3A5D98 , 32'hEAA2FD60 , 32'h089DF700 , 32'hF1E6B6E0 , 32'hF2B99980 , 32'h04831810 , 32'h04DF3130 , 32'h030A62E8 , 32'hF8A1DFD0 , 32'hF2320DB0 , 32'hFE66C3DC , 32'hEA844B20 , 32'hF6A0EC50 , 32'h034EA914 , 32'hF3797D00 , 32'h3C56D400 , 32'h09715130} , 
{32'h08735260 , 32'hFD205384 , 32'hFBF99248 , 32'hFD61FA28 , 32'hF6EB1170 , 32'hD59FFF00 , 32'h00C07976 , 32'h1D05DA60 , 32'hE69EC2A0 , 32'h14C048A0 , 32'h1C2146A0 , 32'h19425780 , 32'hF6ABBD00 , 32'h0EE192A0 , 32'h0FE0E390 , 32'h147F6320 , 32'hE15E7040 , 32'h0AA2B0D0 , 32'hFB2DC690 , 32'hEF182DC0 , 32'hEABFA4A0 , 32'hF33CEB10 , 32'hF7EF2A90 , 32'hEE876180 , 32'hF6E45EC0 , 32'h07A4C620 , 32'h002536CD , 32'hFFB8F613 , 32'hF3D5D630 , 32'hF8CE69C0 , 32'hF0B82350 , 32'hF0A1B100 , 32'hF5C8F0C0 , 32'hF2CF0FB0 , 32'hFB2B57D0 , 32'h1F628340 , 32'hF4F11840} , 
{32'h006E15F6 , 32'hFF62211D , 32'h009FE2E9 , 32'h00C5A8D8 , 32'hFFB8C6AB , 32'hFFFB7C72 , 32'hFFE20CE0 , 32'h0086DB4B , 32'h0055ED7E , 32'h006C436B , 32'hFFEBE203 , 32'hFFF76958 , 32'h007F5446 , 32'h002B0253 , 32'hFFE2AD47 , 32'h00BC1573 , 32'h000FF9E8 , 32'h008A68A7 , 32'hFFEAD106 , 32'hFFCBBA74 , 32'h00025A51 , 32'h005EA377 , 32'hFF6AEB0C , 32'hFF8F3023 , 32'hFF8816A7 , 32'hFFE8E04C , 32'hFEF85D70 , 32'h006E9DF5 , 32'h00270BC1 , 32'hFF8F4583 , 32'hFF2DBA78 , 32'hFEAC6360 , 32'hFFC86155 , 32'h00290908 , 32'hFFA34A76 , 32'hFF8CBA64 , 32'h00D6EC99} , 
{32'h0068504B , 32'hFF58D9F8 , 32'h00DD0BE1 , 32'h00F29FE2 , 32'hFF8C30EB , 32'hFFFD31E3 , 32'hFFEA3DAC , 32'h00AE233A , 32'h00631D8A , 32'h009C410C , 32'hFFF9235C , 32'h0007709B , 32'h00AC9CED , 32'h003209EF , 32'hFFEF0DED , 32'h00EFAB9C , 32'h001B77D5 , 32'h00BDE577 , 32'hFFFB194D , 32'hFF9DDF9C , 32'h000BAEAC , 32'h0075CAE4 , 32'hFF7651ED , 32'hFF963D46 , 32'hFF346AA1 , 32'hFFAE4AFB , 32'hFEDF0124 , 32'h00E681C6 , 32'h002007A3 , 32'hFFAA3878 , 32'hFF0DF552 , 32'hFEA1F94C , 32'hFFA8FD3B , 32'h003A12BC , 32'hFFA31086 , 32'hFF6ED33D , 32'h00FD057D} , 
{32'h00647FA5 , 32'hFFA929F2 , 32'h007C22EC , 32'h005C1456 , 32'hFFA7DB12 , 32'hFFEE7951 , 32'h00124F56 , 32'h0073FCA8 , 32'h004D3B71 , 32'h00510087 , 32'hFFAA69E7 , 32'h0008675B , 32'h002F9989 , 32'hFFF2C476 , 32'hFFF34A67 , 32'h005FABAB , 32'hFFAB0BC0 , 32'h00478534 , 32'h001BAD48 , 32'hFF8AA878 , 32'h0034CC6D , 32'h0044C9B2 , 32'h00085208 , 32'hFFA0F85C , 32'hFF926D47 , 32'hFFEB550D , 32'hFF75A650 , 32'h0064B493 , 32'h0025355F , 32'h0000C239 , 32'hFF6A7324 , 32'hFF0F7F19 , 32'hFFFF1BC6 , 32'h0063FDF1 , 32'hFFD4AA91 , 32'hFF6DBB25 , 32'h0055783A} , 
{32'h00053C78 , 32'hFFFE5630 , 32'h0000A738 , 32'h000720FB , 32'h00098656 , 32'hFFFFE12F , 32'hFFFD2C39 , 32'h0000B3DB , 32'hFFF8C3E7 , 32'hFFFBB2CD , 32'hFFFE5D05 , 32'hFFFDA2B1 , 32'h00080545 , 32'h0007223F , 32'hFFFEA202 , 32'h00013C5F , 32'hFFF93CA5 , 32'h0009600F , 32'h000141E6 , 32'hFFFA4A0B , 32'h0000F8D3 , 32'h0004A5AB , 32'h00046F52 , 32'h0001C7E8 , 32'h00047E73 , 32'hFFFD8ADC , 32'h000222E1 , 32'hFFFF3968 , 32'hFFF54C9F , 32'h0000A6BC , 32'h0003CAE3 , 32'hFFFCFDEF , 32'hFFFDA9E0 , 32'h00011D2F , 32'h00070DCC , 32'h0006C38A , 32'hFFFA1FC9} , 
{32'hFFFA5B9C , 32'h00011DA7 , 32'h000AB665 , 32'h00038317 , 32'hFFFDC1C2 , 32'hFFF98A16 , 32'h000541B3 , 32'h000037E8 , 32'h0000BAD8 , 32'hFFF89C62 , 32'hFFF9D94B , 32'hFFFB34AD , 32'h00010526 , 32'hFFFEF004 , 32'hFFF98524 , 32'hFFFC9FE3 , 32'hFFF533BF , 32'hFFFEF3D0 , 32'hFFFD01DB , 32'hFFF75159 , 32'h0000CA91 , 32'hFFFD3988 , 32'hFFFEF207 , 32'h000183DB , 32'hFFFF1B20 , 32'hFFFCC8C2 , 32'hFFFD15F3 , 32'hFFFE5CFE , 32'h0009D988 , 32'hFFFFC6D6 , 32'hFFFF960C , 32'hFFF9C906 , 32'hFFFA9097 , 32'hFFFDB2FB , 32'h000485B6 , 32'hFFFDB355 , 32'hFFFBA0EB} , 
{32'hFFFA91F3 , 32'hFFFC0DA9 , 32'hFFFE6F3D , 32'hFFFD93BE , 32'hFFFD32A8 , 32'hFFFB2A00 , 32'hFFFB177C , 32'h0007A31B , 32'hFFFAA8FA , 32'h0000A1AD , 32'h00082C68 , 32'hFFF84051 , 32'h0000E636 , 32'hFFFF2DB8 , 32'h00046087 , 32'h00009447 , 32'h000994AA , 32'h000130F3 , 32'h00083A1F , 32'hFFF34679 , 32'h0008B64F , 32'h00056007 , 32'hFFF9915E , 32'hFFFC0AE6 , 32'h000156FA , 32'hFFF6E36E , 32'hFFFBB905 , 32'h000B659E , 32'h000579FE , 32'h0002056D , 32'hFFFD51E7 , 32'h0001E00F , 32'h00044ED0 , 32'h00082B06 , 32'h00048D29 , 32'hFFF92173 , 32'hFFFFF264} , 
{32'hFFFCDA02 , 32'hFFFD45D3 , 32'hFFFAE8D7 , 32'hFFFABC72 , 32'h000738C1 , 32'h0004D68F , 32'hFFFF470E , 32'h0004BAD8 , 32'hFFFD3CD4 , 32'hFFFFB00E , 32'hFFFB9911 , 32'h000B3ECD , 32'hFFFD6D3E , 32'hFFFCFA3D , 32'hFFF81AFB , 32'hFFFE9E35 , 32'hFFFFFBCB , 32'hFFF8EF4C , 32'h00035FA5 , 32'hFFFD6725 , 32'h0005BF0B , 32'h00092849 , 32'hFFFE14EF , 32'hFFFF1B8F , 32'h0003237F , 32'h000241DC , 32'hFFFF0B6A , 32'hFFFC33EC , 32'hFFFE00EB , 32'hFFFA8605 , 32'h0003E8F4 , 32'h0002CD84 , 32'hFFFE9065 , 32'hFFFDBC5B , 32'h0001A8C6 , 32'h0001CBB6 , 32'h0001DC4B} , 
{32'h000137F3 , 32'h00007E98 , 32'hFFFB7C14 , 32'hFFFF587E , 32'hFFFC1588 , 32'h00064FDA , 32'hFFFE311B , 32'hFFFDF707 , 32'hFFFEDDF8 , 32'h00002675 , 32'hFFFF062E , 32'h00035B28 , 32'h0002149E , 32'hFFFD0A7C , 32'hFFFB82F8 , 32'hFFFCC23C , 32'hFFFC9E13 , 32'h000638DD , 32'hFFFF3D26 , 32'hFFFEED3D , 32'h0002B7A4 , 32'h0001BB11 , 32'hFFFEAF97 , 32'h00026E6E , 32'h00016A56 , 32'h00045D65 , 32'h00041338 , 32'hFFFF72C3 , 32'h00055237 , 32'h0001C360 , 32'hFFFD624E , 32'hFFFF9D6A , 32'hFFFC725A , 32'hFFFB84FC , 32'h00088691 , 32'h00062848 , 32'hFFFA68B6} , 
{32'h0003E025 , 32'hFFFFAE78 , 32'hFFFC9FA1 , 32'hFFF9EB95 , 32'h000368D6 , 32'h00076568 , 32'h0003B7F4 , 32'h0000750F , 32'hFFFEC5BF , 32'h00048772 , 32'hFFFD7667 , 32'hFFFC2656 , 32'h0008DB45 , 32'hFFF485D4 , 32'hFFFCB767 , 32'hFFFDF315 , 32'h00098DFC , 32'hFFFFE429 , 32'hFFFD0142 , 32'h00094C55 , 32'hFFFDB3D4 , 32'h00076321 , 32'h00054829 , 32'hFFFAF36D , 32'h000A67CD , 32'h00056FE9 , 32'h0000E664 , 32'h0002DEEA , 32'hFFFDD65E , 32'hFFFFBF52 , 32'h000075BC , 32'h000B0315 , 32'h00031642 , 32'h0000AAED , 32'h0004B5FB , 32'hFFFEE0F9 , 32'h000376C4} , 
{32'h03B833E4 , 32'h0303F8B0 , 32'hFA605370 , 32'hFC91FEBC , 32'hFF1175C0 , 32'h019D1550 , 32'hFC8BDC54 , 32'h0187ED14 , 32'hFC3795F4 , 32'h004A4B78 , 32'hF3A0D3E0 , 32'h016D7E9C , 32'h06F807B0 , 32'h055FF818 , 32'h0509B598 , 32'hFEC16768 , 32'h05775A20 , 32'h05DB8B68 , 32'h0283149C , 32'hF8EE5B90 , 32'h03F20F5C , 32'hFE3ECFC4 , 32'hF6C16EF0 , 32'hFDDE0180 , 32'h00C3EA06 , 32'h03E741E0 , 32'h10437DC0 , 32'h04AA91F0 , 32'h065030F0 , 32'hFC82A8C8 , 32'hFA9BE338 , 32'h0711F1E0 , 32'h06508DA8 , 32'hFCD30988 , 32'h037E7354 , 32'h01B80070 , 32'h06CA1F00} , 
{32'h012BAA98 , 32'h0F537CD0 , 32'h1B83C020 , 32'h0776ABE8 , 32'h19311F00 , 32'h01C80744 , 32'hF60670A0 , 32'h17368160 , 32'h1486C180 , 32'h01C42DF8 , 32'hF1762430 , 32'hF97EEB20 , 32'h22397780 , 32'h0BCF3A50 , 32'h040B9DA8 , 32'h11E858A0 , 32'hFD3B547C , 32'h009322C0 , 32'h039398D4 , 32'hF3909750 , 32'h038C6134 , 32'hF8A967E8 , 32'h06E703B0 , 32'hFBF89E50 , 32'h09A19120 , 32'hF459DAC0 , 32'h09A97E00 , 32'h18FAB920 , 32'h02C9F048 , 32'hFEE73484 , 32'hF7AF1260 , 32'hFBAE5EF0 , 32'h1C7ADD20 , 32'h07575BF0 , 32'h054E54E8 , 32'h05D09170 , 32'h03D07524} , 
{32'h09A2A500 , 32'hFCC724F0 , 32'h054C3DD0 , 32'h03B3479C , 32'h052A60D8 , 32'h05D2F5C0 , 32'hFB688F48 , 32'hFE94E020 , 32'h0C6D2B50 , 32'h0087D5D1 , 32'h0A871E50 , 32'h18949EE0 , 32'h090ECDE0 , 32'hF6F2D130 , 32'hED292700 , 32'hFD2527C0 , 32'h1E87D4C0 , 32'hF44D0280 , 32'hEE3CCC60 , 32'h0F781A60 , 32'h01B25D10 , 32'h16656E80 , 32'hFE0CC830 , 32'h03B85424 , 32'hF3F5B320 , 32'hF234B820 , 32'hFF5A78BC , 32'h06582E90 , 32'h0EAC3660 , 32'h094AA840 , 32'h0937D6F0 , 32'h11B0CCC0 , 32'h042F19D8 , 32'hFCDD8910 , 32'h0DEE69D0 , 32'hEA8F4F40 , 32'hF76E9250} , 
{32'h035411E4 , 32'h16030200 , 32'hFF6CB4BA , 32'hF4038110 , 32'hE6102BE0 , 32'h359733C0 , 32'h1DA578E0 , 32'hFE3A4920 , 32'h2BCA9E00 , 32'hFA8F4E08 , 32'h1588D0A0 , 32'hF55F8320 , 32'h042C2FA0 , 32'hFD5A131C , 32'h20972100 , 32'h11F78320 , 32'hF5E579B0 , 32'h13049660 , 32'h1ED7E3E0 , 32'h1C953B00 , 32'h002A7C1F , 32'h25BFFE80 , 32'hF4E48CD0 , 32'h05F395A0 , 32'h0A877C40 , 32'h09A3DEE0 , 32'h136D52A0 , 32'hFAC2A4A8 , 32'h139BE400 , 32'hDDDFF080 , 32'h25FC7480 , 32'hEF06EC00 , 32'h00848907 , 32'h00AE9348 , 32'hEB852440 , 32'hD9E4D400 , 32'hF3FB8E50} , 
{32'hEF2B51E0 , 32'h0D1EDEC0 , 32'h09A445D0 , 32'hF097DF20 , 32'h0887AE80 , 32'h02E565B8 , 32'hF5BC0400 , 32'hF83B80E0 , 32'h23DB8640 , 32'h021EACE8 , 32'hFD424354 , 32'hF8B66938 , 32'h156776E0 , 32'hE803ACE0 , 32'h1F300900 , 32'h1EEF2A00 , 32'hEC85A5A0 , 32'hEF7B27E0 , 32'h1187AD00 , 32'hE7AC35C0 , 32'hFE1FC8A8 , 32'h20274FC0 , 32'hD83BEAC0 , 32'hE4A8C480 , 32'h031D16B4 , 32'h0CFE6610 , 32'h211067C0 , 32'hF8DA52E0 , 32'hFCAA3D84 , 32'h0015C3DB , 32'h0F950130 , 32'hFB8040C0 , 32'hF36350A0 , 32'hF3701040 , 32'hEF135280 , 32'hF00EEF90 , 32'h0803AC80} , 
{32'hEDD37320 , 32'h289D4A40 , 32'h23F52880 , 32'hC2F6DF80 , 32'hF7329460 , 32'h161F2A60 , 32'hBF0B4080 , 32'h4AD52500 , 32'hF4CAAC50 , 32'h00DB8B55 , 32'hF50A3040 , 32'h154B1500 , 32'h2975D940 , 32'hF4A62B60 , 32'h2D853F80 , 32'h1BA08660 , 32'hC930A740 , 32'hD9507F40 , 32'hD4ACE540 , 32'hFF19FFBC , 32'hF8103BB0 , 32'h067098F8 , 32'hCE31E8C0 , 32'hF0A42A40 , 32'h23F47DC0 , 32'hCAB80540 , 32'h1F2A6E20 , 32'h0BF90990 , 32'h06D26E90 , 32'h3680BC00 , 32'h25387D80 , 32'hC5924FC0 , 32'hE7D61B00 , 32'hFE8E0404 , 32'hCE3D7380 , 32'hF0D5F790 , 32'hF7E92620} , 
{32'hE2877400 , 32'h0073A67E , 32'h2052F7C0 , 32'hE00D4320 , 32'hF854C468 , 32'hD7113680 , 32'hF0635790 , 32'h2A7F98C0 , 32'h197A6FC0 , 32'h0C551A00 , 32'hF9741258 , 32'h1EC41EA0 , 32'h18A90CC0 , 32'hDEDDFC40 , 32'h4184E800 , 32'h1A30F660 , 32'hF9C67740 , 32'hF31D5480 , 32'h0316ED00 , 32'h03A6EE84 , 32'hDFC53C80 , 32'h0B6AA350 , 32'hC75AAAC0 , 32'hEC393CE0 , 32'hFB0E6D88 , 32'h03508938 , 32'h13872C40 , 32'h0A1EE1D0 , 32'hF0435840 , 32'h11466DE0 , 32'h12601140 , 32'hFFC55E9F , 32'h0239ACB4 , 32'hF8B939A8 , 32'h048537E8 , 32'h01244CA0 , 32'hF4F9F670} , 
{32'hE9E97620 , 32'h0AA48EA0 , 32'h1D10F960 , 32'hDE4D7CC0 , 32'h09FA50F0 , 32'hDDCAC600 , 32'hE2695B60 , 32'h215ED4C0 , 32'h08B7D480 , 32'h1EF0E5A0 , 32'h09939650 , 32'h0EF061C0 , 32'hF38EDC70 , 32'hCBD5DDC0 , 32'h26D3C800 , 32'h110D3680 , 32'hFF2CB4AB , 32'hF310E6B0 , 32'h0F3F84B0 , 32'hED2F2B00 , 32'hF42D2870 , 32'h074325A8 , 32'hDFA92840 , 32'hF71BBA90 , 32'hF5525FB0 , 32'hF273A6C0 , 32'h136F6620 , 32'hFE80E6E0 , 32'hFCCF04EC , 32'h1A614220 , 32'h2BDD6640 , 32'h0ABE39A0 , 32'hF67BFD40 , 32'h05475020 , 32'h1E4E1D00 , 32'hEE356FE0 , 32'h0BE08200} , 
{32'hF255CBA0 , 32'h14F770A0 , 32'h1E1A1EA0 , 32'hC3E1D080 , 32'hEED42420 , 32'hA623BA00 , 32'hF3E642A0 , 32'h28DA2380 , 32'hA4BD2300 , 32'hE4184DA0 , 32'hF08742C0 , 32'h0AB16460 , 32'hE81AAB60 , 32'hC3904180 , 32'h3A2C1600 , 32'hE8AF1380 , 32'h33ED5900 , 32'hDD017780 , 32'h05FF3120 , 32'h13901AC0 , 32'hF35CA750 , 32'h208DE740 , 32'hEE67AA00 , 32'h17368F80 , 32'hEFCC9E00 , 32'h001F4127 , 32'h1BC2F380 , 32'hE9AC9B00 , 32'h19C2E760 , 32'hFC0FB440 , 32'h16CDBF60 , 32'h02888104 , 32'h0B37DA90 , 32'h285868C0 , 32'hF4530E30 , 32'h010B7E90 , 32'h01E50588} , 
{32'hCE4B5C40 , 32'h25A02640 , 32'h25880F00 , 32'hED196F00 , 32'h032400AC , 32'hBF13F400 , 32'h04311C28 , 32'h167F7DA0 , 32'hCAAD0380 , 32'hC97AC900 , 32'hF1A8E4B0 , 32'hFD566320 , 32'h0325FC60 , 32'hC6A78140 , 32'h0DDC0F70 , 32'hE30A7CC0 , 32'h1966E560 , 32'hF99C8F90 , 32'h16A24D40 , 32'h11769000 , 32'h0601B7B0 , 32'h0178BF1C , 32'hF20863D0 , 32'h0CD84090 , 32'hEB232180 , 32'hFCF70520 , 32'hD9B3D3C0 , 32'hF75A1870 , 32'h0618D5E8 , 32'h09A45880 , 32'h0D348850 , 32'hFBBC77E0 , 32'hFA8C7D88 , 32'hEED96180 , 32'h182DE5C0 , 32'hF9FE1F90 , 32'h1C50B600} , 
{32'hC9629CC0 , 32'h1A4221C0 , 32'h016C2400 , 32'hE09DF0C0 , 32'hF7AB53C0 , 32'h065233F0 , 32'h08EAF990 , 32'hF5C83570 , 32'hD7753A00 , 32'hD4E29540 , 32'hEDA44B80 , 32'h0586CD48 , 32'h09F028E0 , 32'hD87F8A80 , 32'hFADA4E10 , 32'hDB6BD0C0 , 32'h0AAC1D60 , 32'h00D5899D , 32'h1FA8AEC0 , 32'h5945B600 , 32'h0E0C8BD0 , 32'hF47E8B20 , 32'hF89E3100 , 32'h0FCD2760 , 32'hC2436480 , 32'h287A2CC0 , 32'hE3B959A0 , 32'hEC5AE5C0 , 32'hF850E4A8 , 32'h14EF9BC0 , 32'hFED64CE4 , 32'hFAF4EB68 , 32'hCCE7ED40 , 32'hDE98BD80 , 32'hF0E11D10 , 32'h090C5D00 , 32'h1A069A80} , 
{32'hDC96D1C0 , 32'h2B9642C0 , 32'hFA269E10 , 32'h096DAB20 , 32'hE6F03040 , 32'h14D197C0 , 32'h118A0840 , 32'hED958240 , 32'hFAAEA8E8 , 32'hE39027A0 , 32'hE344D800 , 32'hF6981530 , 32'h230FE5C0 , 32'h0B3A58D0 , 32'hE9C87580 , 32'hDFCC85C0 , 32'hEA68BE20 , 32'h0D63D6A0 , 32'hF95D77A8 , 32'h1D7D0480 , 32'hE7E86C80 , 32'h1A1D0B80 , 32'h0140EA9C , 32'h20605E80 , 32'hE6DB1700 , 32'h20417B40 , 32'hE6C1ADC0 , 32'hFE2D770C , 32'h0E08EED0 , 32'hF71BAD20 , 32'hF841AAB0 , 32'hE6230520 , 32'hFECFDBC4 , 32'hFCFBF478 , 32'hFAAAE460 , 32'h0403AF68 , 32'h19FA3F20} , 
{32'hE2F09EE0 , 32'h11379860 , 32'hF1A9F960 , 32'hF0601F40 , 32'h07A7A1C8 , 32'h1F4D7A20 , 32'h03DB74DC , 32'hC8753B00 , 32'h0B6B8FE0 , 32'h01C4D718 , 32'hF0199E00 , 32'hEFAC0B00 , 32'h12C739C0 , 32'hCC0E97C0 , 32'hF46B6DF0 , 32'hF8A25618 , 32'h097302E0 , 32'h147A3360 , 32'h01DC14D0 , 32'h1D3032C0 , 32'hFDF1C81C , 32'hE2905EA0 , 32'h1957AFA0 , 32'h21272A00 , 32'h05727FB0 , 32'h0D81DA60 , 32'h09090F20 , 32'h1E78BF60 , 32'h0D44E0B0 , 32'h0CD048C0 , 32'h074D8988 , 32'h0BF9C4C0 , 32'h070D3158 , 32'h02AB2254 , 32'hF4CBC5A0 , 32'h1F0FB360 , 32'h014D4CB0} , 
{32'hE09C05C0 , 32'h2E5E52C0 , 32'h06B5CFB8 , 32'hE08E8900 , 32'h0BDAF4F0 , 32'hFC921150 , 32'h10C3AB20 , 32'hC6EE4DC0 , 32'hFB7CF4A0 , 32'h34171A40 , 32'h095AD080 , 32'hEB113560 , 32'h0F39CA90 , 32'h0CEC8310 , 32'hEEA544A0 , 32'hE6551CE0 , 32'hFC7DFC44 , 32'hF955C4E0 , 32'h1B704D20 , 32'h21BE8180 , 32'h018256AC , 32'h1F4215A0 , 32'h152A95C0 , 32'h1F69C0E0 , 32'hEC6ECCA0 , 32'h10FF7000 , 32'h18B22F40 , 32'hF2942CE0 , 32'hE9345620 , 32'h014CDF60 , 32'hDF5C0280 , 32'hE9017CC0 , 32'hEF7F27E0 , 32'h0CE17140 , 32'hEC6E2280 , 32'hE8C69140 , 32'h0E59FEA0} , 
{32'h0AC787D0 , 32'h37689500 , 32'hF34B9AE0 , 32'hAA70A580 , 32'hF1EB5A10 , 32'h097A9B30 , 32'h0D8E1C10 , 32'hAF95A600 , 32'hF7E4B970 , 32'h3AF5CD80 , 32'hE276E100 , 32'hDAE2F900 , 32'hF4F29A40 , 32'h16FD0CA0 , 32'hF8AD9C30 , 32'h0FD56C40 , 32'hE77CD400 , 32'hFD3C82DC , 32'h41F25A00 , 32'h22B60300 , 32'hF5F22230 , 32'hFD0C983C , 32'h2B8D4940 , 32'h088BADB0 , 32'hF6A49470 , 32'h1F9ACE20 , 32'h37E39180 , 32'hF9E13E08 , 32'hCDDD8440 , 32'hFDD7EE30 , 32'h2A860CC0 , 32'h0E51A420 , 32'h39B20000 , 32'h054A1898 , 32'hCE8F7A40 , 32'h12325340 , 32'h19BE6F80} , 
{32'h097AB9C0 , 32'h22BC6F40 , 32'h0441A6D0 , 32'hC8814A40 , 32'h02200E08 , 32'h155FD340 , 32'hF69B34C0 , 32'hBA746100 , 32'h0D24C930 , 32'h25133840 , 32'h2BDE3FC0 , 32'h1222D460 , 32'h0F58B710 , 32'h029DA1FC , 32'h107690C0 , 32'h09C7F7E0 , 32'h216FC240 , 32'h14D3FE00 , 32'h03AB4EFC , 32'hFAF22778 , 32'h1021E6C0 , 32'hFB1BAC08 , 32'hF1BD70D0 , 32'h14F9AA80 , 32'hEB3D2300 , 32'hEC1D0860 , 32'hF0F6DBF0 , 32'h20446FC0 , 32'hEA3ECEA0 , 32'h13F88700 , 32'h190FB8A0 , 32'h20204A80 , 32'hF58A8740 , 32'h16AAA640 , 32'hF60AEB90 , 32'h4ADD6280 , 32'hD93E5000} , 
{32'h00A7C1CC , 32'h1598E480 , 32'h118239E0 , 32'hD15AF980 , 32'h0E7BD5C0 , 32'hF8F66B70 , 32'hFB7C4BD0 , 32'hFC9D4FB8 , 32'hF684A440 , 32'h239A2CC0 , 32'h0CD82AF0 , 32'hE91E30E0 , 32'hFC3881C0 , 32'hFC714D30 , 32'hFDC9560C , 32'h0CB99000 , 32'hEB04AF60 , 32'hFC319020 , 32'h20DBC9C0 , 32'h18167D20 , 32'hDC98AF80 , 32'h1C802580 , 32'hE01F1EE0 , 32'hEF3C6360 , 32'h08298B40 , 32'hECE9F320 , 32'hF280DAF0 , 32'h0D897460 , 32'hEF542A40 , 32'hFCEC5C9C , 32'h05081D20 , 32'h1964BCA0 , 32'h09E23B30 , 32'hFCFAAA08 , 32'h236AD640 , 32'h081C03F0 , 32'hFD4FFEF0} , 
{32'h03A8AF90 , 32'hFD8D1A00 , 32'h09DC7F60 , 32'hF3E26C60 , 32'h055C07C8 , 32'hFE65A750 , 32'hF072E0F0 , 32'h0EC8D6E0 , 32'hF8402C80 , 32'h08A84980 , 32'h246FFD40 , 32'h1BAEDDE0 , 32'h414CEC00 , 32'h0DABD1F0 , 32'h0C4D5F40 , 32'h06C7A980 , 32'hED028F00 , 32'h0A1BC8D0 , 32'hFF34D60D , 32'hFF223772 , 32'h0AF5C630 , 32'hF9D13AB0 , 32'h07D06C20 , 32'hF36BE220 , 32'hF057C920 , 32'h124FE000 , 32'hF3514560 , 32'h14F49580 , 32'h06F0FFF0 , 32'h02629DE4 , 32'hF2E88360 , 32'hFC0F8AA8 , 32'h0100F60C , 32'h0FB9ED00 , 32'hFFBE3484 , 32'hF9DFE7B8 , 32'h091D4720} , 
{32'h076933E8 , 32'h16F23BA0 , 32'h1EF0F100 , 32'hD4D585C0 , 32'h10DC19C0 , 32'hEC8CEA20 , 32'hFDA2AC78 , 32'hDD6FA3C0 , 32'hB7391B80 , 32'h1179F060 , 32'h307E46C0 , 32'h05A43720 , 32'h0CF21880 , 32'h09262E20 , 32'h0D0BDCC0 , 32'h23C07E00 , 32'h05A2BD40 , 32'hF687B610 , 32'h0279AFCC , 32'h00BF0325 , 32'hEDAE3AA0 , 32'hF31CF4F0 , 32'h0D73CA00 , 32'hC61076C0 , 32'hFE2B0BB4 , 32'hE58B32A0 , 32'hECF08FE0 , 32'hF63958F0 , 32'hE61733C0 , 32'hF7AA13B0 , 32'hEAECBDC0 , 32'h0D880AE0 , 32'h142C6A60 , 32'hFCA7B204 , 32'h04D28E70 , 32'hF7578DD0 , 32'h000E4DC9} , 
{32'h04FD1BF8 , 32'hFE43D814 , 32'hFF0B823A , 32'h02EF6A90 , 32'hFE251E5C , 32'hF9A892F8 , 32'hFB143530 , 32'h12FE9140 , 32'hF9C60FF8 , 32'h0860BAF0 , 32'h0B5A4230 , 32'h0E0D40A0 , 32'h11384120 , 32'h04CBCE78 , 32'h0A1043D0 , 32'h08B4F530 , 32'hF28C3480 , 32'h03F5E3A4 , 32'hF1BF2FE0 , 32'h00521949 , 32'hFF531F48 , 32'h02E54430 , 32'hFAA5ADA8 , 32'hF52CB800 , 32'hFBE12038 , 32'h0BCB29B0 , 32'hF8136488 , 32'h08FEFC20 , 32'hFB6BF620 , 32'hFD99826C , 32'hF66B8340 , 32'hFB131D30 , 32'h067AF7F0 , 32'hFE666A50 , 32'h01009510 , 32'hFCCB0B80 , 32'hFE06D178} , 
{32'h0068D050 , 32'h004357C6 , 32'h009B8F40 , 32'hFF795E33 , 32'h0094FFA9 , 32'hFFD50A6E , 32'h00047C61 , 32'hFF9A24EB , 32'hFEFB8DCC , 32'h00441226 , 32'h0134AC8C , 32'h00DCDC74 , 32'h00A169C3 , 32'hFFD43ACE , 32'h001BB98C , 32'h008ABEB7 , 32'hFF8AFFE0 , 32'h0070F5C1 , 32'hFF5F870E , 32'hFFC57C86 , 32'hFFC49917 , 32'hFF5BE239 , 32'hFFF8A2E5 , 32'hFED769F0 , 32'hFFD76916 , 32'hFFD6AE73 , 32'hFF797D25 , 32'h00939D20 , 32'hFF8EC911 , 32'hFFEDAA96 , 32'hFF083A47 , 32'hFFC92F46 , 32'h013A39B8 , 32'hFF6E6AE4 , 32'hFF9CB8FE , 32'hFF3B9376 , 32'hFF4E6324} , 
{32'h000153C4 , 32'h0000B645 , 32'hFFF53691 , 32'h000185BB , 32'h0004A9FA , 32'h00014B16 , 32'hFFFB63AC , 32'h0002A23A , 32'hFFFD2863 , 32'hFFFA5018 , 32'hFFFE2A5B , 32'hFFFEF5C6 , 32'hFFF9814C , 32'hFFFFEE00 , 32'hFFFBE575 , 32'h0001EB44 , 32'hFFF8D374 , 32'hFFFF00A5 , 32'hFFFC73DF , 32'hFFFB37E9 , 32'hFFFE393B , 32'hFFFF848B , 32'h0006613A , 32'hFFFCA26B , 32'hFFFD268C , 32'h0004A1F5 , 32'hFFFCAC9A , 32'hFFF7E897 , 32'h000165C6 , 32'h000CCB9B , 32'h0000567C , 32'hFFFDA486 , 32'hFFF8118E , 32'hFFFC497F , 32'h0001112A , 32'h0001C76B , 32'h00048C82} , 
{32'hFFFB174D , 32'h00008FB8 , 32'h0000F167 , 32'h000139EC , 32'hFFFDF663 , 32'hFFFFB295 , 32'h0001C812 , 32'h0001D908 , 32'h000136D6 , 32'hFFFB7202 , 32'hFFF93846 , 32'h00007492 , 32'hFFFF99E8 , 32'hFFFF3320 , 32'h000176D6 , 32'h0005D7BF , 32'h0000728C , 32'hFFFFCB2E , 32'hFFFB5FFB , 32'hFFFFE87C , 32'hFFFF0AC1 , 32'hFFF8BE14 , 32'h00054C14 , 32'hFFFE27A5 , 32'hFFFAE48A , 32'h00004073 , 32'hFFF4AC27 , 32'hFFF54AFB , 32'hFFFDB4AE , 32'h00046FB1 , 32'h0002BDD1 , 32'h00075AD8 , 32'h000A5BBC , 32'h0001A060 , 32'h00085237 , 32'h0000D661 , 32'hFFFDDE0B} , 
{32'hFFF9EB46 , 32'h0001E34D , 32'hFFF4E21A , 32'hFFFA110D , 32'h0001F6E0 , 32'h00017307 , 32'h0001DB80 , 32'hFFF91CA8 , 32'hFFFC2AB7 , 32'h00007714 , 32'h0000DC4B , 32'hFFFEEAC7 , 32'hFFFDBB51 , 32'h0001D37C , 32'hFFFA3482 , 32'h00080DCF , 32'hFFFACBC5 , 32'hFFFBCDC2 , 32'hFFFFA977 , 32'h0000593E , 32'h00002F83 , 32'h000083A9 , 32'hFFFB8972 , 32'h0000332D , 32'h0007AF15 , 32'h0006C43F , 32'h0009FF57 , 32'hFFFF4EF5 , 32'h000412B9 , 32'h00040DBA , 32'hFFFEFF4D , 32'hFFFC487A , 32'hFFFDC5E8 , 32'hFFF9B394 , 32'h00003818 , 32'hFFFC68E7 , 32'hFFFD7810} , 
{32'hFFF9E442 , 32'h000B5637 , 32'h0002BEE5 , 32'hFFFEEAD7 , 32'hFFFE067C , 32'h0006F88A , 32'hFFFFE1AE , 32'h00004411 , 32'h00014908 , 32'h000124EB , 32'h0007C795 , 32'h0003A86B , 32'h0003A41B , 32'h0000CF8E , 32'h00067254 , 32'hFFF49554 , 32'hFFFF9B54 , 32'h0003E2D3 , 32'h00034152 , 32'h00011AF6 , 32'hFFF9FDEB , 32'hFFFFCF23 , 32'hFFF8C0BF , 32'hFFFEEECF , 32'hFFFE3CC8 , 32'h0004FD31 , 32'hFFFCB57C , 32'h000159A7 , 32'h00017A39 , 32'hFFFBEB94 , 32'hFFF9AE21 , 32'h0003BB64 , 32'h0004B789 , 32'hFFFF37A1 , 32'hFFFC89FC , 32'h000637D4 , 32'hFFFA5520} , 
{32'h0001D35C , 32'hFFFD09B0 , 32'hFFF6C461 , 32'hFFFF81FA , 32'h0003D94D , 32'hFFFF3802 , 32'h0005A25B , 32'h00094851 , 32'hFFF53B0D , 32'h00074535 , 32'h0006CACE , 32'hFFFF24BF , 32'hFFFF3703 , 32'hFFFB37BE , 32'hFFFEC273 , 32'h00069242 , 32'h00003592 , 32'h0004D20F , 32'h0000600F , 32'h0009CA5A , 32'hFFFC6369 , 32'hFFFDE50D , 32'hFFFC1214 , 32'h00028B6B , 32'h000215C2 , 32'h0005D6EC , 32'hFFF716B6 , 32'hFFF90452 , 32'hFFF4B07A , 32'hFFF8E38D , 32'hFFFE9601 , 32'h00027430 , 32'hFFFF3C51 , 32'h000AE5E4 , 32'h00060CEE , 32'h000826FE , 32'hFFFC4042} , 
{32'h00065442 , 32'hFFFF758A , 32'h0002779F , 32'h0002974D , 32'h00002580 , 32'h00009F57 , 32'h0004FF92 , 32'h00027F67 , 32'hFFFD1E44 , 32'h00001D2B , 32'h00041ED9 , 32'h00003CEB , 32'h00005A08 , 32'hFFFD3674 , 32'h0000A8BD , 32'hFFFD99AE , 32'h00035562 , 32'h0003D41F , 32'hFFFD6614 , 32'h00019A7E , 32'hFFFC2F05 , 32'hFFF98BB6 , 32'hFFFB7703 , 32'h00014A80 , 32'h00002F4E , 32'hFFFB3358 , 32'hFFFD10FA , 32'hFFFE8ECB , 32'hFFFDD15D , 32'hFFFBFC10 , 32'h00060B49 , 32'hFFFB2EB0 , 32'h000104A9 , 32'h0002625B , 32'h0005F679 , 32'h00000AFB , 32'hFFFB99D9} , 
{32'h00F492FC , 32'h07D08200 , 32'h046D47A0 , 32'h064C1560 , 32'h04BF5118 , 32'h03A215C4 , 32'hF47A81A0 , 32'hFDE3AB18 , 32'h05482438 , 32'hFF901F99 , 32'h016F7F4C , 32'h03DD8BF0 , 32'hFBA6BB28 , 32'h0D819260 , 32'hF83EFF50 , 32'h02ED0B94 , 32'h08BC7F80 , 32'hF0AF7C80 , 32'h090407E0 , 32'h054B6658 , 32'hF88FA5D0 , 32'hF8D25078 , 32'h00445386 , 32'h00473BCF , 32'hFE775D08 , 32'h052F1D90 , 32'h0C0C8BA0 , 32'h054802A0 , 32'h054548F0 , 32'hF1274A00 , 32'hF9740958 , 32'hFE303D80 , 32'h0257DBAC , 32'h03952478 , 32'hFC44BE1C , 32'h00BDBDD7 , 32'h001F4D99} , 
{32'h006F20D7 , 32'hFE9D3DC4 , 32'hFC7048F4 , 32'hFF9196CD , 32'h0377261C , 32'h14A85D60 , 32'hFC4BD230 , 32'hF94AB960 , 32'h140F17E0 , 32'h056B0618 , 32'h04070F50 , 32'h025E2974 , 32'h01EE7DA4 , 32'h01AFB99C , 32'hFF1D8275 , 32'h0CDBFE20 , 32'hF703B210 , 32'h00B5A005 , 32'hF7B181B0 , 32'hFF84A154 , 32'h002386F3 , 32'hF3577E80 , 32'hFDB420E4 , 32'hFA1D0CA0 , 32'hF6134620 , 32'h031A90B4 , 32'hFF71FC71 , 32'hFAA41FD8 , 32'h0073C9A9 , 32'h02AD2D20 , 32'hFD0C5808 , 32'hFBF884D0 , 32'hFC5E9408 , 32'hF934E090 , 32'h0D1EDF60 , 32'h045501A8 , 32'h023F2AF4} , 
{32'h0EC7A6B0 , 32'h020D39F0 , 32'hF8AFAC20 , 32'h011D7E4C , 32'h016B069C , 32'h0DE24E90 , 32'hF08F2C80 , 32'h023A3FF0 , 32'hF65F8D20 , 32'hFF9A37D8 , 32'hF4327B70 , 32'h0728AF38 , 32'h0D4A1D60 , 32'h006C9B81 , 32'hFC9D0798 , 32'hF765BD00 , 32'h15F76320 , 32'hFE06AF74 , 32'hFF92F12E , 32'h05838880 , 32'h0320DB64 , 32'h0015F53F , 32'hFC1C68DC , 32'hF85CE5E8 , 32'hFEA1CDEC , 32'h06573B38 , 32'h1BD90740 , 32'h08E1C840 , 32'h0D7A3310 , 32'hF8A72568 , 32'hFB1253D0 , 32'h0DE0BD30 , 32'h08F20950 , 32'hFE63623C , 32'h00D3D88C , 32'hF6744580 , 32'h0659E238} , 
{32'h0ADA1010 , 32'h11B57F20 , 32'h060FC590 , 32'hE2E93540 , 32'h001C0688 , 32'h17FAB6E0 , 32'hFB40D050 , 32'h170823E0 , 32'h0E2B3440 , 32'hFA680AF8 , 32'hFD46CC8C , 32'hF141A180 , 32'h08801F80 , 32'h120DBCC0 , 32'hF33C4F00 , 32'h0A681D10 , 32'hF55452F0 , 32'hF2BC1F20 , 32'hED8FEC60 , 32'h000615A2 , 32'h1691A340 , 32'hE67C68A0 , 32'hF232B0B0 , 32'h10377560 , 32'hFFBEEC21 , 32'hE6447C40 , 32'h054D9758 , 32'hF9A3ABC0 , 32'hE923E660 , 32'hF6BB5840 , 32'hFAAC3648 , 32'hFDE8F5E0 , 32'hF7F9F770 , 32'hE8B80C40 , 32'hF7B6C510 , 32'hF3AD2110 , 32'hFF5277EA} , 
{32'h0ABE78E0 , 32'h065B8960 , 32'hF9EC8698 , 32'hEF6DA700 , 32'hFB995728 , 32'h437A8300 , 32'h10F29160 , 32'h146E4480 , 32'h1BE30F40 , 32'hB078AE80 , 32'hFC989980 , 32'h098D7690 , 32'h2F7ECA40 , 32'hFA898B98 , 32'hFA7DB8F8 , 32'hDB9730C0 , 32'h0C526990 , 32'hF5007B10 , 32'hF02811A0 , 32'h3B83F9C0 , 32'h04F51490 , 32'h40757B00 , 32'hE1F240E0 , 32'hD1D7F380 , 32'h06BDEC28 , 32'hDDCCF680 , 32'h14892EE0 , 32'h1687E780 , 32'h03B20B18 , 32'h08CB5CF0 , 32'hE521CA80 , 32'h079DBCD8 , 32'hFD762E34 , 32'h17BC7EE0 , 32'h187601E0 , 32'h1AA07080 , 32'h1563C8E0} , 
{32'h0AD20310 , 32'hFF66D8CE , 32'hFAD1A770 , 32'hE4BE1A80 , 32'hF3791960 , 32'h29A6C500 , 32'hE471EF80 , 32'h08EE47F0 , 32'h1F153120 , 32'hF9755540 , 32'hF366DD50 , 32'hFEAFB0F0 , 32'h041829D8 , 32'hEED9CB80 , 32'h17229FE0 , 32'h29156A80 , 32'hE5032A60 , 32'hF90204C8 , 32'hF41C01F0 , 32'h0D1ADA60 , 32'hEBDE9080 , 32'hF182FE10 , 32'hD87FA1C0 , 32'hFD577978 , 32'hD9FD79C0 , 32'h0C739020 , 32'h0B493D80 , 32'hE5D5F240 , 32'hFAE95010 , 32'h20526B40 , 32'hF969BCE0 , 32'hFC402090 , 32'hFCBFA8A0 , 32'hFADEE208 , 32'hF9124910 , 32'h1C956E40 , 32'hF67280D0} , 
{32'h03CC5AB8 , 32'h1A0A8FA0 , 32'h1AD88780 , 32'hEE66CCC0 , 32'h07805DA0 , 32'h192D7840 , 32'hE26692A0 , 32'h0F5DCE10 , 32'h2D1C7A80 , 32'hFC404F14 , 32'hE62F1DE0 , 32'hFE78D088 , 32'hFB39B268 , 32'hD4D27A00 , 32'h27B46740 , 32'h30DC7CC0 , 32'h01BB5D14 , 32'h06BCB240 , 32'hCCC7A8C0 , 32'h152F8140 , 32'hF32BBD40 , 32'h0C263150 , 32'hDCA39840 , 32'hDB99F440 , 32'hD81A0400 , 32'h13B41D00 , 32'h0BA47660 , 32'h08493940 , 32'hE3347940 , 32'hFC127C48 , 32'h091CC850 , 32'h1D2B0800 , 32'h0A397C70 , 32'hF667A240 , 32'hD1DCCF40 , 32'h0EEA1F30 , 32'h1C73B240} , 
{32'h03FDC75C , 32'hFBF3E9B8 , 32'hF317C790 , 32'hE27FA0E0 , 32'h06C77268 , 32'h04CAE390 , 32'hD1928B40 , 32'h050BE218 , 32'hEB3B51E0 , 32'hE6E02CA0 , 32'hFF0D55B9 , 32'hFE2E51A4 , 32'hF1769AB0 , 32'hEB020380 , 32'h10533D60 , 32'hFE7D9B64 , 32'h03015E38 , 32'hF95B9BA8 , 32'hF19D7660 , 32'h0FD6B3B0 , 32'hFE99C4B0 , 32'h02FA8FF8 , 32'hF6BAE9F0 , 32'h102A6820 , 32'hFD7A6590 , 32'h0B6C59E0 , 32'h03E96EDC , 32'hD929B040 , 32'h1D5D2E40 , 32'hFFEBB278 , 32'hF74E9240 , 32'hF82E7908 , 32'h11D576A0 , 32'h06033550 , 32'h13F0FC00 , 32'hFD27052C , 32'hF7758510} , 
{32'h11E743E0 , 32'h0923D740 , 32'hFAC7AF60 , 32'hE7638180 , 32'hFC5C6D5C , 32'hFE0818D4 , 32'hE63037A0 , 32'h134087C0 , 32'hDDD5A500 , 32'h1230E100 , 32'h0B6D7D40 , 32'hFDF18BF8 , 32'hF21E2C50 , 32'hDB7FD940 , 32'h133ECC60 , 32'h1C4F0420 , 32'hFDD87E88 , 32'hFD2EEB30 , 32'hFCB4A6AC , 32'hF372DCC0 , 32'hE7CE0680 , 32'h0371C924 , 32'hF8A9C218 , 32'h092BF8F0 , 32'hE4571280 , 32'hE52DA1C0 , 32'hF74200F0 , 32'hCDBB0E00 , 32'h01CCA220 , 32'h171C41C0 , 32'hF80D5D88 , 32'h09DAC560 , 32'h0D044700 , 32'h1492DE20 , 32'h22FBE580 , 32'hEE0034A0 , 32'h0A10EA10} , 
{32'h25D01280 , 32'hEBEE2C20 , 32'h02BC7E38 , 32'hDB3A9600 , 32'hEB3F6500 , 32'hCA7186C0 , 32'hFDD4D7F8 , 32'h1849C3A0 , 32'hC2CBC900 , 32'hE3D976C0 , 32'hFCDA02D0 , 32'h08EF2A50 , 32'hED476220 , 32'hEA24C820 , 32'hFC24447C , 32'h0C485000 , 32'h131D2240 , 32'h045382D0 , 32'h229C9E40 , 32'h1349A400 , 32'hE8226B80 , 32'h1185DDA0 , 32'hF32F7190 , 32'h107888A0 , 32'hF3117D50 , 32'h0A03A240 , 32'h00B9786D , 32'hF75BE990 , 32'hED79A380 , 32'h012B3798 , 32'hD5763200 , 32'h00006F25 , 32'h10895BC0 , 32'hE7C16300 , 32'hF5984C70 , 32'h14AA3A20 , 32'hFD988DB4} , 
{32'h04BE9E88 , 32'hEF6BA7C0 , 32'h1DAECE20 , 32'hF9855F78 , 32'hFBC460C0 , 32'hD3802180 , 32'hFFA978B3 , 32'h30E9FD80 , 32'hBCDA2880 , 32'hAD4FB000 , 32'hF0092E80 , 32'h0222FA88 , 32'h13434980 , 32'hF6969710 , 32'h01C22534 , 32'hE3E9B8A0 , 32'h24881A40 , 32'h0FE88650 , 32'h00DECCB1 , 32'h24AFEE80 , 32'h0E495B10 , 32'h06FA46B0 , 32'hEFF0EB80 , 32'h02F53E30 , 32'hF55A6A50 , 32'hECAF2560 , 32'hC8A62700 , 32'h080BC830 , 32'h0936C2B0 , 32'h1FA85F00 , 32'h21363680 , 32'h0BC0D600 , 32'h1E54F7C0 , 32'hDE712580 , 32'h14709DA0 , 32'h08DB9E60 , 32'hFB098928} , 
{32'hFF8F69C6 , 32'h02A0BB9C , 32'h1DC55720 , 32'hD8CBF440 , 32'hFE336294 , 32'h072686C0 , 32'hFDDE14F0 , 32'hD57AEE40 , 32'hDA6F2280 , 32'hA89B2980 , 32'hEB676C20 , 32'h1CAE9180 , 32'h262422C0 , 32'h17EF7420 , 32'hEB61CD80 , 32'hFF8710EA , 32'hE581AD20 , 32'h1C53BE60 , 32'hF9C602F0 , 32'h2BE98D80 , 32'h037952EC , 32'hF91591C0 , 32'hEE149640 , 32'hEB1B5920 , 32'h155BBC80 , 32'h0D822000 , 32'hE3847400 , 32'hEDFCC740 , 32'h04AC3958 , 32'hE5789D00 , 32'h0E98A460 , 32'hEE35E0E0 , 32'h0DEFEDD0 , 32'hEBCF4A60 , 32'hD11BC6C0 , 32'h03AA6530 , 32'h06E702E8} , 
{32'h1A48B760 , 32'hEAA35BC0 , 32'h17DFED20 , 32'hD317E540 , 32'h02F9FF14 , 32'h256E9800 , 32'h1BD149C0 , 32'hB1595A00 , 32'h09E41740 , 32'hBB534200 , 32'hF0AECB60 , 32'h0BACBD70 , 32'h2F65FB00 , 32'h0AD90080 , 32'h04E4A900 , 32'hEE738640 , 32'hCC6DAD40 , 32'h25425500 , 32'h080E8FA0 , 32'h0B4B3DC0 , 32'h133C9C40 , 32'h04CF52E0 , 32'hE54AE420 , 32'h22343F80 , 32'hF9CC2FB0 , 32'h19177A20 , 32'hC216FD80 , 32'h194E4F20 , 32'hE3483BC0 , 32'h16972260 , 32'hF9821DC8 , 32'hEA7923E0 , 32'h1FC95E20 , 32'h0A108000 , 32'h008D5614 , 32'hC5268180 , 32'h24EDC840} , 
{32'h0BABF000 , 32'h12578280 , 32'h1549B4E0 , 32'hB9171980 , 32'h03FBFF84 , 32'h1FE7E320 , 32'hFFCA02A5 , 32'hA6CA6380 , 32'hF6275D60 , 32'hE1A28EA0 , 32'h0CB3F660 , 32'hF7A92610 , 32'hFDFEDA18 , 32'h0A2D6E40 , 32'hFD611A84 , 32'h0514F078 , 32'h002AFDF7 , 32'hF9891DE0 , 32'h1D5F7300 , 32'hF52A64A0 , 32'hF0919E20 , 32'hEA285A20 , 32'h0BABF1A0 , 32'hED9D4560 , 32'h02AE73EC , 32'hE947F6E0 , 32'hF031AA60 , 32'hF5CF5DD0 , 32'hEE80CCA0 , 32'hFD473DDC , 32'hFC012990 , 32'hF36259F0 , 32'h1DAB2C80 , 32'h09AE15D0 , 32'hF2D299D0 , 32'hED6E63E0 , 32'h0E04C5B0} , 
{32'h13D17940 , 32'h201A53C0 , 32'h243A9840 , 32'hA47FBF80 , 32'h202B0F80 , 32'h191E44A0 , 32'hF302F8A0 , 32'h9F7D1D00 , 32'hFBD59E20 , 32'h38450200 , 32'h27F73840 , 32'hF7C55590 , 32'hEF162AC0 , 32'hEA9E65E0 , 32'hFFDDCC3B , 32'hFF564692 , 32'hFB97C1B0 , 32'h01595D08 , 32'h18C73200 , 32'h0AD62520 , 32'h02BEB68C , 32'h0670C228 , 32'hF2B042E0 , 32'hE49A2BA0 , 32'h0C2C29B0 , 32'h011975DC , 32'hFD288828 , 32'h0516DB48 , 32'h07520E80 , 32'hF9F9A2F8 , 32'hE85EFAA0 , 32'hF22FE970 , 32'h0855DC30 , 32'h1536DD20 , 32'hF63C6610 , 32'hF6375F90 , 32'h0B3C80B0} , 
{32'h0A63F060 , 32'h109D5640 , 32'h040C93C8 , 32'hC6E34240 , 32'h077FDF10 , 32'h13A23720 , 32'hF738EFB0 , 32'hDE481480 , 32'h01BD7B90 , 32'h30396F80 , 32'h2EF53AC0 , 32'hFB3AC438 , 32'hFB76E5F8 , 32'h0B0DC380 , 32'h08C43BD0 , 32'hEF079B20 , 32'hEF2425C0 , 32'h03C0E7E0 , 32'h1345C360 , 32'hFEE88FB0 , 32'h14108440 , 32'h2F719C80 , 32'hDA6358C0 , 32'hFCEAC740 , 32'h09D2B780 , 32'h00FB5190 , 32'hFFC38DB8 , 32'h1490D880 , 32'hF5DF37E0 , 32'hFE021300 , 32'hF4C4BE60 , 32'hFC6D6D5C , 32'h1096A420 , 32'h2806DC40 , 32'hF477F1F0 , 32'hF073F680 , 32'hFCCFBFD4} , 
{32'h140B7F40 , 32'h1B1C4680 , 32'h1E742F20 , 32'hD6D43D40 , 32'h1F65C7E0 , 32'h0DBE9450 , 32'hFF640018 , 32'hD61E0B80 , 32'hED8E1700 , 32'hE976A3E0 , 32'h1729ED60 , 32'h2901EBC0 , 32'h08DC4AC0 , 32'h0A6A3650 , 32'h1092F220 , 32'h01A61B20 , 32'hFB0EBC90 , 32'h101AA9E0 , 32'hFFD1FC79 , 32'hF5B65A90 , 32'h14FB4260 , 32'hFDA6648C , 32'hF8636C60 , 32'h03178680 , 32'h1DDE7000 , 32'h0C87DD30 , 32'hF5818A20 , 32'hF1E01730 , 32'h113BBD60 , 32'h072D3710 , 32'hF63E16F0 , 32'h0556D0D8 , 32'hFD416CA8 , 32'h0EA75B50 , 32'hDD4BA580 , 32'hF0F3BE20 , 32'hF71D9F40} , 
{32'h08C54290 , 32'h0427F2C0 , 32'h0834CC10 , 32'hF688EF00 , 32'h0B486010 , 32'hE6D6E9C0 , 32'h15422320 , 32'hEE6D4CE0 , 32'hEE381E00 , 32'h1D1AA940 , 32'h1F0E2E40 , 32'h12E7EBA0 , 32'h1036E7A0 , 32'h15E52C40 , 32'h01FA028C , 32'hFD03B448 , 32'hF75AB980 , 32'h0509D138 , 32'hF363CF90 , 32'hF1B76440 , 32'hF6024E40 , 32'hFB573A90 , 32'h15688880 , 32'hFF98EFF6 , 32'hFBC1CD98 , 32'h10645AC0 , 32'h0DC26530 , 32'h1262C4E0 , 32'hE466E2A0 , 32'hFD36E0BC , 32'hDF22B980 , 32'hFB968308 , 32'hFACC6F70 , 32'h06D1B1A8 , 32'hF3197980 , 32'hFFBC4981 , 32'hFFED4BF7} , 
{32'h0C90EFC0 , 32'h17F66CE0 , 32'h09958B00 , 32'hC700FCC0 , 32'h038E5D38 , 32'hFFA39D6B , 32'hFAB51870 , 32'hF99337D0 , 32'hDB818680 , 32'h0A879120 , 32'hF7CAE250 , 32'hF066C1C0 , 32'h11E205A0 , 32'h14D48000 , 32'hFC535F18 , 32'h089216C0 , 32'hDD7D6740 , 32'hF38C8CB0 , 32'h0E453EF0 , 32'h0B915D20 , 32'hEA89B7E0 , 32'h0893BEC0 , 32'h01411C4C , 32'hFE339840 , 32'hFFFC5014 , 32'hF7F022A0 , 32'h040DC990 , 32'h01EF9C50 , 32'hEF83E260 , 32'h1316CA60 , 32'h0AB3AA20 , 32'h09731A10 , 32'h31A6E1C0 , 32'h065358A8 , 32'h0661F118 , 32'h096C20D0 , 32'hD5B25640} , 
{32'h13043120 , 32'h03A9517C , 32'h131E5220 , 32'hE67C3C60 , 32'h114D2040 , 32'h0737D150 , 32'h02987970 , 32'hE575F180 , 32'hEB30F560 , 32'hFC9F8080 , 32'h2340E600 , 32'h0A7AFE80 , 32'h0F8B2650 , 32'hF59753E0 , 32'h19B02120 , 32'h1261EB00 , 32'hF196E120 , 32'h062D1DB8 , 32'hFD6EC728 , 32'hF3C55340 , 32'h0DB914E0 , 32'h02C53724 , 32'h017B7B3C , 32'hF137D360 , 32'h068DF070 , 32'h07C7AAA8 , 32'hFD89D0DC , 32'h0F8665C0 , 32'h11EE3DA0 , 32'hF9E4F708 , 32'hFBD66DA0 , 32'h0AE8C820 , 32'h02B845D0 , 32'h015DD724 , 32'hECF7DA60 , 32'hF04C0440 , 32'hD8E69D80} , 
{32'h085FEB10 , 32'h02A7B8EC , 32'h0FF8D2C0 , 32'hF376D2D0 , 32'h0D147520 , 32'hFB1FA3D0 , 32'hFC7C21E8 , 32'hF2B968A0 , 32'hEDA7D040 , 32'h03FB9C20 , 32'h3236B380 , 32'h1C634EC0 , 32'h30B23200 , 32'h0D7EB610 , 32'h0D003F00 , 32'h0415A340 , 32'hECA49BC0 , 32'h05DA0D60 , 32'hEBA36FA0 , 32'hF23BEA70 , 32'h04933CC8 , 32'hEC6F1A00 , 32'h031F3220 , 32'hF5570B90 , 32'hF5B4B1F0 , 32'h092547D0 , 32'hF30D1840 , 32'h1F0B8640 , 32'hEC18CF80 , 32'h05B90A48 , 32'hDDEE18C0 , 32'hED29D5C0 , 32'h188FC1C0 , 32'h06DE9248 , 32'hF13C8C90 , 32'hF54A2080 , 32'h0415ABD0} , 
{32'h01FE83EC , 32'h007AEF2F , 32'hFD5AAEC4 , 32'hFDA87894 , 32'hFF4E0F8B , 32'hFCB50BB4 , 32'h060DFEE8 , 32'hFCFE4828 , 32'hFF5F3124 , 32'hFE4D9584 , 32'h0A6C5B90 , 32'h0A989B00 , 32'hFDFB3924 , 32'h0010D9E3 , 32'hF9240A10 , 32'hFF791A01 , 32'hFC25D504 , 32'h084CE390 , 32'hFEA1A168 , 32'hFFB964AC , 32'hF26726B0 , 32'h0153A5C4 , 32'hFE884930 , 32'hFC664BF8 , 32'hFCF15EB0 , 32'h04EA3720 , 32'h01A7EDE0 , 32'hFD31C89C , 32'hFCF00D2C , 32'h03EF7A34 , 32'h045047B0 , 32'hFCB02968 , 32'hFE550D60 , 32'hF62EFCE0 , 32'hFDDC02DC , 32'h096103A0 , 32'hEECAA1C0} , 
{32'h000376AB , 32'h00068A11 , 32'hFFFF3DFF , 32'hFFFFD8C9 , 32'hFFFC8361 , 32'hFFFFEDF3 , 32'h0001C63A , 32'h000766DE , 32'h0004BCF6 , 32'h00017059 , 32'hFFFE83A1 , 32'h00020F57 , 32'hFFFCC22C , 32'h0001A02E , 32'hFFFCE840 , 32'hFFFD63CE , 32'h0000A8BB , 32'h0003872B , 32'h0003C315 , 32'hFFF52626 , 32'hFFFFEB13 , 32'h0002B902 , 32'hFFF31D4E , 32'h00017AA7 , 32'hFFFB9F0B , 32'hFFFDFADD , 32'h00053BBA , 32'h00032B1D , 32'h00029815 , 32'hFFFD7B99 , 32'hFFF86DF8 , 32'h00045C2A , 32'hFFFAD4E6 , 32'hFFFB1D3A , 32'h0000FCDE , 32'h00040216 , 32'h00035660} , 
{32'h0000E98F , 32'hFFFFB70C , 32'hFFFE45F2 , 32'hFFFF954B , 32'hFFFD2C01 , 32'hFFF564D7 , 32'h000B5B8B , 32'hFFFD9DB8 , 32'hFFFE07B6 , 32'h000413D0 , 32'h00001956 , 32'hFFFFFF21 , 32'hFFF9BE44 , 32'h00027632 , 32'h00072F54 , 32'h00038470 , 32'h000550CC , 32'h00040FF3 , 32'hFFFD8B18 , 32'h0004EED3 , 32'h00014AA4 , 32'hFFFAD179 , 32'hFFF4D45E , 32'h0001F262 , 32'hFFF9E4EC , 32'hFFFEFB70 , 32'h000249EA , 32'hFFFD4A22 , 32'h0009E606 , 32'h000550C4 , 32'hFFFBEF66 , 32'h000261E3 , 32'hFFF9FB1B , 32'hFFFEC6D8 , 32'h00082438 , 32'h0005F6C3 , 32'hFFFCE83B} , 
{32'hFFF84CC7 , 32'h000118E9 , 32'h00053CFE , 32'h000691DF , 32'h0002DD19 , 32'hFFFD37B5 , 32'hFFFEE8F3 , 32'h0003606A , 32'h000A9F2F , 32'h000182D1 , 32'hFFFEFAED , 32'h0002938E , 32'hFFFD9095 , 32'hFFFE6F67 , 32'h00020353 , 32'hFFFCB31F , 32'h0002C0FB , 32'h000315ED , 32'h000B3969 , 32'hFFFDDE85 , 32'hFFFEB4A7 , 32'h0005CFA8 , 32'h000456B2 , 32'hFFF652B1 , 32'hFFFFABB1 , 32'hFFFD1405 , 32'hFFF9D230 , 32'hFFFECBE9 , 32'hFFFEBEB5 , 32'hFFF70346 , 32'h00078578 , 32'hFFF53569 , 32'h00061681 , 32'h0002AEF8 , 32'h00093029 , 32'hFFFF83FD , 32'hFFFB74F7} , 
{32'h000795D5 , 32'hFFFD21A2 , 32'h0001EEA7 , 32'h0001BAF8 , 32'hFFFD2A63 , 32'h0000715C , 32'hFFFD2141 , 32'h0001FAC3 , 32'hFFFD3F0F , 32'h0004538D , 32'h00097FEB , 32'h0003709A , 32'h00034961 , 32'hFFFDD1F0 , 32'h0001223E , 32'hFFFCF613 , 32'hFFFE67A4 , 32'hFFFD67B1 , 32'h00069173 , 32'h000D14E0 , 32'h000D2B7B , 32'hFFF60EFF , 32'h000507F1 , 32'hFFFE6765 , 32'h00056E84 , 32'h0002E035 , 32'hFFF9E454 , 32'hFFF925F1 , 32'h00095F70 , 32'h0000AE80 , 32'hFFFF8A3D , 32'hFFFCDCBE , 32'h0000705F , 32'h0004FC00 , 32'hFFFD7FB2 , 32'h000149AF , 32'h00046E64} , 
{32'hFFF9FB8B , 32'hFFFA97B9 , 32'hFFFF193B , 32'h000072D9 , 32'hFFF8FA54 , 32'hFFFF1100 , 32'hFFF79003 , 32'h00015695 , 32'hFFFE6E3E , 32'hFFFA40EF , 32'h00016BD1 , 32'h0002F116 , 32'hFFFF1B5B , 32'hFFF5DB3A , 32'h0004D2A2 , 32'h00013E54 , 32'h00035614 , 32'hFFFCCA40 , 32'hFFFDA752 , 32'hFFFBFA15 , 32'h00060BEE , 32'h0002EA5A , 32'hFFFBED75 , 32'h0000B65F , 32'h0005374E , 32'h000552C1 , 32'hFFFC1C33 , 32'h000124A4 , 32'hFFFC7347 , 32'hFFFC6750 , 32'h0000B784 , 32'hFFFE5B50 , 32'h0000E1AF , 32'h00067FC2 , 32'hFFFD22E3 , 32'hFFFB4BE4 , 32'hFFFE2C12} , 
{32'h0000F09E , 32'hFFFBBF3A , 32'h0000B444 , 32'hFFF84026 , 32'h000904CC , 32'hFFEEC331 , 32'h00041882 , 32'hFFFB8A00 , 32'h000247F6 , 32'h0005675F , 32'hFFFF0C34 , 32'hFFF93F72 , 32'hFFFD346E , 32'hFFF36A43 , 32'h0002AB81 , 32'hFFF64A88 , 32'hFFF9B2EE , 32'h00088A50 , 32'hFFFF4739 , 32'h00042588 , 32'h0002C1CD , 32'h00036FAD , 32'h000109B0 , 32'h0009A9FF , 32'hFFFF8766 , 32'hFFFD1E23 , 32'hFFFB46DB , 32'h000C2D87 , 32'h0003D804 , 32'hFFF87327 , 32'h000CEC99 , 32'h0003263E , 32'h0003ADA1 , 32'h0001EF6F , 32'h000871F0 , 32'h00067E7B , 32'h0007D274} , 
{32'h0045C625 , 32'hFF7F1F1F , 32'hFFFE00DA , 32'h000B27C8 , 32'h00562F81 , 32'hFFF1335A , 32'hFFD00313 , 32'h00397100 , 32'hFFB6B096 , 32'hFF828258 , 32'hFFEEF397 , 32'h005CF486 , 32'hFFFD4355 , 32'hFFC60350 , 32'hFFEA6F3E , 32'hFFC63904 , 32'h009F7B9A , 32'hFFC606D5 , 32'hFF9C4173 , 32'h0022DCD7 , 32'hFFC1EA3A , 32'hFFECC3EE , 32'hFFF049F6 , 32'h006996A8 , 32'hFFC4DFE8 , 32'hFF94B51F , 32'h0005E629 , 32'hFFF18E2D , 32'h002CD15E , 32'h006F18A9 , 32'hFFF0340F , 32'h001C1586 , 32'h005DC929 , 32'h0007CC00 , 32'h003FD79E , 32'hFFE83BC6 , 32'hFFBE6CFE} , 
{32'h0C8F3020 , 32'h10C1D4A0 , 32'h0C38E030 , 32'h084831F0 , 32'h1196A3E0 , 32'hFF607073 , 32'hF1994560 , 32'h049BF3A8 , 32'hFE01E0A0 , 32'hF98C7608 , 32'hFAE96728 , 32'h07506890 , 32'hF8279818 , 32'h0CB03A10 , 32'h020C474C , 32'h05578F68 , 32'h06901A18 , 32'hE5A4D0C0 , 32'h00A362D4 , 32'h0F018350 , 32'hF4E25BE0 , 32'hF7840CC0 , 32'h03CC7790 , 32'h083B0820 , 32'h03E35ABC , 32'h0B845720 , 32'h090AE4B0 , 32'h16834980 , 32'h11D35080 , 32'hEBD2E380 , 32'hF9695898 , 32'hFCC9D524 , 32'h0AFCA090 , 32'h05D6CF10 , 32'h03AA74F4 , 32'hF8BDFA20 , 32'hF5213C40} , 
{32'h0785EFB0 , 32'h061930E8 , 32'hFF4DFDB6 , 32'hF7791BF0 , 32'h018011D0 , 32'hFA336A08 , 32'h0084E865 , 32'h09102580 , 32'h005008D0 , 32'hF8665938 , 32'h07DAA8D0 , 32'hF8B108D8 , 32'h06054130 , 32'hFEBED94C , 32'hF6BCB5D0 , 32'hFF7EF2EC , 32'hF9CBDC78 , 32'hF6D0C4B0 , 32'hFA10C790 , 32'hFB8991D0 , 32'h00C54FE3 , 32'hFCE78188 , 32'h02C6A5C0 , 32'h01439918 , 32'hFB3619D0 , 32'h049537C0 , 32'h040B5AF8 , 32'h0AE83760 , 32'h1695FB40 , 32'hF0D6CBA0 , 32'h094CCB90 , 32'hF4653C80 , 32'h04E84E50 , 32'h01B43B80 , 32'hFBD2B818 , 32'h01B36EE4 , 32'hFED59360} , 
{32'h16FAF6A0 , 32'h131D5BE0 , 32'h05312D60 , 32'hFB8B6500 , 32'hFB015968 , 32'h1151B740 , 32'hFE9576A4 , 32'h07E3BD10 , 32'h1162F060 , 32'hE7202220 , 32'h064A5998 , 32'h132D1580 , 32'hF985D2B8 , 32'hFFDD5181 , 32'hEAFD2920 , 32'h1C13CB20 , 32'h16107A00 , 32'hEAB01300 , 32'hF58B0460 , 32'h0FBCB3F0 , 32'hFCFC8E70 , 32'h35E117C0 , 32'h02F5CF34 , 32'h05C08678 , 32'hFF860E6A , 32'hF25254F0 , 32'hFC3FE360 , 32'h11A5A9C0 , 32'hFF99D115 , 32'h04AC6C80 , 32'h0089109F , 32'hE7C63D60 , 32'h123B2120 , 32'hFFD39C73 , 32'h0E2DF530 , 32'h0B701640 , 32'h070C09C8} , 
{32'h0459B390 , 32'h084BD890 , 32'hF7EAFE80 , 32'hF63E41F0 , 32'hF4D31050 , 32'h1EE34460 , 32'h006825BF , 32'h06146E68 , 32'h0D29B510 , 32'hE83F92A0 , 32'hEF74ED80 , 32'hF6A5C790 , 32'h100A7A40 , 32'h065DB448 , 32'hFF3D2C20 , 32'hF56A64D0 , 32'hFE16AFD0 , 32'hFD1E00BC , 32'hF8208BD8 , 32'h0E3A99E0 , 32'h11B6F300 , 32'hFF1386AD , 32'hE34BB560 , 32'h10D126E0 , 32'h065E7920 , 32'h025E36DC , 32'hF616DD70 , 32'h078E2FC8 , 32'h0974C750 , 32'hFC486214 , 32'h05442478 , 32'h01892910 , 32'h014CE514 , 32'hFCBA3968 , 32'h0655BB10 , 32'hFB5129A8 , 32'hFE18BAF0} , 
{32'h11A6EA40 , 32'hF9229748 , 32'hF34D7C90 , 32'hFA883440 , 32'hF96405C0 , 32'h2BEC7880 , 32'hEDD29DE0 , 32'h02EABFD8 , 32'h0AFE12D0 , 32'hFF8F3A6C , 32'h0AA2DBD0 , 32'h04916708 , 32'hFF6C50A6 , 32'h024FB968 , 32'hF98C4970 , 32'h0752E088 , 32'hF24D65E0 , 32'hFA648A38 , 32'hF43974F0 , 32'h0C8E67D0 , 32'h009CC31E , 32'hF9A22C68 , 32'hF9BCDBF0 , 32'hEC1C6320 , 32'hEE91C2E0 , 32'hF862DC50 , 32'hF52DBA40 , 32'hFB1F1BC0 , 32'h06A00F48 , 32'h09168A00 , 32'h0D28F1F0 , 32'hF8C74618 , 32'hEF0B2600 , 32'h0375E090 , 32'h09ABE8E0 , 32'h07C98488 , 32'h0536D680} , 
{32'h48C09A00 , 32'hE5035500 , 32'hECC24920 , 32'hEB0709E0 , 32'hD4FA9CC0 , 32'h48829500 , 32'hED1E14E0 , 32'h2DE7F040 , 32'hF97EF920 , 32'hF8A13F38 , 32'h2EDCE180 , 32'h0B638AB0 , 32'hEF0E5BA0 , 32'hF50CF540 , 32'h330D94C0 , 32'h179172A0 , 32'hD6CB0000 , 32'h03788B60 , 32'hDCBD7280 , 32'h2EDBEC80 , 32'h09040F50 , 32'h294B5E00 , 32'hEE4486E0 , 32'h0F559D40 , 32'h0425C328 , 32'h04BF6748 , 32'hD3006080 , 32'hF3E8D210 , 32'h2F638D80 , 32'hFF542582 , 32'h2AF0C300 , 32'hD7D14F40 , 32'h03C9C504 , 32'h1A2EAE00 , 32'hD88A2380 , 32'hF13C4210 , 32'h0DE7CF00} , 
{32'h2A137040 , 32'hF78BEDC0 , 32'hE0734C80 , 32'hF974B9B0 , 32'hF09A4D50 , 32'h31521400 , 32'hDB297C40 , 32'h0B116930 , 32'hE1786620 , 32'h31F5F700 , 32'h0D8B7120 , 32'hFAB5A238 , 32'hFE8667A4 , 32'hFDC11DE0 , 32'h1F2DC000 , 32'h378B1300 , 32'hD31D8A40 , 32'h16C9A660 , 32'hEC0181C0 , 32'hF8193270 , 32'h00DE89DC , 32'h0D3344A0 , 32'hE8C95660 , 32'hF25CB540 , 32'hF5ABEED0 , 32'h40202280 , 32'h0DE32E60 , 32'h13011660 , 32'h12B06720 , 32'hF4609E60 , 32'h1A6F8380 , 32'h17B64560 , 32'hFD3E6828 , 32'hF345CB20 , 32'hDE393680 , 32'hFE48FCC8 , 32'h17D28F40} , 
{32'h53648000 , 32'hFFD53412 , 32'hFA7FFE38 , 32'hFC4EF0F0 , 32'hF8709788 , 32'h2B57A640 , 32'hC9CB0440 , 32'h294B67C0 , 32'hC2029C80 , 32'h2E51AE40 , 32'hF1E7AF10 , 32'hF1F58610 , 32'hF41A6FF0 , 32'hFCD9DAD8 , 32'h3616FB00 , 32'h0855CB50 , 32'hF8551868 , 32'h104EAB40 , 32'hF2AD9A70 , 32'hD7F7B2C0 , 32'hECCE4EE0 , 32'h1FDEAC20 , 32'h0B2E0E30 , 32'h453CD800 , 32'hEB2FC8C0 , 32'hFC3106AC , 32'h393B62C0 , 32'hF1E77CD0 , 32'h2D440F80 , 32'h2B984440 , 32'h0739AEE0 , 32'h02068AFC , 32'h051BD7C0 , 32'h045F3FF8 , 32'hF96690A0 , 32'hDCA6E840 , 32'h4F2CC280} , 
{32'h737C2F00 , 32'hC63A8E40 , 32'h148F4760 , 32'hFD32E640 , 32'hFEE781E4 , 32'hF3CC02A0 , 32'hE3015D60 , 32'h3185E000 , 32'h9D9C5880 , 32'hF3FA1CC0 , 32'h152CC100 , 32'hF14CEE80 , 32'hEA151B80 , 32'hE6AADA80 , 32'h174DE500 , 32'hFEF6C7E8 , 32'h19DE1280 , 32'h1B54EE00 , 32'h20FCAD40 , 32'hE7B72060 , 32'h1B042280 , 32'h1662C5C0 , 32'h06BCB868 , 32'h1E3D6DE0 , 32'h1AB25D20 , 32'h0D79A700 , 32'h0B7B2950 , 32'h1CC3ADC0 , 32'hFFD735BC , 32'hFF2AA322 , 32'h1D57C620 , 32'h2A2EC040 , 32'h04EE7480 , 32'hF247ECE0 , 32'hFA917248 , 32'h000F3818 , 32'h0B667F70} , 
{32'h78C8DB80 , 32'hC3960E00 , 32'h320AE740 , 32'hFF3AF308 , 32'h0AA8CBC0 , 32'hC5218BC0 , 32'hE9CF9CC0 , 32'h2303DF80 , 32'hC2422800 , 32'hC38AFD80 , 32'h08C97A10 , 32'h057937B8 , 32'h1A16EE00 , 32'hEC6209A0 , 32'h1C0D4780 , 32'h16D12960 , 32'h1530EBC0 , 32'h1D48E260 , 32'h04BD4EA0 , 32'h0D884BC0 , 32'h242BC540 , 32'hD33F5800 , 32'hE5D6FFC0 , 32'h0230DE3C , 32'h0DAC8B30 , 32'h20581E80 , 32'hFA28B270 , 32'h3704F640 , 32'hECAE7F40 , 32'h1498AE80 , 32'hFA3A2730 , 32'hFBA986E8 , 32'h200B2AC0 , 32'hE69AD120 , 32'h11696560 , 32'hF503FDC0 , 32'hFB7DC270} , 
{32'h3DF4B300 , 32'hCD96C400 , 32'h0E261310 , 32'hEF7E9760 , 32'h0CFE2A90 , 32'hF4BDC4E0 , 32'h1AC7E7E0 , 32'hF4A9AF50 , 32'h03E141CC , 32'hA0CB5200 , 32'hEC2B6D60 , 32'h0816CCB0 , 32'h03E7F44C , 32'h004C4FCD , 32'hFDD92D88 , 32'h141F5F80 , 32'hFC6E8BE8 , 32'h0FA6E7A0 , 32'h208D9580 , 32'h1F71D4A0 , 32'h0A6C0AD0 , 32'hD149C880 , 32'hEC732E60 , 32'h121EC020 , 32'h1A0D2E40 , 32'h1503EB80 , 32'hFCFCD938 , 32'h073C1098 , 32'hE7053EC0 , 32'hF9A5F930 , 32'hF66F6A90 , 32'h195DDF00 , 32'hFB05DFA8 , 32'hE16BAFA0 , 32'hCFBC01C0 , 32'hFC1DE530 , 32'hEEFAB5E0} , 
{32'h56A48F80 , 32'hBAFCE280 , 32'h3082A300 , 32'hB5160880 , 32'h0FD2B4A0 , 32'h04361FD0 , 32'h1E2A2A80 , 32'hC8E2B140 , 32'h401B1B80 , 32'hB5501A00 , 32'hE342AD60 , 32'hE7D88580 , 32'h05507370 , 32'hED67CAA0 , 32'hDE992B00 , 32'h18DADE60 , 32'h0BC84FC0 , 32'h0C01AA30 , 32'h43F13880 , 32'h003925C0 , 32'h33FFB0C0 , 32'hBF982200 , 32'h1679E560 , 32'hFF320E3A , 32'h0A32F980 , 32'h313ED0C0 , 32'h1F3C3620 , 32'h09BE2FD0 , 32'h08B4D240 , 32'h102EA0A0 , 32'h22586DC0 , 32'h0C386B70 , 32'hEA98AFA0 , 32'hFC6C9794 , 32'hFC4CD3A4 , 32'hFF019FEB , 32'h0A2BE1C0} , 
{32'h7FFFFFFF , 32'h984EA680 , 32'h4AC46E80 , 32'hBAB0DB00 , 32'h0D5CD170 , 32'hD971D3C0 , 32'h042DBE00 , 32'hB7DD6600 , 32'h44E18700 , 32'hCF95FD00 , 32'hEB37A760 , 32'hEEB6C080 , 32'hEFE4DB60 , 32'hEAC54B60 , 32'hFB884F08 , 32'h0DAD2460 , 32'h20C65200 , 32'hF0513650 , 32'h1B7D4F00 , 32'hEB975B80 , 32'hF4DE2ED0 , 32'hC1068200 , 32'h0C53AB30 , 32'h0BBBCC80 , 32'hEDCEA380 , 32'h0B6AC930 , 32'h10F1CFA0 , 32'hCD414240 , 32'h23FC14C0 , 32'h0B29BD20 , 32'h04D8EE28 , 32'hF0D6E470 , 32'hDDA541C0 , 32'h014F3C58 , 32'hE8F92E80 , 32'h0916CEE0 , 32'h0E70BEC0} , 
{32'h5AE7EB80 , 32'hC1B95900 , 32'h329F4140 , 32'hC0056280 , 32'h0D219ED0 , 32'hD6178200 , 32'hFD7368D8 , 32'hDD0CD3C0 , 32'h3677B880 , 32'h14EE9EE0 , 32'h08B6E240 , 32'hF73255F0 , 32'hE2437300 , 32'hFE68F794 , 32'hF413BFA0 , 32'h0152C530 , 32'h2CE16180 , 32'hFB9D9F90 , 32'h29B66740 , 32'hF36B5830 , 32'h10D89480 , 32'h01932778 , 32'h0D112610 , 32'hECF58A40 , 32'h05F4FF50 , 32'h00E35AB8 , 32'hFD2A3DE4 , 32'hED26A0C0 , 32'h0749F7F0 , 32'h1C36B5C0 , 32'hF5CDF2F0 , 32'hDBBD5F00 , 32'hFC8EDF94 , 32'h221503C0 , 32'hF6C2B690 , 32'hEC7A79E0 , 32'h29D62B80} , 
{32'h5EF12280 , 32'hAE0BA980 , 32'h3B396400 , 32'hB4553980 , 32'h1697F560 , 32'hD501C8C0 , 32'hF3F14600 , 32'hF1D79B60 , 32'h4FB39780 , 32'h39E43BC0 , 32'h11CCD5C0 , 32'hF0215890 , 32'hF482A420 , 32'h2861AFC0 , 32'h05911950 , 32'hBE4D6280 , 32'h1A41F960 , 32'h14678140 , 32'hF591B150 , 32'h2969C180 , 32'h2472A080 , 32'h2AF6F080 , 32'hD7DD9AC0 , 32'hFC3B9968 , 32'hE5BD8660 , 32'hF8AF97B8 , 32'hFAE6E590 , 32'h0E4DAD10 , 32'hF0994230 , 32'hF21A1C90 , 32'hE607A7C0 , 32'h014629E8 , 32'hEEF74AE0 , 32'hEECD41E0 , 32'h1A1977E0 , 32'hFDE6D940 , 32'hFAA4FF48} , 
{32'h653DD480 , 32'hCA6B1440 , 32'h223AFDC0 , 32'hD27C1040 , 32'h07E8C3C8 , 32'hD761F000 , 32'h07C3E200 , 32'hE24629E0 , 32'h28EC8500 , 32'h4689E380 , 32'h20397340 , 32'hEF42FD20 , 32'h0CF528A0 , 32'h433B9600 , 32'h04990330 , 32'hC296CA40 , 32'h117C13E0 , 32'hFAA393C0 , 32'hE2D8DC00 , 32'h2477AE80 , 32'hFEBDC568 , 32'h342BE100 , 32'hE5EEDC00 , 32'h0E744F90 , 32'hFB990D70 , 32'hE8A13F80 , 32'h00D2A6B9 , 32'hEF885B20 , 32'h113E9E40 , 32'hFC0A63C0 , 32'h18AA9340 , 32'h0C0DA710 , 32'h02E471A4 , 32'h0CC3C9B0 , 32'h19EBF460 , 32'hFAF10868 , 32'hF29EE3D0} , 
{32'h64970D00 , 32'hC7E5B8C0 , 32'h2413E480 , 32'hDDF629C0 , 32'hFEF128DC , 32'hD5F57A80 , 32'h0FD10CD0 , 32'hF61765A0 , 32'h2721E2C0 , 32'hF91E0C10 , 32'h02F20F1C , 32'h019506A8 , 32'h0F72E340 , 32'h3549AB40 , 32'h136694E0 , 32'hF12C97B0 , 32'h1BE60440 , 32'hF9B9D5C0 , 32'hFF8B6B3B , 32'h1754B8A0 , 32'h01A7D250 , 32'h18803FC0 , 32'hFEBB2214 , 32'hF642FFF0 , 32'h186417A0 , 32'h0B9A2030 , 32'h06CD9CE8 , 32'hE1C50F80 , 32'hF5535FA0 , 32'h0EEEEC00 , 32'h0B7CA7C0 , 32'hF841F608 , 32'h052F52C0 , 32'h0A0D3490 , 32'h034AACA0 , 32'hFC2F0300 , 32'h100ECB60} , 
{32'h42598A00 , 32'hCFC04840 , 32'h1A94F0A0 , 32'hE2136AA0 , 32'hF8DAE768 , 32'hEA0D28E0 , 32'hF6BA0710 , 32'h04DEA910 , 32'h244FC440 , 32'h0031DD91 , 32'hF23FEA60 , 32'h04DCCEF0 , 32'h09719130 , 32'h1EFFD0E0 , 32'h13362460 , 32'h13226300 , 32'h13573D20 , 32'h092D8810 , 32'h024DCAF0 , 32'h04DF9AB8 , 32'h00495061 , 32'h091FF1D0 , 32'h001D593D , 32'hF3976860 , 32'h12191560 , 32'h1B2E12C0 , 32'h147311A0 , 32'hF91106F0 , 32'hE1DD66A0 , 32'h0994BF80 , 32'h027D2590 , 32'h07E6E808 , 32'hFE103264 , 32'hF383E060 , 32'hE8096D00 , 32'h15CCB100 , 32'hF3368FA0} , 
{32'h25AD6800 , 32'hEEF61860 , 32'hFD19E6E8 , 32'hFDD3C5E0 , 32'hF6534820 , 32'hE065D180 , 32'h091A1500 , 32'h181E70A0 , 32'h0DEF0270 , 32'h11520760 , 32'h1A4AD8E0 , 32'h22ADCB00 , 32'h1A034EA0 , 32'h27432900 , 32'h08F3F7A0 , 32'hEF354E00 , 32'hEB570880 , 32'h1FEDA4E0 , 32'hCD60F2C0 , 32'h0281A88C , 32'hD16562C0 , 32'h152CE680 , 32'hF4527190 , 32'hF0AD1E60 , 32'h013B69A8 , 32'h01358770 , 32'h0CC3B420 , 32'hF3B71230 , 32'h115CDB20 , 32'h04A5DA58 , 32'hFDF1E718 , 32'hF6A55F90 , 32'h04FC0C30 , 32'hF26D7620 , 32'hEED0C2C0 , 32'hFD98CA4C , 32'hE51CC460} , 
{32'h1CD1A680 , 32'hF9094FE8 , 32'h08503450 , 32'hF2C02EC0 , 32'hFE33E294 , 32'hEE3BB200 , 32'h08A0F240 , 32'hEB199CE0 , 32'hF0565010 , 32'hFFAEFBC0 , 32'h1AC863A0 , 32'h1D8D2F40 , 32'hFD9F16D0 , 32'hF0D17D20 , 32'hF722F080 , 32'hF1617F30 , 32'hF4BB9F90 , 32'h13D65100 , 32'hDEB92F40 , 32'h0991FF50 , 32'hDDCE47C0 , 32'hE4C986E0 , 32'hEAD318C0 , 32'h06249C48 , 32'hE64A06E0 , 32'hF2739BA0 , 32'h0493D798 , 32'h1E2ED2C0 , 32'h08D48B80 , 32'h0D8A76E0 , 32'hF330A6D0 , 32'hEC01CD40 , 32'h0D1AB250 , 32'hD4549780 , 32'h01787700 , 32'hFF28EF9A , 32'hF1936060} , 
{32'h0001DB49 , 32'h0003611B , 32'hFFFBEF3E , 32'h00008FA2 , 32'hFFFF7800 , 32'hFFFE92B8 , 32'h0001C2F3 , 32'hFFFBBBF5 , 32'h0000F8DE , 32'hFFFA791D , 32'hFFFE1627 , 32'hFFFE7BFD , 32'hFFFCE253 , 32'h00002661 , 32'hFFFFCC7D , 32'hFFF7249C , 32'h0003C319 , 32'hFFFF8728 , 32'h00072597 , 32'h000144C5 , 32'hFFFF87C1 , 32'hFFFFE644 , 32'h00052E07 , 32'h00043B83 , 32'h00029917 , 32'hFFFBBD8F , 32'hFFF91C51 , 32'hFFFED483 , 32'hFFFB1A8B , 32'h00059ADF , 32'h000302D8 , 32'h000018FB , 32'hFFFD5B3D , 32'hFFFF4351 , 32'h00021F2E , 32'h0002D3A1 , 32'h000009E3} , 
{32'h0000BAD9 , 32'hFFF9BC14 , 32'h00032BAA , 32'h0001FC57 , 32'hFFFEB12B , 32'hFFFDA9E4 , 32'hFFEF941D , 32'h0000D34A , 32'h0008FEE3 , 32'hFFFDBC8E , 32'h0002364B , 32'hFFFBCD2A , 32'hFFFF7C66 , 32'h00047924 , 32'h00013A4C , 32'hFFFBEA9C , 32'hFFF8D72E , 32'h00023961 , 32'hFFFCA4FB , 32'hFFF9C1F2 , 32'hFFFD7FFE , 32'hFFFEEFB4 , 32'hFFFE5053 , 32'h000576ED , 32'h00037CC4 , 32'hFFFDCC9B , 32'hFFFB6485 , 32'h00025502 , 32'h00004561 , 32'hFFF6D271 , 32'h0002AE05 , 32'hFFFEAC94 , 32'h000464FD , 32'hFFF092BC , 32'h0001A7F0 , 32'hFFFC0478 , 32'hFFFDCFE7} , 
{32'hFFFBC968 , 32'h00040686 , 32'hFFFD40CD , 32'h0001D248 , 32'h00025F32 , 32'h000030D9 , 32'h000158D4 , 32'hFFFEE230 , 32'h00032048 , 32'hFFFEF581 , 32'hFFFF055C , 32'h0001E001 , 32'h00010F78 , 32'hFFFE73B3 , 32'h0001DC6E , 32'h000687FB , 32'h0005A6AA , 32'hFFFD376F , 32'hFFFE4D67 , 32'h00013AFC , 32'h0008057D , 32'hFFFFB345 , 32'h00008637 , 32'hFFFD7495 , 32'h0007CC8E , 32'hFFFFE539 , 32'h0001586A , 32'h00005833 , 32'hFFFC1A03 , 32'h00022EC6 , 32'h00000C4A , 32'h0003C43A , 32'h00048A15 , 32'h000179AE , 32'h0002493E , 32'h0003A3C5 , 32'hFFFA5640} , 
{32'hFFFEC5CA , 32'hFFFF4989 , 32'hFFFC4037 , 32'hFFFC1DEC , 32'h00088D61 , 32'hFFF64BB6 , 32'hFFFB35C6 , 32'h000562BC , 32'hFFF7D442 , 32'hFFFDF2BF , 32'h00023C1F , 32'h0000D757 , 32'h00029B9C , 32'h000597A2 , 32'h0000D1CD , 32'h00055A53 , 32'hFFFAB08B , 32'h00012387 , 32'h0000747E , 32'h0000804C , 32'h000000CC , 32'h0000D217 , 32'hFFFD672F , 32'h00013FAF , 32'h00020C28 , 32'h00039572 , 32'hFFFBFC75 , 32'h0004ED6A , 32'h00000B39 , 32'hFFFEED04 , 32'hFFFE2181 , 32'hFFFA8C5F , 32'h000655D4 , 32'h0003FF89 , 32'hFFFF80F3 , 32'hFFF8B210 , 32'hFFFC7EBF} , 
{32'h0003EC32 , 32'hFFF91BF2 , 32'h00066559 , 32'h0006928D , 32'hFFFE33D6 , 32'hFFFD8E46 , 32'h0000E591 , 32'h0007BCD0 , 32'hFFFF934F , 32'hFFFAAF45 , 32'h00039762 , 32'h0003CA98 , 32'hFFFC20B8 , 32'hFFFBEFEF , 32'hFFFF66B9 , 32'hFFFA33F6 , 32'h0001DA9B , 32'hFFFE45D3 , 32'h00011F8B , 32'hFFFDD64E , 32'h0006EF22 , 32'h00048AA4 , 32'h00009725 , 32'hFFFD580B , 32'h0009152A , 32'h00007CDD , 32'h0005D870 , 32'h00006E74 , 32'h0007C4F5 , 32'hFFFD9FCC , 32'h00072FD8 , 32'hFFFC7866 , 32'h0006ED18 , 32'h0003F798 , 32'h00015CD3 , 32'h00054628 , 32'hFFFB9B1C} , 
{32'h0001812A , 32'hFFFFD8AD , 32'hFFF9D0E2 , 32'hFFFAF863 , 32'h00029F9C , 32'h0005AC5C , 32'h000248A6 , 32'h000255E4 , 32'hFFFD8F4E , 32'hFFF8B8C3 , 32'h000BED76 , 32'h00004033 , 32'h00009832 , 32'h000302C6 , 32'hFFF4F7CA , 32'hFFF8530B , 32'hFFF87D1D , 32'h000191B3 , 32'hFFF9B0AC , 32'h0005E6B0 , 32'hFFF89EA0 , 32'h000B0C34 , 32'h00014AAC , 32'h0007E886 , 32'hFFFE8520 , 32'h00025175 , 32'hFFFEEE90 , 32'h00027101 , 32'h0001D9F3 , 32'hFFFE1BF5 , 32'h00030B9E , 32'h0001EB74 , 32'hFFFC8703 , 32'h0005B7DD , 32'hFFFCFB7F , 32'h00053E5E , 32'h00078DDC} , 
{32'h0000DD80 , 32'h000237F2 , 32'hFFFC5BC1 , 32'h000C29AF , 32'h00020194 , 32'hFFF70488 , 32'h0002F678 , 32'h00085937 , 32'hFFFC2444 , 32'hFFF812DA , 32'hFFF9F480 , 32'hFFFD8E10 , 32'h0005EDB4 , 32'hFFFD899C , 32'hFFFEF89A , 32'h0003EBAF , 32'hFFF59F1D , 32'h00038DFF , 32'h00086D34 , 32'hFFF5B694 , 32'hFFFD0E39 , 32'h0004A7B4 , 32'hFFFF09C4 , 32'hFFF6EF2E , 32'hFFFCF3E4 , 32'h000894A4 , 32'hFFFFAFB5 , 32'hFFF636C1 , 32'hFFFA8AC4 , 32'h00090AA6 , 32'h0005A8BD , 32'hFFF9B9AA , 32'hFFFA3815 , 32'h00055DF7 , 32'hFFFCDDD8 , 32'h0007AEB8 , 32'hFFF91A27} , 
{32'h01B537BC , 32'hFF0A29C7 , 32'hFFAEFE83 , 32'hFF7197AF , 32'h00701170 , 32'hFF88C00E , 32'hFF79FC50 , 32'h00B300F3 , 32'hFE548C78 , 32'hFFCEF399 , 32'hFF8C788A , 32'h0003A27E , 32'h0029E306 , 32'hFF1F1396 , 32'h00B6AFB9 , 32'hFED17708 , 32'h00B786C4 , 32'hFFC3C2EC , 32'hFF7B081B , 32'h00C12BCB , 32'hFF0A71CD , 32'h01608384 , 32'hFEBB6D78 , 32'h02B4C248 , 32'h0003B876 , 32'hFDBBAE24 , 32'h013F89F0 , 32'h008F4836 , 32'h0202A160 , 32'h010BDAC8 , 32'hFF888767 , 32'h004E03AF , 32'h0108FF34 , 32'hFFB1C2C4 , 32'hFE97D250 , 32'hFEA62D20 , 32'h00C14EAA} , 
{32'h0C47C380 , 32'hFF017D53 , 32'hF5A1B800 , 32'hFF256713 , 32'hFCD6684C , 32'h07DD23C8 , 32'hFC8CF7D8 , 32'h003E064C , 32'hF5333BF0 , 32'h012F5C58 , 32'hF59EAA20 , 32'hFEFB9074 , 32'h03DD2468 , 32'h08DC37A0 , 32'hFF6ADCF1 , 32'hFB52E578 , 32'h06318FB8 , 32'h071AAC08 , 32'hFFD02AE4 , 32'hFAD348B0 , 32'h067E5128 , 32'hFF63AA71 , 32'hFDE897C4 , 32'hFFA584D9 , 32'h02710270 , 32'h02965AD0 , 32'h0E534DB0 , 32'h03A1CC90 , 32'h093F3A10 , 32'hF9DE6E58 , 32'hF6A2A980 , 32'h04FBB698 , 32'h04C540D8 , 32'hFE855598 , 32'hFFAF154F , 32'h0354E65C , 32'h07B884B0} , 
{32'h64272200 , 32'hF41FF290 , 32'hDB17F380 , 32'h0BEEE9A0 , 32'hECD2FA20 , 32'h237BDB40 , 32'hEA4E9020 , 32'hFF0AFB30 , 32'hDEBDF540 , 32'h054F6F58 , 32'h05E79708 , 32'h0AFB1320 , 32'hF0A737B0 , 32'h25B9C640 , 32'hF420D480 , 32'hD53830C0 , 32'h150A41A0 , 32'hF769DA80 , 32'h0AC153B0 , 32'h0A3D8450 , 32'hE71FF140 , 32'h14AF7280 , 32'h25C88480 , 32'h195048A0 , 32'h04A30C70 , 32'hE8E82CC0 , 32'hE420D360 , 32'hD52B6200 , 32'hF6C121A0 , 32'hEF2E2460 , 32'hE99E1440 , 32'hE724E1C0 , 32'hFC4A665C , 32'h160B1200 , 32'hE700F440 , 32'h0C2665B0 , 32'hEA087780} , 
{32'h22636380 , 32'hEBA4C800 , 32'hED3BC120 , 32'hFFB80767 , 32'hEFB61500 , 32'h2BE5CF00 , 32'hE7F32980 , 32'h09DEB700 , 32'hD97BF1C0 , 32'hFE8E0F90 , 32'h14A0B740 , 32'hFB03D518 , 32'hE8A94540 , 32'h01B74BE4 , 32'hF2A3DEF0 , 32'hEE644C60 , 32'hF7D55EF0 , 32'h00D64703 , 32'hFD9D31C8 , 32'h15DCCF60 , 32'h079A3D30 , 32'h04872A30 , 32'h1562FA80 , 32'hF67029C0 , 32'hFC3BD320 , 32'hF6D85990 , 32'hE68DA1C0 , 32'hFBFB6448 , 32'h04C032F8 , 32'h03CBB2F0 , 32'h146181A0 , 32'hFB9DD878 , 32'hE1E63780 , 32'h00176498 , 32'hF7FCDE90 , 32'h085821B0 , 32'hFA85A830} , 
{32'h299C4000 , 32'hF5957D30 , 32'hEA563520 , 32'hFB17D598 , 32'hF17A2700 , 32'h3B99DD80 , 32'hF980BD90 , 32'h08183540 , 32'hE2C3A400 , 32'h0AE0ACC0 , 32'h23B41240 , 32'hF6BEFD00 , 32'hE28201E0 , 32'hFCDB6E64 , 32'hF342C270 , 32'hEABCF1E0 , 32'hEAD12060 , 32'hF8B83390 , 32'h0326B17C , 32'h253B9FC0 , 32'hFDF828A8 , 32'h07218578 , 32'h17C284A0 , 32'hE8EDBD80 , 32'h0CD9ED00 , 32'hEFFF88C0 , 32'hF14543B0 , 32'h03B3EB4C , 32'hF5BCBB30 , 32'hFD8B1BA0 , 32'h103D83E0 , 32'hF54149F0 , 32'hCDDC0C00 , 32'h0DB260A0 , 32'hE6A78E20 , 32'h061A7A10 , 32'hFEA26528} , 
{32'h5C5EFD80 , 32'hE0574200 , 32'hDC78AC00 , 32'h06760FD8 , 32'hEBE52CA0 , 32'h72027900 , 32'h0635CFF8 , 32'h1294F8C0 , 32'hF241BF60 , 32'hE2C06B20 , 32'h3FC942C0 , 32'hF871B780 , 32'hCCA42480 , 32'hF0DBBF50 , 32'h076C4088 , 32'h0862CCF0 , 32'hE8A8D120 , 32'h03271204 , 32'hF4744100 , 32'h22021B00 , 32'h0061B01A , 32'hEA8168E0 , 32'h1D993320 , 32'h02479F50 , 32'h02F07324 , 32'hE5F279A0 , 32'hEE73C960 , 32'hF8C3CB78 , 32'hFD28515C , 32'hEDC45D20 , 32'hFF5A338A , 32'h03AA4440 , 32'hE91E9EE0 , 32'h1CA5A000 , 32'h0611A6D0 , 32'h15385340 , 32'hED1CFCC0} , 
{32'h62C67B00 , 32'hF2B79100 , 32'hD5D7FDC0 , 32'hF458C620 , 32'hE98DA980 , 32'h66D48400 , 32'hE4397340 , 32'hF8FDA480 , 32'hE3448180 , 32'h17FF2BC0 , 32'h0CD6EE80 , 32'hFE1A4740 , 32'hF2F68290 , 32'h1E0B6DC0 , 32'hF94CF190 , 32'h22419000 , 32'hCCECFB00 , 32'hFC49F7C8 , 32'hEB0ED320 , 32'h178F5520 , 32'hF9598138 , 32'hF7397630 , 32'h17C0FD20 , 32'hDFBFE540 , 32'h01EB2F4C , 32'hF2DE74D0 , 32'hE7846AE0 , 32'hFB748498 , 32'hF9A78788 , 32'h2440F680 , 32'h1328A120 , 32'hF9EEE488 , 32'hDF8AB800 , 32'hE828D7E0 , 32'hEDF63140 , 32'h1BCC02A0 , 32'h04FA6768} , 
{32'h61732D80 , 32'h10329020 , 32'hCE4868C0 , 32'h2D6B48C0 , 32'h0B253F30 , 32'h63F75800 , 32'hEBC28200 , 32'hE4A371C0 , 32'hEF870100 , 32'h25CB6780 , 32'hF7BAF2C0 , 32'hF2284370 , 32'hF308C970 , 32'h2D25F280 , 32'h0252D554 , 32'h249F9280 , 32'hF169F6B0 , 32'h21B1C9C0 , 32'hE4748BA0 , 32'hC5310FC0 , 32'h0EB23340 , 32'hF4035E00 , 32'h3EB43480 , 32'h04252D68 , 32'hE884DAA0 , 32'hF7B25AE0 , 32'h1A9FC320 , 32'hDDE2D100 , 32'hFE2DF438 , 32'h1DF3F6A0 , 32'h009AA1E3 , 32'hF87F50F0 , 32'h1D22D700 , 32'hD34A2A40 , 32'h26D219C0 , 32'hFFCBAFFA , 32'hF916E898} , 
{32'h365AA500 , 32'hE88E4D40 , 32'hD6F9BBC0 , 32'h0CB743C0 , 32'hF24483E0 , 32'h29189540 , 32'hE67677A0 , 32'h02296F7C , 32'hCB5D3940 , 32'h161E9940 , 32'h08EB0CF0 , 32'hE7646900 , 32'hF7169310 , 32'h17AFAEC0 , 32'hF4076B70 , 32'h111C0DA0 , 32'hFECB8368 , 32'h1B9B1180 , 32'h03725038 , 32'hDD7E3D00 , 32'h08BF18E0 , 32'h09CFD370 , 32'h2DE5DA40 , 32'h081C7D00 , 32'hDF3F9E80 , 32'hFF746B80 , 32'h13AFA0E0 , 32'hFD3DF4A8 , 32'h0C2FDE30 , 32'h10162920 , 32'h1B58A860 , 32'h0B236650 , 32'hF2621830 , 32'h04B9CA98 , 32'h120A8CA0 , 32'hECAABC20 , 32'h13383440} , 
{32'h51BCBB00 , 32'hF974F4E8 , 32'hFF744736 , 32'h5B112380 , 32'h3279AD40 , 32'hE531ABE0 , 32'h0B9E4B20 , 32'hF83B3918 , 32'hA7AFF200 , 32'h081474B0 , 32'hDDF2BC00 , 32'hE7505820 , 32'hEFE8CBC0 , 32'hFC2F5040 , 32'hE42A3C60 , 32'h1CDE6900 , 32'hFB309CA8 , 32'h174B7740 , 32'hFD64BA6C , 32'hEE53EF00 , 32'h16195C20 , 32'h1C1B6C40 , 32'hDB006E80 , 32'hD9F635C0 , 32'h16E05580 , 32'hEB832B00 , 32'hF6642E50 , 32'hFC34FAC4 , 32'hE5921CA0 , 32'h13EDA5C0 , 32'hDDFDDA80 , 32'h21F18300 , 32'hEC777820 , 32'hFA2D9A10 , 32'h1C5EE320 , 32'h0EA9C4D0 , 32'h0E172DC0} , 
{32'h28B5E300 , 32'hC822B900 , 32'hE42A0F20 , 32'h6634B780 , 32'hF2ACA980 , 32'hCDAF2B00 , 32'h52500B00 , 32'hF8F551D0 , 32'hCF70FB40 , 32'hC51DC440 , 32'hFC79CDF0 , 32'hB5E66B80 , 32'hEAFBDB00 , 32'h156A1D20 , 32'hEED59FA0 , 32'h13CDF960 , 32'h09126380 , 32'h081897F0 , 32'h0D92F2E0 , 32'h175B5680 , 32'h121B0FE0 , 32'h23CA9DC0 , 32'hBE178700 , 32'hF5CCB9B0 , 32'h0A6D4F80 , 32'hE2939920 , 32'h1C788B80 , 32'h36222500 , 32'hDF725440 , 32'hEAACDCE0 , 32'h1E9E6740 , 32'h03DA1774 , 32'h17873020 , 32'hE35997C0 , 32'hDEDB82C0 , 32'h097A5970 , 32'hE0B80EC0} , 
{32'h2CC6A9C0 , 32'hC2D662C0 , 32'hE9140D80 , 32'h254541C0 , 32'hF2B0DC40 , 32'hFEACB960 , 32'h136067C0 , 32'h184760C0 , 32'hF8C7F908 , 32'hBF785100 , 32'hE99BFAC0 , 32'hDC134940 , 32'h0605BF78 , 32'hEB4A3B80 , 32'hCC0D1E00 , 32'h4E45A300 , 32'hDD744900 , 32'hF09494F0 , 32'h1D2D0A00 , 32'hF6854AE0 , 32'hB3851C80 , 32'h0460CB48 , 32'hFB5AFEE0 , 32'h2A526380 , 32'h16B91D40 , 32'h10BCD240 , 32'h07EA2C80 , 32'h1D3188C0 , 32'h02504434 , 32'hE4206A60 , 32'h05D4F860 , 32'h099428E0 , 32'h0B7367B0 , 32'h143F3FA0 , 32'h0317D09C , 32'hEC0BBD00 , 32'h04ADB708} , 
{32'h34A11EC0 , 32'hD798E040 , 32'h01F48778 , 32'hFBD3C8A0 , 32'h04502338 , 32'h1CBD2E00 , 32'h0A9B0B50 , 32'hD5122500 , 32'h2F4CA880 , 32'hD574E7C0 , 32'hCBCB1440 , 32'hC71A2A40 , 32'hC8495F00 , 32'hDCAEC940 , 32'hE561DF20 , 32'h165ECF20 , 32'hF74EEBC0 , 32'hE9FFFF80 , 32'h1BB6FE20 , 32'hF1A264F0 , 32'hE00951E0 , 32'hFACAD9C8 , 32'hE0A59B60 , 32'h1BCFF380 , 32'h22408400 , 32'hDED1ED80 , 32'h09D2C990 , 32'hE2A5C200 , 32'h242BCA00 , 32'hF6C117D0 , 32'h027AB8A0 , 32'h038B3A8C , 32'h0DECD230 , 32'h1F1549C0 , 32'hE382A0A0 , 32'hE7F8D380 , 32'hF9D46C58} , 
{32'h09EC04F0 , 32'hFC0A56F0 , 32'hF771B4F0 , 32'hFC49D15C , 32'h0274C988 , 32'h13293CE0 , 32'h07DA4798 , 32'hEEF8F3A0 , 32'h3B109300 , 32'h018D8920 , 32'hCA291280 , 32'hE2496940 , 32'hE5558300 , 32'hE2170160 , 32'hE7B72EA0 , 32'hFF5B975D , 32'h0EC72CE0 , 32'hF5E3AB50 , 32'h28ADCE40 , 32'h06FB0A20 , 32'hE860C700 , 32'hD0830DC0 , 32'h05F73EC8 , 32'h05C54450 , 32'h0708ADD0 , 32'hDDD76B00 , 32'h167F8860 , 32'hE6417FC0 , 32'h1501C320 , 32'h13C5A900 , 32'h078B32B0 , 32'hF9841810 , 32'hF6A0EE60 , 32'hF9B03F60 , 32'hF7709150 , 32'h04FC1E80 , 32'h0D5F2690} , 
{32'h3F705040 , 32'hC8852100 , 32'h0F9B0C60 , 32'hE2638FC0 , 32'hFF0E1A29 , 32'hD3BD3C80 , 32'hFBB6D628 , 32'h224227C0 , 32'h46AEA180 , 32'h120D02C0 , 32'hDDA25F00 , 32'hE511FE80 , 32'hD8F613C0 , 32'hEA279440 , 32'hEAB7BAC0 , 32'hF68AD570 , 32'hFF1B8848 , 32'h002BE9C4 , 32'h27F8D900 , 32'h0811BDC0 , 32'h16FE7F40 , 32'h094AAB10 , 32'hF539AAA0 , 32'hD1848B00 , 32'hF7D4D550 , 32'hF513A770 , 32'hFE1570E8 , 32'h0DC59640 , 32'hFF791D29 , 32'hFA21C440 , 32'hD71F0600 , 32'hEC5857C0 , 32'hF2E81020 , 32'hDF0E8F40 , 32'h0621EDD8 , 32'hFB53D890 , 32'h052E4600} , 
{32'h4FAF5100 , 32'hB8B90700 , 32'h1D7C91A0 , 32'hED077920 , 32'h10545320 , 32'hC27A3C40 , 32'hF3E91800 , 32'h274DF800 , 32'h3CA4A480 , 32'h3087F0C0 , 32'hF43188A0 , 32'hEE7DE240 , 32'hF9588668 , 32'h0747DF38 , 32'hEEF44D40 , 32'h01F391C0 , 32'h05F3C2D8 , 32'hFCC48DE8 , 32'h22065600 , 32'h0C2372D0 , 32'hF7374F60 , 32'h06CFEEF8 , 32'h0AEE6A10 , 32'hED4702C0 , 32'h01FC6B00 , 32'hF2615550 , 32'h098AE4E0 , 32'hE7C648C0 , 32'hF594F110 , 32'hFCB96BDC , 32'hF6D24370 , 32'hF7AF7F30 , 32'hE8637860 , 32'hF0461A80 , 32'hFDDAF3B8 , 32'h09ABA8E0 , 32'hFE5BA1F4} , 
{32'h44337380 , 32'hCAC4B500 , 32'h1C0F1F00 , 32'hFA0BDC30 , 32'h04173E78 , 32'hCFA0CA80 , 32'hF6876430 , 32'h2CCF1740 , 32'h2688E7C0 , 32'h2A5F22C0 , 32'h0FB1D630 , 32'h1DF2AAC0 , 32'h52D02200 , 32'h2FC49AC0 , 32'h0B1D1C00 , 32'hF6732E50 , 32'hD76EE3C0 , 32'hFA39E068 , 32'hFDFF7B18 , 32'h12C5FB40 , 32'h044B1AB8 , 32'h1B248D40 , 32'h123C8D40 , 32'h0BE7CA90 , 32'hF1821210 , 32'h0D748660 , 32'hE6F917E0 , 32'hEF724720 , 32'hE9930D40 , 32'hE75E5960 , 32'hF03C8260 , 32'hF899B288 , 32'h1F50E2E0 , 32'h0AFDC6A0 , 32'hFA1BBFD8 , 32'h069E1968 , 32'h282AD180} , 
{32'h3FDCDC80 , 32'hE575EE80 , 32'h15745760 , 32'hF4AC0130 , 32'h02FEB638 , 32'hD79220C0 , 32'hFA8B5B00 , 32'h307055C0 , 32'h0FBC0F50 , 32'h0BF64540 , 32'h0E88D980 , 32'h1F628AA0 , 32'h1FE30280 , 32'h260104C0 , 32'h290C5AC0 , 32'hFE1C9EA8 , 32'hF7F89A10 , 32'h0CD49340 , 32'hE06F72C0 , 32'h16DB3020 , 32'hFF1CAA5B , 32'h2054B900 , 32'h0D9CCB80 , 32'hFEF42894 , 32'h05B7C4C0 , 32'h35369280 , 32'hF8FA6430 , 32'h0A04B320 , 32'hE55EFA20 , 32'hEFE69380 , 32'hF58914C0 , 32'h04157CA0 , 32'h03F870A8 , 32'hFD83B4C8 , 32'h06E9CFF8 , 32'hF8A63B40 , 32'hF2671D20} , 
{32'h27FE1E00 , 32'hE63CD640 , 32'h04C3D560 , 32'h1607F900 , 32'h023DD6C8 , 32'hD3E7A100 , 32'h00B7B344 , 32'h16C5CF60 , 32'hFFA3A462 , 32'h09B2C630 , 32'hD36B9DC0 , 32'hEE46EAE0 , 32'h00D8EBFE , 32'h16077660 , 32'hF16AC8A0 , 32'hDF507140 , 32'h079D4EC0 , 32'hECC8AEC0 , 32'hFDABFBA0 , 32'h03B4AB1C , 32'hF0B3B610 , 32'h1DF98B40 , 32'hF5C2FB20 , 32'hFDBE58D4 , 32'h0D802C40 , 32'hF4A0F4C0 , 32'hF66A65F0 , 32'hF20EA7C0 , 32'h0BC0A150 , 32'h0F12E8A0 , 32'hFDAB49CC , 32'hFB3AC850 , 32'h0CF095F0 , 32'h0D542840 , 32'hFA64FAC8 , 32'hFEDCBFA0 , 32'h0BD91000} , 
{32'h2DF3D880 , 32'hFE721318 , 32'h0DA52420 , 32'hECB0CE00 , 32'h10EA83C0 , 32'hEC651360 , 32'h0B040D30 , 32'h09BA3460 , 32'hFC9D2E90 , 32'hFB59D480 , 32'hFD040688 , 32'h031CF1CC , 32'h214E9FC0 , 32'h2C7EBDC0 , 32'h03C2C1BC , 32'h07711B78 , 32'hF6706780 , 32'hF6DC68D0 , 32'hE7D625E0 , 32'h10A419A0 , 32'hC530B500 , 32'h19C8FA20 , 32'h037AAA38 , 32'h150C00C0 , 32'h1BB5D580 , 32'hF10CBE80 , 32'hFE7FFA24 , 32'hF152B830 , 32'h0E1D2910 , 32'h0AC8EB70 , 32'h20FA5C80 , 32'h238C50C0 , 32'h098E9810 , 32'h1AB194C0 , 32'h188D2900 , 32'h13A5FBC0 , 32'hEF9F8620} , 
{32'h0D54D7B0 , 32'hF71AF700 , 32'h011ED978 , 32'hFE352D04 , 32'h0663CCC8 , 32'hF67F65A0 , 32'hF48B0960 , 32'hEFC60FE0 , 32'hF5C77930 , 32'hFEC0F9BC , 32'hF5118CD0 , 32'h07835F58 , 32'h03609EA8 , 32'hFE4DA5D8 , 32'hF11B16E0 , 32'hFB740BB0 , 32'hEDCF75C0 , 32'hF81F7C90 , 32'hEFB64F80 , 32'hF3DBF7B0 , 32'hF1FB0670 , 32'hEE419DE0 , 32'hEF6133C0 , 32'hF86DF3B0 , 32'hF2F2BEE0 , 32'h0A126E70 , 32'hF9F91140 , 32'h105A94C0 , 32'hF80CD1D8 , 32'h18787B40 , 32'hE9539060 , 32'hFEE0F3C0 , 32'h06834C50 , 32'hF5BF30D0 , 32'hF3560A10 , 32'h0691DA78 , 32'h050AE7B0} , 
{32'h0674C748 , 32'hFBC68E70 , 32'h03F872E0 , 32'hFE2685E8 , 32'h01BEA860 , 32'hFE63F9FC , 32'hFFB62599 , 32'hFB3B1F48 , 32'hFF2F81EA , 32'hFACCE148 , 32'h02C0F5B8 , 32'h01A0E1AC , 32'hFF3DC176 , 32'hFAFE1358 , 32'hFFDAE163 , 32'h009372D6 , 32'hFC777A8C , 32'h02C50D64 , 32'hF8F7DE20 , 32'hFE9D972C , 32'h003075F6 , 32'hF33978D0 , 32'hFC11F444 , 32'h01472468 , 32'hFB0FD668 , 32'hFE226188 , 32'hFC8B7C40 , 32'h08D67E30 , 32'hFAE8B678 , 32'h03ABA25C , 32'hF6CAA780 , 32'hF72F6D00 , 32'h094FDDF0 , 32'hFF3A74E3 , 32'hFF8E86CE , 32'hFDA4E1B8 , 32'h02DAB61C} , 
{32'h0007D67D , 32'h0002FAC6 , 32'h0002933C , 32'hFFFD20ED , 32'h0000A3D6 , 32'h0002BEF4 , 32'h0000445B , 32'hFFFF2041 , 32'h00027231 , 32'hFFF90178 , 32'h00015EAC , 32'hFFF94175 , 32'h0000CCF3 , 32'h0002C20B , 32'hFFFFE3F2 , 32'h000140E5 , 32'h00075E13 , 32'h000638BC , 32'hFFFE5DAC , 32'hFFFCD8AD , 32'hFFFF28C7 , 32'h00007C2E , 32'h0004E4FD , 32'hFFFFA2DA , 32'hFFFBE3CA , 32'hFFFB0000 , 32'h0000873F , 32'h00010C31 , 32'h0001C60D , 32'h0001A38B , 32'h000040B5 , 32'hFFFBA415 , 32'hFFFE8FE9 , 32'hFFFDCA7E , 32'h00004AFA , 32'h00070EE6 , 32'h0002E982} , 
{32'hFFF69493 , 32'h0000AA0B , 32'h000188E0 , 32'hFFFA0A4F , 32'h0005C946 , 32'hFFFE957E , 32'h00071A5D , 32'hFFFD103B , 32'h00018B40 , 32'h0004043B , 32'hFFFD6EB4 , 32'h0000D05E , 32'hFFFF1D56 , 32'h00066F28 , 32'hFFFE1C5C , 32'hFFFD83F7 , 32'hFFFEE336 , 32'hFFF710C2 , 32'h000061DB , 32'hFFFE78CC , 32'h00019690 , 32'h00055C75 , 32'hFFFB1179 , 32'hFFFEFA7D , 32'hFFFC978F , 32'hFFFE274A , 32'h00003D82 , 32'h00017662 , 32'hFFFE8E75 , 32'hFFFDE0DA , 32'hFFFB93D0 , 32'hFFFA8ECF , 32'h00052A16 , 32'hFFFD731F , 32'hFFF73F4F , 32'hFFF74312 , 32'h0003EF5C} , 
{32'h00063764 , 32'h000318D6 , 32'h000526CA , 32'h000B979A , 32'h00065D80 , 32'h0003A7C8 , 32'h00099CF8 , 32'hFFF39B57 , 32'h0003B615 , 32'h00084DC5 , 32'h00012545 , 32'hFFFED700 , 32'h00074839 , 32'hFFFB7D37 , 32'hFFF8308C , 32'h0000EA55 , 32'h0009A3DE , 32'h0009BC2F , 32'h000856D6 , 32'h00072B06 , 32'h0003EF19 , 32'hFFF88312 , 32'h000166A2 , 32'h00041461 , 32'hFFFD2117 , 32'hFFFAAC2A , 32'hFFFAA867 , 32'hFFF697BC , 32'h000210CC , 32'hFFFC0A80 , 32'hFFFB1CD8 , 32'h0003CE3B , 32'hFFFDADD2 , 32'hFFFC2BCC , 32'h000A3773 , 32'hFFF95148 , 32'hFFF7183A} , 
{32'hFFF69A6D , 32'h00033CDD , 32'hFFF72B01 , 32'h0000AEA6 , 32'h0003B19C , 32'h00007B92 , 32'h0001FE0E , 32'hFFFB77A4 , 32'hFFFD0D5F , 32'hFFFE28FF , 32'hFFF9DA58 , 32'hFFFB9F26 , 32'h00009ADA , 32'h00049256 , 32'hFFFFA842 , 32'hFFFB287B , 32'hFFFE5921 , 32'hFFFA32E7 , 32'h000A19C9 , 32'h0003CBFC , 32'hFFFBAE3E , 32'h0006559A , 32'h0001F712 , 32'hFFFFCA6F , 32'hFFFD5E58 , 32'h0000C95C , 32'h00015E40 , 32'h00026EA7 , 32'h00015858 , 32'hFFF7F831 , 32'h00034895 , 32'hFFFE7009 , 32'hFFFAC0F5 , 32'h0005A459 , 32'hFFFC4660 , 32'h0002BB9C , 32'hFFFB525C} , 
{32'h00085C18 , 32'h0005E231 , 32'hFFFCAFBA , 32'hFFFF79F6 , 32'h000108B2 , 32'hFFFB579D , 32'hFFFD29B2 , 32'hFFFEC7AF , 32'hFFFECFA5 , 32'h0006FC46 , 32'h000097D4 , 32'hFFFD3594 , 32'h0002355B , 32'hFFFE55CB , 32'h0003A4A1 , 32'hFFF780D4 , 32'hFFFBF1B0 , 32'hFFF876E4 , 32'hFFF7BD84 , 32'h000307DD , 32'hFFF45698 , 32'hFFFF7704 , 32'hFFFE0902 , 32'h00007FC0 , 32'hFFFFFCD0 , 32'h00013956 , 32'h0001CC2C , 32'h0002CC1A , 32'h000425D1 , 32'hFFFD0C62 , 32'hFFFDFF40 , 32'h0004C20E , 32'h0001FC28 , 32'h00006BE3 , 32'h0000156E , 32'hFFFA79A9 , 32'hFFFC6219} , 
{32'h065818E8 , 32'hFBDE5F00 , 32'h037B0CEC , 32'h010AE600 , 32'h034460F4 , 32'hFC64C948 , 32'h012867D4 , 32'h02F206A8 , 32'h052A6AB0 , 32'hFF85D01B , 32'hFD022058 , 32'hFB8A9050 , 32'hFDCCCAE8 , 32'hFE1E7950 , 32'hFB361D50 , 32'h0054B565 , 32'hFA8149F8 , 32'h001ACD01 , 32'hFFFC05DD , 32'hF9CC1120 , 32'hFC3DBAEC , 32'h02F7D0B8 , 32'h00761D38 , 32'hFCCAA884 , 32'hFEBB2CCC , 32'hFECAF938 , 32'hFCAD484C , 32'hFF921D8B , 32'h02859884 , 32'hFEE4FBF4 , 32'hFB0F8D48 , 32'hF8312298 , 32'h00ECA62D , 32'h0168C7A4 , 32'h047910B0 , 32'hFBF14C98 , 32'h02843A48} , 
{32'h125FEF80 , 32'h0A06D6C0 , 32'hFDE0610C , 32'h15CBE020 , 32'h0774C1B8 , 32'h0A70D6E0 , 32'hF57CB320 , 32'hFB253318 , 32'hFCF0F524 , 32'hFE25F934 , 32'h019ED534 , 32'h04FEA7F0 , 32'hF84F1258 , 32'h2331F300 , 32'hED5A8820 , 32'h018523D0 , 32'h141511A0 , 32'hF0F18A20 , 32'h046ECF98 , 32'h07631898 , 32'hFD8EF8B4 , 32'hF49107D0 , 32'h101E3B20 , 32'h0932E2C0 , 32'hFE4520EC , 32'h066C3938 , 32'h0C1F1560 , 32'h03344B4C , 32'h0D0AE0C0 , 32'hEBE8FB60 , 32'hE89FB060 , 32'hFC0C0CB0 , 32'h0ECE6410 , 32'h027B3EFC , 32'hF8FAE4D8 , 32'h08B1A880 , 32'hFD62A0F4} , 
{32'h35D24240 , 32'hF3A0AEF0 , 32'hE753C4A0 , 32'h1C0DE820 , 32'hECB2CC00 , 32'h1D4E7B80 , 32'h08C8EDE0 , 32'hF7B00310 , 32'hD8D6B4C0 , 32'h001153A9 , 32'h1545F820 , 32'hEC9D2100 , 32'hF61F1120 , 32'h0E18BEA0 , 32'hEE2B3CA0 , 32'hE7A5A300 , 32'h006E6F1A , 32'hF27FEAE0 , 32'hFAC57420 , 32'h201D54C0 , 32'h15007880 , 32'h07570250 , 32'h0D0E5460 , 32'hF204C510 , 32'hFFF77D93 , 32'hFA764670 , 32'hF5FFBC10 , 32'hFBC48F00 , 32'h09DD0020 , 32'h08D8A420 , 32'h008C92AE , 32'hE5500E60 , 32'hF46EF380 , 32'h0A58F220 , 32'hFA00AC60 , 32'h07D19A40 , 32'hFEEF11D0} , 
{32'h2B9D66C0 , 32'hEDD10DC0 , 32'hEC8416E0 , 32'h04BA1158 , 32'hF74275C0 , 32'h2DB40000 , 32'hEF3D4C40 , 32'h0A24F4D0 , 32'hD809EF80 , 32'h02AE3854 , 32'h13FA05C0 , 32'h05B07D40 , 32'hEC90DB80 , 32'h03C6254C , 32'hF92BB5A8 , 32'hEF1E4DA0 , 32'hF04C8DE0 , 32'hF8F5DD28 , 32'h073C02C0 , 32'h0E488A90 , 32'hFEE04BB8 , 32'h04269B50 , 32'h178926E0 , 32'h0608F9F8 , 32'hFADB5CD0 , 32'hED8A4D00 , 32'hF121E000 , 32'hEFC5D7E0 , 32'hF98045A8 , 32'h0F23A050 , 32'h05BE2AB0 , 32'hFCC6BCA4 , 32'hEB41D320 , 32'h063822B8 , 32'hF7B11050 , 32'h09FD30A0 , 32'hE9D92CE0} , 
{32'h47191A80 , 32'hF7D97910 , 32'hDD24BEC0 , 32'h1CEF4200 , 32'hED73BFE0 , 32'h2A852D40 , 32'h02510F04 , 32'hF462D8E0 , 32'hD1AEDA00 , 32'h06ECA200 , 32'h1C80B560 , 32'h03521830 , 32'h04B83820 , 32'h0171150C , 32'hE72B3AE0 , 32'hE3D8CB60 , 32'hFD29A76C , 32'hF6E1AFA0 , 32'hF959E5A8 , 32'h24E64240 , 32'hFBED9230 , 32'h0770CE80 , 32'h0A1741A0 , 32'hDD1671C0 , 32'hF6735A80 , 32'hF73CA220 , 32'h15386E40 , 32'hF63B09E0 , 32'h04F9D4A8 , 32'h293F3A40 , 32'h140BC740 , 32'hEB116540 , 32'hF0D0A540 , 32'hE452D020 , 32'hFF9E7D58 , 32'hF45AC3D0 , 32'hDCAB4B00} , 
{32'h1F090580 , 32'h0B5BD3D0 , 32'hE00D7FA0 , 32'h16D06000 , 32'hEA9E0F20 , 32'h27A03040 , 32'h08FBC120 , 32'hEBBB1380 , 32'h0B5D7B80 , 32'hFB0EBFE8 , 32'hFF988D13 , 32'hFEBAE8F0 , 32'h0F3FD310 , 32'h10D9EFA0 , 32'h016189FC , 32'hE62573C0 , 32'hFB5BFCC8 , 32'hEBBE08E0 , 32'h0BFC9E30 , 32'h0FCA73F0 , 32'hF956EEE0 , 32'h0082BEC8 , 32'hF68D5BF0 , 32'hFC2FE9B0 , 32'h027B2A30 , 32'hFB4B1C38 , 32'hF3189880 , 32'h03707DA4 , 32'hFD7AB25C , 32'h0F66AE90 , 32'h12686200 , 32'hEDC824C0 , 32'hF9C40E28 , 32'hF01BF870 , 32'h03E6A734 , 32'hFF7BE2F4 , 32'hE354BDA0} , 
{32'h255EF580 , 32'h149DBC40 , 32'hECF05020 , 32'h25AAA500 , 32'h09342A30 , 32'h25B61E40 , 32'h1E4E96E0 , 32'hFEEDFB9C , 32'hFE0A667C , 32'hFBC3E710 , 32'h0AE81C60 , 32'hFF790167 , 32'hF2D32D70 , 32'h03D419F0 , 32'h05E12020 , 32'hDF3B77C0 , 32'hF1D20690 , 32'hDE5B17C0 , 32'hF45D60C0 , 32'h1C9A1680 , 32'h09B879D0 , 32'hFF0A67A6 , 32'hF1FA2B30 , 32'hE5BC18A0 , 32'h0EE3BBD0 , 32'hF88AA240 , 32'hFB0A7328 , 32'h0AC33420 , 32'hF05D31E0 , 32'h01EA3AA0 , 32'h1107C100 , 32'hF65AB8A0 , 32'h1BBFA9A0 , 32'h03667320 , 32'h0CD350C0 , 32'h0D895EB0 , 32'hDD57BE00} , 
{32'h2B4D5AC0 , 32'h1744BB80 , 32'hEA5D5240 , 32'h2DA09FC0 , 32'hFDE321CC , 32'hFD264F7C , 32'h38586E00 , 32'hEB6066A0 , 32'hFD5DBFD0 , 32'h0EB6BDD0 , 32'h0C31F9C0 , 32'hF66BA2C0 , 32'h0915A0F0 , 32'h048165C8 , 32'h091C4060 , 32'hFB7DCA10 , 32'h07304F78 , 32'hF9169E08 , 32'h040C5748 , 32'h049F7B98 , 32'h09FCF380 , 32'hFD6FF90C , 32'h01069B04 , 32'hF8FB42F8 , 32'hFFBDBA76 , 32'h052A5F80 , 32'h092C52C0 , 32'hF9248228 , 32'hFDD35D70 , 32'h039F32A4 , 32'hF9D3F7C0 , 32'hE9E213E0 , 32'h051C0CA8 , 32'h00D9E728 , 32'h043A05D0 , 32'h03E97B6C , 32'hFCE1B2A8} , 
{32'h4A50FB80 , 32'h3838E9C0 , 32'hFA1A3018 , 32'h48073300 , 32'h248D4080 , 32'hF0952F20 , 32'h511B0880 , 32'hD603E600 , 32'hE470D6A0 , 32'h17BC52A0 , 32'hFB075DD8 , 32'hFBECAD70 , 32'hE1E382E0 , 32'hFC250C08 , 32'h136097E0 , 32'h01917E2C , 32'h01C0AD34 , 32'h0400DD68 , 32'hEE2652E0 , 32'hFF35B589 , 32'h14B52600 , 32'h12C87320 , 32'h0566C0D8 , 32'h0CEFADE0 , 32'h093E9710 , 32'h1F6AAAE0 , 32'hF5A9F2D0 , 32'hE302F500 , 32'h05CFFCA8 , 32'h20C931C0 , 32'hFC597D3C , 32'hF8F3CBF8 , 32'hFCA1DC3C , 32'hDAF04EC0 , 32'h03E992C4 , 32'h0977D660 , 32'hF29DF680} , 
{32'h1A328540 , 32'h35D73340 , 32'hE683F280 , 32'h6493E800 , 32'h202427C0 , 32'hDE806580 , 32'h63772900 , 32'hD4FFA140 , 32'hEC3DCDC0 , 32'h194864C0 , 32'hFBE2E658 , 32'hD8A77100 , 32'h1F1F5FC0 , 32'hFD324A34 , 32'h1D084740 , 32'h24962300 , 32'h02063638 , 32'hF5D37570 , 32'hFEEF1BA0 , 32'hFDC311FC , 32'h07D1D928 , 32'h07EEC550 , 32'hE8657240 , 32'hFF93AFD1 , 32'hE3576A20 , 32'h26ABC3C0 , 32'h15325940 , 32'hE25B8140 , 32'h219F7BC0 , 32'h2604FD00 , 32'h05FB28F0 , 32'h01A5F160 , 32'h171AE760 , 32'hE47CB000 , 32'h0BE36A00 , 32'h0C528800 , 32'h0658CC10} , 
{32'h1DF92E20 , 32'hE576AAA0 , 32'hE7C2D7A0 , 32'h584FA400 , 32'h0BEFDF40 , 32'hF3D334F0 , 32'h35FB6100 , 32'hE0205940 , 32'hE2DC3840 , 32'hEEBB88A0 , 32'hFDDFB1EC , 32'hCD222A40 , 32'h12573280 , 32'h124B1880 , 32'hF0E40D50 , 32'h29E5C4C0 , 32'h0B4BF530 , 32'h0BC00E30 , 32'hCD829600 , 32'h100D7600 , 32'h25C72680 , 32'hEEDBE0C0 , 32'hF2964140 , 32'hED2CC820 , 32'hCC14EB80 , 32'hDDE12740 , 32'h257873C0 , 32'h05D97D98 , 32'h0C7AB8F0 , 32'hF7BDDFC0 , 32'hE02F23C0 , 32'h15412C00 , 32'h11AE1C80 , 32'h20B7F400 , 32'hE96432C0 , 32'hEF916DE0 , 32'h0DB1E030} , 
{32'hFC516E2C , 32'hCAD08780 , 32'hDC428D40 , 32'h31CC9AC0 , 32'hDA1EF6C0 , 32'hE9D709A0 , 32'h202C3C40 , 32'hE00E8F40 , 32'hF654D720 , 32'hD1F948C0 , 32'hF0AFBD20 , 32'hC1B95840 , 32'h256874C0 , 32'h0FAF46C0 , 32'h14531E00 , 32'h043BDBA0 , 32'hEDA73E80 , 32'hE84FDF00 , 32'h04921488 , 32'h2E36BF40 , 32'hF36545B0 , 32'hEE1493E0 , 32'hE625E020 , 32'hE2C38BA0 , 32'hF3579E60 , 32'hD50F4740 , 32'h2D0197C0 , 32'h113BC440 , 32'h1389A300 , 32'hF94B1EF8 , 32'hFC3241C8 , 32'hE215A280 , 32'hF6FFA9D0 , 32'h29DE1600 , 32'h040A9318 , 32'hEDC120C0 , 32'h079B1640} , 
{32'h03B84168 , 32'hDEC32A80 , 32'hCD005480 , 32'h15911260 , 32'hEB0A2C00 , 32'h05302460 , 32'h03F933E4 , 32'hD18BE280 , 32'h16D16A60 , 32'hC7C43140 , 32'hD5F4F380 , 32'hCD267A40 , 32'hED9BDB60 , 32'h0DB2A720 , 32'hD6B6FF80 , 32'h156E6240 , 32'hFD4AC8D8 , 32'hD8547B40 , 32'hD4DF0980 , 32'hF98050A0 , 32'hF3DD0D90 , 32'h145C2FA0 , 32'h0DA04930 , 32'hFB4ABC90 , 32'h0CF8D040 , 32'h10415FE0 , 32'hF4153D10 , 32'hFFF2C27D , 32'hEC0BDA80 , 32'hDEA2E900 , 32'hEF78BDC0 , 32'hFF43A889 , 32'h150595C0 , 32'hFFBF1842 , 32'hFBC493B0 , 32'hF311DA50 , 32'hEF35F800} , 
{32'hE655DB80 , 32'h03ABBB18 , 32'hE899E400 , 32'h10CED980 , 32'hF71B91E0 , 32'h065BFA80 , 32'h134F1400 , 32'hEBE0E520 , 32'h0C3B8D90 , 32'hE3FAD6A0 , 32'hDC8466C0 , 32'hE25E67C0 , 32'hBC7CC480 , 32'hEDF7A3A0 , 32'hF8966090 , 32'h0A9009E0 , 32'h14063980 , 32'hE6B4DDA0 , 32'hE97A3160 , 32'hFFC1BFE9 , 32'hEBC29AC0 , 32'h04DEFBD0 , 32'hFE928748 , 32'h030A0354 , 32'h09F590A0 , 32'hE90FA160 , 32'h0464F9E0 , 32'hDD2A4180 , 32'h0B7BCB40 , 32'hFA6199D0 , 32'h03E75B80 , 32'h0248FFE8 , 32'hFA45ABE8 , 32'hE357FDC0 , 32'h00655EF5 , 32'h15682660 , 32'hE8DBBC60} , 
{32'hF3839A20 , 32'hFF12FEA6 , 32'hEF3CDD80 , 32'h1ACA4860 , 32'hEE1DC780 , 32'h06402CC8 , 32'hEA4752C0 , 32'h24FD6E40 , 32'h29E63D00 , 32'h2BDE8380 , 32'hDF89EC80 , 32'hD2DBB440 , 32'hCE6D1E00 , 32'hE23C7880 , 32'h0CD9AC10 , 32'hF7460B30 , 32'h1FEB4640 , 32'hE6C2AB80 , 32'h02918F54 , 32'h035F3F80 , 32'h2C432500 , 32'h0A316310 , 32'hF08DAB10 , 32'hDD77E1C0 , 32'h04686750 , 32'hF406A910 , 32'hEBD96960 , 32'hFF185A1F , 32'hF20F6F00 , 32'hF7389860 , 32'hED056EE0 , 32'hFD19D34C , 32'h1BB00B20 , 32'hEBE294C0 , 32'hF9319960 , 32'h13580100 , 32'h0EFCE400} , 
{32'h08311D80 , 32'hEABE7360 , 32'hF12F3B00 , 32'h1B488B60 , 32'hD942C0C0 , 32'hE314EDA0 , 32'hEAE94780 , 32'h2BF15640 , 32'h40DF5600 , 32'h5565A780 , 32'hBB5F6780 , 32'hE0F7B360 , 32'hB953D500 , 32'hD2DF76C0 , 32'hF6CFCF20 , 32'hF459F610 , 32'h04E818A8 , 32'hF1355C20 , 32'h0544A6A8 , 32'h1B04E380 , 32'h403E5800 , 32'hED9FD040 , 32'h0D4F55D0 , 32'hE16186A0 , 32'hD5A56880 , 32'hF325F3D0 , 32'hE2B749C0 , 32'h0CA29C50 , 32'h16BC55C0 , 32'h0850C4C0 , 32'h0352F534 , 32'hF60AA740 , 32'h19F5BE20 , 32'hE73AF880 , 32'hF93AD230 , 32'hECDB10C0 , 32'hED327DC0} , 
{32'h1F3B35E0 , 32'hE2D06A60 , 32'hE1FE7A80 , 32'h23D90C80 , 32'hF5F7A730 , 32'hE0B76520 , 32'h0236C1C4 , 32'h5CD9AD80 , 32'h2E27DD40 , 32'h2FD09780 , 32'hC1674F00 , 32'hEE3A1160 , 32'hFBA656D0 , 32'hEA72FA80 , 32'hE3677BA0 , 32'h0A8E8EF0 , 32'hE0BD02E0 , 32'h1DD1A900 , 32'h1BEE7540 , 32'h250019C0 , 32'hDCD8C4C0 , 32'hFE7F30B8 , 32'h05680500 , 32'h0B66E3B0 , 32'hF23CC2E0 , 32'hF5B41B80 , 32'hE3791080 , 32'h09F1A2D0 , 32'h03676E80 , 32'h026AE540 , 32'h12693520 , 32'hFD8C890C , 32'hF59DDAE0 , 32'hED582580 , 32'h030399F4 , 32'hF381A780 , 32'h003840E9} , 
{32'h1EC11CC0 , 32'hE4983740 , 32'hEC8CAC40 , 32'h28F03E40 , 32'hF56CDA90 , 32'hF46632D0 , 32'hEBDACE00 , 32'h5E867F80 , 32'h256F5040 , 32'h34523100 , 32'hE160D960 , 32'hFEEB6D94 , 32'h1CDF4AE0 , 32'hFA1B4C10 , 32'hDF1D0940 , 32'h0610AC88 , 32'hD48D5DC0 , 32'h0E229DE0 , 32'h25A65F40 , 32'h30E9A240 , 32'hEF1B1F00 , 32'hF92D0F90 , 32'h10BF2140 , 32'h09CC5960 , 32'hFE685840 , 32'h0A009500 , 32'hE52C1520 , 32'h22838000 , 32'h06381F78 , 32'hF740E420 , 32'hEE904C60 , 32'hFB2D4188 , 32'h02E2B7D0 , 32'h00244EEF , 32'hFF40BFD9 , 32'hED076520 , 32'h0B682BB0} , 
{32'h08A539D0 , 32'h074175C0 , 32'hF4F10150 , 32'h0DF9F160 , 32'hFDA486A8 , 32'hFE905CA0 , 32'h0D1F0270 , 32'h15923E00 , 32'h0E815710 , 32'h2A50F780 , 32'hE6971D20 , 32'hEFD42E80 , 32'hFB26FE40 , 32'h07746120 , 32'hF729B380 , 32'hF82B2630 , 32'hDE392800 , 32'hFEDB61CC , 32'h07293B98 , 32'h0FAB2150 , 32'hF6664EC0 , 32'h0BE90DD0 , 32'h03FE3FB0 , 32'h1929D2C0 , 32'h10FB7B40 , 32'hF48F9CB0 , 32'h12504F80 , 32'h10242CC0 , 32'h00055EF1 , 32'h0E5C50D0 , 32'h013BD8B0 , 32'hF3B100E0 , 32'h019724E0 , 32'h0000DDC1 , 32'hEBDD81E0 , 32'hF8259D50 , 32'h0EDFD300} , 
{32'h10769FE0 , 32'hF8B2DD40 , 32'hFE70F204 , 32'h09AD7650 , 32'hF5505A30 , 32'hF0B460D0 , 32'hFB1F1DE0 , 32'h23236C80 , 32'hFA129890 , 32'h0918BD70 , 32'hFC123AE8 , 32'h01B215E4 , 32'h1AFE19C0 , 32'h01DCA064 , 32'h13E111C0 , 32'hF8FAEA40 , 32'hD7312080 , 32'h050DA5D0 , 32'hEB35C480 , 32'h072316C8 , 32'hF4B2EDA0 , 32'hFCB38890 , 32'hF77FB1A0 , 32'hF0CBD2B0 , 32'hFD98F31C , 32'h0CD95440 , 32'h05E828B0 , 32'h07A2C9A0 , 32'h04633060 , 32'hF7A6BD30 , 32'hDF6A4600 , 32'hEBCE7920 , 32'h00B0566A , 32'hFE205E5C , 32'h027FF5B0 , 32'hE49275A0 , 32'h0E103B80} , 
{32'h3FD5E440 , 32'hEB1ABC20 , 32'h166A5B80 , 32'hEC66A460 , 32'h0F694620 , 32'hD9DA05C0 , 32'h1BC1FB20 , 32'h04A11680 , 32'h1961D700 , 32'h00932EC1 , 32'h0001DD24 , 32'hF1CE3020 , 32'h0C7CE3B0 , 32'h1FCC9F80 , 32'h017DD0FC , 32'hF2FD77D0 , 32'hF0BEB900 , 32'h040B65F8 , 32'hEE6A0C40 , 32'hFF4EA75E , 32'hD49C0380 , 32'h1D89EFA0 , 32'h0A117050 , 32'h01D838A4 , 32'h07C122D0 , 32'h08301030 , 32'h029FA1E0 , 32'hFC2EBAAC , 32'hF7931C30 , 32'h02C176C4 , 32'h05D6FA10 , 32'h134D5B80 , 32'hFBFD2918 , 32'h027C7434 , 32'h18222CA0 , 32'h0712C538 , 32'h01CF01D8} , 
{32'h12B6E240 , 32'hF0DEDBB0 , 32'h06E67408 , 32'hFB131038 , 32'h11025CC0 , 32'hE9F174C0 , 32'hF421D560 , 32'hF905ED40 , 32'hFF468C38 , 32'h09C5AC50 , 32'hE13E5F00 , 32'hF5FAFFD0 , 32'h00F8E9F1 , 32'h18CEE780 , 32'hE95E3CC0 , 32'hEF4C2720 , 32'hEEBE95A0 , 32'hECEFBCA0 , 32'hEFABC1E0 , 32'hE8FE8EA0 , 32'hEF8908E0 , 32'h0B8F5BC0 , 32'hF96046A8 , 32'hF60AA600 , 32'h055284D0 , 32'h0468B1A0 , 32'hEDA1B460 , 32'h0110FA88 , 32'h05EDCFE0 , 32'h17837B40 , 32'hFC9B7BD4 , 32'h10193160 , 32'h0073092D , 32'h09AAD9E0 , 32'h099487D0 , 32'hFD187FE4 , 32'h0F385810} , 
{32'hFFFF6B8F , 32'hFFFF3F1F , 32'h000484AC , 32'h000013AE , 32'hFFFAA083 , 32'h0000C109 , 32'hFFFEC00A , 32'hFFFC3793 , 32'h0001603E , 32'h00034860 , 32'hFFFCC3B7 , 32'hFFFBF07D , 32'hFFFB93BE , 32'hFFFE503F , 32'hFFFB72AF , 32'h00002A90 , 32'hFFFEB169 , 32'hFFFD5BB4 , 32'h00040F42 , 32'h00015A9F , 32'h00024FEE , 32'hFFFDC35B , 32'hFFFF05B1 , 32'h0002119B , 32'h00063E49 , 32'h0002C04F , 32'h0001CD77 , 32'hFFFD3DDD , 32'hFFFC0723 , 32'hFFFC9442 , 32'h0001EC05 , 32'h00043649 , 32'hFFFED703 , 32'h0000E3CB , 32'h00010AD3 , 32'hFFFB8553 , 32'hFFFEAD70} , 
{32'h00022333 , 32'hFFFC27F1 , 32'h0005D66C , 32'h000121D9 , 32'h000691D3 , 32'hFFFB29AF , 32'h00018675 , 32'hFFF7CC2C , 32'hFFFF76F0 , 32'h00008C97 , 32'h00059E02 , 32'h0001516F , 32'h00007DBA , 32'h00017883 , 32'h00015172 , 32'h00031E3E , 32'hFFFD196A , 32'hFFFC80AD , 32'hFFFE87B6 , 32'hFFFC321A , 32'h000816B5 , 32'h000131CD , 32'h00015049 , 32'h000A1052 , 32'hFFFF4322 , 32'hFFFBAFA0 , 32'h00007E58 , 32'hFFFD83EF , 32'h000590B2 , 32'h00069B48 , 32'hFFFDAAEB , 32'hFFFF7C6D , 32'h00002A25 , 32'h00024F34 , 32'h0007DFED , 32'h0000AB24 , 32'hFFFB8B5E} , 
{32'h000CAC84 , 32'hFFFCCD34 , 32'h0006E8B1 , 32'h0002A22C , 32'h000075D4 , 32'hFFF8F2DC , 32'h0000A3B4 , 32'h00038F7B , 32'hFFF9B594 , 32'h000912FE , 32'h00049362 , 32'hFFF220AB , 32'hFFFAFAE3 , 32'h0001E767 , 32'hFFFB95D4 , 32'hFFF66B3E , 32'h0003F222 , 32'h0001D7E6 , 32'h00024C5D , 32'h0005A595 , 32'h00077043 , 32'hFFF8EC15 , 32'hFFF60C96 , 32'hFFF99BF4 , 32'h000029AD , 32'hFFF54E76 , 32'hFFFFA895 , 32'h0005C1DB , 32'hFFFE49DB , 32'hFFF93D8B , 32'h000095B8 , 32'hFFFA5B18 , 32'hFFF8813F , 32'hFFFB2C31 , 32'h0001E33C , 32'h00005ADE , 32'hFFFDF1F4} , 
{32'hFFFF9128 , 32'h00063C2F , 32'h0004A1CB , 32'h00011B3F , 32'hFFFA33D5 , 32'hFFFE23C0 , 32'h0001FB9B , 32'hFFF4819D , 32'hFFFE9A94 , 32'hFFFD6848 , 32'hFFFCEB5C , 32'h0003C5C1 , 32'h0007FE61 , 32'h0000C06A , 32'hFFFDBA80 , 32'h000030D5 , 32'hFFFC314F , 32'hFFF9810E , 32'h00017882 , 32'hFFFF1C3F , 32'h000290A2 , 32'h000098B3 , 32'h0004A1C8 , 32'hFFFE31FA , 32'h000011E7 , 32'hFFFE1008 , 32'hFFFA11D1 , 32'h0009AE18 , 32'hFFFB7323 , 32'h0001CE8B , 32'hFFED6446 , 32'h0004C422 , 32'h00088735 , 32'hFFF95BBD , 32'h0006B44A , 32'h0003D8B6 , 32'hFFFD3BF8} , 
{32'h0000D111 , 32'h0007CC2D , 32'hFFF9743E , 32'h00020E5D , 32'h00047EBF , 32'hFFFCE459 , 32'hFFF7EF19 , 32'h00068963 , 32'hFFFC1674 , 32'hFFF924CF , 32'h00012F8C , 32'h0000D2E2 , 32'h000112C3 , 32'hFFFDD687 , 32'hFFF9B091 , 32'h000178B4 , 32'h00071209 , 32'h0000F846 , 32'hFFFFA22C , 32'h0001C7DA , 32'h0001D7AD , 32'h0003FADB , 32'hFFFDC480 , 32'hFFFDF15B , 32'hFFFFDF3E , 32'hFFFBB327 , 32'hFFFDF17D , 32'h000023D5 , 32'hFFFF94A2 , 32'hFFF5FF7E , 32'h0004FF3D , 32'hFFF2E594 , 32'hFFFEDB27 , 32'hFFFF49D1 , 32'h00032389 , 32'h0000B77E , 32'hFFFB77EA} , 
{32'hFFFC5D65 , 32'hFFFF0700 , 32'hFFF9F72C , 32'hFFFF7D8A , 32'h0002B2D6 , 32'hFFFDA645 , 32'hFFFCC480 , 32'h000A6800 , 32'hFFF880AC , 32'hFFFE074D , 32'hFFFEF68A , 32'hFFF90457 , 32'h0002523F , 32'hFFFDB22B , 32'h00084CE4 , 32'hFFF95772 , 32'h0005AA0E , 32'hFFFE8452 , 32'h00003D56 , 32'hFFFF718A , 32'h0003B4F5 , 32'hFFFC8B68 , 32'hFFFEF02F , 32'hFFFF61D0 , 32'hFFF97986 , 32'hFFF79F85 , 32'hFFF59A57 , 32'hFFFEAB8C , 32'hFFFBDC4A , 32'h00013A09 , 32'hFFFF98DD , 32'h0001B3DF , 32'h00035455 , 32'hFFF5D3A1 , 32'hFFFE2908 , 32'h0000A0EE , 32'hFFF5CFCC} , 
{32'hFFF7C028 , 32'hFFF66011 , 32'hFFFFEF55 , 32'hFFFEB1B8 , 32'hFFF7F8CA , 32'hFFFD9F1A , 32'hFFFB8021 , 32'hFFFED5AE , 32'h0005F56B , 32'hFFFAA548 , 32'h0005FCB9 , 32'hFFF6FD97 , 32'hFFF9E393 , 32'h00065F6E , 32'hFFFDB46F , 32'h000C8F0C , 32'h00025073 , 32'h00070DBF , 32'hFFFF3354 , 32'h000708F2 , 32'h00047F5D , 32'hFFFB7105 , 32'hFFFDE91C , 32'h00013023 , 32'hFFFF7138 , 32'hFFFC0104 , 32'h00033B5C , 32'h00040E68 , 32'hFFFD9324 , 32'h0000F6F0 , 32'h00046A0D , 32'hFFFC3E7B , 32'h0008E689 , 32'h0007BAA2 , 32'h00040522 , 32'h00018EFC , 32'h000022EA} , 
{32'h1E656A40 , 32'h0E977240 , 32'hF8793A50 , 32'h0CB6EB20 , 32'hF4BBD290 , 32'hFAA23EA0 , 32'h137CFF20 , 32'hFD696430 , 32'hEEA70DE0 , 32'h07408B20 , 32'h033EDE14 , 32'hEB88F220 , 32'h140C9EC0 , 32'h060E68E8 , 32'h04419320 , 32'h03F0D98C , 32'h05CDB1C8 , 32'hE1AC3860 , 32'hF8817B10 , 32'h0A98DE90 , 32'h17C12FA0 , 32'hF8FCECD0 , 32'hDF91BDC0 , 32'h009E6797 , 32'h041E60E0 , 32'hF9FDAFB8 , 32'h0FFC1800 , 32'hFD46D9E8 , 32'hFEF03AAC , 32'h0E476A80 , 32'h04AD25C0 , 32'hED894CA0 , 32'hFF5CD05F , 32'hF78B88F0 , 32'h05E46F18 , 32'hF40C35C0 , 32'hFA57E6C8} , 
{32'h2568E840 , 32'h14735880 , 32'hFB8F2BD8 , 32'h1030A180 , 32'h10FB9600 , 32'h09C7E1B0 , 32'h32C73800 , 32'h032287C8 , 32'h05DFD518 , 32'h065D2148 , 32'h1E550CA0 , 32'hE991AA00 , 32'h129255A0 , 32'hF2351B60 , 32'h0E68BC00 , 32'hF034C630 , 32'hF0E24590 , 32'hD213F9C0 , 32'h1B6385A0 , 32'h0707F5C0 , 32'h0F195250 , 32'h030F6404 , 32'hEDC6F440 , 32'hEBFDAAC0 , 32'hF500ACA0 , 32'hFE3A4FA0 , 32'h10E76800 , 32'hFD44BF08 , 32'h13D51280 , 32'h07F5AFE0 , 32'h14EC8420 , 32'hF278E5A0 , 32'h0F43EB40 , 32'h0E425970 , 32'hEEDD1F60 , 32'h05315080 , 32'hF3E72C30} , 
{32'h257351C0 , 32'h025C452C , 32'hF0C9D2D0 , 32'h141340C0 , 32'hFD0D7B28 , 32'h1390AB00 , 32'h18F28380 , 32'h01A719B8 , 32'hECF21FE0 , 32'h022B4AC4 , 32'h1A3A1120 , 32'hF5A89AC0 , 32'hF662AB40 , 32'hF6F0B520 , 32'hFFBDABB5 , 32'hDFA84FC0 , 32'hFB4EBC58 , 32'hDF705480 , 32'h005917A6 , 32'h0E80CD00 , 32'h0BA77C50 , 32'h008E033C , 32'h07059D50 , 32'hF1E274A0 , 32'hFBD6C980 , 32'h04503600 , 32'hFC919B58 , 32'h09750270 , 32'h0A089B60 , 32'hFD1CBF54 , 32'h17291BC0 , 32'hF7E5BC00 , 32'hF06C5350 , 32'h0D4EDB40 , 32'hF4A05B90 , 32'h092B47B0 , 32'h16457B20} , 
{32'h3ACAC400 , 32'h25AE1580 , 32'hE6386BE0 , 32'h2D0ADF40 , 32'hF502CBA0 , 32'hF5264550 , 32'h275C0480 , 32'hEFD1C260 , 32'hFD3D1578 , 32'h0F94B040 , 32'h0FF35E80 , 32'h1089F4A0 , 32'h17306BC0 , 32'hF0B743C0 , 32'h078507D0 , 32'hE4C6C820 , 32'h022FD6C4 , 32'hF6306EA0 , 32'h0AB5FFA0 , 32'hFC1DEC6C , 32'hEA812340 , 32'hF4876DA0 , 32'hDE1C1E40 , 32'hEEE92580 , 32'hF6690990 , 32'hF91DDEF0 , 32'h0C2BEB10 , 32'hEF317500 , 32'hF9053860 , 32'h1DEC8F40 , 32'h1B573F00 , 32'hE7BA76C0 , 32'hF6194CD0 , 32'hF1B5DD00 , 32'hFE540510 , 32'hF5693100 , 32'hF6227CD0} , 
{32'h47DDCA80 , 32'h22A42240 , 32'hE0EECAE0 , 32'h41B2DD80 , 32'h0FFC3310 , 32'hEE4DA900 , 32'h575C4E00 , 32'hE563D940 , 32'h012F93E4 , 32'h16F52300 , 32'h168DEA80 , 32'hF999F950 , 32'h1CAD95C0 , 32'hF77C7220 , 32'hF7E72240 , 32'hEB890EA0 , 32'hF8091230 , 32'hE4D7FB40 , 32'h0937FF70 , 32'hEE272CC0 , 32'hF2D86F90 , 32'hF67FC6C0 , 32'h05900558 , 32'hFC7C146C , 32'h007604FD , 32'h11340AC0 , 32'hFE584F80 , 32'hFF87A1D3 , 32'h08393840 , 32'h06AFB6C8 , 32'hFAA67898 , 32'hE5492E60 , 32'hF6941890 , 32'hFA6E5580 , 32'hFC4982CC , 32'h044B5A60 , 32'h09BAA8A0} , 
{32'h366EDB80 , 32'h301797C0 , 32'hFDD9E9C0 , 32'h46E69480 , 32'h170096C0 , 32'hF6FC9740 , 32'h764A9780 , 32'hEB0A26C0 , 32'h0EE18CF0 , 32'h0FEA1990 , 32'h234B0C40 , 32'h0FCF91D0 , 32'h0823C500 , 32'hDABFE740 , 32'h216E7640 , 32'hE2CF2160 , 32'hF0B6E080 , 32'hDF5A1740 , 32'h0F556E10 , 32'h0AE68420 , 32'h08503CB0 , 32'hFFD81553 , 32'hF8250FD0 , 32'hFC481890 , 32'h0F8927D0 , 32'h0A121090 , 32'hF5EF7E30 , 32'h08686D30 , 32'hF3812510 , 32'hF57D3C70 , 32'h0585AA68 , 32'hECA0E2E0 , 32'hDED9E2C0 , 32'h101DD820 , 32'h1BF96A80 , 32'h0E8E92B0 , 32'h0605E748} , 
{32'h08292910 , 32'h36782940 , 32'h14398F80 , 32'h31575980 , 32'h2C2D8D40 , 32'hD2772A00 , 32'h5354AE80 , 32'hE308E3A0 , 32'h147B76E0 , 32'h2766F100 , 32'h10940EA0 , 32'hFAF14A90 , 32'h09494B00 , 32'hE920E920 , 32'h2D7B4380 , 32'h021B4F08 , 32'hFDA9AFA4 , 32'hE0F9D980 , 32'hEDB11BA0 , 32'hDC5401C0 , 32'h07557D70 , 32'hFAA4F598 , 32'h0A148AD0 , 32'h10E82780 , 32'hF868B8D0 , 32'h2E43F840 , 32'h0CAB2DF0 , 32'h007687ED , 32'h0AA37D10 , 32'hF8303910 , 32'hFD3B3EA8 , 32'hF9CA9658 , 32'h04BEFF68 , 32'h13F1D760 , 32'h10214EE0 , 32'hEB2E3FC0 , 32'h21A7F7C0} , 
{32'hF2286C70 , 32'h29013840 , 32'h030861FC , 32'h51089C00 , 32'h3E078B40 , 32'hD4636600 , 32'h306F1880 , 32'hD8D92A40 , 32'h1292C2A0 , 32'h1E1706A0 , 32'h2C3B4700 , 32'hDB49F340 , 32'h070CD9D8 , 32'hEE026C80 , 32'h2B638500 , 32'h49592480 , 32'h09524110 , 32'h30653080 , 32'hFDDBC1A4 , 32'h091045B0 , 32'hEA477300 , 32'hF9B32B78 , 32'h08BF4070 , 32'h432BE480 , 32'hFACF9920 , 32'h058DFEF8 , 32'hEBA9A0E0 , 32'hD9DD0380 , 32'h07C85178 , 32'h13D2E120 , 32'h10BCAAA0 , 32'h0B0522B0 , 32'hE8C54540 , 32'hEB8E3940 , 32'hF725AC60 , 32'hED197B80 , 32'h1785F020} , 
{32'hB060C200 , 32'hF26310E0 , 32'h215C87C0 , 32'h1D92A920 , 32'h0D386F60 , 32'hA3E2A480 , 32'h152150E0 , 32'hF79F71F0 , 32'h2242DF00 , 32'hFACF8B10 , 32'h4BB6A400 , 32'hCD25E200 , 32'hDE339400 , 32'hFECC19F4 , 32'h28B71D00 , 32'h5FCBA480 , 32'h05B78040 , 32'h33759900 , 32'hFCE912E4 , 32'h30C32EC0 , 32'h16A78560 , 32'hFE09E808 , 32'h162DCC20 , 32'h21266600 , 32'hEE041F40 , 32'hF6AE24E0 , 32'h064D59A8 , 32'hDC87B500 , 32'h20512680 , 32'hEE101DA0 , 32'hE50024C0 , 32'hDC463180 , 32'h0B5015C0 , 32'hECF38660 , 32'hF30308E0 , 32'h1341DF00 , 32'hD5FE8880} , 
{32'h9A75F380 , 32'h7FFFFFFF , 32'h09756FD0 , 32'h125B6760 , 32'hD4F69700 , 32'hBDFF0B80 , 32'h14D00160 , 32'hE5468120 , 32'hFB20D238 , 32'hFB43EE90 , 32'h4104D480 , 32'h9AF24100 , 32'h1AC80080 , 32'h0EA5C830 , 32'hE89CF940 , 32'h20438280 , 32'h02885300 , 32'hE72DBA00 , 32'hE8C0CB00 , 32'h1B9BAFA0 , 32'hFC600EB8 , 32'hFE21A0C8 , 32'hED5AFE20 , 32'hE3966BE0 , 32'hCD74DBC0 , 32'hF6045F80 , 32'hFD0BAA88 , 32'hF6871AA0 , 32'h05C7A298 , 32'h02339140 , 32'h03C5CF64 , 32'hF79C63C0 , 32'hF6621540 , 32'h312C8E40 , 32'h0B92B6B0 , 32'h2782E840 , 32'hF3FE69F0} , 
{32'hE6C06C40 , 32'hB3185400 , 32'hC2178F00 , 32'h142F81C0 , 32'hCC0FA180 , 32'hDE97CCC0 , 32'hF41FD940 , 32'hD79890C0 , 32'h0028F21E , 32'hE8A636E0 , 32'hE7C51800 , 32'hEB636EA0 , 32'h0CAEB050 , 32'h0D910440 , 32'h11240FE0 , 32'h12E2D700 , 32'hF55633D0 , 32'hE4B851E0 , 32'hDD38AC40 , 32'hDE4CCD80 , 32'hF6132BE0 , 32'h135F7780 , 32'h016AA0A0 , 32'h085D20C0 , 32'hE47795A0 , 32'h01857B64 , 32'h03BAB4B4 , 32'h19AD62C0 , 32'h0B323CB0 , 32'h0B2B9570 , 32'h08660110 , 32'h272C6980 , 32'hF3D69F30 , 32'h153ED240 , 32'hF3874C50 , 32'hEE6F98A0 , 32'h02699534} , 
{32'h04D2DAC0 , 32'hF0D0F5C0 , 32'h07F1A7F8 , 32'h164F02E0 , 32'hEA4AA780 , 32'hF8BBE378 , 32'hD35E5D00 , 32'hC27B6500 , 32'hF11795E0 , 32'hE5554380 , 32'hA1487600 , 32'hFB8D6E20 , 32'hEE2B5DA0 , 32'hE9A5DD60 , 32'hF84FB7D0 , 32'h3B69FE40 , 32'h14524B40 , 32'hBD164100 , 32'hA25C3C00 , 32'hF83831E8 , 32'hC0BD1540 , 32'h1D377700 , 32'hFCF1E8BC , 32'hD0201A40 , 32'hF9A27A30 , 32'h321A4100 , 32'hED505F60 , 32'h0180FD98 , 32'hDF563340 , 32'h08822110 , 32'hEC520080 , 32'h0D85FA10 , 32'hD8B3B7C0 , 32'h123D9900 , 32'hE862E040 , 32'h06787030 , 32'h0B0BDA10} , 
{32'hEDC450C0 , 32'h02556A60 , 32'hD4FD3380 , 32'h10C7B040 , 32'hCD50A3C0 , 32'hFF184A38 , 32'hF8581C10 , 32'h007C13EE , 32'hF797C260 , 32'h1933C8A0 , 32'hD43C3A00 , 32'hF37AC5A0 , 32'hA5801E80 , 32'hF49CB640 , 32'h074A2DF0 , 32'hE8428F60 , 32'h1E219BE0 , 32'hF1FCE6F0 , 32'hD1692800 , 32'h08386C20 , 32'h10393760 , 32'h39BC6280 , 32'hF7E4FA90 , 32'hECF8DEA0 , 32'h077B2F28 , 32'h1C14F840 , 32'hE32D6060 , 32'h070540E0 , 32'hE8805700 , 32'hE2CE0280 , 32'hEA076380 , 32'hB72D8E00 , 32'h05038448 , 32'hD41802C0 , 32'h00C007D0 , 32'hF11532F0 , 32'h23B92FC0} , 
{32'hF4876DF0 , 32'h06B4B640 , 32'hE8D211C0 , 32'h1722E600 , 32'hE6C1DE80 , 32'h1BC3F160 , 32'hE3805FA0 , 32'h24D0DD80 , 32'h0BF7D830 , 32'h20E1B100 , 32'hE415F180 , 32'hF4554ED0 , 32'hCCEFA600 , 32'hE34F9A00 , 32'h11AB3520 , 32'h0F65BD40 , 32'h25615D00 , 32'hD30387C0 , 32'h13511920 , 32'h01B7D434 , 32'h52DDD500 , 32'h00F0783D , 32'hD5222F40 , 32'hD6E3F500 , 32'h2B353B40 , 32'hEBF569C0 , 32'hE7EC7480 , 32'hF7B583B0 , 32'hED5AAE40 , 32'h052F0318 , 32'h02558D94 , 32'hE708C300 , 32'h3662A5C0 , 32'h30671900 , 32'h040F8020 , 32'hFE220120 , 32'h15172DC0} , 
{32'hEB0F9EC0 , 32'h09C39A20 , 32'hF0E4EE70 , 32'h145F7580 , 32'hF934BE08 , 32'h11AB3D80 , 32'hF36EB650 , 32'h052B7460 , 32'hFE7E2004 , 32'h08397050 , 32'hFD83BB5C , 32'hFBA2BB18 , 32'hF94A0020 , 32'hEAA85E80 , 32'h0876C720 , 32'h09C01030 , 32'h10C5B480 , 32'hF176A800 , 32'h147AF4A0 , 32'hFF6A26B6 , 32'h20C9DC80 , 32'hEC7E73C0 , 32'h0A217800 , 32'hF3D29E80 , 32'h08D765C0 , 32'hFC92ACC4 , 32'hFAA873C8 , 32'hEA6C2A60 , 32'hFACEF958 , 32'h007B8A3A , 32'hF8168A30 , 32'hE5954B20 , 32'h24B26A40 , 32'h03F53D1C , 32'hD5A65740 , 32'h116183C0 , 32'h0AB24BA0} , 
{32'h1D86B3E0 , 32'h0354000C , 32'hE81C3320 , 32'h461A3D80 , 32'hE537D400 , 32'hE9B4ED60 , 32'h1750F4E0 , 32'h5F7F0100 , 32'h0FD1C810 , 32'h332422C0 , 32'hE9D79080 , 32'h1365DB20 , 32'h286C6940 , 32'h04812770 , 32'h1DF67CE0 , 32'h1FA9D080 , 32'hE69AD9A0 , 32'hF9802480 , 32'h05C18CB0 , 32'h2BDFC580 , 32'h1B0B5280 , 32'hFD954578 , 32'h049F5440 , 32'hF75AE810 , 32'hEF0828A0 , 32'h53297000 , 32'hDC2284C0 , 32'h07381EA8 , 32'hF9472B90 , 32'h2C2445C0 , 32'hFC7CA2E4 , 32'hECE7BDE0 , 32'h173B22C0 , 32'h1CBB7FA0 , 32'hF804D210 , 32'h133EE4A0 , 32'h03C31954} , 
{32'h00B90A74 , 32'hE43DC640 , 32'hE6D750E0 , 32'h3CFD6840 , 32'h137F87A0 , 32'h008698FA , 32'hF6322CA0 , 32'h5F118600 , 32'h262BA4C0 , 32'h308B3F40 , 32'hDEBE3280 , 32'hEE4B2660 , 32'h477C9D00 , 32'hCEE77600 , 32'hC802FA40 , 32'h17E7C640 , 32'hF13AA1A0 , 32'h0B40D350 , 32'h203A6540 , 32'h2F401080 , 32'hE3A13E20 , 32'hE4435520 , 32'h29484300 , 32'h0F21B3B0 , 32'h0FF27CC0 , 32'hDC7C9780 , 32'hFDF00DC0 , 32'h0D0D8B00 , 32'h0F940DD0 , 32'h00B70763 , 32'hF994A3E0 , 32'h259CF900 , 32'hFC0F5448 , 32'hE8A2FD00 , 32'h00DAC5FD , 32'h1354B9C0 , 32'hEEE1A140} , 
{32'h10ECB820 , 32'hFAA23310 , 32'hF537DA50 , 32'h13EBCA00 , 32'hF20F2A10 , 32'hF7D734C0 , 32'h06016DB0 , 32'h2BEAFA00 , 32'h13B7B520 , 32'h080DA3E0 , 32'hD9D2F800 , 32'hF4AE69B0 , 32'hF5679080 , 32'hEB694AC0 , 32'hF35F9600 , 32'hF60178F0 , 32'hEC3351E0 , 32'hF32CA3A0 , 32'h08B72E00 , 32'h113A69E0 , 32'hEDE9B120 , 32'hF73A7500 , 32'hFD77C9B4 , 32'h0C588AB0 , 32'hF7E5C650 , 32'hF7235AE0 , 32'h0745E4D0 , 32'hFD42C59C , 32'h0F0C99C0 , 32'h0218DDC0 , 32'hF9F459D8 , 32'h015DE134 , 32'h001276BA , 32'hF096FA20 , 32'hFD9835FC , 32'hF1773170 , 32'h152578A0} , 
{32'h244DC280 , 32'hF129C6C0 , 32'h05D9E770 , 32'h06C881D0 , 32'hEDB7CEE0 , 32'hF2988780 , 32'h004AD94B , 32'h22A4F840 , 32'h1482D020 , 32'h01056084 , 32'hE7784260 , 32'hFB4ACBC0 , 32'hFF0419D8 , 32'hF4F28130 , 32'hFCB0145C , 32'hFB9B4738 , 32'hEBE3F360 , 32'hEF6F59A0 , 32'h0DA7FCD0 , 32'h254AF5C0 , 32'hEDEE8980 , 32'hEE62CB00 , 32'hFBF9FB60 , 32'h0E6B48E0 , 32'h135B39E0 , 32'hFC5FD310 , 32'h14A7B5A0 , 32'h06D7ECC0 , 32'h030A88A8 , 32'h0C360B30 , 32'hFE3E895C , 32'h159FF940 , 32'hF2EF1790 , 32'hEB3E7600 , 32'h0537B1A0 , 32'h01CBBFA8 , 32'h14A19A40} , 
{32'h08FE41D0 , 32'h1468F200 , 32'h0FD64F20 , 32'hE426D5E0 , 32'hE81FEC20 , 32'h06C6FCF8 , 32'h1A43D800 , 32'h1F6A6F00 , 32'hF075E850 , 32'h0CF2C7A0 , 32'h050A99D0 , 32'hED1DDC60 , 32'h13F11780 , 32'h0C6ADAE0 , 32'hDEC08AC0 , 32'h01FA3FB4 , 32'hECD030A0 , 32'hC9FA4000 , 32'hDD2A9A80 , 32'hF8E1E920 , 32'hFCEC5BB0 , 32'hF10DCCD0 , 32'hEE899A00 , 32'h2648C7C0 , 32'h186ADAC0 , 32'hF1C95770 , 32'h0C262210 , 32'hF243BE00 , 32'hE836D020 , 32'hF4488640 , 32'hF7D7DEB0 , 32'h2189C2C0 , 32'hF568CFC0 , 32'hECDE3360 , 32'hFBE0A718 , 32'hFE6B2BD8 , 32'hFC0825E0} , 
{32'hF6996340 , 32'hF127F7A0 , 32'h0650A760 , 32'h039AEA1C , 32'h01C899F8 , 32'h0224C2CC , 32'h02B4067C , 32'h045BAD10 , 32'hF11EA660 , 32'h040DD9F0 , 32'hEB38C5A0 , 32'hDEDA7D80 , 32'h074FCDE0 , 32'hF91AA518 , 32'h1C4D0A40 , 32'hDD895640 , 32'hDE54B240 , 32'h18A498A0 , 32'hF4BB57E0 , 32'h05BAC920 , 32'hF72CF550 , 32'hDC319180 , 32'h0258D844 , 32'hE92A6D60 , 32'h1A0AC080 , 32'h08F5FB90 , 32'h14200420 , 32'hF21891D0 , 32'hF797A370 , 32'hE797D880 , 32'hF159FB50 , 32'hF6CF7B00 , 32'hF15BC4B0 , 32'h12348A80 , 32'hFE6A57B4 , 32'hEC312AC0 , 32'hF9980BA8} , 
{32'h0000FADB , 32'h0001DB7A , 32'h00024378 , 32'h0004F084 , 32'hFFFF3A93 , 32'hFFFC7F1F , 32'hFFFCC904 , 32'h00004A96 , 32'hFFFD692A , 32'h00003E96 , 32'h000256EC , 32'hFFFFF918 , 32'hFFFEA7B7 , 32'h0001118B , 32'h0001B8C6 , 32'h000058FF , 32'hFFFCA1AB , 32'hFFFF0A3C , 32'hFFFF0E93 , 32'hFFFCAC48 , 32'hFFFC98B6 , 32'hFFFB227E , 32'hFFFF1EFA , 32'h00062AC3 , 32'h00007FB5 , 32'hFFFD2866 , 32'hFFFC35FE , 32'h000532F1 , 32'hFFFD572B , 32'h000117CC , 32'hFFFF9A12 , 32'h0001A72B , 32'hFFFDDE61 , 32'h0006D84E , 32'h00039075 , 32'hFFFA4586 , 32'h00013E9E} , 
{32'h00105F7C , 32'h00063A6C , 32'hFFECA2DA , 32'h001022EA , 32'hFFF9CFC7 , 32'h00037012 , 32'h0003EF63 , 32'hFFEE37B0 , 32'hFFFAD84C , 32'hFFF6E445 , 32'hFFFE2B1E , 32'hFFF4B899 , 32'hFFFD1152 , 32'h0009CE26 , 32'hFFED6B7C , 32'hFFFA2721 , 32'h0002A8AD , 32'h00059FAB , 32'hFFF5CEB0 , 32'hFFFFA476 , 32'h0002F984 , 32'hFFFB2CA4 , 32'h001494A5 , 32'hFFFA684A , 32'hFFFECDB1 , 32'h00018C2E , 32'hFFFE3BF4 , 32'hFFF2F670 , 32'hFFF8F4D4 , 32'hFFFD2E47 , 32'hFFE95816 , 32'h0000D854 , 32'h000D2E69 , 32'h0001B64C , 32'hFFFA1A1C , 32'h000627B0 , 32'hFFF92235} , 
{32'h000197A3 , 32'h00012B0B , 32'hFFFA0B97 , 32'hFFFE1A70 , 32'h00002FCB , 32'hFFFD8AB9 , 32'hFFF9A454 , 32'hFFFCCDF2 , 32'h00011ADB , 32'h0006281F , 32'h00032D5D , 32'h0007BAC6 , 32'h00062C7C , 32'hFFFD83E4 , 32'hFFFFFF31 , 32'hFFFDAF38 , 32'h0003B404 , 32'h00054E24 , 32'hFFFECACC , 32'hFFF962D0 , 32'h000235C7 , 32'hFFFE9B63 , 32'hFFFBFF14 , 32'h0005D182 , 32'h0007946D , 32'hFFFB0401 , 32'h0004CD2A , 32'h0000C47B , 32'hFFFA5859 , 32'h00052D1D , 32'h000059C5 , 32'hFFFE83CA , 32'hFFFF2B29 , 32'hFFFFC318 , 32'hFFF9A0AE , 32'hFFFBD2EA , 32'h0005EA58} , 
{32'h00015468 , 32'hFFFF5914 , 32'h0002510B , 32'h00077EF5 , 32'hFFFE8505 , 32'h00025CAF , 32'hFFFF1E9C , 32'h0000E1F9 , 32'hFFFC90C5 , 32'hFFFC15DD , 32'hFFF8D5E9 , 32'h0002D2DA , 32'hFFF86B67 , 32'hFFFFFEFA , 32'h0003E8E8 , 32'hFFFAC65F , 32'hFFFDE47D , 32'hFFFB5D0D , 32'hFFF83C97 , 32'h0009827F , 32'h000BC560 , 32'hFFFD7EFD , 32'hFFFCA92E , 32'h00078903 , 32'hFFF9978A , 32'h00079EBA , 32'h0000A6C6 , 32'hFFF2674B , 32'h00008ADD , 32'h00058440 , 32'h0004A34C , 32'hFFFD95E8 , 32'h00020666 , 32'hFFFE6A65 , 32'hFFFF722A , 32'hFFF187DB , 32'hFFFB763B} , 
{32'hFFFE9D1A , 32'hFFFF7BBA , 32'h0002A889 , 32'hFFFEC897 , 32'h0004F6AA , 32'hFFF95272 , 32'hFFFEDBCD , 32'hFFFF66F3 , 32'h0001893C , 32'h000A3F3F , 32'hFFFFEDA0 , 32'h0001F021 , 32'hFFFA0E24 , 32'hFFFD7089 , 32'hFFFD0D79 , 32'hFFFF91D2 , 32'hFFFE2781 , 32'h0000E51F , 32'hFFFC1B27 , 32'hFFFAB354 , 32'h0002D439 , 32'hFFF2C95F , 32'h000418A3 , 32'h0004FEE2 , 32'h0005F43B , 32'h0008C52C , 32'hFFFD4B25 , 32'hFFFCD794 , 32'h00037D9F , 32'hFFFF3E04 , 32'h0001ED20 , 32'h00041348 , 32'h000D883B , 32'hFFF9FCFA , 32'h00007012 , 32'h00027952 , 32'hFFFFEBBA} , 
{32'h00080EB4 , 32'h0008BDCB , 32'h000D7881 , 32'h0001BBF2 , 32'h00114EBD , 32'hFFFD295D , 32'hFFF9C46F , 32'hFFFF5921 , 32'hFFFE9957 , 32'hFFFE4F3B , 32'hFFFA6819 , 32'h000BF4FF , 32'h000260FF , 32'hFFFF529F , 32'h00007D33 , 32'hFFFFACB9 , 32'h00024694 , 32'h000680AB , 32'hFFFC8EEF , 32'h0004D34B , 32'hFFF8798D , 32'h000392BC , 32'h0004A3FF , 32'h000ABC08 , 32'h00073C67 , 32'hFFFA2B86 , 32'h000518C5 , 32'hFFFB875E , 32'h00005930 , 32'hFFFB8031 , 32'hFFFD1B01 , 32'h00020830 , 32'h0002FF1D , 32'h0000F766 , 32'h000129D6 , 32'h0003CC39 , 32'hFFF62ADB} , 
{32'hFFF7B3D3 , 32'hFFF27960 , 32'hFFF52AFA , 32'hFFFE0E31 , 32'hFFF2D4C3 , 32'hFFFACF35 , 32'hFFF469A9 , 32'h000079BD , 32'hFFF5CAA4 , 32'hFFF9E89E , 32'hFFFDB818 , 32'hFFF9D53C , 32'h0004C53F , 32'h00010CDA , 32'hFFF5875F , 32'hFFFBC981 , 32'h0003BD21 , 32'h00040AAF , 32'hFFFFE567 , 32'h000930D5 , 32'h000532FC , 32'hFFFE0121 , 32'h00051472 , 32'h00016840 , 32'hFFF63E21 , 32'hFFFB38D7 , 32'h000274F0 , 32'h0007CEAE , 32'hFFFFFD65 , 32'h00039D70 , 32'h0000CF87 , 32'hFFFE32D1 , 32'h0001AA6B , 32'h0004630E , 32'h0004AA26 , 32'hFFF751EF , 32'hFFF64545} , 
{32'h03FFC9A4 , 32'h02F8A6C4 , 32'hFF9508BF , 32'hFD0A8454 , 32'h0628A5C8 , 32'h01374248 , 32'h07A4BA40 , 32'h06DFB360 , 32'h037AC964 , 32'hFE7E19DC , 32'h0CD1B020 , 32'hF27EF0A0 , 32'h069C8510 , 32'hFAC01E50 , 32'h04C13A68 , 32'hF8DA7EF8 , 32'h03CBC610 , 32'hF5D95F40 , 32'h046F2008 , 32'hF6AA1010 , 32'hFE979B18 , 32'hFDF6850C , 32'h04FE55B8 , 32'h05DC2120 , 32'hFFC39785 , 32'h028D39A4 , 32'hFD24B4E8 , 32'h062A45F8 , 32'h0FAAB9B0 , 32'hFDC00220 , 32'h093E6AD0 , 32'hF4F362C0 , 32'h0A6D1810 , 32'hF714B290 , 32'hF8390DE8 , 32'h02ACB2A8 , 32'h011976A0} , 
{32'h3585E5C0 , 32'hFFC8BB53 , 32'hF28553B0 , 32'h2E353700 , 32'h0A440450 , 32'h0FC33DE0 , 32'h2B2DFBC0 , 32'h02A7C2B4 , 32'hEC74EC20 , 32'h0C842430 , 32'h3D50AB80 , 32'hF4747CB0 , 32'hF241E270 , 32'hE5C845E0 , 32'hF9F66518 , 32'hEEAF0C20 , 32'hF073C6C0 , 32'hE5ED3860 , 32'hF8DBC900 , 32'hF6BAEDC0 , 32'h10081E80 , 32'h02B3E5B0 , 32'h115316E0 , 32'h03996E68 , 32'hFE2854AC , 32'h1DEAD300 , 32'hD617DA80 , 32'h20B1D180 , 32'h1ACECD00 , 32'hD8656CC0 , 32'h1FE38960 , 32'h0B5A6B00 , 32'hDA1F0100 , 32'h108E04A0 , 32'hF4B42FE0 , 32'h02EAFBC4 , 32'h24A364C0} , 
{32'h2656BE00 , 32'h2A62A180 , 32'h00AF14E2 , 32'h1E442C60 , 32'h30BB4580 , 32'hFEF63A30 , 32'h53135A00 , 32'h06953ED8 , 32'h0F0E1B10 , 32'h03B04DF0 , 32'h0A9A58A0 , 32'h1FA2C900 , 32'hF055E3A0 , 32'hE83B8040 , 32'h0D748420 , 32'hE4AF3C00 , 32'hE2348180 , 32'hDF736740 , 32'hFBEF8D30 , 32'hF5FF2DB0 , 32'h0E3CBAA0 , 32'h004BB670 , 32'h01A9F0B4 , 32'hFFF6DFBC , 32'hF9B81D28 , 32'h09AD4E00 , 32'hE8E32E00 , 32'h01207F88 , 32'h0D4DB4F0 , 32'hE941B620 , 32'hFCE307F4 , 32'h2B89C340 , 32'hD99DF1C0 , 32'h07DA2CB0 , 32'hE2375360 , 32'h0EAB5EF0 , 32'h2A8A1580} , 
{32'h0596A5C0 , 32'h213FE340 , 32'h0FF78140 , 32'h2E876D00 , 32'h145984A0 , 32'hDB31E940 , 32'h4C59F800 , 32'hF20A1660 , 32'h26A790C0 , 32'h05180988 , 32'h1CE3BA40 , 32'h0A014110 , 32'h02E65EFC , 32'hDDEF1240 , 32'h045A9FA8 , 32'hE05444C0 , 32'hED5CC4E0 , 32'hD431C440 , 32'hF8979D68 , 32'h02320994 , 32'hFD7A2A70 , 32'hF28B56A0 , 32'hFFF72054 , 32'h01316BF8 , 32'h0C82DB50 , 32'h0E6A5630 , 32'hF55A41A0 , 32'h0EA468E0 , 32'hF096D4B0 , 32'hF1E5B740 , 32'hF2C5C990 , 32'h1A245C60 , 32'hED230220 , 32'h28ABDE00 , 32'hF14AD0D0 , 32'h07DF69B8 , 32'h25623B00} , 
{32'h0B28BBA0 , 32'h2AB55380 , 32'h2492CEC0 , 32'h1FB2C000 , 32'h25FC6780 , 32'hFD4DC478 , 32'h45BD6A00 , 32'h0A293CB0 , 32'h1B413C00 , 32'hFED8293C , 32'hF91F9858 , 32'h2D5C86C0 , 32'hFB5251C8 , 32'hE8A7D7C0 , 32'h07EBB458 , 32'hEC1C01A0 , 32'hF62DD1A0 , 32'hE7C26860 , 32'hF8C7DE68 , 32'h043504D8 , 32'h039788F8 , 32'hF7205520 , 32'hEB958420 , 32'hF6CB2EA0 , 32'h04805878 , 32'hF8DBEA90 , 32'hFA360948 , 32'hFC59525C , 32'hFDFB1D70 , 32'h0F7D3190 , 32'hF1327DA0 , 32'h15D6A600 , 32'hF8AB7148 , 32'h16DAE9E0 , 32'h065ACEA8 , 32'h1BB90160 , 32'h011FF21C} , 
{32'hF01F97D0 , 32'h1AA2DD60 , 32'h1FFF7CC0 , 32'h1D1286A0 , 32'h000B9167 , 32'hE5041AE0 , 32'h2A0F47C0 , 32'hFBFBA510 , 32'h2C852BC0 , 32'hF4AA28D0 , 32'h2C434500 , 32'h0CF58180 , 32'hEA6A9F80 , 32'hDF3E2DC0 , 32'h15F22880 , 32'h0914AC40 , 32'hF7F77BB0 , 32'hF636EBB0 , 32'hFA3C55E8 , 32'h19970FC0 , 32'hEBA15AE0 , 32'hEF18A380 , 32'h0CA7F000 , 32'h05FC8BC8 , 32'h193A4F60 , 32'hF0888100 , 32'hEB5D3EC0 , 32'h030327AC , 32'hFB574BB8 , 32'hF5039DE0 , 32'h0AFD6240 , 32'hE7E21120 , 32'h04795120 , 32'h10724AC0 , 32'hFCCBEE90 , 32'hEC911A60 , 32'hF6AC42B0} , 
{32'hE9B5D400 , 32'h0A3D5240 , 32'h45298F80 , 32'h21A38B40 , 32'h19B7F0C0 , 32'hDB6F7600 , 32'h04186938 , 32'hF47123F0 , 32'h1AEEDC80 , 32'h05923150 , 32'h03BB03F4 , 32'hF2CE5AF0 , 32'hF6B8D7A0 , 32'hDA46F0C0 , 32'hFE473204 , 32'h14EA6480 , 32'hF42FA1B0 , 32'hE3311460 , 32'hF9B7D1A8 , 32'h04544460 , 32'hEA535340 , 32'h036221E8 , 32'h06A416C8 , 32'h142BACC0 , 32'h01BFA11C , 32'h08A61C90 , 32'hE769E900 , 32'hFB312338 , 32'hEC26FEE0 , 32'hFF4AE0A4 , 32'h12EB5C40 , 32'hD7C8F580 , 32'hFC140228 , 32'h081C7EB0 , 32'h04A14030 , 32'hFFFA5C42 , 32'hEA10DA20} , 
{32'hBED5A300 , 32'hEBF9D1E0 , 32'h3F6A4F40 , 32'h31550500 , 32'h067848F8 , 32'hD34C8800 , 32'hFF7200F8 , 32'hE7E805A0 , 32'h05B39BE8 , 32'h0D5BCDE0 , 32'h27823840 , 32'hC0B56E00 , 32'hFB5BBAE8 , 32'h12A37860 , 32'h06BD3508 , 32'h2B3D0280 , 32'hF89C4E18 , 32'h184A4F60 , 32'hE8AD72A0 , 32'h2E027A40 , 32'h113F39C0 , 32'h004D13A9 , 32'h09C90C60 , 32'h0AB46730 , 32'h155DF140 , 32'h1FC5BB20 , 32'h04863498 , 32'hF6535E40 , 32'h25C818C0 , 32'h05FB8190 , 32'hE98DE740 , 32'h063ECD50 , 32'hF3B0CD60 , 32'hDF8FC240 , 32'hF3AA5E70 , 32'hF9F333A0 , 32'h153619C0} , 
{32'hCA1C57C0 , 32'hCB3AED80 , 32'h342E46C0 , 32'h11C15480 , 32'hF5415140 , 32'hDAFBA2C0 , 32'hDC357040 , 32'hF548BA90 , 32'hEC37A240 , 32'h0B152AC0 , 32'h184444C0 , 32'hD2312300 , 32'hEC6936A0 , 32'h11A1D8A0 , 32'h25386C40 , 32'h17EE0060 , 32'hD92C6B80 , 32'h29E60940 , 32'hFC2E612C , 32'h12F32C40 , 32'hF5246310 , 32'hF755B870 , 32'hF26940D0 , 32'hF9BD1070 , 32'h171AA920 , 32'h1AD8B460 , 32'h003AA1BF , 32'hF8DBDD98 , 32'h1E37EB00 , 32'h12733580 , 32'hF73C51C0 , 32'hEA9C9600 , 32'hEC1A4420 , 32'hF3C82920 , 32'h08E7D670 , 32'hFD521E68 , 32'h055C7628} , 
{32'hD8AE3B80 , 32'hC85E8600 , 32'hB3C4E900 , 32'hF121AAC0 , 32'hA62EAE80 , 32'hCAF4E600 , 32'hF5DD9C70 , 32'hF999F780 , 32'h14D841C0 , 32'hED513980 , 32'h0A6F10C0 , 32'hD56CCC00 , 32'h0D187F90 , 32'h265ADFC0 , 32'h1FA11CC0 , 32'h09373A30 , 32'hF83177D8 , 32'hF3E9E730 , 32'h0C424A60 , 32'hEA176A80 , 32'h044D1ED0 , 32'hFA0CE050 , 32'h03598B2C , 32'h197CC180 , 32'hD860FF00 , 32'hF0B9BE20 , 32'hFF1BA229 , 32'h1BF75220 , 32'hFF25246B , 32'h1C20F7A0 , 32'h02FC247C , 32'hF5D4ACA0 , 32'hE27C67E0 , 32'h2B0716C0 , 32'h00001018 , 32'h3C35B680 , 32'hF3093D20} , 
{32'hD9996F40 , 32'hD27BAC80 , 32'hD5FBBD00 , 32'hF86DE858 , 32'hA6993000 , 32'hEA166740 , 32'hFD7F3904 , 32'hBC901E80 , 32'hFD0C8F60 , 32'hFE92E0D0 , 32'h011050EC , 32'hF5698120 , 32'h0FBB1B40 , 32'h1E187DA0 , 32'h44EC7280 , 32'hDFF16880 , 32'h07883078 , 32'hC4D9BEC0 , 32'hF4D4D000 , 32'h19013A00 , 32'hE72474E0 , 32'h05E643C8 , 32'h06A58F70 , 32'hF5FD5F30 , 32'hE089B360 , 32'hFF80BFC3 , 32'hFFCE770A , 32'h303A9300 , 32'h13172200 , 32'hF226F080 , 32'hD148E380 , 32'h027BDC94 , 32'hEF4F8D20 , 32'hDE1EE000 , 32'h0393A118 , 32'hF0D05DB0 , 32'hFCC921F0} , 
{32'hEEF76220 , 32'hFC9E9620 , 32'hE982AC60 , 32'hFDFAD590 , 32'hD7CFC340 , 32'h0E051F30 , 32'hFD533D1C , 32'hE74663E0 , 32'hF7630990 , 32'h0EE06D00 , 32'hEE4CDCC0 , 32'h0B70A050 , 32'hF43F00F0 , 32'h015D0150 , 32'h3E25E900 , 32'h053801E0 , 32'h12CDF500 , 32'hFD4D3384 , 32'hEB851FE0 , 32'h09BD3D50 , 32'h022AA550 , 32'h139C02A0 , 32'hFB79CD30 , 32'h0F8F7EA0 , 32'h036D92B0 , 32'h1B29E6C0 , 32'h085D9050 , 32'h0D4132C0 , 32'hE32BFFE0 , 32'hF7894D50 , 32'hF24AAC80 , 32'h14064760 , 32'hEFAEEC40 , 32'hD74E6380 , 32'hEECA5B00 , 32'h06400730 , 32'hF6B70DA0} , 
{32'h008876B3 , 32'hFEA0F79C , 32'hEE5C8E20 , 32'h1EABC0E0 , 32'hF4EA6760 , 32'hFFD176C7 , 32'hEAE67BA0 , 32'hD1A21100 , 32'hF862B978 , 32'hED580D60 , 32'hE8ADFFA0 , 32'h0C726A40 , 32'hDB3F0B80 , 32'hFA0112A0 , 32'h1A162AE0 , 32'h0C934090 , 32'h2183A5C0 , 32'h08400130 , 32'hFD98E770 , 32'h0A4883C0 , 32'h09C49DF0 , 32'h0D594370 , 32'hE8080560 , 32'h1338E760 , 32'h294F4980 , 32'h16324D40 , 32'h0486E358 , 32'h0347BC68 , 32'hDB315B40 , 32'h02E4FAA4 , 32'hFB93DAE0 , 32'h00A804DF , 32'hEB9E4F40 , 32'h067D5AA0 , 32'h100E0CC0 , 32'hEB046620 , 32'hF1663CF0} , 
{32'hE95FCB20 , 32'hFFC62F80 , 32'hFA517008 , 32'h0D69D1D0 , 32'hEED09BA0 , 32'h172D1440 , 32'hF5461640 , 32'h0553D350 , 32'hF644FE30 , 32'h159BAD20 , 32'hF1BF8710 , 32'hFBEC8B28 , 32'h018C76B4 , 32'h00A93A00 , 32'h2958B980 , 32'h16044B80 , 32'h288C2FC0 , 32'hE35C9560 , 32'h08E0AC20 , 32'h0C6B18B0 , 32'h38E463C0 , 32'hFC091298 , 32'hF2113750 , 32'h174DFF20 , 32'h36DC2400 , 32'h04B85A60 , 32'hE36A6600 , 32'hFA360AA0 , 32'hF2AF1220 , 32'hFBFCEE68 , 32'h071F8B00 , 32'h19DCBCC0 , 32'hFC774E04 , 32'hFB3B9D70 , 32'hFE252EB4 , 32'h06E112D0 , 32'h111DBC40} , 
{32'hF806FDE8 , 32'hFE201764 , 32'hFFC97E5B , 32'h1728D260 , 32'hFE852298 , 32'h042A2CE0 , 32'hF58ED4D0 , 32'h086A6BE0 , 32'hFCCC1ED8 , 32'hFF43BA5F , 32'hFCF295C0 , 32'h02E87B64 , 32'h0CFF5570 , 32'h06179550 , 32'h11F8D880 , 32'h15061920 , 32'h0972D1A0 , 32'h061CFC28 , 32'h0F7E0510 , 32'h093B3330 , 32'h16276C00 , 32'h09D16260 , 32'h05C747E8 , 32'hFAC48BC8 , 32'h148BB160 , 32'h11BBEA20 , 32'hF5B7C270 , 32'hF5E69370 , 32'hF0D06FC0 , 32'hFF5EC22D , 32'hF83CCA88 , 32'h0292C0A0 , 32'hF98A1DC8 , 32'h03078EA0 , 32'h078C4B28 , 32'h041379C0 , 32'hF6BC8810} , 
{32'hFC9482E8 , 32'h08A6FC70 , 32'hF255BE70 , 32'h1CFF1AA0 , 32'hF4BFC600 , 32'h0B7795B0 , 32'hE58950E0 , 32'h50983600 , 32'hFB431970 , 32'h03C40070 , 32'h1ACA7E00 , 32'h0B8E88D0 , 32'h650D8980 , 32'h246F0EC0 , 32'hFCC12500 , 32'h24E1AC80 , 32'hF21D21B0 , 32'hD4F359C0 , 32'h39838000 , 32'h12F49B40 , 32'h1371D9A0 , 32'hDF543000 , 32'h10520BA0 , 32'h1C6E6700 , 32'h0A906390 , 32'h102D0AA0 , 32'hFFDE1EC6 , 32'h04752740 , 32'hEA4477E0 , 32'hFD5FD4B8 , 32'hDCF230C0 , 32'hF77E6740 , 32'h065F12C0 , 32'h19BB00E0 , 32'hF4654AF0 , 32'hF936B3A0 , 32'h0DF41560} , 
{32'hFD296D80 , 32'hF445E470 , 32'hF9027898 , 32'h2875AD80 , 32'hF18900C0 , 32'hFB857040 , 32'h12E3BC20 , 32'h0C91CC10 , 32'hE63321A0 , 32'hD6188900 , 32'hFA881448 , 32'hF1ACDB50 , 32'h1B24DC00 , 32'h0F052F40 , 32'h042C8860 , 32'h11CB40E0 , 32'hFFF2382F , 32'hF15CEA90 , 32'hFD6965A0 , 32'h01A256A4 , 32'h04D01C30 , 32'hF7099F40 , 32'h0EDE2860 , 32'hF9A3CC50 , 32'hF8741118 , 32'h0DD26700 , 32'h0D3FB940 , 32'hF25DFBA0 , 32'hF272C360 , 32'h1115E120 , 32'h09724D50 , 32'hF837C938 , 32'h1338EB60 , 32'h00A01B45 , 32'hFE9868A8 , 32'hFD51D704 , 32'h0925B2C0} , 
{32'h0778BCC0 , 32'h110C6C20 , 32'h0C6CDE70 , 32'h0595A4A8 , 32'h01F463F8 , 32'hFFF32981 , 32'hFAE33928 , 32'h1658D160 , 32'h048DE488 , 32'h0EA652A0 , 32'h04F9B1D8 , 32'hF0623D10 , 32'h1B721440 , 32'h0F8A30A0 , 32'hF9FE6810 , 32'hE5BC8E60 , 32'h00A3E10D , 32'hE78CDA40 , 32'hF1F58BF0 , 32'h0B09FFC0 , 32'h19947C20 , 32'hECA0FAA0 , 32'h09C36E00 , 32'h16F9F8A0 , 32'hFE4E8A68 , 32'hD60E9E80 , 32'h07B31B80 , 32'h05264E68 , 32'hF30D9D00 , 32'h079579B0 , 32'hFDCA7278 , 32'h039D1F90 , 32'h0301E508 , 32'hFBC2B1E8 , 32'h038478F4 , 32'hF4AFD2C0 , 32'hF3CFF6A0} , 
{32'h05BF1E68 , 32'hFBEF8630 , 32'hFBFF5200 , 32'hF7BEEEF0 , 32'hFDACD860 , 32'h07B9EC80 , 32'hFC8B0FA8 , 32'h10906260 , 32'h072718B0 , 32'hF61E5070 , 32'h07471FB0 , 32'hFCF8ECFC , 32'h02F7308C , 32'hEF830360 , 32'hEFEDD5A0 , 32'hF790D5D0 , 32'hF985BA10 , 32'hE51E0D40 , 32'hEF4CC0A0 , 32'hF0ABBC10 , 32'hEF904700 , 32'h0E84E660 , 32'h0041C289 , 32'hFF73EDF5 , 32'h097A9B50 , 32'h08EC7B30 , 32'hFF2ABEC5 , 32'h0EDA2BE0 , 32'h0247D044 , 32'hF75F03A0 , 32'hFC6B1E88 , 32'hE9013720 , 32'h09744880 , 32'h027EA1F4 , 32'hF8276008 , 32'hFC40CB80 , 32'h0BFCE460} , 
{32'hFE1D42C8 , 32'hDAD2DE00 , 32'hFB82D818 , 32'h17E7F3E0 , 32'hF5178EE0 , 32'h1565A3E0 , 32'h0FEB8540 , 32'h3B6EF240 , 32'h19873840 , 32'hF99194B0 , 32'hC925FC00 , 32'hF2E82660 , 32'hE98F5C00 , 32'hE1601560 , 32'h003A77CB , 32'hBC363B00 , 32'hD6B26140 , 32'hF5FCE890 , 32'hED2CB2A0 , 32'hEE987C20 , 32'hEC29E520 , 32'hD7550280 , 32'hF46E5040 , 32'hE8D0E1E0 , 32'h175F8900 , 32'hF79880C0 , 32'h3BFF08C0 , 32'hFD5DAF8C , 32'hFBA46C90 , 32'hDAC70340 , 32'hF89AFB88 , 32'hFC171414 , 32'hE8EB36A0 , 32'h26B79B00 , 32'hFDBD88B4 , 32'hFB429F90 , 32'h0572D0A0} , 
{32'hFCBDA764 , 32'hF5C4B7E0 , 32'hF9B4CF20 , 32'h0B47A630 , 32'hFD9EC2F0 , 32'hFF2ED2B1 , 32'hFCBD0EC0 , 32'h05F2B620 , 32'h0D024340 , 32'hFD34B2C8 , 32'h018D68D0 , 32'h0A5497F0 , 32'hFDB4E194 , 32'hFCD1710C , 32'h02230438 , 32'hF56D9930 , 32'h042A51C0 , 32'h023202D8 , 32'hF6677DA0 , 32'hF2B5BBA0 , 32'h0ACA9840 , 32'h0175998C , 32'hFE4F78C4 , 32'h0FECC280 , 32'hFFC13D4E , 32'h077771B0 , 32'h0F992540 , 32'h043FABC8 , 32'h03878984 , 32'h015968C0 , 32'h00C77200 , 32'hF9D4F480 , 32'hF69730A0 , 32'h05EBE610 , 32'hF7B08D40 , 32'h057C2AF8 , 32'hFB208E40} , 
{32'h0020628B , 32'h001A1AE4 , 32'hFFC08EB0 , 32'h005BEEB9 , 32'h0040B127 , 32'h00609C66 , 32'hFFD8F801 , 32'h00274F9D , 32'hFFED8437 , 32'h00430329 , 32'hFFCC98D3 , 32'hFFC00F74 , 32'h00538223 , 32'hFFE54436 , 32'hFFC9326A , 32'h00298ECB , 32'h0066CFFA , 32'hFFAA8AD5 , 32'hFFD8D4CE , 32'hFFD6B182 , 32'h00424B4F , 32'h00A0A6D8 , 32'h00500C4C , 32'hFFFDF0EC , 32'hFFDDA2FF , 32'hFF94994B , 32'h003E2665 , 32'h0049DF72 , 32'h0017A39C , 32'hFF93760F , 32'hFFFB4357 , 32'h0049409F , 32'h00440385 , 32'hFFF2A212 , 32'hFF882612 , 32'h001A1623 , 32'h002092C6} , 
{32'h0032F6EE , 32'hFFE44B16 , 32'hFFAA8D7E , 32'h0089FD7A , 32'h002FE071 , 32'h00301AF6 , 32'hFFF7DC48 , 32'h002172F5 , 32'hFFC20D09 , 32'h000FE91F , 32'hFFD4884F , 32'hFFD0F740 , 32'h003E7EF0 , 32'h001AAF70 , 32'hFFD0E701 , 32'hFFECB278 , 32'h0095B92A , 32'hFFB61FE0 , 32'hFFBC7EE8 , 32'hFFB25A1E , 32'h0049AEDF , 32'h00D3D1E8 , 32'h005DFF71 , 32'hFFF82527 , 32'h0007B328 , 32'hFF87BD61 , 32'h002E2931 , 32'h003F0731 , 32'h002B6ED0 , 32'hFF7D732C , 32'hFFD802E7 , 32'h0028E505 , 32'h005E8191 , 32'h0004B517 , 32'hFF6EDDBC , 32'h00147584 , 32'h00031BA0} , 
{32'hFFF705D5 , 32'h00009D68 , 32'hFFF3F97F , 32'h0002AA79 , 32'h00047C2A , 32'h00057C69 , 32'hFFF7B25A , 32'h00031B54 , 32'h0008A295 , 32'hFFFB3C54 , 32'h0001243D , 32'h0001AC92 , 32'h00077BE1 , 32'hFFF6C3CA , 32'h0004861F , 32'h00019593 , 32'h00088B78 , 32'h0004B6EC , 32'h00030CE3 , 32'h0003B202 , 32'hFFFDDD43 , 32'hFFF60084 , 32'h0003FC02 , 32'h00005A56 , 32'hFFFE4567 , 32'h0000297B , 32'h00094554 , 32'h0001839A , 32'h000C868D , 32'hFFF8D3A4 , 32'h0002A964 , 32'hFFFFAA4A , 32'h0003A0BB , 32'hFFF561EC , 32'h0003F8B9 , 32'h000BB0F7 , 32'h0008058B} , 
{32'h00013E8D , 32'h000DC001 , 32'hFFFCCF48 , 32'h0006A0CC , 32'hFFFCC592 , 32'h0004AFF4 , 32'h0005A5CA , 32'h0000286F , 32'hFFFF067A , 32'hFFF47B0D , 32'hFFF83EAF , 32'hFFFA5A83 , 32'h0007BDED , 32'h000557CF , 32'h0008B887 , 32'h00044AE6 , 32'hFFFBB317 , 32'hFFFFE3DA , 32'h000409FA , 32'h0001FDC8 , 32'h0000A51E , 32'h0008286A , 32'hFFFC2824 , 32'h0000A9E6 , 32'h00042953 , 32'hFFFCBD6E , 32'hFFFE1824 , 32'h0000F0F9 , 32'hFFFD9AE0 , 32'h00004601 , 32'hFFFEA52E , 32'hFFF263E6 , 32'hFFFA4863 , 32'hFFFA37EF , 32'h000115B8 , 32'hFFF88512 , 32'h0000F87B} , 
{32'hFFF8B06B , 32'h00060100 , 32'h00015754 , 32'hFFF973CD , 32'hFFFA326C , 32'h00060215 , 32'h00065CCF , 32'hFFFD3AE4 , 32'hFFF72CFF , 32'h000038D8 , 32'h00044C67 , 32'hFFFBEA84 , 32'h00063740 , 32'hFFFF9336 , 32'h00001863 , 32'hFFFE1649 , 32'hFFF92A44 , 32'h00031A85 , 32'h00090786 , 32'hFFF8E635 , 32'hFFF9B378 , 32'h0003125F , 32'hFFFCBF98 , 32'h0008591F , 32'h000649E7 , 32'h00023D9C , 32'h000411A5 , 32'hFFF77780 , 32'h00059C03 , 32'hFFFCE8D9 , 32'h00009ECC , 32'h000A1359 , 32'hFFFF52C8 , 32'h0005CEFF , 32'h0001DE0A , 32'hFFFF91D2 , 32'hFFFC688D} , 
{32'hFFFA0348 , 32'hFFF7264D , 32'hFFEECB49 , 32'hFFF59882 , 32'hFFF05721 , 32'hFFF80325 , 32'h00027C6E , 32'hFFFB5221 , 32'hFFFEF479 , 32'hFFF96EA4 , 32'h0004C0B5 , 32'hFFF75A8A , 32'h00046210 , 32'hFFFAE238 , 32'h00009357 , 32'hFFF795E0 , 32'h0012A927 , 32'h0002B492 , 32'h00063D77 , 32'hFFF90F8F , 32'hFFF31C47 , 32'h00011EFA , 32'hFFFDCB9A , 32'hFFFEB878 , 32'hFFFA328D , 32'hFFF4E129 , 32'hFFFF9903 , 32'hFFFB9EC8 , 32'hFFEBBA37 , 32'h00088273 , 32'h00107FCC , 32'hFFF9CCDC , 32'h0005C6EE , 32'hFFFCD704 , 32'h00007387 , 32'hFFF5B26B , 32'h00013829} , 
{32'hFFFC35CF , 32'h00087A7B , 32'h00030881 , 32'h0002D7DD , 32'hFFFF7C01 , 32'h0002023C , 32'h0001CA7F , 32'hFFFE0C8A , 32'h0006E598 , 32'hFFF8E7EE , 32'hFFFA26D8 , 32'hFFFB43C7 , 32'hFFF92A2D , 32'h00017E23 , 32'h000382AD , 32'hFFFE0B17 , 32'h0000B16E , 32'h0001F37B , 32'hFFF85B08 , 32'h000107F9 , 32'h00032FE3 , 32'h00016A60 , 32'h00014D81 , 32'hFFFFCC3D , 32'hFFFA5C85 , 32'hFFFD6735 , 32'hFFFFCE1D , 32'h000598B5 , 32'hFFFEE9C7 , 32'h00077FF8 , 32'hFFFBD2FA , 32'hFFFC2B07 , 32'h0000C7F6 , 32'h0002A365 , 32'h0003058D , 32'hFFFFD25B , 32'hFFFC7D15} , 
{32'h000BC009 , 32'h001814DA , 32'hFFF8D0CD , 32'h003522A9 , 32'hFFA47D92 , 32'hFFAC3124 , 32'hFFDA6277 , 32'hFFFBCA50 , 32'h001E005F , 32'hFFE17E20 , 32'h00348350 , 32'hFFFB3A4B , 32'hFFBF1EAC , 32'h000C2108 , 32'h002C9ED1 , 32'hFFF37501 , 32'hFFBF5775 , 32'hFFE3B919 , 32'h0000F589 , 32'hFFDF24D3 , 32'hFFDD1E7C , 32'hFFDD5A02 , 32'hFFFB338F , 32'h002D127E , 32'h00655410 , 32'hFFD3EF8A , 32'h001FABEA , 32'h000E1180 , 32'h0010C638 , 32'h0049E9C7 , 32'hFFDC1010 , 32'h002BD37A , 32'h000E076D , 32'hFFFA6B73 , 32'hFFC6DEAD , 32'hFFED49AE , 32'h004121D6} , 
{32'hE76B43A0 , 32'hE23BE080 , 32'h1D7DE960 , 32'h1A1F44C0 , 32'h24E13740 , 32'h0452B5A8 , 32'h6994B480 , 32'h0191BFF4 , 32'h12A61740 , 32'h1BCD1380 , 32'h265CD5C0 , 32'h23DC6980 , 32'hE7342840 , 32'hF51301A0 , 32'hE6041E80 , 32'hF8BE7FF0 , 32'hE28E78E0 , 32'hBC2F4A00 , 32'hF9CAD7B8 , 32'h0466DF48 , 32'hEA97D640 , 32'hFE770274 , 32'h109A8400 , 32'hFBC0B560 , 32'h0FE1F020 , 32'h0092F2D4 , 32'hE8895AA0 , 32'hF21A8550 , 32'hD33B12C0 , 32'h176562A0 , 32'hF62B4800 , 32'hF3614020 , 32'hFDE28A0C , 32'hFF26F730 , 32'hEA3ACBC0 , 32'hE5797260 , 32'hF2D7C110} , 
{32'hD97851C0 , 32'hEF7CDA20 , 32'h294AA700 , 32'h1533C360 , 32'h0189D5B8 , 32'hF7855340 , 32'h28257500 , 32'hFCF98608 , 32'h13F1C800 , 32'h063E3670 , 32'h0EB63CA0 , 32'h1632A9C0 , 32'hF5BB99F0 , 32'hF8EAD680 , 32'hEE042820 , 32'hFED1C11C , 32'hF765D4B0 , 32'hFC1AAF2C , 32'h00F9024E , 32'hFBC77BF8 , 32'hEC4D6EE0 , 32'h07298908 , 32'h0CA43520 , 32'hE14F41E0 , 32'h08556E20 , 32'h0A31DAA0 , 32'hF2463840 , 32'hF6C688D0 , 32'hFD96D9A8 , 32'h0739F190 , 32'h10004080 , 32'hFCEFEDC8 , 32'h11992B00 , 32'hF0181320 , 32'hFF2DA538 , 32'hF32F4E90 , 32'h02221034} , 
{32'hC42C2880 , 32'hF02FB140 , 32'h35A1FA00 , 32'hEECC02A0 , 32'h1F4787C0 , 32'hF9C36F40 , 32'hFD4503EC , 32'h13D07E00 , 32'h2FB11140 , 32'hECAAEEA0 , 32'h234DE180 , 32'h13C8CB40 , 32'hE4C185E0 , 32'hD4426A40 , 32'h02B05790 , 32'hF6DD2650 , 32'hDD83A040 , 32'hFCE54380 , 32'h0B0C8DD0 , 32'h00F5B492 , 32'hCD0F3040 , 32'h12868FC0 , 32'h19FA76E0 , 32'h01C8D0A4 , 32'hF5637EA0 , 32'hFA97B108 , 32'hD12218C0 , 32'hFA3A5B80 , 32'hE3109480 , 32'h09C6A1A0 , 32'h33991900 , 32'h18E2A3E0 , 32'hF5702E60 , 32'h0F630FE0 , 32'hF349AA10 , 32'h11ADBDC0 , 32'hF4263650} , 
{32'hE17B8560 , 32'h0A3E6AF0 , 32'h35D10E40 , 32'h1043B8C0 , 32'hF7EDE4E0 , 32'hEBD7D2A0 , 32'hFD2F67BC , 32'hF724FDA0 , 32'h23613240 , 32'hE118C800 , 32'h2F3C2040 , 32'hF491BBC0 , 32'hE35C1920 , 32'hE69A2740 , 32'hEADF8540 , 32'hE28DA8C0 , 32'hEB26FF20 , 32'hDE8A3E40 , 32'h0BDE2C80 , 32'h0D8F3910 , 32'hF0B88580 , 32'hF6AC5BF0 , 32'h14741600 , 32'h1B50DFE0 , 32'h10123C60 , 32'hE1A93380 , 32'hE22458C0 , 32'hF1253D80 , 32'hE0DF3BE0 , 32'h2AEE5240 , 32'h190F9420 , 32'hFFFB8176 , 32'h0242035C , 32'hFB03EC18 , 32'h06C6C3D0 , 32'hEF09DFA0 , 32'hF5D892E0} , 
{32'hBEEA2080 , 32'hF98600A8 , 32'h47FF6D00 , 32'hF1CA05F0 , 32'h28263B00 , 32'hE662DF80 , 32'hF8180918 , 32'h1C0D1220 , 32'h28C8A800 , 32'hF0B8B950 , 32'h226D8340 , 32'h114793A0 , 32'hE49E3140 , 32'hD7310B00 , 32'h189DF520 , 32'hF63C1870 , 32'hE3ADC040 , 32'hE1267A20 , 32'hF4884A60 , 32'h0C25DB10 , 32'hE89BCA60 , 32'hFD6EDF94 , 32'h0A551B60 , 32'h11580A20 , 32'h067ACA30 , 32'hF9182120 , 32'hD63F9B00 , 32'h047B4C98 , 32'hF9E5FD08 , 32'hEFA106C0 , 32'h25B10740 , 32'h0C2DDE90 , 32'hEBDF77A0 , 32'h1C616460 , 32'h1DF08D80 , 32'hCF477580 , 32'hE7AB67E0} , 
{32'hC37C9D00 , 32'hDC900780 , 32'h4934B580 , 32'h23DAC900 , 32'h0E961F80 , 32'h034D0A98 , 32'hF3ADBCA0 , 32'hF7916010 , 32'hFB4A3A78 , 32'hF445CB80 , 32'h4731E800 , 32'hD374A600 , 32'hEF1FA7A0 , 32'h12E89D20 , 32'h0C87DE40 , 32'hF9D1E6F8 , 32'hDDD6D240 , 32'h045DCD00 , 32'hEFC51680 , 32'h1D66E940 , 32'h0EFDCE30 , 32'hF5B1C240 , 32'hFEC339D0 , 32'h11FF72A0 , 32'h3E1E5F40 , 32'h0DD07870 , 32'h01D48C98 , 32'hF6E4B240 , 32'h020C0FF0 , 32'h13EFD240 , 32'hE45D7320 , 32'hFF9FA441 , 32'hED2C57C0 , 32'hF15E6900 , 32'h04091CC0 , 32'h0EFD8100 , 32'h0ACED4B0} , 
{32'hC00EBC80 , 32'hDB0CDA80 , 32'h4A95C980 , 32'hEC5D80C0 , 32'h09E93690 , 32'h115F7940 , 32'hC0EE26C0 , 32'h08BC2B30 , 32'h079E40E0 , 32'hEA834320 , 32'h338A0BC0 , 32'hDD324E80 , 32'hDE732980 , 32'h05911BA8 , 32'hF393AE00 , 32'hFBC6E688 , 32'hEC8D9580 , 32'h0DF7D240 , 32'hDE44BDC0 , 32'hFFBD66E0 , 32'h15113C60 , 32'h20AD2640 , 32'h1C5A8A40 , 32'h226A0440 , 32'h2B892CC0 , 32'hFDE89854 , 32'h1D5642A0 , 32'h09D63140 , 32'hFE1721E8 , 32'h046F7930 , 32'hD67773C0 , 32'hFE4ECDE4 , 32'h0669B9B0 , 32'hE95AF260 , 32'hFAAB4368 , 32'h0317730C , 32'h181B60C0} , 
{32'hD5C46C80 , 32'hBE396580 , 32'hF755CB90 , 32'h06C02D40 , 32'hAEDB3980 , 32'hF53B5A60 , 32'hEFA4AB80 , 32'hF13EBE00 , 32'h01661058 , 32'hFBB85CB0 , 32'h2B39E340 , 32'hAD904980 , 32'h18428180 , 32'h0679F4E0 , 32'h03A06C14 , 32'hFF426171 , 32'hF211D650 , 32'h0E481960 , 32'hFC9994D8 , 32'hF165D550 , 32'hE531DF80 , 32'hFAFF47A8 , 32'h03D60A28 , 32'h0BE3D370 , 32'h040791F8 , 32'hF8EF5C38 , 32'h08933560 , 32'hEE963500 , 32'hBF9AEE00 , 32'h2772AE00 , 32'h27B10B00 , 32'hEF651780 , 32'h0C3FC760 , 32'hE8F45F20 , 32'h066E3118 , 32'hEFD7F0C0 , 32'h13AEF4A0} , 
{32'hC140F280 , 32'hB95D5400 , 32'hD8477E00 , 32'hF4AAFB20 , 32'h901EF100 , 32'hD6387A00 , 32'hEDC235A0 , 32'hEF774420 , 32'h1FABB320 , 32'h0DFDD410 , 32'h29D6F8C0 , 32'hF5547BB0 , 32'h01C5734C , 32'h17A06D00 , 32'hF99E5518 , 32'hE35B5120 , 32'h0360ED20 , 32'hE8320540 , 32'hFD698668 , 32'h01AACFC0 , 32'hFCC8E014 , 32'h0BDF97C0 , 32'h0174F120 , 32'h051AA598 , 32'hF77F0BB0 , 32'h0B2D4480 , 32'h099F5480 , 32'h14D746A0 , 32'hD26A1E00 , 32'h0C375630 , 32'h1CE13640 , 32'hEF822680 , 32'hFBED1910 , 32'hE5C51580 , 32'h0B6387F0 , 32'h0BA37AE0 , 32'h36DA7580} , 
{32'hDF572140 , 32'hE834F060 , 32'hEAD8B560 , 32'hF41AFA30 , 32'hB5F89A80 , 32'hF6744190 , 32'hF5D98460 , 32'hDBF0B9C0 , 32'h08652B20 , 32'h0D9EE630 , 32'hED54FC40 , 32'h304FBE00 , 32'hF5610880 , 32'h18E11500 , 32'h1BE55160 , 32'h0F1425F0 , 32'h0FB6B1B0 , 32'hFDAB9CE8 , 32'h0DD80EB0 , 32'h1A640A40 , 32'h14600680 , 32'hDD1975C0 , 32'h179D71E0 , 32'hF10E3850 , 32'hFE78E31C , 32'h11B65980 , 32'hF36032E0 , 32'h1BFC6860 , 32'h120BCB20 , 32'h155969E0 , 32'h01EF0F64 , 32'h0ED7EF20 , 32'hE2CD1260 , 32'h0A5766A0 , 32'hFE934494 , 32'hC39EDE80 , 32'hFD26E818} , 
{32'hFCD0B690 , 32'hF78FD3A0 , 32'h08831D40 , 32'h0CA117B0 , 32'hE92061C0 , 32'h057447A8 , 32'hE8674540 , 32'hE4014500 , 32'h00696D10 , 32'h13790A40 , 32'hE5A2A6E0 , 32'h161DA780 , 32'h037B32B0 , 32'h00FFAA91 , 32'h166E3860 , 32'h178D2E60 , 32'h069ED1B0 , 32'hF2592640 , 32'hF3471650 , 32'h12CB1CC0 , 32'hE683F3C0 , 32'h073C62B8 , 32'hFFC392EE , 32'hFA5EEDB8 , 32'h001CA624 , 32'h12634FC0 , 32'h00308153 , 32'h060B8C18 , 32'hED1C44A0 , 32'h0266DA10 , 32'hF7568460 , 32'hFD797EA4 , 32'hF11BB4B0 , 32'h0DDC79F0 , 32'h07C91DE0 , 32'h0C08AFC0 , 32'hFF1A7413} , 
{32'hF76D3390 , 32'hEFA12840 , 32'h07FBBA00 , 32'h076E10A0 , 32'hE96EF800 , 32'h04DA58B0 , 32'hF1A22470 , 32'hFCF008F0 , 32'hF91BBCB0 , 32'h065D9DD8 , 32'hF81D4970 , 32'h25B11B00 , 32'hF51FAFB0 , 32'h0DFD8C50 , 32'h16C86460 , 32'hFFDFEB02 , 32'h13C6C540 , 32'hFAD60398 , 32'h24E05D00 , 32'h03455CB4 , 32'h09063A50 , 32'hF563E990 , 32'h04C41F10 , 32'h1FD3D5C0 , 32'h2D3EEE40 , 32'h1CC7AD60 , 32'h1176E780 , 32'h058A8698 , 32'hE775B560 , 32'h0DB53330 , 32'hEBF32F20 , 32'hEA0EB5A0 , 32'hE116E200 , 32'h08DC0380 , 32'h2CCC7940 , 32'h0D243F60 , 32'hF636C4B0} , 
{32'hF1CDA7F0 , 32'h03378D04 , 32'h037FC8EC , 32'h16F31660 , 32'hFE8AB0B4 , 32'h0E351590 , 32'hEA84AA20 , 32'hFA335950 , 32'hFFB197D0 , 32'h0B808EB0 , 32'h041FFBA0 , 32'hFD75C06C , 32'h01358A3C , 32'h02A3445C , 32'h0DB26850 , 32'h07C37640 , 32'h26E92380 , 32'hF59A31F0 , 32'h0D6B5850 , 32'h14FD4C40 , 32'h1F507C80 , 32'hEACACF60 , 32'hFFF51A02 , 32'hF5A3B430 , 32'h1549A0A0 , 32'hF94D5DB0 , 32'hFEE46D64 , 32'hF72B3100 , 32'h001B7EB2 , 32'h0B13D920 , 32'h09689950 , 32'h06CC4710 , 32'hFC044944 , 32'hFF30657A , 32'hFCB5F89C , 32'h107924A0 , 32'hF8266C00} , 
{32'hF7994BD0 , 32'hF0928480 , 32'h03D527B8 , 32'h2A9B5B80 , 32'h034E7D1C , 32'h208F7D80 , 32'hDD519980 , 32'hF8D98B60 , 32'hF13C3370 , 32'h04FE1AA8 , 32'h15DE0DA0 , 32'hFDE1486C , 32'h11A696E0 , 32'hE933D3C0 , 32'hEE8C3400 , 32'h07A89B28 , 32'h204F0840 , 32'hEE588020 , 32'hFB9B7130 , 32'h1C6572A0 , 32'h0CF92110 , 32'h09456CD0 , 32'h0DB8D1A0 , 32'hFE66653C , 32'h11AEB140 , 32'hF87A2388 , 32'hF07727A0 , 32'hF430CA20 , 32'h076D8578 , 32'hF3C93A60 , 32'hFDBB6908 , 32'hF4257A90 , 32'hE3AC0380 , 32'h088E2000 , 32'hEE612860 , 32'hFEC4D44C , 32'h100189E0} , 
{32'hF5B15E60 , 32'h04734390 , 32'h043327F0 , 32'h0EBF4160 , 32'h1C66D5E0 , 32'h237FA300 , 32'hE58B22A0 , 32'h1E388020 , 32'h04467698 , 32'hF712B940 , 32'h2906A8C0 , 32'hFCA905A0 , 32'h541E6680 , 32'hDF57B480 , 32'hE93B2FC0 , 32'hFEE723F8 , 32'h2176DD80 , 32'hDF03FD80 , 32'h2B458000 , 32'h0C226660 , 32'hFDB1D020 , 32'h05F44A50 , 32'h12E62E40 , 32'hEFDF4480 , 32'h0B628A40 , 32'hFD22C258 , 32'h2F006500 , 32'h0BF966A0 , 32'h012D5AC0 , 32'h26049FC0 , 32'h0ECC6C80 , 32'h1C4E8540 , 32'hE0B09AE0 , 32'h012C24DC , 32'hF63C5760 , 32'h071BC350 , 32'hF405E1C0} , 
{32'hF7D1ED90 , 32'h11BE5FA0 , 32'h02347440 , 32'hFD4A1F6C , 32'h0CEE21A0 , 32'h118A6B80 , 32'hF3DDF470 , 32'h253D4D00 , 32'h0056564B , 32'h02F30950 , 32'h14335C00 , 32'hE99A3BA0 , 32'h42990D80 , 32'hF460B020 , 32'hF6889B30 , 32'h0118FB6C , 32'hF7907F70 , 32'hE3D6E4E0 , 32'h17908640 , 32'hF77DC930 , 32'h1F02D140 , 32'hE7B4CB80 , 32'h0D82A840 , 32'h06403E80 , 32'hF73DBDC0 , 32'hF0130280 , 32'hFB7316C0 , 32'h0C247E50 , 32'hFEE5A194 , 32'hFBC357F0 , 32'hF57C8620 , 32'hFCFCCC90 , 32'hF9398CF8 , 32'hF58B5B20 , 32'hFB018778 , 32'hFCCAB098 , 32'h094F6D00} , 
{32'hFB8D2F40 , 32'hF8CF2510 , 32'hFE4EA528 , 32'h13559780 , 32'hFD0B1984 , 32'hFA415AE0 , 32'hFD658494 , 32'h1B642D40 , 32'h0091BD0A , 32'hCE456640 , 32'h155E91E0 , 32'hEE5F83C0 , 32'h2015F580 , 32'h04A5C9F0 , 32'hEF8D0CC0 , 32'hF5336220 , 32'h010F18B8 , 32'hF0D08BD0 , 32'h017A1648 , 32'hDD67BD80 , 32'h0BB13700 , 32'h098BFB80 , 32'h12ED99C0 , 32'hF70E8F10 , 32'hE9F2B980 , 32'hFBB74060 , 32'hFF89113C , 32'hF606D500 , 32'hEED6F840 , 32'h053A9EB0 , 32'h07B5BB38 , 32'hEDD5FF00 , 32'h068B9228 , 32'h004D4E6D , 32'h1022DEC0 , 32'h13EFD260 , 32'h0DC38C40} , 
{32'hFD7A43A0 , 32'hF5586760 , 32'hFA590AA8 , 32'h105458A0 , 32'hFF8A2CCB , 32'hFE3F5644 , 32'h0245C6A8 , 32'h0F1865D0 , 32'h0F991610 , 32'hEE02DC20 , 32'hFDE11C5C , 32'h14156C60 , 32'hFC8A1870 , 32'hFEC05480 , 32'h012877E0 , 32'hE85F98E0 , 32'h080FD440 , 32'hFD212E1C , 32'hEE717580 , 32'hEF8B6A60 , 32'h0AA18320 , 32'hFA069210 , 32'h03C55070 , 32'h0FA92650 , 32'hFA9F9850 , 32'h0079AFCF , 32'h0D44A2B0 , 32'h06C7F6B8 , 32'hFDCD3418 , 32'h0937FBE0 , 32'hFF023B26 , 32'hFE3D9A80 , 32'hF708E7E0 , 32'h092880B0 , 32'h0066B51A , 32'h107EDCA0 , 32'h01BE9250} , 
{32'hF9CEFFD8 , 32'hF1FC94E0 , 32'hFF747C1E , 32'h11522100 , 32'h16398320 , 32'h082C9F20 , 32'hFE9266A0 , 32'hF2A289A0 , 32'h06E027B0 , 32'hE9A3A080 , 32'h05D55518 , 32'h10C2EF00 , 32'hF3004940 , 32'hEE17F6E0 , 32'h0D667310 , 32'hE554E8C0 , 32'hF2F8B170 , 32'h0F838FE0 , 32'h18F82720 , 32'hF4E982A0 , 32'hE6FF4B80 , 32'h24169F40 , 32'h0ADF04A0 , 32'hD8CE34C0 , 32'hF41510B0 , 32'h06E72A90 , 32'h0EF29520 , 32'hFF67C6B4 , 32'h0B83E990 , 32'h06E64690 , 32'hFEC8DD88 , 32'h0CE04F60 , 32'h0EC49BA0 , 32'h0D2C0CE0 , 32'h038AEB84 , 32'h23BF7F40 , 32'h0BE75900} , 
{32'hFE3A83C8 , 32'hF64BE7E0 , 32'h05BA75B8 , 32'h051F0560 , 32'h061CE1A0 , 32'h0A887700 , 32'hF82BA190 , 32'h00468B2C , 32'h0656A0C0 , 32'hFF3CD673 , 32'hF842ADD8 , 32'hF2B79800 , 32'hFD5862AC , 32'h0124CE7C , 32'h0D05BBF0 , 32'h0A18CA10 , 32'h07F14C48 , 32'hF6027AC0 , 32'hFD5EEAC0 , 32'hF431F640 , 32'h119FA820 , 32'h00BCC025 , 32'h00CAEF7C , 32'h03AC2CD4 , 32'h0FCC4950 , 32'hF847DB88 , 32'hEF8A22A0 , 32'h0350D818 , 32'h03FFA530 , 32'hF6F6ABF0 , 32'h09CEA840 , 32'h0B7249D0 , 32'h0623A6E8 , 32'h109D4840 , 32'h028065C0 , 32'h01AFE954 , 32'h0A44CB80} , 
{32'hFFF18F65 , 32'h00157B17 , 32'h00108308 , 32'hFFF7B7D2 , 32'hFFF54FC5 , 32'hFFFC3634 , 32'h000619E6 , 32'hFFF101EF , 32'h0003D20F , 32'h000F05B2 , 32'hFFFFCD1D , 32'hFFF3AC02 , 32'hFFFFF21A , 32'h0008DA14 , 32'h000760E1 , 32'h00226CCB , 32'h00028DAA , 32'h00075BF3 , 32'h000C8D80 , 32'hFFFF00D1 , 32'hFFF6F8E9 , 32'h00173344 , 32'hFFF41657 , 32'h000C7338 , 32'hFFF0AB43 , 32'hFFFCD43A , 32'hFFF4ADE6 , 32'h00053DBE , 32'h001CFD99 , 32'h000CCF1E , 32'hFFF187B1 , 32'hFFF6ACEE , 32'hFFF51128 , 32'hFFF225F4 , 32'hFFFFBD90 , 32'h0008E903 , 32'h00059037} , 
{32'hFFF9125F , 32'hFFF3DC46 , 32'hFFFC453E , 32'h00009A22 , 32'h00089049 , 32'h000239E2 , 32'hFFFD6D64 , 32'hFFF1CB80 , 32'hFFF452E8 , 32'h0002CDAD , 32'h00048091 , 32'hFFFBEB68 , 32'h00007E9D , 32'h000A2F29 , 32'h000818B4 , 32'h00000802 , 32'hFFFE0CD1 , 32'h0002F7CC , 32'h000261C6 , 32'hFFFF5DD2 , 32'hFFFA099D , 32'h000D6C23 , 32'h00016F1E , 32'h0009EC81 , 32'hFFFB24DA , 32'hFFF9030B , 32'h00048556 , 32'hFFF5A246 , 32'hFFFCF3E9 , 32'h0002ECAA , 32'hFFF71445 , 32'hFFFDC8EF , 32'hFFFE4EFC , 32'hFFF59263 , 32'hFFFCD9FA , 32'hFFFA6580 , 32'h00022D0B} , 
{32'h0001A479 , 32'h0002A83E , 32'hFFFE29B0 , 32'h0002B548 , 32'h0001B716 , 32'h0007A7CE , 32'hFFFEF519 , 32'h0000A3FE , 32'h00075C85 , 32'h000827F2 , 32'hFFFD9B28 , 32'h00008AD4 , 32'hFFF86368 , 32'h0006C5B8 , 32'hFFFF8331 , 32'h0007EF09 , 32'hFFFBCAA6 , 32'h0004909D , 32'hFFFAEDED , 32'hFFFDE603 , 32'hFFF885DB , 32'hFFFF2510 , 32'hFFFD4327 , 32'h0003609B , 32'hFFFE211A , 32'h000625E6 , 32'h0008A1B0 , 32'hFFF91423 , 32'hFFFDD91E , 32'hFFFF2701 , 32'h0004FEF5 , 32'h00021E3D , 32'h0004555A , 32'hFFFA7143 , 32'hFFFF48DB , 32'h00005837 , 32'h00001F3C} , 
{32'h000024C4 , 32'hFFF562AF , 32'hFFF60607 , 32'h0003006B , 32'h0001C69E , 32'h00060C6B , 32'h0001E7FA , 32'h000072A7 , 32'hFFFB4DBF , 32'h0004B837 , 32'hFFFDCEB8 , 32'hFFFC7149 , 32'hFFFC3210 , 32'hFFFA5666 , 32'hFFFA7F76 , 32'h000630AF , 32'h0006803B , 32'hFFF3BA35 , 32'h000980F0 , 32'h00005E96 , 32'hFFFA01C6 , 32'hFFFDA571 , 32'hFFFA38C9 , 32'h000175E8 , 32'hFFFC1FD8 , 32'hFFFAFA8C , 32'hFFFF97D1 , 32'h00017A0A , 32'h00051C46 , 32'hFFF9FD55 , 32'hFFFACF37 , 32'hFFFA99C3 , 32'hFFFED39E , 32'h00018C5A , 32'hFFFE234E , 32'h0001D453 , 32'hFFF9427D} , 
{32'hFFFE0C80 , 32'h0002EC8D , 32'hFFF6577D , 32'hFFFFB2AF , 32'h00010708 , 32'h0006F370 , 32'h000468BA , 32'h00056E86 , 32'h001274F0 , 32'hFFFE2D27 , 32'hFFFDDBD4 , 32'h0001B73A , 32'h00087B70 , 32'h00019D8D , 32'h00068D30 , 32'h000957C6 , 32'hFFF92814 , 32'h0000F1EB , 32'hFFFFFF98 , 32'h00006935 , 32'hFFFDDC36 , 32'hFFFE1D7E , 32'h0002D7D2 , 32'hFFFB6FAA , 32'h0000C63E , 32'h00010C20 , 32'hFFFD2F76 , 32'h0004AA82 , 32'hFFFE6FE4 , 32'h000702EC , 32'h00034BD0 , 32'h00059381 , 32'hFFF89B50 , 32'h00066293 , 32'h00040639 , 32'hFFFFE4E1 , 32'hFFFE7CB3} , 
{32'h000406D6 , 32'hFFFC6EC1 , 32'hFFFDF10B , 32'h000D5AA2 , 32'h000A4F71 , 32'h0000EEA1 , 32'h00018077 , 32'hFFF8E272 , 32'h00014989 , 32'hFFFEF271 , 32'h000B8475 , 32'hFFFF8184 , 32'hFFFDC5F6 , 32'hFFF89CD6 , 32'h00052E4A , 32'hFFFFD169 , 32'hFFF96F19 , 32'hFFFA14E6 , 32'h00052112 , 32'h00028603 , 32'h00091AE1 , 32'h00068861 , 32'h0005D182 , 32'h000AFB7C , 32'hFFFEF181 , 32'h000135CB , 32'hFFFAC675 , 32'h0002EBC4 , 32'h0005D4D9 , 32'h000107B3 , 32'h00055C16 , 32'hFFF75067 , 32'hFFFB3D1D , 32'hFFF93CCD , 32'hFFF7B397 , 32'h00087DE3 , 32'hFFFF5DD1} , 
{32'h00016DFE , 32'h00017C64 , 32'h0002DFF7 , 32'h0005004C , 32'h00007AC4 , 32'h0008DEE5 , 32'h00045CFE , 32'h00034D67 , 32'hFFF797EE , 32'h00020200 , 32'h000573F7 , 32'hFFFF8156 , 32'h0002D0A4 , 32'hFFFB7C5C , 32'hFFFF9E34 , 32'hFFFF6F51 , 32'hFFFA5935 , 32'hFFFB96AF , 32'h000320FF , 32'h00053E20 , 32'hFFFCCBB8 , 32'hFFFC7E44 , 32'h000B0C98 , 32'hFFFCD805 , 32'h0003270D , 32'hFFFC4697 , 32'hFFF40E64 , 32'h0005B53E , 32'hFFFFDA66 , 32'hFFF9381D , 32'h0002DF4C , 32'hFFFB684E , 32'hFFF666E1 , 32'hFFFCC762 , 32'hFFF5406C , 32'hFFFBF3C3 , 32'hFFFD4498} , 
{32'h02B19B58 , 32'h0016DD07 , 32'h06344520 , 32'hFFAD113B , 32'h087E0A30 , 32'h01C4F708 , 32'h038CFFA0 , 32'h08B5A530 , 32'h0527AB90 , 32'hFC3699F8 , 32'h074D9DC8 , 32'h028E935C , 32'h06DF3C88 , 32'hFC70C14C , 32'hFB558888 , 32'hF75FC620 , 32'hF9892BC8 , 32'hF7904980 , 32'h05153948 , 32'hFFD61514 , 32'hFE630230 , 32'hFA730B30 , 32'h059F3668 , 32'hFCE725E8 , 32'hF865E7C0 , 32'hF45EF490 , 32'hFF69B485 , 32'hFADFAFE8 , 32'h0029095B , 32'h043D2388 , 32'h08B8BD70 , 32'h067BA2B0 , 32'h0172F0F4 , 32'h0BD28CF0 , 32'hFD003DC0 , 32'h023F7FA4 , 32'hF62E3940} , 
{32'hE2A7FA80 , 32'hEC708920 , 32'h306296C0 , 32'hFB422A48 , 32'hF100C7B0 , 32'h047787E0 , 32'h18A8B3E0 , 32'h0EC8C8F0 , 32'h0E2BC740 , 32'hFEC9BF1C , 32'h29444140 , 32'hFF11597D , 32'hEA4BE620 , 32'hF0BE9DF0 , 32'hE8E997A0 , 32'hF56C6660 , 32'hDD89B380 , 32'hDD3F3D00 , 32'hF6700990 , 32'h02FC1828 , 32'hE6758AC0 , 32'h0EEA9AF0 , 32'h0B3A30E0 , 32'h116E7FE0 , 32'h106C5940 , 32'h0CEBB090 , 32'hE1D36020 , 32'hEF7D77E0 , 32'hE6DA0F80 , 32'h18AC4DC0 , 32'h06AB9300 , 32'hF452DA00 , 32'h0C3873C0 , 32'hDA0C9A80 , 32'hF19E8370 , 32'hF9EC41E8 , 32'h05154F70} , 
{32'hE8FD18C0 , 32'hE35BF360 , 32'h29171B40 , 32'hFA9A94F0 , 32'hFCAE7C58 , 32'h1785FF40 , 32'h15C85780 , 32'h139C46C0 , 32'hF3B8D390 , 32'hFB856250 , 32'h11384300 , 32'h03B51308 , 32'hF9034DA0 , 32'h0B0A4790 , 32'hE5A081E0 , 32'h09AF9EC0 , 32'hF093B040 , 32'hEB5AA860 , 32'hF4EF2B20 , 32'h08F16270 , 32'h01835328 , 32'h0D5BB4C0 , 32'hFCEFC508 , 32'hFBB177F8 , 32'h0AC356C0 , 32'h0E64E7E0 , 32'h0B16B2E0 , 32'hF8FF4828 , 32'h0963A580 , 32'h0BBB6700 , 32'h05737100 , 32'h0F093570 , 32'h0E46CF50 , 32'hFD6C0DE4 , 32'hFDECD2A8 , 32'hFF4CEE40 , 32'h070C3FC8} , 
{32'hE8AA0CE0 , 32'hE9E242A0 , 32'h50A2AD00 , 32'hF4DF4210 , 32'h0105F6A0 , 32'h322FD840 , 32'h2C8A4740 , 32'h1CA54B80 , 32'hEF72CC60 , 32'hFB610D70 , 32'h1E99C900 , 32'h10686A40 , 32'hE6B57340 , 32'h0403E5B8 , 32'hE4EBFEE0 , 32'hEB3C9A00 , 32'hE54739A0 , 32'hDB602880 , 32'hEF4C0740 , 32'hF35FB8F0 , 32'h023869A8 , 32'h0D95C1F0 , 32'h04C76050 , 32'hF7672B40 , 32'h0C832EA0 , 32'h140EA660 , 32'h1BE708E0 , 32'hF2208F50 , 32'hEC9E9C00 , 32'h078BC880 , 32'hF67B0C60 , 32'h0FA09CD0 , 32'h1DAF9EE0 , 32'hD8755180 , 32'hEFC5E060 , 32'hFDE4D19C , 32'h18641160} , 
{32'hD43A1200 , 32'hC92860C0 , 32'h76EF6480 , 32'h10F3EE00 , 32'hF1521110 , 32'h36EB1340 , 32'h3DE7D2C0 , 32'h293C0040 , 32'hE620DD40 , 32'h0EC17B80 , 32'h12929660 , 32'h07395A50 , 32'hEAFAF2C0 , 32'h0EA8A7E0 , 32'hE4A8D1A0 , 32'hDB1ACB00 , 32'hECCFAD00 , 32'hE13B4A80 , 32'hEF6EEFA0 , 32'h0A5717E0 , 32'h0BDF5A60 , 32'hFEE81D38 , 32'hFA1D7838 , 32'hF52A4490 , 32'hFCCB686C , 32'h0232EDB0 , 32'h214FB600 , 32'hE55EF3E0 , 32'h17A2B860 , 32'h09C642E0 , 32'hFF4F549D , 32'h13DE76A0 , 32'h1725B440 , 32'hF7A64B80 , 32'h14787B80 , 32'hEB7DE820 , 32'hF3E82440} , 
{32'hB7967E80 , 32'hC498D980 , 32'h7FFFFFFF , 32'hFB2F6DD8 , 32'hE0A10600 , 32'h35D8B2C0 , 32'h283F8380 , 32'h25455EC0 , 32'hEA9CC780 , 32'h0F8CA370 , 32'h06FEEC60 , 32'hF219CD60 , 32'hE4E94360 , 32'h19AEFF00 , 32'hE3D0B300 , 32'hFFD07C9F , 32'hEA5F4DE0 , 32'h02B9B4CC , 32'hE863C960 , 32'h12230E20 , 32'h0F92E4A0 , 32'h0DB35530 , 32'h08C1EA00 , 32'hFAE07B00 , 32'h09A29BE0 , 32'h12233580 , 32'h2473F600 , 32'h07219310 , 32'h0FAC7310 , 32'h179CEBA0 , 32'hEDDF5400 , 32'h174C95C0 , 32'h152AA5C0 , 32'hED57DAC0 , 32'hE9C79E20 , 32'h00866FE1 , 32'h0DCFAAD0} , 
{32'hD4A97A40 , 32'hD92345C0 , 32'h554BC000 , 32'hFB91F438 , 32'hD1B70FC0 , 32'h32478C40 , 32'hF9744770 , 32'h1894DA80 , 32'hE1BDD360 , 32'h046213F8 , 32'h204F87C0 , 32'hE6907C40 , 32'hD9B0FC00 , 32'h12610EA0 , 32'hFC5886B0 , 32'hE278D6E0 , 32'hDDE9DD80 , 32'hFDF2EBA8 , 32'hDF9EB3C0 , 32'h0B1A4940 , 32'hFFDDF585 , 32'hE39D6960 , 32'h16B90D20 , 32'hF9464918 , 32'h0958D0E0 , 32'h1106B620 , 32'h1E371EC0 , 32'hDF9CF400 , 32'h0E1375A0 , 32'hFAE9E840 , 32'hFC52CA3C , 32'h2C288440 , 32'h0337BB88 , 32'hFD07C558 , 32'hFD1B366C , 32'hFAF3EEF8 , 32'h0CEF4E70} , 
{32'hF58E65C0 , 32'hF63FF160 , 32'h0017A4AF , 32'h1107B940 , 32'hCA79C600 , 32'h03A004F4 , 32'h0FF83850 , 32'h0626AC98 , 32'h0DC1ED10 , 32'hF1126930 , 32'h2A0FB640 , 32'hE46B4600 , 32'hFF6545D7 , 32'hF32CBD90 , 32'h08079E80 , 32'hF4794880 , 32'h11BFDA00 , 32'h1B06BEE0 , 32'h0978DE50 , 32'hFBB4A478 , 32'h038A4FC8 , 32'h028191DC , 32'h0D246470 , 32'h0C01D0E0 , 32'hF14597D0 , 32'hEEB66B00 , 32'h13545C40 , 32'hF38C9870 , 32'hEF4588C0 , 32'hE8A15460 , 32'h1B4817A0 , 32'hEE4CBAC0 , 32'h0C112CB0 , 32'h050FB9C8 , 32'h1A4FBF40 , 32'hFCA66D14 , 32'hFBB63AB0} , 
{32'hF376E410 , 32'hAD510E80 , 32'hD61095C0 , 32'h109074C0 , 32'h9DAF2080 , 32'hEBF154A0 , 32'h05B24270 , 32'hE998ADC0 , 32'hFD82C11C , 32'hF9C09258 , 32'h41625900 , 32'hCEE55940 , 32'h0C4D7100 , 32'hEE3D09C0 , 32'hEB519BA0 , 32'hF8ECCF38 , 32'hFEFEC1B4 , 32'h0ED26270 , 32'h121E5AE0 , 32'hF08292F0 , 32'hEC40CFE0 , 32'hFC94FDBC , 32'h07C8A0D8 , 32'hF0A3DA30 , 32'hF66BF390 , 32'hF4D0C570 , 32'hF73B6510 , 32'h002EB023 , 32'hDDE55B40 , 32'h14DB9A00 , 32'h0F6AB9C0 , 32'h2EF70F40 , 32'hFE112784 , 32'h1ED382E0 , 32'h11AF1180 , 32'h03EFCAB8 , 32'h24AEE400} , 
{32'hE1A8DE40 , 32'hEC0D25A0 , 32'hCF420800 , 32'h14CC6D20 , 32'h7FFFFFFF , 32'hE817D440 , 32'hF37CF1C0 , 32'hE1307BE0 , 32'h0C405D10 , 32'h090A8CC0 , 32'h1201D860 , 32'h2E7A3C40 , 32'hE58D9140 , 32'h07D80798 , 32'h06D87258 , 32'hF4BD2730 , 32'h07FAEAD8 , 32'hEEA8A460 , 32'h02A48638 , 32'h1D914440 , 32'h14C2CCC0 , 32'hB8549380 , 32'h01941D60 , 32'h1CC063E0 , 32'h1525B140 , 32'h1022D020 , 32'h0BEE05E0 , 32'h070F4610 , 32'hEFDE2D60 , 32'h1386DBC0 , 32'h1F6E5900 , 32'h2C669A00 , 32'h179C4CA0 , 32'h30AA02C0 , 32'hEDED61A0 , 32'hD4452D80 , 32'h220AA300} , 
{32'hEB8E15E0 , 32'h083A8400 , 32'hFA0FAF98 , 32'h1470DAE0 , 32'hD8BF76C0 , 32'hFF8BC65C , 32'hECFBC800 , 32'h04CFD5C0 , 32'hF77266B0 , 32'h281FD7C0 , 32'h05C254F0 , 32'h2147FDC0 , 32'hEBD5E940 , 32'h224326C0 , 32'h1B341B40 , 32'h111C0680 , 32'h248A9280 , 32'hEF13DC20 , 32'hFC1CBAF4 , 32'h2A021B40 , 32'hE4683740 , 32'hE99F51C0 , 32'h10A25FC0 , 32'h08048360 , 32'hF9129F60 , 32'h047D5FC0 , 32'h033B13D0 , 32'h12BCB280 , 32'h07F702F8 , 32'hE81C7200 , 32'hF69EF3A0 , 32'h152D73C0 , 32'hF3A701C0 , 32'h01399710 , 32'hFBBE7000 , 32'hEDB91A40 , 32'hE813E020} , 
{32'hF2CCF690 , 32'hFBB0CCC0 , 32'h0736F730 , 32'h14E5AA60 , 32'hF65979E0 , 32'h0748FD48 , 32'hF281DC00 , 32'hE6A0E1C0 , 32'hF4F29E80 , 32'h055FEF10 , 32'hE507E680 , 32'h10E005E0 , 32'hF2098AB0 , 32'h14487440 , 32'h076D1920 , 32'h09B1EFE0 , 32'h04EFBE00 , 32'hF3AC8920 , 32'hF9582460 , 32'h13FD5180 , 32'hE4860940 , 32'h06490D80 , 32'hF85A90C8 , 32'hFD64E8BC , 32'hFF9C44F5 , 32'hFA3EBB08 , 32'h0145EED0 , 32'hF3154A80 , 32'hEA2F3860 , 32'h00FA4065 , 32'hF6F39F10 , 32'h139D2A20 , 32'hEA5850A0 , 32'h13ECCE20 , 32'h07A5BBE0 , 32'hF35067B0 , 32'hFD3E3FB4} , 
{32'hEBFE0D20 , 32'hF5B15040 , 32'h0AE5AD80 , 32'h17B45F00 , 32'hFD2304CC , 32'h02B0C62C , 32'hE73715E0 , 32'hEE239820 , 32'hFED13840 , 32'h10C83540 , 32'hE630F7A0 , 32'hFF50C284 , 32'hFE42E6B8 , 32'h085343D0 , 32'h0201B708 , 32'h245C3680 , 32'h26C31AC0 , 32'h00D0C1C3 , 32'h08E91A50 , 32'h0AFF9C30 , 32'h289CB980 , 32'hFFD10C4A , 32'hFF21BABD , 32'hF7C31CC0 , 32'h280C7880 , 32'h01C3111C , 32'hE7F41E40 , 32'hFC408504 , 32'hF03A0CC0 , 32'h05577500 , 32'h1257B080 , 32'hFADC74F8 , 32'h00786881 , 32'h162D5A20 , 32'h222BF8C0 , 32'hFF14ECF1 , 32'hF90CF640} , 
{32'hF6A1A4B0 , 32'hE5230340 , 32'h08065C40 , 32'h289AFCC0 , 32'h0C50AEB0 , 32'h2B39C700 , 32'hDAF76B80 , 32'hE6C522A0 , 32'hF8881FE8 , 32'h0590BAE0 , 32'h0F896F10 , 32'hF266EEC0 , 32'h0E4C6D20 , 32'hF84C80E0 , 32'h28F9C840 , 32'hE0BC76E0 , 32'h194264A0 , 32'hE573F5A0 , 32'h06AA0CD0 , 32'h0848E760 , 32'h043456F0 , 32'hFFFBDDC2 , 32'hFB68C988 , 32'hED1D9700 , 32'h080779F0 , 32'hDFD45B80 , 32'hE8030D60 , 32'hE6C1B7C0 , 32'h05E10CE8 , 32'hF5A93AC0 , 32'hF4B7F820 , 32'h05155740 , 32'hE7B74240 , 32'hE58E1620 , 32'hE726F160 , 32'h0CE94D10 , 32'h0BE3D470} , 
{32'hF588B090 , 32'hF0A92D80 , 32'h09F9E230 , 32'h0DFB0A70 , 32'h1C7744E0 , 32'h1ACB4A00 , 32'hD9A4B940 , 32'hF6F64D30 , 32'h03A88B24 , 32'h01156980 , 32'h2AA9B700 , 32'h0AA64630 , 32'h35BD7700 , 32'hECDE36E0 , 32'hFE5F8D78 , 32'hF6C5E2E0 , 32'h08215270 , 32'hFE0405BC , 32'h214C2A40 , 32'hF5B12330 , 32'h157139A0 , 32'h088918C0 , 32'hF2CD4C60 , 32'hF199E670 , 32'hFFAD6688 , 32'hEDE69C00 , 32'h0E185D90 , 32'hFA554AA0 , 32'hF8F525A8 , 32'h075E7FA8 , 32'hE2716120 , 32'hF881CAB8 , 32'h0826E260 , 32'h08FCA320 , 32'hFC467E28 , 32'h05507C40 , 32'hFC3C918C} , 
{32'h03DD08A0 , 32'hE776C4A0 , 32'hF6448F80 , 32'h1413CE60 , 32'h09805710 , 32'h236D1800 , 32'hDFC26080 , 32'h18ACFF60 , 32'hFB7E4FD0 , 32'hFBF10ED0 , 32'h41F5C180 , 32'hD53D7740 , 32'h30290040 , 32'hFAA1FCC8 , 32'h0310D12C , 32'h01176FD4 , 32'h246AB580 , 32'hD76CD080 , 32'h24050880 , 32'hE0542BA0 , 32'hD97E5540 , 32'hF62D4660 , 32'hEC4627C0 , 32'h1521DD00 , 32'hE3B248C0 , 32'h1519B380 , 32'h034FC598 , 32'h162FD000 , 32'hFC847C64 , 32'hCF144F00 , 32'hE8775FE0 , 32'hE7E68240 , 32'h1EEEFC80 , 32'hF6ED8190 , 32'hEE2419C0 , 32'h045E5558 , 32'h09A7C540} , 
{32'hF8B2DF18 , 32'h02501BFC , 32'hFD1895C8 , 32'h16EC5F80 , 32'h15025900 , 32'h2AE80E00 , 32'hF5AFE430 , 32'h16CC4E60 , 32'h1361F340 , 32'hD6BD2BC0 , 32'hF8B3A030 , 32'hD0822500 , 32'h30562BC0 , 32'h083F4090 , 32'h11EFD720 , 32'hF0DB8770 , 32'hEA583F80 , 32'hE97542E0 , 32'h29727600 , 32'hF56CF950 , 32'h1443BD20 , 32'h4B955880 , 32'hFE87A630 , 32'h0F99EEE0 , 32'hF9A439E8 , 32'h15E1CA80 , 32'h03FC8CBC , 32'hB4CF1B80 , 32'hEE284100 , 32'hFAB3E130 , 32'h059D7CA8 , 32'h1EB97540 , 32'hEBD66AE0 , 32'h06D862B0 , 32'h045F6138 , 32'hFBC16778 , 32'hE964D460} , 
{32'h020E5F04 , 32'hFFFBEB99 , 32'h0172CEB0 , 32'h08DFB1A0 , 32'h017E5FEC , 32'h0A15A800 , 32'hFB8EF318 , 32'h080625F0 , 32'h08FADEA0 , 32'hF6BE2F20 , 32'hFC5C10A8 , 32'hEED84D80 , 32'h12FA4F80 , 32'hFC6B5288 , 32'h03D5C848 , 32'hFD77D768 , 32'hFE76651C , 32'hF54CD290 , 32'h013E5190 , 32'hFD2D0E98 , 32'h149CDE60 , 32'h05442888 , 32'h06825B48 , 32'hFEA26258 , 32'hF9EE2D68 , 32'h025E42C4 , 32'h0410C840 , 32'hD7513580 , 32'hEDE8DEE0 , 32'hFB57C5A8 , 32'hF3AEB340 , 32'h18C05900 , 32'hFDB054E8 , 32'h066EED70 , 32'h0213ACB0 , 32'hF3D6F800 , 32'hF30F9BF0} , 
{32'h05857E90 , 32'hFAA55030 , 32'hFC091DE0 , 32'hFE2EE720 , 32'h09DA8970 , 32'h118F8C80 , 32'h067393B8 , 32'hFE340FD4 , 32'h03BAAFF4 , 32'h05BAD1F8 , 32'hFAB94028 , 32'h0728EF60 , 32'h1B6882E0 , 32'hD6193DC0 , 32'hF251F150 , 32'hF108D9C0 , 32'h1520ED20 , 32'hF77B6B20 , 32'hEA21A9E0 , 32'h15535EA0 , 32'hF90674A8 , 32'h05D978E8 , 32'h15C8EBE0 , 32'hF96A4608 , 32'h0B3D5950 , 32'h004CFCF0 , 32'h106A4840 , 32'h06C79AE8 , 32'hFC4A370C , 32'h03E66E50 , 32'h031EE3C8 , 32'h128AF560 , 32'h06686EB8 , 32'h083DB940 , 32'h017F6554 , 32'h035284D0 , 32'hFD4F92A0} , 
{32'hF15F0580 , 32'h056AD4F8 , 32'h04750EC0 , 32'h07B4F4A0 , 32'h10EA5100 , 32'hF58D0B50 , 32'h0F401D20 , 32'hFBEE0E68 , 32'h19382D00 , 32'hF433B3B0 , 32'hF0E443E0 , 32'h123DB640 , 32'hFEC6AB9C , 32'hFB9AD120 , 32'h0F667EB0 , 32'hFBAF9A00 , 32'hFEB4210C , 32'h076DA1A8 , 32'h0903B420 , 32'hF2159F00 , 32'hEE422560 , 32'h056EAA98 , 32'hFAE11EC0 , 32'hED6BB1A0 , 32'hF6EA86E0 , 32'h04F8B1D8 , 32'h159D3FA0 , 32'h03BFF11C , 32'h01C035AC , 32'h06B02938 , 32'hF8EA4D80 , 32'h0F679A90 , 32'h1B6B07C0 , 32'h0AC33BE0 , 32'h09AA1AC0 , 32'h118746E0 , 32'h05854E98} , 
{32'hF6AD2570 , 32'hEBD80280 , 32'h003E6DDD , 32'h165444E0 , 32'h0AF4A190 , 32'hFD7EEFFC , 32'hF8F7A378 , 32'hEF999FC0 , 32'h05B1AAD0 , 32'hF7A17610 , 32'h0264CBD8 , 32'h15197AA0 , 32'hE8C468E0 , 32'hF639E8F0 , 32'h0CA74460 , 32'hF1B8A860 , 32'hF96DD1C0 , 32'h23DF3D00 , 32'h17F80720 , 32'h00D27137 , 32'hE1E20FA0 , 32'h1506F0E0 , 32'h10528D60 , 32'hDE056C40 , 32'hF1179260 , 32'h123C4760 , 32'hFF8CD9E9 , 32'h00F6ECB8 , 32'h164633C0 , 32'h0C0EDF50 , 32'h04D4A540 , 32'h06C779D8 , 32'h1A96EFA0 , 32'h0C5D80D0 , 32'hFF7A4130 , 32'h1267E660 , 32'h010E1890} , 
{32'hFFE66E67 , 32'h0011B100 , 32'h00041D06 , 32'h0004979B , 32'h0001289E , 32'hFFF06B03 , 32'h000A81B0 , 32'hFFE88219 , 32'h0012CD2E , 32'h00050C71 , 32'hFFF4F5B5 , 32'hFFFA804D , 32'h00042F7D , 32'h000604A7 , 32'h0004D92F , 32'h0024FD63 , 32'h000CFE1E , 32'hFFFF9E71 , 32'h00101216 , 32'hFFF355A6 , 32'hFFF569A8 , 32'h001A8375 , 32'hFFE88D77 , 32'h0012A488 , 32'hFFF9CB86 , 32'h00071D6E , 32'h00014E36 , 32'hFFFCCD19 , 32'h00113887 , 32'h0007DC8F , 32'hFFF2199A , 32'hFFFFEDD7 , 32'h0004D45D , 32'hFFF25FB1 , 32'hFFF6EB38 , 32'h000C135B , 32'h00012D50} , 
{32'h00076717 , 32'h000310BF , 32'hFFFE64E9 , 32'h00034B97 , 32'h00063686 , 32'h00000911 , 32'hFFF3CAF1 , 32'hFFFE3E8A , 32'h000752BB , 32'hFFFFFE8B , 32'h0000DE08 , 32'h0005A29C , 32'hFFF80604 , 32'hFFFF3244 , 32'hFFFE0F69 , 32'h0004F517 , 32'h00028F51 , 32'hFFF9CB3B , 32'hFFF35FE7 , 32'hFFFCAFCC , 32'h0003DD92 , 32'hFFFC937D , 32'h00014D7D , 32'hFFFAEE03 , 32'h0000312C , 32'hFFFCA1FF , 32'hFFF9709B , 32'hFFFA6B75 , 32'hFFFBF159 , 32'h00080A99 , 32'hFFFD4266 , 32'hFFFFED96 , 32'hFFFF7242 , 32'hFFFAAD0D , 32'hFFFFC302 , 32'h00082C9A , 32'hFFFE614A} , 
{32'h0008A47C , 32'h0000BABC , 32'h00074280 , 32'h00086637 , 32'hFFFE5592 , 32'hFFFBA524 , 32'h0002AF67 , 32'h00040691 , 32'h000B74B1 , 32'h00027299 , 32'hFFFFCF05 , 32'h0007CFF0 , 32'hFFFFDCA0 , 32'hFFF7ED06 , 32'hFFFF4FDD , 32'h00090E5E , 32'h0007F41B , 32'h00010A55 , 32'hFFF8E4E0 , 32'h0001E307 , 32'hFFFFCBD9 , 32'hFFFD78C8 , 32'h0000EF22 , 32'hFFF7C1F7 , 32'hFFFBF08F , 32'h0002332A , 32'hFFFE2FAA , 32'h000340C9 , 32'h0006E88B , 32'h0001778B , 32'h0001523D , 32'hFFFC6CCB , 32'hFFFDD537 , 32'h000250B8 , 32'hFFFBBF60 , 32'hFFFBDB9C , 32'hFFFCB821} , 
{32'hFFFF624C , 32'hFFFD5F6D , 32'h0007C92E , 32'h0002B942 , 32'h00011661 , 32'h00025B29 , 32'h00022B56 , 32'hFFFB4459 , 32'hFFFC6928 , 32'h000A752E , 32'hFFF81CD4 , 32'h0006C593 , 32'h000513B6 , 32'h00063E39 , 32'hFFFE06E6 , 32'hFFFF328C , 32'hFFF98722 , 32'hFFFECF53 , 32'h0001CEE5 , 32'hFFFD39F8 , 32'hFFF826F8 , 32'h00026B2A , 32'h0002F8D6 , 32'hFFFDE669 , 32'h0001C1F3 , 32'h0002C5F5 , 32'hFFF8EA09 , 32'h00048C14 , 32'hFFF2E210 , 32'hFFFE8F6F , 32'hFFFC0EDE , 32'h0003BA02 , 32'hFFFC80B6 , 32'hFFFF0AAA , 32'h0008250B , 32'h0006FCDF , 32'hFFFF1178} , 
{32'hFFFAF245 , 32'hFFFA6E5A , 32'h00063307 , 32'hFFF608BC , 32'hFFFBCAB8 , 32'h0005C4C0 , 32'hFFF2D8FF , 32'h00019A0B , 32'h000194AB , 32'hFFFDA433 , 32'hFFFF1EC9 , 32'h00068E63 , 32'hFFF93370 , 32'hFFFEDF8C , 32'h0007C2BE , 32'hFFFCA5CC , 32'h0000B8E9 , 32'hFFFE75E1 , 32'hFFF9DD86 , 32'hFFFC1309 , 32'h00005CB8 , 32'hFFFB9AEF , 32'hFFF250EB , 32'h0001CFBA , 32'hFFF9A948 , 32'hFFFDEBB0 , 32'hFFF7DAEE , 32'hFFFD7B73 , 32'hFFFCDA7D , 32'h00047A3B , 32'h0003009E , 32'hFFFCD751 , 32'hFFFEE4FB , 32'hFFF8C3DD , 32'hFFFD6524 , 32'hFFF97E2C , 32'hFFFEAC5E} , 
{32'h000E153B , 32'hFFFBFF30 , 32'hFFFA86A9 , 32'h000C6A96 , 32'hFFF89FCA , 32'h0010A5A1 , 32'h0002FDFB , 32'hFFF2E0FA , 32'hFFF890BE , 32'hFFFD960A , 32'h00071FF6 , 32'hFFFC0C17 , 32'hFFF88BDD , 32'h0003530C , 32'hFFF0671A , 32'h000132FB , 32'hFFFE5522 , 32'hFFFADA6F , 32'hFFFA22CA , 32'h00057DC5 , 32'h00002777 , 32'h00081D9F , 32'h00023B5A , 32'hFFF79CEF , 32'hFFF9B7C9 , 32'h00034386 , 32'hFFF0137A , 32'h00037965 , 32'hFFFDE9E2 , 32'h00004FE6 , 32'h00030571 , 32'h000530BF , 32'hFFEB67F5 , 32'h0005098F , 32'hFFFE3F2D , 32'hFFF95DBC , 32'h0000FA57} , 
{32'h0074BA92 , 32'hFFB93F10 , 32'hFFC45C16 , 32'hFFEB673E , 32'hFFB6871D , 32'h008CF723 , 32'hFFBC73EC , 32'h00295271 , 32'hFF660C6B , 32'h0016888A , 32'h0091E2C8 , 32'hFFCEAA71 , 32'hFFA19438 , 32'hFFEC403A , 32'hFFB6C388 , 32'hFF7EC55D , 32'hFFE7C7DB , 32'hFFCF6494 , 32'hFFFCD0BA , 32'h005F5036 , 32'h00268F30 , 32'h0002B98B , 32'h008A1CFE , 32'h00028C20 , 32'h0002A212 , 32'h0004CACF , 32'hFF71DBF2 , 32'h00079558 , 32'h002B4FDB , 32'hFFDA2CE0 , 32'h005009D4 , 32'hFFE1F2B0 , 32'hFF768A84 , 32'h001CB17F , 32'hFFACDE13 , 32'h00068AE7 , 32'h00276D0A} , 
{32'hE4801F20 , 32'hE6A3BF80 , 32'h19EEE240 , 32'h0188DA54 , 32'h0A7C2BE0 , 32'hFDA9E298 , 32'h049F4978 , 32'h0897EB00 , 32'hF64A6C30 , 32'hFAB4AD10 , 32'h0CBE9EA0 , 32'hE9FD7740 , 32'hF1E13420 , 32'h0EEF7E50 , 32'hFA29DB58 , 32'h1233DB60 , 32'hF6071680 , 32'hFBD235A0 , 32'hEABAAD60 , 32'h177A5320 , 32'h15A115C0 , 32'h063CD738 , 32'h02295568 , 32'h004B2863 , 32'hFD50B01C , 32'h093F9460 , 32'h134C06E0 , 32'h06A68C00 , 32'h1908BB80 , 32'h055D07D8 , 32'hF51D0420 , 32'h0C41C420 , 32'h04724E68 , 32'h0C2B23D0 , 32'hFEAAE1FC , 32'h056889D8 , 32'h0A7E0290} , 
{32'hD65C53C0 , 32'hC6A4ED40 , 32'h1A2220C0 , 32'hF91D0C18 , 32'h3F19B500 , 32'h0438AE68 , 32'h011E3238 , 32'h0EC1C490 , 32'hECDA2FA0 , 32'h08E1E2D0 , 32'hF070E5B0 , 32'hDC791D00 , 32'hFB255060 , 32'h1EAA2BA0 , 32'hF1D612A0 , 32'h1601D060 , 32'hF8F262A0 , 32'hE3FBF180 , 32'hEB273A80 , 32'h095A9CB0 , 32'h243EA080 , 32'h0CF10CC0 , 32'h049AAB98 , 32'hFF6504E1 , 32'hEEAE0F20 , 32'h03EA4598 , 32'hFCB536C8 , 32'h0FA24100 , 32'h1620FFC0 , 32'h08F07720 , 32'hFC151D6C , 32'h193B91E0 , 32'hFC547128 , 32'h1C3916E0 , 32'hFCF8AA74 , 32'h060A9980 , 32'h14C650A0} , 
{32'hB6F4AA00 , 32'hAB58F000 , 32'h15149060 , 32'hD30E1700 , 32'h6D744000 , 32'h26D1D240 , 32'h15A6C680 , 32'h22F2B200 , 32'hF6C06D10 , 32'h0C0BB390 , 32'hE3489AE0 , 32'hEFD8C0E0 , 32'hF1586770 , 32'h21531AC0 , 32'hFFF2C445 , 32'h333A6280 , 32'h196F6FE0 , 32'hF7C201E0 , 32'hF0AD5600 , 32'h01C9D07C , 32'h2E845B80 , 32'h12BA1C00 , 32'h1EF58AC0 , 32'h0D600500 , 32'hE7485BC0 , 32'hFF147188 , 32'hE0F58B60 , 32'h1116F3C0 , 32'h0179251C , 32'hDECA6C80 , 32'h1CCCEBA0 , 32'h0DD5DE30 , 32'hF3413A40 , 32'h2B56D140 , 32'hFED92C1C , 32'h106B4AC0 , 32'h07198338} , 
{32'hCCF9BC40 , 32'hB5A17A00 , 32'h1D77E280 , 32'hF4A29740 , 32'h62F45800 , 32'h20584D00 , 32'h3600E880 , 32'h0ADFE6E0 , 32'hD7C328C0 , 32'hF4448640 , 32'hF0831DE0 , 32'h083DD5E0 , 32'hD09E4740 , 32'h231A29C0 , 32'hFB50EBA0 , 32'hF7AC0BC0 , 32'hFB318578 , 32'hEA1376A0 , 32'h13A569C0 , 32'h171D9580 , 32'h14B55640 , 32'h009BD3BC , 32'h0C238290 , 32'h0A761BC0 , 32'hF4F6E3A0 , 32'h080DA130 , 32'h14E9B100 , 32'h14966B60 , 32'h24C79500 , 32'h12138620 , 32'hFE8717C0 , 32'h0567FE58 , 32'h01A50FE4 , 32'h04E6AF08 , 32'h0FA71420 , 32'hFC44D220 , 32'h075D9690} , 
{32'hD455A0C0 , 32'hBC94A580 , 32'h227651C0 , 32'hF44320A0 , 32'h41759200 , 32'h27DEEEC0 , 32'h2D21DC40 , 32'h1F2B21E0 , 32'hE05F1500 , 32'h05380ED8 , 32'hF1E68AB0 , 32'h04D6AD58 , 32'hE94C6B40 , 32'h2E5C68C0 , 32'h04B9A550 , 32'h12A10080 , 32'hFFA75D30 , 32'hD0E3FAC0 , 32'hF3881DC0 , 32'h215BC300 , 32'h093F2230 , 32'hF964F960 , 32'hF6BB4130 , 32'hF74B30F0 , 32'hE5464AA0 , 32'h117144C0 , 32'h216C7940 , 32'hFE5DBA70 , 32'h0D42E250 , 32'h04518D10 , 32'h1391C1E0 , 32'h00B1EEE8 , 32'hFE4C5248 , 32'h0AE1E5A0 , 32'hFF4194EB , 32'hF81FBD98 , 32'hF7B805D0} , 
{32'hF13B5F50 , 32'hD94FA580 , 32'h142CB7C0 , 32'hF4BA19D0 , 32'h0788BDE8 , 32'h310E6D00 , 32'h195207A0 , 32'h15DC7040 , 32'hD6DE87C0 , 32'h11A66C80 , 32'hE280E600 , 32'hF6783500 , 32'h083B7F60 , 32'h176ED740 , 32'h1FC85DE0 , 32'hDB7DB140 , 32'h081A5870 , 32'hFF047951 , 32'h0656D598 , 32'hF7E83710 , 32'hF42FB980 , 32'hE8C1D440 , 32'hF077A000 , 32'hF4A6BA40 , 32'h0BA3DB10 , 32'h19DCB4A0 , 32'h1FD93960 , 32'hF4A771B0 , 32'h085E4840 , 32'hF2279980 , 32'h012C9D9C , 32'hFC7DDD40 , 32'hF531A990 , 32'hF1AAFBD0 , 32'h161995E0 , 32'hF90F90C0 , 32'hF34894B0} , 
{32'hE6248C60 , 32'hC6A48B00 , 32'h36F88E80 , 32'h05CB7A70 , 32'hC2AAC600 , 32'h2AC1C0C0 , 32'h20335D80 , 32'h0B294540 , 32'hE1C73820 , 32'h10A26D20 , 32'h037008C8 , 32'hEDDBB2C0 , 32'h09570700 , 32'hFE081650 , 32'hFA302CD8 , 32'hF40244D0 , 32'h02A907D0 , 32'hFD7A4328 , 32'hFD506558 , 32'hE71ECEA0 , 32'hEE8EDCE0 , 32'hE8E3FEA0 , 32'hEE9D50E0 , 32'hF9877AF8 , 32'hDB5D3A80 , 32'h011BD91C , 32'h182115C0 , 32'hFD008770 , 32'hDBF47800 , 32'h10C0FD60 , 32'hE9F87FA0 , 32'hEB959C00 , 32'h2902E500 , 32'h0A78CAB0 , 32'h0A4A8FD0 , 32'h0A456A90 , 32'hF0564E20} , 
{32'hF4843F50 , 32'hA3E39C00 , 32'h1F438D80 , 32'hF5288A50 , 32'h9216C680 , 32'h30301840 , 32'h5A673700 , 32'h1DCF1560 , 32'hFB023C00 , 32'h2CBA8340 , 32'h2ACE7400 , 32'h00A706B7 , 32'h242B1440 , 32'hA3278D80 , 32'hE661B520 , 32'hF1F44440 , 32'h11B3E860 , 32'h3E7A5A80 , 32'hEE68E800 , 32'hE4F8E4C0 , 32'h187A4D40 , 32'h13476360 , 32'h20BFF880 , 32'h058EC1A8 , 32'h0F662170 , 32'hF755C2C0 , 32'h166A9DC0 , 32'hDAC886C0 , 32'hE78F2DC0 , 32'h0A80F7E0 , 32'h02B14F9C , 32'hFAAF7B48 , 32'hFDC760E4 , 32'hEBAB53C0 , 32'hEE4176E0 , 32'h264E4EC0 , 32'h03235FF0} , 
{32'hE0316820 , 32'hDFF214C0 , 32'h1046B920 , 32'hF201BCD0 , 32'h88B96780 , 32'h0FBE52F0 , 32'h241BF1C0 , 32'hF3302CC0 , 32'hEDE589E0 , 32'h1DBBBB80 , 32'h09137880 , 32'h21541BC0 , 32'h106A3F00 , 32'h0A936070 , 32'hE530F6C0 , 32'h0B20EF60 , 32'h01FE2C64 , 32'h04B65E50 , 32'h2B39B880 , 32'hC47986C0 , 32'hEE60F6E0 , 32'hF55C4CF0 , 32'hE070DD80 , 32'h0667E460 , 32'h1B0483E0 , 32'h04BC64B0 , 32'hF2453F80 , 32'hD3C71080 , 32'h19E13140 , 32'h0A1457B0 , 32'hF7FEF270 , 32'hED9FA1A0 , 32'hF7A74D90 , 32'hF892A280 , 32'h0EBA74E0 , 32'hF40CFB00 , 32'hEFE5E3E0} , 
{32'hF89599B0 , 32'h05B27718 , 32'hDE9B50C0 , 32'hF33616A0 , 32'h909E7C00 , 32'h1CAB6340 , 32'h20300480 , 32'hF17292E0 , 32'hFA88BBB8 , 32'h0F8B7ED0 , 32'hFF4B0633 , 32'h4DB81680 , 32'h0BCEBCA0 , 32'h08869090 , 32'h1AD8DDE0 , 32'h003B5579 , 32'h279BE500 , 32'hE266F5A0 , 32'h2FF5E880 , 32'h0452FE10 , 32'hFCEF1624 , 32'h0E7B2A20 , 32'h030CDA6C , 32'h03BEE86C , 32'h0C8F04C0 , 32'h0D0164F0 , 32'h113FB940 , 32'h083B04D0 , 32'h22CE8200 , 32'hF7CB3840 , 32'hFC62F11C , 32'h30858AC0 , 32'hFE4F9284 , 32'hDD11A500 , 32'h01F2EA7C , 32'hFAE44C40 , 32'hEEC26100} , 
{32'hF256EC30 , 32'h11D63B40 , 32'h03D04A04 , 32'h1491ABE0 , 32'hF718ADC0 , 32'h029C7290 , 32'hF267B740 , 32'h0145879C , 32'hFDDDAC50 , 32'h047E67D8 , 32'h025A95AC , 32'h1272BF20 , 32'hEFAD5DA0 , 32'h2B82B380 , 32'h018632E8 , 32'hF9D5CE20 , 32'h02AC1A90 , 32'hF309D5B0 , 32'h177E9800 , 32'h070E2F08 , 32'h018A8B68 , 32'h11C0FF20 , 32'hF386A1E0 , 32'hFAD11B80 , 32'hEAA6AAC0 , 32'h02F86E18 , 32'h0099B153 , 32'hF517F3D0 , 32'h06BCEB20 , 32'hEE31CD80 , 32'h006F67DA , 32'h047C2940 , 32'hF23452E0 , 32'hFDDFE774 , 32'h05647688 , 32'hF9E864F0 , 32'h03D447E0} , 
{32'hE59E8F40 , 32'hF6CC4EE0 , 32'h05AB7EC8 , 32'h28506000 , 32'hFDAA6024 , 32'h0CA7D240 , 32'hF6E94140 , 32'hE6303340 , 32'hFA33E100 , 32'h0199D590 , 32'hF6C98580 , 32'h24464780 , 32'hEBAE5880 , 32'h0E0CCAE0 , 32'h1351AC40 , 32'h0453F5C0 , 32'hF2BDB0D0 , 32'h0CE99C10 , 32'h16C2B9E0 , 32'hFD96E958 , 32'hD6FF1900 , 32'h0AB456A0 , 32'h09C87300 , 32'hEC816220 , 32'h06362898 , 32'hF1FD8C20 , 32'hFCF57BA0 , 32'hF7689410 , 32'h01C7190C , 32'hFB4E7928 , 32'hF8202FB0 , 32'hFB076500 , 32'hF4775300 , 32'h10CE7000 , 32'h16FE5B20 , 32'h115EF120 , 32'hFA1A39C8} , 
{32'hE72F6CC0 , 32'h05F80770 , 32'h11F0D960 , 32'h26455A40 , 32'h02A5FF84 , 32'hFF2E9635 , 32'hDC22A280 , 32'hE527C440 , 32'h07C99670 , 32'h0F9F1930 , 32'hF5FC8650 , 32'h0742E600 , 32'h066991E0 , 32'h2ACE5540 , 32'hF88BA638 , 32'h1BFDA780 , 32'h33B78040 , 32'hFC863DB4 , 32'h133E6EA0 , 32'h05FAE600 , 32'h1D9618A0 , 32'hEA52FF00 , 32'h0C70BED0 , 32'hE97201A0 , 32'h2236E800 , 32'h0293E02C , 32'h01ACEC4C , 32'h1493D380 , 32'hFD06B088 , 32'hEA32C540 , 32'h1A249360 , 32'hF7C5F910 , 32'h071EE518 , 32'hF83B7AD8 , 32'h101D5580 , 32'hFF106527 , 32'hEDBE1B60} , 
{32'hF8FA0050 , 32'hEF9192A0 , 32'h0BDB4620 , 32'h28906240 , 32'h14194B60 , 32'h116F6960 , 32'hE28121A0 , 32'hEA142760 , 32'h12B69A60 , 32'h08CC5F10 , 32'h08F93C10 , 32'h1284A3E0 , 32'h0F3BEC20 , 32'hF79377A0 , 32'h0A8E6050 , 32'hFCEC62AC , 32'h1441C180 , 32'h0017D6C3 , 32'h2263B380 , 32'h0F5A2A90 , 32'hDD7370C0 , 32'hFC5966F0 , 32'h187EB720 , 32'hE6BCD340 , 32'hEBB6B8C0 , 32'hFB06D058 , 32'h0DA56DA0 , 32'h09876770 , 32'h24C50680 , 32'hF98BD6A0 , 32'hF965B0B8 , 32'h0A2A2A40 , 32'h12F0E1C0 , 32'h0014D71B , 32'hE4A8EF40 , 32'hF9079E48 , 32'h0EC29D10} , 
{32'hEB3BE840 , 32'hE23F6080 , 32'h0A7D1D30 , 32'h12DA4480 , 32'h191D65C0 , 32'h06087918 , 32'hCD63CC00 , 32'h19F06EA0 , 32'h015F1B04 , 32'h09952110 , 32'h1AB961A0 , 32'hDEDA2080 , 32'h481CBE80 , 32'h121703C0 , 32'hECE91E00 , 32'hE48DB1E0 , 32'h02560BA0 , 32'hF04C0040 , 32'h1DAE13E0 , 32'hE17BDBE0 , 32'hEE1AD0E0 , 32'hFB73CE60 , 32'hFCBB452C , 32'h034B56B4 , 32'hEE5A3960 , 32'hDC7D9480 , 32'hEA1524E0 , 32'h10DEAE60 , 32'h16FAC8E0 , 32'h11F8A3A0 , 32'h00474899 , 32'h0238F1B4 , 32'hFD231DB8 , 32'hF80E5600 , 32'hF11C0040 , 32'hE93789C0 , 32'h1F0EFC60} , 
{32'hEDBBAEC0 , 32'h052AEEB0 , 32'hF79ACA40 , 32'hDEF99BC0 , 32'h1C157EA0 , 32'h15334280 , 32'hE2596880 , 32'h1AA52AA0 , 32'h14E5D8A0 , 32'hE500A680 , 32'h10182100 , 32'hBD03E680 , 32'h0CD580F0 , 32'h08ACA040 , 32'h01A72A50 , 32'hF524ABF0 , 32'h1A34E640 , 32'hECD54200 , 32'h0C00BB50 , 32'hD6D55240 , 32'hF5636970 , 32'h0F7C1600 , 32'h15F84D20 , 32'hE9DD41E0 , 32'h099893D0 , 32'h0C8F8CB0 , 32'h08FB4800 , 32'h085DCE10 , 32'h0AD69620 , 32'hFB4A2330 , 32'hFA57A4B8 , 32'hFA689F00 , 32'hEF2C6020 , 32'hF566E8C0 , 32'h0039B5B9 , 32'hE455ADC0 , 32'hFB9B3470} , 
{32'hF132AC80 , 32'h178AEB00 , 32'hE5B4EBE0 , 32'hFA26A8C8 , 32'h12C69860 , 32'h281FC400 , 32'hE8766220 , 32'h29DD9600 , 32'h18FBAB00 , 32'hBD61AB80 , 32'h04945EC0 , 32'hBE591980 , 32'h2060E800 , 32'h0575C830 , 32'h0ABF4A20 , 32'h08291460 , 32'h0F062400 , 32'hF24E7560 , 32'h2AA5AAC0 , 32'hD5BBCCC0 , 32'hFCFD9958 , 32'h2C147180 , 32'h052B5970 , 32'hE1B28220 , 32'h1BE2F7A0 , 32'h2DAF4D00 , 32'hFCE04174 , 32'hED6234A0 , 32'hF741D360 , 32'h38CD5F80 , 32'hF4537930 , 32'hE77E6100 , 32'hF83959F8 , 32'hFACDDA18 , 32'hEA3825C0 , 32'hEF3989A0 , 32'hD7E60F40} , 
{32'hE5769A80 , 32'h0E6DA750 , 32'hF40CD5D0 , 32'h0E982120 , 32'h0D6767C0 , 32'h16D3D3C0 , 32'hFA460150 , 32'h2869FC40 , 32'h0A4917F0 , 32'h005457FB , 32'hF930F890 , 32'hDDF63440 , 32'hFEEEFA54 , 32'h2B105380 , 32'h04BDE058 , 32'h1D614B00 , 32'h226CAEC0 , 32'h065A5DE8 , 32'h1E397C60 , 32'hDC066180 , 32'h175EA840 , 32'h233532C0 , 32'h1BD6FF20 , 32'hDF601500 , 32'h20DE1540 , 32'h245399C0 , 32'hF6A36C10 , 32'hE57AFD40 , 32'hF3DCC350 , 32'h11EE9180 , 32'h1F3978E0 , 32'h20B731C0 , 32'hEA8D23C0 , 32'h1DE8D1A0 , 32'hF25B6200 , 32'h086B9930 , 32'hE2E914A0} , 
{32'h0047D021 , 32'h0D2CDC00 , 32'hFB864D10 , 32'hFBD8B8F0 , 32'h02F40260 , 32'h0A02E0A0 , 32'h0C7B11C0 , 32'h20F6A4C0 , 32'h07EAE0B8 , 32'hF4056410 , 32'h096ED6B0 , 32'hE8F0B540 , 32'hFFAA9779 , 32'h0C252A60 , 32'hFFCF7D11 , 32'h056A90D0 , 32'h0ACBC650 , 32'h07CFB6E8 , 32'hFF8FECE0 , 32'hEBCA3A40 , 32'hEBBE5C80 , 32'h0937CE20 , 32'h0C852FB0 , 32'hEAAA7AE0 , 32'h079752E8 , 32'h132A38E0 , 32'hFC898C98 , 32'h0C08F450 , 32'hFD3E4F44 , 32'h14023E00 , 32'hEE91AFE0 , 32'h02E79014 , 32'hEE1C1520 , 32'h07C6F3B0 , 32'hF84B4510 , 32'hF50CE1E0 , 32'hF3A65B20} , 
{32'h047A8378 , 32'hF5A24390 , 32'hF4FBA680 , 32'h0FE74440 , 32'hF50DC600 , 32'hFC043214 , 32'hFD9740F0 , 32'h1B14E480 , 32'h11BEE000 , 32'h06658BE0 , 32'hE17242C0 , 32'hF78ED760 , 32'hF0FAA920 , 32'hF6392890 , 32'hF1F2D480 , 32'hFE5A9CA8 , 32'hFCD63C18 , 32'h00B2DAA2 , 32'h095F5BE0 , 32'h0A2BF270 , 32'hF7750730 , 32'hF8B51460 , 32'hFEA89910 , 32'h04110560 , 32'h01F38730 , 32'hFA3A74B8 , 32'h01B13390 , 32'hFFB4A00A , 32'h0260CDA0 , 32'hFE539E04 , 32'h0712CF98 , 32'h02EC68B0 , 32'hFD51EE18 , 32'hF8A429D0 , 32'h0833F9D0 , 32'hFF7AA89D , 32'h058F6C80} , 
{32'hF7CCA9E0 , 32'hEEB2B580 , 32'hFAB45398 , 32'h1418F360 , 32'h019AE454 , 32'h000C5F5F , 32'hF8D0C7E0 , 32'hFFF1A4C1 , 32'h0CBF5570 , 32'hFA761F98 , 32'h04582DF0 , 32'h11F97E60 , 32'hF706C970 , 32'hF5FDF680 , 32'h06779C20 , 32'hF25D7770 , 32'h02760EE8 , 32'h0E8F7170 , 32'h0243DC74 , 32'hF3EAA720 , 32'h01C118C0 , 32'h0629AFE8 , 32'h03228E94 , 32'h02667B2C , 32'hF8BBF9D8 , 32'h0D575170 , 32'h0CCEFA20 , 32'h0251811C , 32'h09F04600 , 32'h03789A70 , 32'hFD2B8B3C , 32'hF9C51050 , 32'h00456C83 , 32'h08C92980 , 32'hF46F38B0 , 32'h0C251D00 , 32'hFAF4E750} , 
{32'hFFA8D2EE , 32'hFE4E5380 , 32'hFECD992C , 32'hFEEF8988 , 32'hFCB5E690 , 32'h011192A8 , 32'hFD89AD9C , 32'hFFF3184A , 32'h008720F7 , 32'hFEA73220 , 32'hFF721E82 , 32'h02AFD730 , 32'hFEC8E088 , 32'h012D839C , 32'hFDAFBE84 , 32'hFE92CBF4 , 32'h00FC9BC3 , 32'h00848A1A , 32'hFFBFE31E , 32'hFEBE7AEC , 32'hFF3F0CBE , 32'hFE0770E4 , 32'h0035EA75 , 32'h0032F1C6 , 32'h01E7BA74 , 32'hFD178000 , 32'h00CC1A9F , 32'h00C927DE , 32'hFD225888 , 32'h0042C9FD , 32'h01B29284 , 32'h01ECE8C0 , 32'hFFD8F911 , 32'h0032DDDD , 32'h00B8A4CA , 32'hFE6175C8 , 32'hFFAE92F5} , 
{32'hFFFFFA4C , 32'hFFFBDCD8 , 32'hFFFD8BFD , 32'hFFF8618D , 32'h00006A36 , 32'hFFFCCA46 , 32'h00038E02 , 32'h00075137 , 32'h000095CC , 32'h0003B11E , 32'h00052B51 , 32'hFFFD902F , 32'hFFFDE3C0 , 32'hFFF0717E , 32'hFFFFB124 , 32'hFFFC07D0 , 32'h0003CAA2 , 32'h000716BA , 32'h0002DE4B , 32'hFFF7EBA5 , 32'hFFFD8EC1 , 32'hFFFEC3E6 , 32'hFFFD3B0D , 32'h00064FDF , 32'h0001D3BC , 32'h0008F203 , 32'hFFFCB988 , 32'hFFFEAA9A , 32'h00013034 , 32'hFFFE9CB9 , 32'hFFFF94E0 , 32'hFFFEDD14 , 32'h0006038D , 32'h00053710 , 32'h0003D548 , 32'h0000FA5D , 32'h00014A82} , 
{32'h0008AD51 , 32'h0007F44E , 32'hFFFB9CC2 , 32'hFFFF8831 , 32'hFFFEB0FF , 32'h00014DB0 , 32'hFFFAA22B , 32'hFFF71718 , 32'hFFFCE17B , 32'hFFFB085C , 32'hFFF74109 , 32'hFFFC0A00 , 32'hFFFECCDC , 32'h0004E9CD , 32'hFFFA3EE6 , 32'hFFFE1A3D , 32'hFFFE8B7B , 32'h00062399 , 32'h0004CE58 , 32'hFFFCE4B9 , 32'h00039DF8 , 32'hFFFF8FF2 , 32'hFFF77F5B , 32'hFFFAC850 , 32'h000A74A5 , 32'h000272BC , 32'hFFFBEE58 , 32'hFFFEF4CE , 32'hFFF3663C , 32'hFFFDD9C5 , 32'h00093C0B , 32'h000D73B4 , 32'h0000A4B5 , 32'h0000158E , 32'h000006C2 , 32'hFFFD2EA9 , 32'h000161D6} , 
{32'h00054DC8 , 32'hFFFF53A8 , 32'hFFFD7708 , 32'h0003AF3F , 32'hFFFD9E1C , 32'h0000FD0B , 32'hFFFF94D1 , 32'hFFFD99BF , 32'hFFFE38BE , 32'h00020F8E , 32'h00018426 , 32'h0001BA83 , 32'h00034F38 , 32'hFFFD823B , 32'hFFF8727A , 32'h00025358 , 32'h00003D99 , 32'hFFF38361 , 32'hFFF724C9 , 32'hFFFCEBBE , 32'h000224A9 , 32'hFFFECA09 , 32'h0002FEC6 , 32'hFFFF981D , 32'h0008CBF4 , 32'hFFF95C23 , 32'hFFF946E3 , 32'hFFFEEC24 , 32'h000681D0 , 32'hFFFE18E2 , 32'hFFFBCB8F , 32'hFFFC6BA9 , 32'h000613E9 , 32'hFFFE3DE0 , 32'hFFFD2362 , 32'h00039BFA , 32'hFFFE1860} , 
{32'hFFFDB919 , 32'hFFFF5231 , 32'h0000D2D3 , 32'h00042DFA , 32'hFFF8BD54 , 32'h00026575 , 32'hFFF9C17A , 32'hFFF9F14D , 32'hFFFA50BE , 32'h0005ABAE , 32'h0002E5BD , 32'h00088A1C , 32'hFFFE71B0 , 32'hFFF4087B , 32'h0002DD53 , 32'hFFFFBD87 , 32'hFFF65FA1 , 32'h000C18C9 , 32'h0001B72C , 32'hFFFBEA94 , 32'h00082D1E , 32'hFFFE24FF , 32'hFFFCC0C2 , 32'h00036E6D , 32'h00028C72 , 32'hFFFDC6B7 , 32'h00067D59 , 32'h0006D3CD , 32'hFFFE185B , 32'hFFFF0C25 , 32'hFFFFC05A , 32'hFFFB6BA6 , 32'hFFF6464F , 32'hFFFA9E90 , 32'hFFF9A767 , 32'hFFFA34EC , 32'h0001E558} , 
{32'h005047D5 , 32'hFFB95D3A , 32'hFFE1B08E , 32'hFFFBEF89 , 32'hFFD34E6B , 32'h00654DA5 , 32'hFFCEB0C9 , 32'h000DC369 , 32'hFF9E2E54 , 32'h0017C763 , 32'h0058F069 , 32'hFFE24322 , 32'hFFAAD244 , 32'hFFDFEDC2 , 32'hFFCDCBDE , 32'hFF9BCDC8 , 32'hFFD07ABA , 32'hFFFC908D , 32'h0010390E , 32'h0054EC26 , 32'hFFFD7F2F , 32'h001E55DD , 32'h005B4474 , 32'hFFEE079B , 32'hFFEC35D5 , 32'h00055222 , 32'hFF7D0125 , 32'h0010B3E6 , 32'h0022AEFA , 32'hFFE63B8C , 32'h00342D6D , 32'hFFDB202F , 32'hFFA67B88 , 32'h00253C43 , 32'hFFBA9330 , 32'h0014EBDD , 32'h001C0C10} , 
{32'h0069C884 , 32'hFFC041D0 , 32'hFFC61A05 , 32'hFFEBD8F2 , 32'hFFB35F95 , 32'h008F281F , 32'hFFC08FB5 , 32'h00260F72 , 32'hFF642E21 , 32'h001A63C7 , 32'h0095C6B4 , 32'hFFC1386B , 32'hFF9E98E1 , 32'hFFE39F53 , 32'hFFBF1E89 , 32'hFF7F4347 , 32'hFFEDAB48 , 32'hFFDBAEC5 , 32'h00020E30 , 32'h006E1387 , 32'h0020F27F , 32'h0008D8DA , 32'h007EE564 , 32'h000952DA , 32'h000591F8 , 32'h00015B47 , 32'hFF6F2017 , 32'h00103DEE , 32'h0035091A , 32'hFFD48AE8 , 32'h0054C28F , 32'hFFD37BDB , 32'hFF7DDF0F , 32'h001C28E3 , 32'hFFAAF17E , 32'h00138F26 , 32'h00374D06} , 
{32'hFE4B57CC , 32'hF8541898 , 32'hFF19D237 , 32'h0318C950 , 32'h0C2A86F0 , 32'hF8883978 , 32'hEEFB21C0 , 32'hF6DE24C0 , 32'hF2E4D5E0 , 32'h05B71AF8 , 32'hEBBABFC0 , 32'hFDF00DD0 , 32'h03AB3AB8 , 32'h06E75968 , 32'hECEEC4A0 , 32'hF40D06F0 , 32'hF5DC0C70 , 32'hEE477A60 , 32'hFB37C3F0 , 32'hEDE0DAA0 , 32'hFF3758AA , 32'hFE483BB0 , 32'hF6EB7CB0 , 32'hFA635D40 , 32'hFF5FFD36 , 32'h07C00D58 , 32'hF34F0AD0 , 32'h06C901D0 , 32'h0038E7BF , 32'h131190C0 , 32'hF6B0FDD0 , 32'h113C3DA0 , 32'hFA5F6460 , 32'h013F9D80 , 32'hFBE2CA48 , 32'h045C36B8 , 32'h0856D8E0} , 
{32'hD2FE5C80 , 32'hBCF4EF80 , 32'h0BD45FE0 , 32'hF93E63B0 , 32'h3FABB900 , 32'h06B67D68 , 32'h0F2901D0 , 32'h05C44738 , 32'hE25CEDC0 , 32'h04B246D8 , 32'hF4D318B0 , 32'hFD184674 , 32'hED79F320 , 32'h19BBF5C0 , 32'hFA63B688 , 32'h1576DE40 , 32'hFAB69F48 , 32'hF58EE220 , 32'hF2DCF8C0 , 32'h0F3769F0 , 32'h112EBCA0 , 32'h0DC455F0 , 32'h0148FBB8 , 32'hF28DF440 , 32'hE80273E0 , 32'h12BC6C40 , 32'h0B63BC60 , 32'h12928B40 , 32'h20F91900 , 32'h137A59A0 , 32'hFC75DB78 , 32'h0AF23700 , 32'h04FF3970 , 32'h11655040 , 32'hFEC134CC , 32'h0BE3A880 , 32'h08E652C0} , 
{32'hE48D18C0 , 32'hDF2C7100 , 32'hE243B9C0 , 32'hE341D0E0 , 32'h3B3FC7C0 , 32'h1511F780 , 32'h11C0E6E0 , 32'h0C587B30 , 32'hECC0DCE0 , 32'h019CCDB8 , 32'hEB2A90A0 , 32'h11AECA80 , 32'hFB894228 , 32'hFEBFEA38 , 32'h02932424 , 32'h11F44560 , 32'h08E071A0 , 32'hF6EC5170 , 32'h066143D0 , 32'hFE83020C , 32'h0412DD88 , 32'hFC60E20C , 32'h08CCF450 , 32'h00F77490 , 32'hEE619280 , 32'h04BDE9E0 , 32'hFD45B7A8 , 32'h08F632B0 , 32'h00136741 , 32'hEE292D20 , 32'h104B2AC0 , 32'hEE40C520 , 32'hF6468570 , 32'hF30FA7C0 , 32'h0AF305B0 , 32'hFBF61DE0 , 32'hFFBCCFA4} , 
{32'hE535C860 , 32'hCB40AC40 , 32'hF67C52C0 , 32'hF7F787A0 , 32'h3B4E2840 , 32'h35BC7E40 , 32'h23797E40 , 32'h10EE0B00 , 32'hE7AA0EA0 , 32'h0C2380D0 , 32'hF285EF40 , 32'hE56ADA40 , 32'h17CC41A0 , 32'h197C5100 , 32'h0E3BA6F0 , 32'hF71A05B0 , 32'h2F23A640 , 32'hF7604060 , 32'hFE18C7A8 , 32'hF49EBCF0 , 32'hCAC6BE00 , 32'hF243B320 , 32'hDE7CB740 , 32'h01EB4BE0 , 32'hD4511040 , 32'h15AEACA0 , 32'hFEF48EB0 , 32'hFEE33464 , 32'hCDE4D140 , 32'hCAFCEF80 , 32'h35AD5080 , 32'hD8C8AAC0 , 32'hF8FAFFA8 , 32'h119A49E0 , 32'h1306D3E0 , 32'h29022240 , 32'hFC46DEDC} , 
{32'hE6B29220 , 32'hBEDD8780 , 32'hFD931394 , 32'hF8611C38 , 32'h5A0B7500 , 32'h3222BC80 , 32'h1E2E9480 , 32'h0DD9F510 , 32'hDB42A5C0 , 32'h115DC900 , 32'hD78813C0 , 32'hFFF04B0F , 32'hF7AFD0F0 , 32'h33059480 , 32'h353CFF80 , 32'hE7F73960 , 32'h0858BE30 , 32'hF4BB4DB0 , 32'h10CC3900 , 32'h23797500 , 32'hFFCD51B6 , 32'hDD35F580 , 32'hF733F4F0 , 32'h021345D8 , 32'hD18D3900 , 32'h066E4C70 , 32'h0DA55950 , 32'h01796F70 , 32'hE6C94920 , 32'h105E0480 , 32'h3130E3C0 , 32'hEFA16800 , 32'hE9A17820 , 32'hF64F3B40 , 32'hFE519DB4 , 32'hF32F3350 , 32'hDFCD7000} , 
{32'hD8B2F980 , 32'h9FC79880 , 32'hD7C74240 , 32'hE6049100 , 32'h46BB0C80 , 32'h20BA8C80 , 32'h3569A240 , 32'h08AAF950 , 32'hE2ED9E60 , 32'h1518FC80 , 32'hDDCC5D80 , 32'hE99919A0 , 32'h08DA6520 , 32'h0203F05C , 32'h38C41B40 , 32'hF5187910 , 32'hFD169E04 , 32'hFCB78F20 , 32'hF8B2BF50 , 32'h057AC3A0 , 32'hF7381CC0 , 32'hF5A22E80 , 32'hFAFA6608 , 32'hFBB920D0 , 32'hF36C9BB0 , 32'hFB4D75E0 , 32'h05E4E770 , 32'hFEE7D5E4 , 32'hD4E6A880 , 32'h0B315790 , 32'h127BA3C0 , 32'hD724E180 , 32'hFB7640C8 , 32'hFEBB22FC , 32'h03783EA4 , 32'hE8FD1C20 , 32'hEDB5D6A0} , 
{32'hD9290F00 , 32'hB5E6A800 , 32'hE7E03580 , 32'hBCD0C680 , 32'h28C9E880 , 32'h2411FF00 , 32'h3EC9DAC0 , 32'h07C5A740 , 32'hDE4EF5C0 , 32'h3A7C6F80 , 32'hC68F1800 , 32'hF095DFF0 , 32'h23505300 , 32'hAC2C0B80 , 32'h0CAD2C50 , 32'h01D0FB34 , 32'hFD25316C , 32'h44FA7380 , 32'hE46D64E0 , 32'hF3A451C0 , 32'h0539CF20 , 32'hF4F7FA10 , 32'h249C05C0 , 32'h06798D70 , 32'h1E55FDC0 , 32'h02E608E8 , 32'hF0E889F0 , 32'hF73B5FC0 , 32'hFF045857 , 32'hD41E55C0 , 32'h0177FBA0 , 32'hE84A1A20 , 32'hFB567F58 , 32'h003AD09A , 32'hFE556B84 , 32'h12728A00 , 32'hFA30D568} , 
{32'hD5CA8C80 , 32'hA3468C00 , 32'hC6F10940 , 32'hB45C3C80 , 32'hE70E2280 , 32'h1C18EB00 , 32'h63C23880 , 32'h0D869850 , 32'hE32861E0 , 32'h1CD33080 , 32'hE0A69540 , 32'h2BAA2180 , 32'h1F772DC0 , 32'hC961E540 , 32'hE7504760 , 32'h0EF36DD0 , 32'h099927C0 , 32'h357D2500 , 32'hFDB8232C , 32'hC579F780 , 32'h1D752B40 , 32'h145D0900 , 32'hF9BD51A0 , 32'hE6AC9D60 , 32'h00B68D9B , 32'hF2F70610 , 32'hD26FCBC0 , 32'hDAD8DBC0 , 32'h1560A620 , 32'hF9C08668 , 32'hFB0F7A88 , 32'hF8B393B0 , 32'h04E4E768 , 32'hFF30B4C3 , 32'h031C2404 , 32'hD97DA4C0 , 32'h1AD32B40} , 
{32'hDE6BC4C0 , 32'hAACB3300 , 32'hCDEF1B80 , 32'hC8273A80 , 32'hA74C0F00 , 32'h0D4AFF60 , 32'h618C0400 , 32'h016BF9A8 , 32'hECDF7440 , 32'h01BA44C8 , 32'h0C353970 , 32'h4A576400 , 32'h1191F780 , 32'h08F3F810 , 32'hB5A47280 , 32'h277B6140 , 32'h16B31120 , 32'hD4CD4800 , 32'h29E20780 , 32'hE13A1960 , 32'hDFE30C40 , 32'h1FD8EA40 , 32'hCB38FC80 , 32'hE5280000 , 32'h149D2AE0 , 32'h19512820 , 32'hF529EAC0 , 32'hEAC6ED60 , 32'h3C80B540 , 32'hDDD4A140 , 32'hF37E7050 , 32'hF2DAB970 , 32'hF9D8B290 , 32'hEAF1F180 , 32'h14101B80 , 32'h0C777E10 , 32'h0AD35050} , 
{32'hF5A0CF00 , 32'hF6987090 , 32'h198C44C0 , 32'h13811FC0 , 32'hF4E6D0F0 , 32'h203CF2C0 , 32'h2263C140 , 32'h1E922560 , 32'hE2197320 , 32'hF6257A30 , 32'hE0E40780 , 32'h314F44C0 , 32'h109DA980 , 32'h22280D80 , 32'hF1CC3B00 , 32'h08B5EEB0 , 32'h1D9A4440 , 32'hDA7DC000 , 32'h07F13B38 , 32'hF9CA2BC8 , 32'hEF51ED40 , 32'hEF7B29E0 , 32'h0EF2A500 , 32'hFA4A2CD0 , 32'h02E98718 , 32'h0711C8E0 , 32'h11847760 , 32'hE8321000 , 32'h2254C400 , 32'hE6ECB080 , 32'h06A99EF0 , 32'h0BCB2A80 , 32'h0A100250 , 32'hF6B7C6E0 , 32'h03AEDC44 , 32'hEFA3CFE0 , 32'hFCFC2760} , 
{32'hF2FCE8B0 , 32'hFB7646D8 , 32'h0FED74E0 , 32'h05EBF830 , 32'hF0EF3730 , 32'h19AC8600 , 32'h04C58A40 , 32'h190A8C60 , 32'h01A4F6E4 , 32'hF4BE1B00 , 32'h0A8BEA60 , 32'h16224760 , 32'hEA0DAC80 , 32'h293595C0 , 32'h0075D2A7 , 32'h0C846AF0 , 32'h0918F250 , 32'h0C894F70 , 32'h10D9BAC0 , 32'hFF1DEDA8 , 32'h03CA65C4 , 32'h0000F801 , 32'hF1EE77F0 , 32'hEE05A660 , 32'h06977C20 , 32'hF616DB60 , 32'h1A16CD00 , 32'hEFB95D00 , 32'hFC184918 , 32'hE37B6400 , 32'h1560AD00 , 32'hFA602888 , 32'h0C867360 , 32'hEBB8E400 , 32'h0931AE40 , 32'hD9CED240 , 32'hEDF7C700} , 
{32'hFECD0FC0 , 32'hF1EE98E0 , 32'h17CC60C0 , 32'h3D85E300 , 32'h10A20C60 , 32'h01A56D88 , 32'hDA6675C0 , 32'hE8AFE060 , 32'hF394D990 , 32'h14887BE0 , 32'hEFFE3840 , 32'h2AA64240 , 32'h0CB797C0 , 32'h17183AC0 , 32'hF1F9CD10 , 32'h3DED6C80 , 32'hFC50E6D0 , 32'h12067FE0 , 32'h1E05B4A0 , 32'h30991600 , 32'hEE860580 , 32'hFD48B55C , 32'hE2C88580 , 32'h1C122680 , 32'h2137D500 , 32'hDACEE140 , 32'h003E569C , 32'hEB35DCC0 , 32'hFFD11807 , 32'hFBD5BAB0 , 32'hFD6D4000 , 32'h037374B4 , 32'hE1F35560 , 32'h03367FE8 , 32'hF92CF1D8 , 32'hE68544E0 , 32'hFBA09330} , 
{32'hE8960D80 , 32'hF3B5E2A0 , 32'h18D85BC0 , 32'h27BC8D40 , 32'h2147DCC0 , 32'h193E3400 , 32'hD41EF900 , 32'hC7224500 , 32'h1569A3A0 , 32'h13715FA0 , 32'h1F756FE0 , 32'h0FF6FFD0 , 32'h36528AC0 , 32'hFE8A98D0 , 32'hF41A3FD0 , 32'hF697F180 , 32'h2FDA97C0 , 32'h106E23A0 , 32'h06028C90 , 32'h10617040 , 32'h039E99BC , 32'hF08861A0 , 32'h185F2E60 , 32'hBC002D00 , 32'h18814B60 , 32'hE9C0F000 , 32'h0DB53A40 , 32'h0DFD0190 , 32'h2A5685C0 , 32'h0DC91790 , 32'h03DEAA88 , 32'hF8712D80 , 32'h11419C20 , 32'h0D4DDF70 , 32'h05CDEC38 , 32'hE9B00560 , 32'h1156DC60} , 
{32'hEE86E8A0 , 32'hF451BC80 , 32'h0B717BA0 , 32'h1F9C3300 , 32'h208C9D80 , 32'h16F66800 , 32'hE96B99C0 , 32'h0CA0A0C0 , 32'h0C581550 , 32'h0FD19B00 , 32'h1B092780 , 32'hF23D9050 , 32'h22230480 , 32'hFE57CD68 , 32'hFABB2988 , 32'h0069A4A2 , 32'h1FA18260 , 32'h13452B40 , 32'h181D7D80 , 32'hF2AE0810 , 32'hFAD5D7E0 , 32'hED5EACE0 , 32'hF3054640 , 32'hF40B33C0 , 32'hFE9FA220 , 32'h090E9A20 , 32'hE4917720 , 32'h019C12C4 , 32'h09D46580 , 32'hEAB5AF40 , 32'h0537AC58 , 32'hED0EA520 , 32'h07FCE6B0 , 32'hFDF82A5C , 32'hF0413FC0 , 32'h0A444B50 , 32'h28ABA380} , 
{32'h00B1183C , 32'hE2A9C560 , 32'h0949B800 , 32'h27C32900 , 32'h175A8640 , 32'h09999670 , 32'hE4D38A60 , 32'hF6FD1990 , 32'h14D93B20 , 32'h081324C0 , 32'h2A1A8F00 , 32'hEF6D9380 , 32'h17976AC0 , 32'hF6B31650 , 32'h02771CB8 , 32'hF8317510 , 32'h22793D40 , 32'h0707D8B0 , 32'h0265E190 , 32'hE53FB400 , 32'hF6746340 , 32'h01633350 , 32'hFF1F03FB , 32'h0B188A30 , 32'hF1C163F0 , 32'hFCEEA4A4 , 32'hF62721D0 , 32'h0C9F2A80 , 32'h149FC6C0 , 32'hE6E57FC0 , 32'h03716ABC , 32'h05733730 , 32'hFA71A3E0 , 32'hDF6291C0 , 32'h0ACE7DF0 , 32'hE21EFD80 , 32'hF8B24D00} , 
{32'h195BE600 , 32'h20D57B80 , 32'hDECDA940 , 32'hFA93E250 , 32'h11749BA0 , 32'hFDF675A4 , 32'h0343C714 , 32'h0823DB70 , 32'h208AE040 , 32'hF2A34B70 , 32'h05F38BA0 , 32'hF3B9BDF0 , 32'h029D2EA8 , 32'hF3AEBF00 , 32'h07158678 , 32'hE9256600 , 32'h0853DE70 , 32'hF85F0788 , 32'h17840E60 , 32'hC13A9440 , 32'hD9C32080 , 32'h013187C4 , 32'h2483C200 , 32'hF33DF9D0 , 32'hD1C28800 , 32'hFC158D20 , 32'hF7F20600 , 32'hF6FD2140 , 32'hC9742E00 , 32'hE3A897A0 , 32'h0B3E5C90 , 32'h1843C7E0 , 32'h01032D04 , 32'hD6E36940 , 32'hF06D0260 , 32'hC7C8EB00 , 32'hFB0A0938} , 
{32'hF337C910 , 32'h0B70D650 , 32'h08DA2F20 , 32'hF703B550 , 32'h00AB0650 , 32'h0B23B690 , 32'hF90824A0 , 32'hE7C31FC0 , 32'hF0D63140 , 32'hD0B44C00 , 32'h15F62280 , 32'h01B85138 , 32'h0BE722D0 , 32'hED16B2E0 , 32'h005D868D , 32'h13D60040 , 32'h02EF7604 , 32'hEA152640 , 32'hF1B4BB20 , 32'hE24AC440 , 32'hFCB21608 , 32'h025104C8 , 32'h02670A6C , 32'hE7B89BC0 , 32'h02FCC23C , 32'h0AC76E70 , 32'h0666C898 , 32'hFDC8BCD8 , 32'h004C351D , 32'hFD2C1C84 , 32'h091129E0 , 32'hF2F22EA0 , 32'hDE7E8540 , 32'hF10E3870 , 32'hF07D27D0 , 32'hE9D04F80 , 32'h0721B898} , 
{32'hF900D420 , 32'h04A863C8 , 32'hF73EEBF0 , 32'h0427D340 , 32'hFE20EEB4 , 32'h0773A588 , 32'h08DE5070 , 32'h12925A20 , 32'h0A6B7EC0 , 32'hEECE4FE0 , 32'h10218260 , 32'h0B018C50 , 32'hFA401EF8 , 32'h065B5BC8 , 32'h00C947A3 , 32'hF0EF61A0 , 32'h15143B00 , 32'h17E25E60 , 32'hF7320D00 , 32'h01A52334 , 32'h02DE4228 , 32'hF8C67540 , 32'h02505E00 , 32'hF7146460 , 32'h01DB4548 , 32'hF9A0AA78 , 32'hFEE20390 , 32'hF12C92D0 , 32'hEECF29C0 , 32'h0FE572F0 , 32'hF2E37490 , 32'h0E697220 , 32'hFD7FBC40 , 32'hF6ED1930 , 32'h0B2AB790 , 32'h0A8B9290 , 32'h17FA6980} , 
{32'hF99B6530 , 32'h14894340 , 32'hFF8AF592 , 32'hF9102A40 , 32'h19CD1020 , 32'h1027C440 , 32'h1674E7E0 , 32'h08B3AF90 , 32'h13C28EE0 , 32'hD8AC4040 , 32'h03DAFC48 , 32'h0261986C , 32'h0F9B9AA0 , 32'hF45122D0 , 32'h144C67E0 , 32'hF837AE78 , 32'h0266BB28 , 32'hF68E3CE0 , 32'h04AC7680 , 32'hED6F1AA0 , 32'hF9359D68 , 32'h2156B480 , 32'hF4F419A0 , 32'hE9C704E0 , 32'h080F00F0 , 32'hE95479E0 , 32'h2C64FAC0 , 32'h039B4CDC , 32'hEC41A0A0 , 32'hFEA926D4 , 32'hE2AE3BC0 , 32'h135F7A40 , 32'hF868F648 , 32'h01AFBEDC , 32'h16B226A0 , 32'h1E3A2980 , 32'h24B56300} , 
{32'h002476F4 , 32'hFED5BD50 , 32'hFD5BDF64 , 32'hFCCD8C48 , 32'hFDF3BFF0 , 32'hFE6F37B0 , 32'h036F4BE4 , 32'hFFF3C23A , 32'hFEAD9C68 , 32'hFD8813D4 , 32'hFF61FCB7 , 32'h011C4710 , 32'hFCDA75EC , 32'h01DDBD88 , 32'hFBB26CC8 , 32'h067B96E0 , 32'hFD62DC2C , 32'h00EF3BBA , 32'h02637344 , 32'hFE0ACC20 , 32'hF8A55268 , 32'h065E3788 , 32'hFAC6FB28 , 32'h045596A8 , 32'h00E58A30 , 32'h04A05B10 , 32'h010CB10C , 32'h0408AF48 , 32'h00D2ED15 , 32'hFD036978 , 32'hFFB9BAFC , 32'hFE344118 , 32'hFD947910 , 32'h00F8C2E0 , 32'h025991D0 , 32'h011CBB08 , 32'h03BFECE4} , 
{32'hFFF92D4D , 32'hFFFFA994 , 32'h000534A6 , 32'h00070321 , 32'hFFFF2E57 , 32'hFFFD1B4F , 32'hFFFF55B9 , 32'hFFFD6875 , 32'h0001A84A , 32'hFFFE4AE6 , 32'hFFFAA63F , 32'h00006BD3 , 32'h00048C87 , 32'hFFFD4CB6 , 32'h0004653C , 32'h0004E9D6 , 32'h00022EAB , 32'h00044C0B , 32'hFFFE7B4D , 32'hFFF8F3E5 , 32'h00026FDA , 32'h00002017 , 32'hFFF941CC , 32'h0005A8FD , 32'h0003FAC2 , 32'hFFFC83C1 , 32'hFFFD7443 , 32'h00005745 , 32'h0007B03A , 32'hFFFDDAF5 , 32'hFFFFFCB0 , 32'h0003E83B , 32'h0001FE6C , 32'h00023F49 , 32'hFFF717E1 , 32'h00021E63 , 32'h000139DB} , 
{32'h00004D97 , 32'h0002401B , 32'h0005818C , 32'hFFF5FB09 , 32'hFFF7EFE6 , 32'h0006BB85 , 32'hFFFC488F , 32'h0002230F , 32'h0002A32E , 32'h0000BD8D , 32'h000069E2 , 32'hFFFDE376 , 32'h0000DFA1 , 32'hFFF9C79E , 32'h0003B7B6 , 32'hFFFFAD80 , 32'hFFFFD64D , 32'h000128F7 , 32'hFFFB783D , 32'h0000863A , 32'h0000DCD7 , 32'h000522BF , 32'hFFF97E22 , 32'hFFFD8714 , 32'hFFFF54F0 , 32'hFFFA307D , 32'h0005D29A , 32'hFFFC18BF , 32'h00064936 , 32'h00093D17 , 32'hFFFCAC51 , 32'hFFFD1355 , 32'h0002F030 , 32'hFFFEF457 , 32'hFFFD8A4C , 32'h00014D36 , 32'hFFFFB87D} , 
{32'hFFF7F6C5 , 32'h00009AA6 , 32'h000B0B4B , 32'hFFFE7857 , 32'hFFFF177D , 32'h0005243E , 32'hFFFE76A6 , 32'hFFFEB19D , 32'h00053C21 , 32'h0008C91D , 32'hFFFE5DE8 , 32'hFFFF0314 , 32'hFFF81913 , 32'h0002E6A0 , 32'h0001964E , 32'hFFFCA468 , 32'h00020191 , 32'hFFFA5838 , 32'h000288DB , 32'hFFFBC6BA , 32'h0003BA9B , 32'h0008E02C , 32'hFFFCE77F , 32'hFFF1D73C , 32'hFFFB7FB2 , 32'hFFFD7E0E , 32'h00018D59 , 32'h00000177 , 32'hFFFB6D4F , 32'hFFFCF6E8 , 32'h0000D770 , 32'hFFFAAE95 , 32'h0006C2D0 , 32'hFFFCEBCF , 32'hFFFF285D , 32'hFFFE9D6B , 32'hFFF96C41} , 
{32'hFFFD600C , 32'h00016598 , 32'h00074920 , 32'hFFF627D1 , 32'hFFFEC874 , 32'hFFFD799E , 32'hFFFF32DF , 32'h0006586F , 32'h0002110A , 32'h000AA72E , 32'hFFFE584C , 32'hFFFFA588 , 32'hFFFCA30A , 32'hFFF81C33 , 32'h00095B26 , 32'h0003B285 , 32'hFFFE8DC0 , 32'hFFFC8CB5 , 32'hFFF8C5C6 , 32'h00033CB5 , 32'h000593CA , 32'hFFF6EEBB , 32'hFFFE2689 , 32'hFFFD2DA1 , 32'hFFFEA678 , 32'h00015E16 , 32'h00014456 , 32'hFFFDEDE5 , 32'h000B5136 , 32'hFFFFB449 , 32'hFFFE3EDD , 32'h00079C0A , 32'h00034787 , 32'h000820AF , 32'hFFFEEE9E , 32'hFFFA3AA1 , 32'hFFFB4077} , 
{32'h0002FD2C , 32'h0000C69A , 32'h0007F121 , 32'h000B1C7F , 32'hFFF86875 , 32'hFFFC719E , 32'hFFFEAEE7 , 32'h000540EC , 32'hFFF95C2C , 32'hFFFA0DAD , 32'h0002DB02 , 32'hFFFE132C , 32'h00063E48 , 32'hFFFC4AE4 , 32'h0005B9AC , 32'h0000E679 , 32'h00023B20 , 32'h0004E357 , 32'hFFFC0158 , 32'h0000684D , 32'h000220A0 , 32'h0002BB7C , 32'hFFFD0F8F , 32'hFFFF0BDC , 32'hFFFB2C24 , 32'h00042A1E , 32'hFFFF0D21 , 32'hFFFC79FD , 32'hFFFE885B , 32'h0005EECC , 32'h00001D9B , 32'hFFFE4EF9 , 32'h0001E3E6 , 32'hFFFE5812 , 32'h00006284 , 32'h001047FA , 32'hFFFF0903} , 
{32'h00032F21 , 32'h000083C1 , 32'h00029377 , 32'hFFFAA90F , 32'hFFFDDA1C , 32'hFFFFAD6E , 32'h000268AC , 32'hFFFB0CDA , 32'h000328A4 , 32'h00043278 , 32'h0005773E , 32'h000120B7 , 32'hFFFF0C0A , 32'hFFFD5301 , 32'hFFFEA652 , 32'hFFFB9AD4 , 32'hFFF7E5DB , 32'hFFFBDE7C , 32'hFFFB6CB5 , 32'h000398CB , 32'h0007E827 , 32'hFFF9D1C6 , 32'hFFFE5651 , 32'h0002DAD9 , 32'h000A5A52 , 32'h0008EC64 , 32'h00023F28 , 32'hFFF6F41D , 32'h00047DA4 , 32'h0006E675 , 32'h0000D70F , 32'h0000F920 , 32'h00032C00 , 32'h0002E006 , 32'h000387C1 , 32'hFFFD0B07 , 32'h00066622} , 
{32'h00056977 , 32'h000C98DA , 32'hFFFA2DAD , 32'hFFFEBB70 , 32'hFFF6F05D , 32'h00038648 , 32'h00100167 , 32'h000ECBCA , 32'h0004EADD , 32'h000A67A2 , 32'h00038337 , 32'hFFFEF4CC , 32'h00124F2F , 32'h00016677 , 32'hFFF44023 , 32'h00085B6B , 32'h00018BB8 , 32'hFFF3DBE4 , 32'hFFFB9FAE , 32'hFFFCCD7D , 32'h000684C6 , 32'hFFFF8CA5 , 32'hFFFDB519 , 32'h000934D3 , 32'h000733E0 , 32'h000128E8 , 32'h00041AAF , 32'h000138BE , 32'hFFFBB919 , 32'hFFFF5AB3 , 32'hFFFEDBB3 , 32'hFFFBD839 , 32'h00061193 , 32'h000372D2 , 32'hFFFDEEC0 , 32'hFFFC95CF , 32'hFFFDD90C} , 
{32'hFE626518 , 32'hFC5C1744 , 32'hFD7343E0 , 32'hFDCD98EC , 32'h00ED3364 , 32'h0332F4D8 , 32'h02EEA814 , 32'hFEF2A6C4 , 32'h0062EB7F , 32'h035AF3F0 , 32'hFCDA8050 , 32'hFD88444C , 32'hFF63B823 , 32'hFEDB4AB4 , 32'h0A47D870 , 32'hFDEBF150 , 32'h035D2D40 , 32'hFC111730 , 32'h0234E9B0 , 32'h01543D1C , 32'hFCA1D0D8 , 32'hFE575F54 , 32'h00489A93 , 32'h0392180C , 32'h06316B60 , 32'hFDE77918 , 32'hFD59FDCC , 32'h012DF094 , 32'hFF1A2AAC , 32'h061F1F70 , 32'hFBA73418 , 32'h037178A0 , 32'h04BD7240 , 32'hFB70DC88 , 32'h00160EDE , 32'h01A2C978 , 32'hFFACC4BA} , 
{32'hF5369C30 , 32'hE95745A0 , 32'hFCE8D404 , 32'h11A8EEA0 , 32'h0A9AA2B0 , 32'h015B6288 , 32'hFD311924 , 32'hEFF2C700 , 32'h05760600 , 32'hFC7B9A34 , 32'hFE92C1A8 , 32'h10029F80 , 32'hEAB59EE0 , 32'hF5FFB320 , 32'h179ADD40 , 32'hF0C88320 , 32'hFE58CFE8 , 32'h1B518060 , 32'h17FD07C0 , 32'h027E6F64 , 32'hE0D60B00 , 32'h110754A0 , 32'h0EEC0330 , 32'hE5EBFBE0 , 32'hF953CEF8 , 32'h0DD646D0 , 32'hFCB98004 , 32'h0234172C , 32'h1259D120 , 32'h121A6020 , 32'hFF4EF05D , 32'h0A3F8FD0 , 32'h1DB0A7E0 , 32'h05A76CE0 , 32'h0029C3DC , 32'h12894D60 , 32'h00D38E3E} , 
{32'hE5FBFD20 , 32'hE7BD58C0 , 32'hD144B140 , 32'hFD60BAEC , 32'h1E4C5020 , 32'h100D8E00 , 32'hE14E1A00 , 32'h00584D48 , 32'hDF817F80 , 32'hEB072260 , 32'h14C6D5A0 , 32'h0A6811F0 , 32'hE059E880 , 32'hEF4B7DC0 , 32'hFF16618D , 32'hF4139E20 , 32'hE71B5900 , 32'h010B35A4 , 32'h239EEE00 , 32'h1559C5E0 , 32'hF58F4A60 , 32'hFA04B630 , 32'h10CEA260 , 32'hEFE83A60 , 32'h059CCA70 , 32'h10865320 , 32'h0763B188 , 32'h06F1C250 , 32'h09229AE0 , 32'h17E1BFA0 , 32'h04C085C8 , 32'hEFE44A80 , 32'h060DD8C8 , 32'hECBE0F00 , 32'h1617FC80 , 32'h054DC9C8 , 32'hFDBDB1D0} , 
{32'hF788A6F0 , 32'hFA9E5C60 , 32'hE298F140 , 32'h055AEBC0 , 32'h2BB65D80 , 32'hEED24BA0 , 32'hD832D300 , 32'hF399F220 , 32'hF3F4E5A0 , 32'hF5A50110 , 32'hFED2D104 , 32'hF0A956B0 , 32'h0149586C , 32'h1C01A0E0 , 32'h1AB472E0 , 32'hE92782A0 , 32'hED201980 , 32'hF047CB90 , 32'h0BE77B30 , 32'h0CAE7630 , 32'hF71715D0 , 32'hE7B48E00 , 32'hFF9FD983 , 32'h0A783CC0 , 32'h0E5DA3F0 , 32'h10D8FBA0 , 32'h02DD3C84 , 32'hFCDD12B0 , 32'h067719C8 , 32'h0B2BF0A0 , 32'h0D47EFB0 , 32'hF723CA10 , 32'hEB9F5D80 , 32'hFDAA561C , 32'h25E79A00 , 32'h0C5618C0 , 32'h06664908} , 
{32'hEC0E9D00 , 32'hE5A63F80 , 32'hD5447300 , 32'hDDDFC9C0 , 32'h4087AF80 , 32'hF493A8F0 , 32'hE01686A0 , 32'hFF8B005D , 32'hEBB814A0 , 32'h04C2F470 , 32'hE8A83F40 , 32'hF7E12D70 , 32'h150F2320 , 32'hF6193810 , 32'hE1CF9220 , 32'hFEEB2330 , 32'hF2327570 , 32'h0451FFC8 , 32'hE798CD00 , 32'hF2A79DA0 , 32'hEF7E95A0 , 32'h057D9F20 , 32'h1EB88CC0 , 32'h147C2660 , 32'h11407940 , 32'h05BEC230 , 32'h07365120 , 32'h0107DD8C , 32'hFDE21704 , 32'hF768E260 , 32'hFC142798 , 32'h20791D00 , 32'hFF5F9957 , 32'hE72BE9C0 , 32'h0B2BFAE0 , 32'h1C2C86E0 , 32'h10BD8F20} , 
{32'hE57A4980 , 32'hD618DE00 , 32'hD4BF7880 , 32'hDFFEA300 , 32'h5C109A00 , 32'hFF9CE63B , 32'hEEC43540 , 32'h0F2FE550 , 32'hFD360224 , 32'h0877C960 , 32'hFAF46E28 , 32'hEC60AC20 , 32'h146139C0 , 32'hEE7A5D60 , 32'hFF0683B0 , 32'hF0F217B0 , 32'hF90F2820 , 32'h15FFC5A0 , 32'hE51A9320 , 32'h0F403060 , 32'hDEE12200 , 32'hE91D03E0 , 32'h173711C0 , 32'h0C8039B0 , 32'h17B67320 , 32'h06F3EF28 , 32'hFE711190 , 32'hF6E58180 , 32'hD81637C0 , 32'hE0E5E480 , 32'h044D9018 , 32'hE6F8DF20 , 32'hF68D96B0 , 32'hFBA36500 , 32'hF4E9EB70 , 32'h0762D7B0 , 32'h06127FD8} , 
{32'hDDF14080 , 32'hC5447F00 , 32'hDB81C980 , 32'hCFE3BF80 , 32'h37023200 , 32'h09A096C0 , 32'h39D44340 , 32'h104E36C0 , 32'hE5B0B800 , 32'h04859748 , 32'hDC9A5F40 , 32'hF40139B0 , 32'h00CF648F , 32'hF263EAC0 , 32'h1F726FA0 , 32'hE4A06FA0 , 32'hEAD8B7C0 , 32'h1CF8EE00 , 32'hF91EE4D8 , 32'hF3F404F0 , 32'h0CAE9D40 , 32'hF8C47480 , 32'h09F9E940 , 32'h0703FEE0 , 32'h0BDCE8A0 , 32'hE7B76BE0 , 32'hF8006818 , 32'hFCFE1364 , 32'hEB3655E0 , 32'hFF5EB75A , 32'hF666D350 , 32'hEB410AE0 , 32'h05679AE0 , 32'h0A606550 , 32'h03F74CD8 , 32'hD3921C00 , 32'hEB9B2BC0} , 
{32'hDA042E00 , 32'h9CFE3380 , 32'h9413B500 , 32'hCB131E00 , 32'h38F37280 , 32'h02F37EE0 , 32'h54FC7380 , 32'h0A0846A0 , 32'hF99F4B90 , 32'h148E7F00 , 32'hF3D9F070 , 32'h1D116980 , 32'h08322820 , 32'hF0AE0290 , 32'h20F107C0 , 32'hF6B284C0 , 32'h0A7E0E50 , 32'h17043500 , 32'hF48B6080 , 32'hF09F6C70 , 32'h210A4780 , 32'hFF995B38 , 32'hEC873820 , 32'h17D9FEA0 , 32'hFC62490C , 32'hE5471540 , 32'hF48E4F40 , 32'h06B2FBB0 , 32'h018CDC88 , 32'h1C171180 , 32'hDF5B1AC0 , 32'hFC1CDE40 , 32'h0D32ACF0 , 32'hFE2F5B60 , 32'hE72DE5E0 , 32'hF3986080 , 32'hFA167978} , 
{32'hD9B51C00 , 32'hA2706F80 , 32'h8EAAE180 , 32'hC9689D80 , 32'h01992E30 , 32'hE8EC8D80 , 32'h41510000 , 32'hF1997CB0 , 32'hFAD3A570 , 32'h1EFA35C0 , 32'h1B377880 , 32'h1B8B0BC0 , 32'h201475C0 , 32'hEA03F6C0 , 32'hFDEF9740 , 32'h29FF5140 , 32'h1B7A0E80 , 32'hECE7A100 , 32'h1124FAE0 , 32'h040ADDD0 , 32'hF5BC38F0 , 32'h0112DDD8 , 32'hFE0C8CB4 , 32'h066F9FE0 , 32'h0F0EF2C0 , 32'hDFEE2640 , 32'hEC0F92A0 , 32'h01A374DC , 32'hF9EB4190 , 32'h33416A00 , 32'hEF5D58A0 , 32'h1F6E3BA0 , 32'h00942F89 , 32'h187E94E0 , 32'hFB3003C0 , 32'hECE0EF80 , 32'h08AFE9A0} , 
{32'hFFB17A64 , 32'hBE11A500 , 32'hD38BF000 , 32'hC110AD40 , 32'h2D0CD900 , 32'hFA185B80 , 32'h2EBEE940 , 32'h1002B120 , 32'hF82A3AD0 , 32'hF99EE068 , 32'h039C9264 , 32'h3CB35A40 , 32'hFF105A7C , 32'h1091E200 , 32'hCEFAA680 , 32'h51079B80 , 32'h1E589C60 , 32'hF960E360 , 32'h238ACF80 , 32'h007CE91D , 32'hEA14FC00 , 32'h29BBA480 , 32'hF7E7C450 , 32'h1EADCF20 , 32'hF4CCCE90 , 32'h00395A58 , 32'hFD211534 , 32'h191A46E0 , 32'hF2B64DB0 , 32'h0AD72AA0 , 32'hFF4FD47F , 32'hEFA12340 , 32'hE7A81C80 , 32'hEF573C20 , 32'hF86D8F40 , 32'h1728FBC0 , 32'h0A332CD0} , 
{32'h1015EF40 , 32'hC8BC5800 , 32'h18CC4800 , 32'h10475CA0 , 32'h1BC10D00 , 32'hFC9CFC18 , 32'h05323458 , 32'h0755FDB8 , 32'hF6240640 , 32'h155EBCC0 , 32'h08C62D10 , 32'h465DCA00 , 32'hEB3806C0 , 32'h214B6C80 , 32'hDF3C5C80 , 32'h14E98520 , 32'h09ED8CD0 , 32'hDEE01800 , 32'h3BA30D00 , 32'h1300AF20 , 32'hFF3BD1CB , 32'hEF823260 , 32'h00F6E8BE , 32'hFF8C3F4D , 32'h226B65C0 , 32'h02B6B6B0 , 32'h1D34FFC0 , 32'h03DCFBD4 , 32'hCD3DAC00 , 32'hDCF73400 , 32'hE9841140 , 32'h041B4E40 , 32'h09C96A40 , 32'hE840E160 , 32'h16D01120 , 32'hF0C0E030 , 32'h098E1C50} , 
{32'hF62B4D50 , 32'hCC16E380 , 32'hF58DD7E0 , 32'h3CE430C0 , 32'h22F65D00 , 32'h12592820 , 32'hED125D80 , 32'hF607ADE0 , 32'h0398C70C , 32'h0B50F4A0 , 32'h0869B3E0 , 32'h1D569D00 , 32'hF35AEEC0 , 32'hFE1892DC , 32'h01052C40 , 32'h18E98B40 , 32'hF54B1940 , 32'h116DB940 , 32'h225C6DC0 , 32'h152D98A0 , 32'hEEF5BFA0 , 32'h10CF0120 , 32'hEBADF7E0 , 32'h05EA89A8 , 32'h022C5414 , 32'hDB769100 , 32'h066F2958 , 32'h05022998 , 32'hD9E1B2C0 , 32'h0FA8E190 , 32'hD9A942C0 , 32'h061B0B70 , 32'hE7766FA0 , 32'hFCF8FBE0 , 32'hE093DD20 , 32'hE26D44E0 , 32'hFDF2A938} , 
{32'hEC0B91E0 , 32'h0071E2B8 , 32'h00D3276F , 32'h3985B840 , 32'h18D09F80 , 32'h13553480 , 32'hD681A540 , 32'hF018F490 , 32'hEF4C7CC0 , 32'h10A8BAA0 , 32'h0B9F6A50 , 32'h09FF55A0 , 32'h1971FE40 , 32'h046C1868 , 32'hDB5A7E00 , 32'h06F7DB20 , 32'h0BCCC780 , 32'h04FB2230 , 32'h04075908 , 32'hF17B8220 , 32'hEAA66280 , 32'hF2D77420 , 32'hD2003900 , 32'h028E4BE4 , 32'h0632FC48 , 32'hF1FFF020 , 32'hEC931740 , 32'hE3C06880 , 32'h0F528E40 , 32'hFA6899F8 , 32'hF116E310 , 32'hFA53F630 , 32'hE853C840 , 32'h0CDB8A60 , 32'hE60A5740 , 32'h0A5E7F80 , 32'h189FF8C0} , 
{32'hEA459360 , 32'hD7B69940 , 32'h0DC63440 , 32'h3F055E40 , 32'h0E0129F0 , 32'h06C17C60 , 32'hDA1AABC0 , 32'hE95C64A0 , 32'h04E0E630 , 32'h0DC82E20 , 32'h1E3B2A80 , 32'h1D157D00 , 32'h19B66860 , 32'hF517E930 , 32'h0294D324 , 32'hFD0F5A2C , 32'h1288F360 , 32'h1C6BEEE0 , 32'h1EC98D00 , 32'h0CD60C20 , 32'h11ECD320 , 32'hFE786338 , 32'hE5E6C020 , 32'hF27E78D0 , 32'hF7C44270 , 32'hF0C88590 , 32'hEC1623A0 , 32'hF08D34E0 , 32'h19399FA0 , 32'hFF71667B , 32'hF7B6AD30 , 32'hFD0F2854 , 32'hF8861750 , 32'hF44974F0 , 32'hDEB50D40 , 32'h22709740 , 32'h054B5058} , 
{32'h0FC0FAC0 , 32'hF34ABAA0 , 32'h12EB10C0 , 32'h0EA3D600 , 32'h20699200 , 32'hF9742AB8 , 32'hE2552840 , 32'h07DF7160 , 32'h19E0A420 , 32'h1501B7A0 , 32'h12299420 , 32'hF9574520 , 32'h29F49140 , 32'h189C2260 , 32'hFACFCC28 , 32'hD95C9800 , 32'h18A6E2C0 , 32'hDD610440 , 32'h0EEB6060 , 32'hFFA9CE31 , 32'hF2E30F20 , 32'hF1652B90 , 32'h13442B40 , 32'h0082ADB2 , 32'hE0679AA0 , 32'hFE52919C , 32'hF46B5F30 , 32'hEFF14C80 , 32'h1E489E00 , 32'hE091C660 , 32'h05A5AF98 , 32'h07FE3120 , 32'h23063C00 , 32'hFBF4C2F0 , 32'hE93A17E0 , 32'hFC77AE34 , 32'hDEFFD200} , 
{32'h02F3B224 , 32'h15BAD9E0 , 32'h04E95FC8 , 32'hFD9CFDF4 , 32'h1B8B8500 , 32'h049B4820 , 32'hFB9D1F00 , 32'h0FB75E00 , 32'h0E0576D0 , 32'hF15BDB00 , 32'h074E24F8 , 32'hE8DEF220 , 32'hFFB152DF , 32'hF9E3DFE8 , 32'hF3745160 , 32'hFCD628A8 , 32'h221C4540 , 32'h0B328540 , 32'hEEF868C0 , 32'hF0682610 , 32'hF67C24E0 , 32'h016AF954 , 32'hF11C8060 , 32'hE8C0B1C0 , 32'hFF45A9D9 , 32'h149A6900 , 32'hF36B2420 , 32'hF920F538 , 32'h045EC8B8 , 32'hFEFA71A8 , 32'h087BFE70 , 32'h0BE04750 , 32'hF57EC3E0 , 32'hFEB88284 , 32'hE6571D80 , 32'hE6B76F60 , 32'hF4B7EC80} , 
{32'hF0A24430 , 32'h0CFE5640 , 32'hEAD26880 , 32'hDD7B9780 , 32'h09D60A90 , 32'h11DCFAC0 , 32'h08867C60 , 32'h2FF1B500 , 32'h1987C1A0 , 32'hF3EC73E0 , 32'h1993F9C0 , 32'hCEF92AC0 , 32'hF0E62460 , 32'h083EB990 , 32'h0C8F88B0 , 32'hEE81B860 , 32'h2F5FB700 , 32'hFA5601C0 , 32'hF7D8D210 , 32'hD4D16EC0 , 32'hD7AAB540 , 32'hFA1FEBC8 , 32'h15062400 , 32'hED477C80 , 32'hF38FAE70 , 32'h1A71BD80 , 32'hE80EB520 , 32'h1A2431E0 , 32'h0D2ACA40 , 32'h0EB76770 , 32'hD091CE80 , 32'h16655BE0 , 32'hE9781AA0 , 32'hE5B36C40 , 32'hDDB06480 , 32'hE2EDC980 , 32'hDFE4E680} , 
{32'hFE0FEC94 , 32'h0B3877F0 , 32'hF0B979E0 , 32'hFAD30F48 , 32'h07BF1168 , 32'h0B50C880 , 32'h1638F840 , 32'h160C9000 , 32'h00363282 , 32'hF25584C0 , 32'h0A6C0CA0 , 32'hEC5B74C0 , 32'hF887A8D8 , 32'h05317788 , 32'h0417BEB0 , 32'h033596B4 , 32'h16BFB740 , 32'h1136D5E0 , 32'hFA5CBB08 , 32'hFAE50650 , 32'hFA9B2E00 , 32'h04550390 , 32'hFB025428 , 32'hF96E01C0 , 32'h073F7398 , 32'hF35F5860 , 32'h02556174 , 32'h0BA90580 , 32'h02447298 , 32'h0FD09D10 , 32'hE406D560 , 32'h07F74080 , 32'hFD165DF4 , 32'h01F6DA3C , 32'hFAA5EDE0 , 32'hF659A330 , 32'hFF26ED38} , 
{32'h05374388 , 32'h259BC140 , 32'hE752C640 , 32'hF53725D0 , 32'hF9119238 , 32'h283FDA40 , 32'h1DAE57A0 , 32'h406D7980 , 32'h1F424EC0 , 32'hC40C16C0 , 32'h210BF100 , 32'hF5F3CFA0 , 32'hEF5CCE20 , 32'hF44FB310 , 32'h39A76840 , 32'h190DCAC0 , 32'h263E36C0 , 32'h1F320B20 , 32'h0AE245B0 , 32'h21305200 , 32'hFD1569A0 , 32'h10CC65C0 , 32'h177A8C40 , 32'hE37AD820 , 32'h08E769E0 , 32'hF74B6410 , 32'h120D7B40 , 32'hFC4AE964 , 32'hF2258920 , 32'hFD891724 , 32'hF0A38980 , 32'h019F545C , 32'hF24B65A0 , 32'h274C33C0 , 32'h12439000 , 32'h0A5C5D10 , 32'h0D2494F0} , 
{32'hEFDD9D40 , 32'h06E14E00 , 32'hFB2E5458 , 32'hFF3C86D2 , 32'h07373AA8 , 32'hF5B0C6C0 , 32'h0F2F02A0 , 32'h08066C50 , 32'h0F1E6880 , 32'hF445C300 , 32'hEC41FDC0 , 32'h03BA0B40 , 32'h1231B4C0 , 32'h01729F54 , 32'h0F078040 , 32'h11DDC840 , 32'hFDBC2680 , 32'h07624860 , 32'h0BF087F0 , 32'hEC62CD00 , 32'h077ECB30 , 32'h03766DE0 , 32'hF7FACEE0 , 32'hFA91EC70 , 32'h07088CB0 , 32'h06DC2618 , 32'h0391EE08 , 32'hEEB659A0 , 32'hF4C6BC20 , 32'h09352360 , 32'hEDD34B40 , 32'h051CFB38 , 32'h18A92660 , 32'h08C749A0 , 32'h0505FBA8 , 32'hF278C6F0 , 32'hFD36588C} , 
{32'hFCAF28A4 , 32'hF733B520 , 32'hFAB043E0 , 32'h0674EEF8 , 32'hFA647EE8 , 32'hFD1FDDF8 , 32'h00B8B9E3 , 32'h08962000 , 32'h0BB2BC20 , 32'hFADA8220 , 32'h078A2C48 , 32'h0F9E5F20 , 32'hF9AC5538 , 32'h0268A26C , 32'hFED667B0 , 32'hF284BA10 , 32'hFD5B5A98 , 32'h0DE83430 , 32'hF2ECF6B0 , 32'hEFE69220 , 32'hF8B7BA60 , 32'h007D9B9D , 32'h04FFD260 , 32'h0CE310E0 , 32'hFEBD5154 , 32'h04D70248 , 32'h145157E0 , 32'h13FE5800 , 32'h01B1CE4C , 32'h08C45710 , 32'h04B95908 , 32'hF8AC8258 , 32'hEF59F900 , 32'h05DD9938 , 32'hF911AB90 , 32'hFD3FCB84 , 32'hF98C13A0} , 
{32'h00ACEE02 , 32'hFE8E23F8 , 32'hFEA19FF0 , 32'hFF509317 , 32'hFAC84618 , 32'h02C30AB0 , 32'hFC20FF48 , 32'h00BEDA62 , 32'h00ACB286 , 32'hFF734C09 , 32'h01D92D84 , 32'h04E3D568 , 32'hFE795ACC , 32'h024DA9D8 , 32'hFCF1622C , 32'h0038DA42 , 32'hFFCE174A , 32'h0271FE34 , 32'hFF664B07 , 32'hFE6A777C , 32'hFDDD4A3C , 32'hFC371410 , 32'h01479FE0 , 32'h006F17EB , 32'h01AB8C08 , 32'hFAE041A8 , 32'h017EE878 , 32'h014D0DD0 , 32'hFD5BB74C , 32'h04B30F20 , 32'h0510D370 , 32'h0342F700 , 32'hFB8F6600 , 32'hFE201A60 , 32'hFFA89664 , 32'h010C6F54 , 32'h030F65A8} , 
{32'h000378D0 , 32'h00037A36 , 32'hFFFA6F66 , 32'hFFFD1964 , 32'h0000A205 , 32'h0003DFAC , 32'hFFFCDE65 , 32'h0001B1CE , 32'hFFFE9D33 , 32'h0004BA7C , 32'hFFFB9A21 , 32'hFFFD0CA4 , 32'hFFFA1F78 , 32'hFFFD9024 , 32'hFFFF81B8 , 32'h00029355 , 32'hFFFD32C5 , 32'hFFFA1977 , 32'hFFFCD5B1 , 32'h00050257 , 32'h0003C52A , 32'h00006C94 , 32'h00050112 , 32'h0002BA21 , 32'hFFFC41C1 , 32'hFFFFE08D , 32'h000642AD , 32'h00040A43 , 32'h0001B9E1 , 32'h00018801 , 32'h00045C51 , 32'h0003364A , 32'h00052F11 , 32'hFFF88575 , 32'hFFFBC117 , 32'h0005FD35 , 32'h0005C8AC} , 
{32'hFFFEF142 , 32'h0009D9A2 , 32'h0001CFF9 , 32'h000605A5 , 32'hFFFACE4A , 32'hFFF8B63D , 32'hFFFF3797 , 32'hFFFF2123 , 32'hFFFFC985 , 32'hFFFEB75C , 32'h000C3558 , 32'h0001C7F7 , 32'hFFF9A026 , 32'hFFFFAC48 , 32'h0009FF2E , 32'h00001777 , 32'h00043972 , 32'hFFFAA482 , 32'h00092B73 , 32'hFFFE9C8D , 32'h0003FC24 , 32'h000AE987 , 32'hFFFAC798 , 32'h0008F8AA , 32'h0004CF18 , 32'h000CA85B , 32'hFFF4F6BA , 32'hFFF7FE4E , 32'h00005223 , 32'h0000B01C , 32'h00047DE0 , 32'h0006BA50 , 32'h0005E479 , 32'h00057F72 , 32'h0007A1AC , 32'hFFF54F2D , 32'h0000345E} , 
{32'h00033D8D , 32'h0000EF42 , 32'hFFFE2FF2 , 32'h00030EB7 , 32'h0001CEC0 , 32'hFFFB9398 , 32'h000584BA , 32'hFFFA2973 , 32'h0002E836 , 32'h0006793F , 32'hFFF90117 , 32'hFFFA531D , 32'hFFFF8598 , 32'hFFFCD22A , 32'h000685AB , 32'h000864D1 , 32'h00051AAD , 32'hFFF5B6FA , 32'hFFEF6F48 , 32'h000026B4 , 32'h00036CD1 , 32'h0000B875 , 32'h00093484 , 32'h000CBC99 , 32'hFFFB1457 , 32'h000775AD , 32'h000120A9 , 32'hFFFE6310 , 32'h00015C7C , 32'hFFFB3FF8 , 32'h00064E37 , 32'h0005F840 , 32'h000584B8 , 32'hFFFC5B39 , 32'h0003AB2C , 32'hFFF4373C , 32'h0006E033} , 
{32'hFFFEB4FC , 32'hFFFD73DC , 32'hFFF97BA4 , 32'hFFFC4FFA , 32'h00019661 , 32'hFFFA94FB , 32'h000C190E , 32'h000AF7CB , 32'hFFFFB288 , 32'h000284EA , 32'h0007079B , 32'h000EC82C , 32'h0001727D , 32'hFFFE20D3 , 32'h000436B3 , 32'hFFFEEAE9 , 32'hFFFDB2CD , 32'h0002D95F , 32'hFFFC7B31 , 32'h00013668 , 32'hFFFFF8C3 , 32'h00045CD6 , 32'h0007ED48 , 32'h0003A267 , 32'h00062B1B , 32'hFFFFAA7B , 32'h0000DEFF , 32'h00004CBA , 32'h0006DB95 , 32'h0006775B , 32'h00095E3B , 32'h00008311 , 32'hFFFE7E6D , 32'h00036816 , 32'hFFFB04FE , 32'hFFFCA46A , 32'h0001286E} , 
{32'h0005195A , 32'h0002B4EA , 32'hFFFD7299 , 32'h0004B3A0 , 32'h0007DF55 , 32'hFFFF1DB5 , 32'h00018EA9 , 32'hFFFD0114 , 32'hFFFFDCC6 , 32'h000433C6 , 32'hFFF8F4C2 , 32'h000A37B2 , 32'hFFF6B3DB , 32'hFFFF6743 , 32'hFFF7C712 , 32'hFFFA4CA2 , 32'h0005201C , 32'h0001E17A , 32'h00002C3E , 32'h000859AF , 32'h0009F628 , 32'hFFFF5851 , 32'h0002A4D1 , 32'hFFFBE8A3 , 32'hFFF8CEEF , 32'h00024201 , 32'hFFFC982F , 32'hFFF8B878 , 32'h0000D315 , 32'hFFFE8568 , 32'h0000F7CB , 32'h000272BD , 32'hFFF81F9C , 32'hFFFECD43 , 32'hFFFBE4D6 , 32'hFFFB9FF2 , 32'hFFFFE2CB} , 
{32'h000201A1 , 32'h00001E6A , 32'h00001006 , 32'hFFF61A15 , 32'h00001C67 , 32'hFFF63F23 , 32'hFFF8E08E , 32'h00007A0B , 32'hFFFF8E91 , 32'hFFFDB227 , 32'h0000345F , 32'hFFF9DEDC , 32'h00018F25 , 32'h0000A02F , 32'hFFFE88B2 , 32'h000BC5C7 , 32'hFFFE91FB , 32'h0008319F , 32'h00060498 , 32'hFFFE3688 , 32'h0005B458 , 32'hFFFD74D0 , 32'h00066AAB , 32'h00024566 , 32'hFFFBC7F1 , 32'h0001B363 , 32'h000168A8 , 32'hFFFF54C2 , 32'h00024289 , 32'hFFFB0361 , 32'hFFFF3DB1 , 32'h00016CF6 , 32'hFFFA557C , 32'h0004065A , 32'hFFFE1398 , 32'h000376F7 , 32'hFFF9176D} , 
{32'h05A3A590 , 32'h0B694240 , 32'hEC967C00 , 32'h0127318C , 32'h0A516B70 , 32'hF0C9F4F0 , 32'hED810C80 , 32'hF62D9990 , 32'h075B9428 , 32'hF8D12518 , 32'hFF2B2A8E , 32'hF40CC660 , 32'h0302B4CC , 32'h0039188C , 32'h0F2AC330 , 32'h04D54070 , 32'h026B93BC , 32'h0B719A50 , 32'hFF99D5FE , 32'h083ACCE0 , 32'h02DD2468 , 32'hFEA4FCD4 , 32'h01A5B2C8 , 32'h07BC8B60 , 32'hFBE65398 , 32'hF8F8A610 , 32'hF88C2420 , 32'h0C2676F0 , 32'hFF44211D , 32'h016D112C , 32'h03D4E5E4 , 32'hFDB45648 , 32'hF616F620 , 32'h0DC58500 , 32'hFFE2CE62 , 32'h09E700F0 , 32'hFEEFD994} , 
{32'hFFA50DEF , 32'h0003662F , 32'hFF3A50AB , 32'hFFD6C8B1 , 32'hFF232FF2 , 32'hFFD00945 , 32'h001D1CA9 , 32'h0031457F , 32'hFFAF81D0 , 32'h003284B6 , 32'h00669967 , 32'hFF762C44 , 32'h0079A5A7 , 32'h000162A1 , 32'hFFA13F8B , 32'h000D55D3 , 32'h004D669B , 32'hFF22EA52 , 32'hFF8FAC2F , 32'h003B37A9 , 32'h002663FD , 32'h004581D9 , 32'hFFE56F77 , 32'h00BD297E , 32'hFF2844DE , 32'hFFAEC5E2 , 32'hFFC32F43 , 32'h0002107D , 32'hFF591A91 , 32'hFFCA8093 , 32'hFFBB6D73 , 32'hFFA6EC00 , 32'hFFD5B398 , 32'hFFD67924 , 32'h007C4641 , 32'hFFAAAD3C , 32'h00ECA2BD} , 
{32'h083C2460 , 32'h03BE7134 , 32'hE3472AC0 , 32'h11B002E0 , 32'h0367EE84 , 32'hECFAF4E0 , 32'hF7D63E00 , 32'h14D9D0A0 , 32'h1046FA20 , 32'h00126BFC , 32'hE77E98E0 , 32'hEC0451C0 , 32'hF1EC8570 , 32'hFB23A7A0 , 32'hF87D6408 , 32'h0E749A60 , 32'hFD989D40 , 32'h14C58160 , 32'h083E64F0 , 32'h0E6BA750 , 32'hE9A671C0 , 32'h06E61F98 , 32'hEA10A820 , 32'h19D866E0 , 32'hFA3FFB60 , 32'hFB2D2888 , 32'hFB9BFE38 , 32'h0DF85DE0 , 32'h04AA7E10 , 32'h02BC915C , 32'h0F5BDA50 , 32'hFB018ED0 , 32'hF132FE40 , 32'h0904D880 , 32'h05EA22C0 , 32'h068E2948 , 32'h11DE4CE0} , 
{32'hFA35CD58 , 32'hF873E2E8 , 32'hF5A3D320 , 32'h017ED350 , 32'h0E99C2C0 , 32'hFF79A3C8 , 32'hF5B6A1B0 , 32'hFFC01290 , 32'hFCCCC7F4 , 32'hFC76932C , 32'h01F372D4 , 32'hF6E8B3D0 , 32'hFDD9413C , 32'h052F7FA0 , 32'h0E8EA1C0 , 32'hF2F60860 , 32'hF87A9E68 , 32'hF696F910 , 32'hFDBBD394 , 32'h087E13D0 , 32'hFA887308 , 32'hF7FA0270 , 32'h03605FA4 , 32'hFDAE1A14 , 32'h03D585E0 , 32'h09284D20 , 32'h073FCF18 , 32'hF4692340 , 32'hFDB99DDC , 32'hFB229AA8 , 32'h0A1D2D90 , 32'hFBA33E88 , 32'h0192EB08 , 32'hF53860C0 , 32'h0D6D3340 , 32'hFC07BFD4 , 32'h04BF68A0} , 
{32'h04E8AB40 , 32'h021A2150 , 32'hC45028C0 , 32'hF46FA390 , 32'h22E95440 , 32'hEDD454A0 , 32'hCBF1B740 , 32'hFEA12A74 , 32'hF7637520 , 32'hEBD99A80 , 32'hF3646AA0 , 32'hE62F68C0 , 32'h049D7130 , 32'h08016260 , 32'h1DC23FA0 , 32'hEC4E00C0 , 32'hF92900D0 , 32'h1080CBA0 , 32'hFE7DD364 , 32'h0FEB0F40 , 32'hFE1ED9F0 , 32'hE73663E0 , 32'hFEF1C5DC , 32'hFB4F0890 , 32'h16FB2BC0 , 32'h0C64DCD0 , 32'h1C169660 , 32'hF7F616A0 , 32'hFE56D7AC , 32'hF6A7A250 , 32'h02BB3114 , 32'hFAD76608 , 32'h06D636B8 , 32'hFFE683AD , 32'h13F14EC0 , 32'hFFF83E0C , 32'h1387B740} , 
{32'h0C9741F0 , 32'hFDF4C2C0 , 32'hA3381600 , 32'hDD143440 , 32'h406DC100 , 32'hD334F900 , 32'hE153D760 , 32'hF950A2B8 , 32'hF2CBD6E0 , 32'hDC784500 , 32'h0860E890 , 32'hD4BB7A80 , 32'h1CA4AE00 , 32'hE24B61E0 , 32'h2C64C680 , 32'hD86C4D00 , 32'hD66335C0 , 32'h1E1A7F00 , 32'hF63FF620 , 32'hF21D0010 , 32'h020ABFF0 , 32'hFABBF958 , 32'hFC8889A8 , 32'hE7756640 , 32'h20A03F40 , 32'hE953A700 , 32'h141AC540 , 32'hE34C44E0 , 32'hE9946140 , 32'hE9B4C760 , 32'hFB15ECD8 , 32'h0C53AEF0 , 32'hECB87020 , 32'hE7B4E480 , 32'h162E7680 , 32'h0465CD90 , 32'h10522A80} , 
{32'hF355BCE0 , 32'hF38C5420 , 32'h8E8B4180 , 32'hE61F7920 , 32'h31827D40 , 32'hC3628C00 , 32'hDAB75340 , 32'hF4C50CA0 , 32'h013D0204 , 32'hE4DAE980 , 32'h1655DC40 , 32'hE66FA3C0 , 32'h03DC3FD8 , 32'hFD91DED0 , 32'h121758C0 , 32'hE6D3B080 , 32'hF089DE40 , 32'h02AE9224 , 32'hF195BFF0 , 32'h1C268280 , 32'h05A69D48 , 32'hDBBB7C40 , 32'h0BC58A50 , 32'hF2A70350 , 32'h29CF8F80 , 32'h0CFD0FC0 , 32'hFE0FDB4C , 32'hE9B39580 , 32'h15831B80 , 32'hE7D34260 , 32'h08DB7120 , 32'hFCB152F8 , 32'hF951B130 , 32'h089DB940 , 32'h1C52CA20 , 32'hEAF4B920 , 32'h107C7D60} , 
{32'hD543F940 , 32'hE8DBB6E0 , 32'h7FFFFFFF , 32'hD5D62A80 , 32'h4139FF00 , 32'hB8E6BB00 , 32'hEF92E980 , 32'h05F3C900 , 32'h12CBDB80 , 32'hF0E0B250 , 32'h46DEE780 , 32'h141DEA60 , 32'hEEB8E9C0 , 32'h15924320 , 32'hF4B7BF90 , 32'hF65BF1E0 , 32'hE750CF80 , 32'hDCCA7380 , 32'hEC92C620 , 32'h392D9DC0 , 32'h041FE188 , 32'hEDF2B3A0 , 32'hFC88B83C , 32'hE7C4CC60 , 32'h1E2420E0 , 32'h0DB78380 , 32'h157C3A20 , 32'hC71992C0 , 32'h17BF7080 , 32'hF2B5DDE0 , 32'h0809D2A0 , 32'h0F0FC0F0 , 32'h0512AFD8 , 32'hCCB059C0 , 32'hF6370710 , 32'hEDB863A0 , 32'hF1125970} , 
{32'hF9AB4C48 , 32'hEBC63780 , 32'h7FFFFFFF , 32'hD3B1E040 , 32'h23575C40 , 32'hBFE67E80 , 32'hEF6A27C0 , 32'h11AC9C00 , 32'h2D4DA600 , 32'hF65FDCA0 , 32'h39AAD580 , 32'h3775EF40 , 32'hF5A26B60 , 32'h01789C20 , 32'hF65D26A0 , 32'h0B3E9580 , 32'hF90D9DE0 , 32'hD7C04F00 , 32'hEE777620 , 32'h0E367CC0 , 32'h232181C0 , 32'h0ED3DB50 , 32'hFF9B60D9 , 32'h0827E2E0 , 32'h03277438 , 32'h1BDB0680 , 32'h09889800 , 32'h090C2D90 , 32'h13DFD020 , 32'h0D513130 , 32'h002634BC , 32'h08D15E00 , 32'h1278EF80 , 32'h03C14F00 , 32'hFECA11F4 , 32'h030A0E6C , 32'hF3186E60} , 
{32'hFFB62381 , 32'h075F4B60 , 32'hDB617240 , 32'hEAFC21C0 , 32'h39AA9B00 , 32'hF1C5BB90 , 32'h0D3FD3C0 , 32'hD72B2FC0 , 32'hFCF6B75C , 32'hEA3DEBA0 , 32'h3E0D0180 , 32'h261D7E40 , 32'h04903DF8 , 32'h09824D50 , 32'hFD091530 , 32'h201ECA00 , 32'h08A07EA0 , 32'hE71A4020 , 32'hF6C2C370 , 32'hF5DC9130 , 32'h2BCA3440 , 32'h35A37880 , 32'h060C9FD0 , 32'h1479EC20 , 32'hF5767230 , 32'hDBDFABC0 , 32'h02FF20E4 , 32'h168844E0 , 32'hFA2D8280 , 32'h1A1D8180 , 32'hF6B332A0 , 32'h0DF07150 , 32'h02603390 , 32'hFB7AB988 , 32'hE58E5B80 , 32'h071F3300 , 32'h06F577E8} , 
{32'hF456BE20 , 32'hEED00700 , 32'hF42443C0 , 32'h03F8B950 , 32'h2B51CF40 , 32'h03246460 , 32'hF8F34CB8 , 32'hFC915118 , 32'h0E832CE0 , 32'hF9D45830 , 32'hF38D9B90 , 32'h2DC71D40 , 32'hE1D4B0A0 , 32'h20508CC0 , 32'hE5D24600 , 32'h2300B140 , 32'hF8795E90 , 32'hE4877060 , 32'h1C096720 , 32'h0B5601A0 , 32'hFA00DFD0 , 32'h0D806090 , 32'h07A43248 , 32'h154FD080 , 32'hE6EBD100 , 32'hDE223FC0 , 32'hF9BEF730 , 32'h10E27E20 , 32'hDE618200 , 32'h01DBD304 , 32'hED999140 , 32'h19088BA0 , 32'hF48AB990 , 32'hF9224098 , 32'hE04C6AE0 , 32'hF09EBDC0 , 32'hFAC4A8F8} , 
{32'hE9CD37C0 , 32'hDB79C300 , 32'hEA2421C0 , 32'h429B0600 , 32'h3DE60CC0 , 32'h1AE75D80 , 32'hE81E94C0 , 32'hFBC940A0 , 32'hFBA88500 , 32'h0F66A4A0 , 32'h1400C420 , 32'h4448DC80 , 32'h0178A320 , 32'hF76AA1C0 , 32'hDBF62F40 , 32'h0DB03640 , 32'hFBBFBCE0 , 32'h2EF66140 , 32'hF0880510 , 32'h0E6450A0 , 32'hFD76E57C , 32'h045C30B0 , 32'hC62CB680 , 32'h047140D8 , 32'hF5E12A40 , 32'hF08CE700 , 32'h17CE6F40 , 32'hE00D1A60 , 32'hDA15B980 , 32'hED6ADD60 , 32'h110030A0 , 32'hE0FFA720 , 32'hFE4EFFD8 , 32'h13A8A6C0 , 32'hF0F4C820 , 32'hE075BB60 , 32'h1FC69220} , 
{32'hDE93CCC0 , 32'hDFB9A5C0 , 32'h030134D4 , 32'h5ED8A080 , 32'h1DF85D40 , 32'h0D3E1090 , 32'hD2F2B580 , 32'hE04CDCA0 , 32'hFA0E7738 , 32'h01ECE20C , 32'h1D29A600 , 32'h1AFCD620 , 32'h05882798 , 32'hF9432678 , 32'hD2614880 , 32'h0378FDC8 , 32'h319D9640 , 32'h60C9DC80 , 32'hFD433FA8 , 32'h13226BE0 , 32'hE5D7B160 , 32'h1B8D4080 , 32'hC13A3780 , 32'hECF7CD80 , 32'hEFD10100 , 32'h0FD2A0E0 , 32'hF4BA71A0 , 32'hDAD18D00 , 32'hECCAD440 , 32'hF4E182A0 , 32'hFC465308 , 32'hFD64A774 , 32'hF35B42B0 , 32'hFE8367B0 , 32'h03C8C504 , 32'hDDC72180 , 32'hFCCAA524} , 
{32'hFADA73D8 , 32'h0C70C970 , 32'h08906D50 , 32'h13711A40 , 32'hFFDC18D9 , 32'hF8484008 , 32'hFBA70310 , 32'h01D9D14C , 32'h08E52830 , 32'hFC3C0F00 , 32'h1464F240 , 32'h01EF61C4 , 32'hEE4C4340 , 32'h1F0BAA60 , 32'h06B304F8 , 32'hE533C6A0 , 32'h05911E30 , 32'h1AE4D720 , 32'h210DBEC0 , 32'hED1F75C0 , 32'h0D7549D0 , 32'hEC0F1F00 , 32'hE8EF0940 , 32'hFAE0A598 , 32'hD5D8F500 , 32'hF70AF0C0 , 32'hF9E5FF70 , 32'hEB60DC80 , 32'hF2E548F0 , 32'hFAF1B558 , 32'h0693D6D0 , 32'h17337480 , 32'hFF2D2741 , 32'h02A069F4 , 32'h07AA7DD0 , 32'hF1C37850 , 32'hFA4BDDB0} , 
{32'hFF60CB5E , 32'hF7167E40 , 32'hF23DB6E0 , 32'hFB54BAD0 , 32'h0F86FB00 , 32'hF6AB0470 , 32'h01368E00 , 32'h0C331D10 , 32'h14E950C0 , 32'h0D9F7EC0 , 32'h1D9124A0 , 32'h034E2370 , 32'hF903FB10 , 32'h01EB9018 , 32'hFAB4E8A8 , 32'hCF693AC0 , 32'h12BF4B60 , 32'h143C3B40 , 32'hE4AA9A60 , 32'hE65952A0 , 32'h062C8680 , 32'hD41D4F00 , 32'hDD0E7D80 , 32'h2359F3C0 , 32'hE7DA5500 , 32'hFCD8E810 , 32'h0D66E000 , 32'hFDBE1868 , 32'h22CB8C00 , 32'h0CC26900 , 32'h133CAB20 , 32'h11DDC500 , 32'hFFF5D733 , 32'hEDC1B0A0 , 32'hF222E370 , 32'h078A94B0 , 32'h04A9C4B8} , 
{32'hFFEC7CB7 , 32'h092B05F0 , 32'hED6EF1E0 , 32'hF1E76450 , 32'h078DDCA8 , 32'h07092538 , 32'h09F3BC00 , 32'h18EE8400 , 32'h10928BC0 , 32'hF9D44738 , 32'h1D8BAC60 , 32'hF0703760 , 32'hFC284144 , 32'h053A84E0 , 32'hFA97CB08 , 32'hF2FAB9C0 , 32'h16A33560 , 32'h02535C9C , 32'h079E9320 , 32'hF03A81B0 , 32'h04B86168 , 32'hFF5AA1A2 , 32'hFB9DBA98 , 32'hFD404C44 , 32'hF5C65D50 , 32'h02F921C4 , 32'hF711BCE0 , 32'h02053C78 , 32'h14518AE0 , 32'h104E4720 , 32'hFB96FD60 , 32'h0BD51250 , 32'h0424E4A0 , 32'hE9212EE0 , 32'hEB469CE0 , 32'h029DC840 , 32'hFB7FD738} , 
{32'hFEA04D50 , 32'h0B55BB90 , 32'hF9885CA8 , 32'h02473588 , 32'hFC1AAE68 , 32'h052ED488 , 32'h06E16AE8 , 32'h071BCB00 , 32'h0809AF80 , 32'h0031D6F3 , 32'h0C8FB2E0 , 32'h0790D808 , 32'hF7176DD0 , 32'hFF9546AB , 32'h004A02BD , 32'h0D3077C0 , 32'h102F9820 , 32'hFB2B39C8 , 32'hFFE1D159 , 32'h035A2FF0 , 32'hFE7C4D58 , 32'h0A428D70 , 32'h01EB49BC , 32'h06C1CA90 , 32'hFF3D5790 , 32'hF3790510 , 32'hFC9E7BC0 , 32'hFF13EDE8 , 32'hFD9D3E28 , 32'hFC190248 , 32'h074E8040 , 32'hFBF38D88 , 32'h106C4AE0 , 32'hF7BF2B20 , 32'hFCF120D0 , 32'h0CA1CBF0 , 32'hFE85D0E0} , 
{32'h0DB64450 , 32'h18D225E0 , 32'hFC04C0D8 , 32'h03443A68 , 32'h0FDEE100 , 32'h0ED3DBB0 , 32'h20B30840 , 32'h0E02EC30 , 32'h07DD9318 , 32'hF25EC1C0 , 32'h033C5110 , 32'h0FD14C30 , 32'hF41605F0 , 32'hF7F0A0F0 , 32'h107B76E0 , 32'hFB531AD0 , 32'h03236A08 , 32'h04127318 , 32'hF80EA538 , 32'h0B319250 , 32'hFC46D504 , 32'h05DD39D0 , 32'h02E53134 , 32'hF1498350 , 32'h093B8720 , 32'hFBD240B8 , 32'h0499E858 , 32'h07FE2980 , 32'hFE77A670 , 32'h0171AE0C , 32'hEA916B40 , 32'h11E40840 , 32'hEC259CE0 , 32'h0BF64680 , 32'h064A11B8 , 32'h0AF6E9E0 , 32'h2075B740} , 
{32'hF693C7F0 , 32'h19554760 , 32'hF067DF80 , 32'hF791F580 , 32'hF2654D30 , 32'h1CA58800 , 32'h19AF8980 , 32'h122729E0 , 32'h04CA7CD8 , 32'hE9E81CA0 , 32'h1D557640 , 32'h0EDCE180 , 32'hF69D1D10 , 32'h06C38488 , 32'h22572900 , 32'h0835C460 , 32'h1FFEB300 , 32'h1BA25FE0 , 32'h035F3DC0 , 32'h248F1180 , 32'h009A87DF , 32'hF7438040 , 32'h05593398 , 32'h098770C0 , 32'h09B802E0 , 32'hF30A58A0 , 32'h1BE9C4E0 , 32'hFBCA9BC0 , 32'hE3E5B160 , 32'hF6DE4340 , 32'h06895908 , 32'h135B9E40 , 32'hFEB8D390 , 32'hFD5B0D70 , 32'hFB29B208 , 32'h05C3A558 , 32'h19FE5720} , 
{32'hFA8F5E48 , 32'h19DE9680 , 32'h0A50FAB0 , 32'hFA1AD150 , 32'h084F2D70 , 32'hFED7D7D8 , 32'hFDE4A024 , 32'h160156C0 , 32'h088F8230 , 32'hF003B220 , 32'hE7596A60 , 32'h0BBE0660 , 32'h02797FA4 , 32'h017F3B68 , 32'h14352180 , 32'h14DA4A80 , 32'hFB324860 , 32'h0691DA80 , 32'h08BA0550 , 32'hF904FB68 , 32'h13F3DD60 , 32'h04C5D750 , 32'hFE270D94 , 32'hF1258E00 , 32'h0FA796A0 , 32'h044DEFE8 , 32'hF185F9B0 , 32'hE3C93180 , 32'h110D39E0 , 32'h01DA07B8 , 32'hF38CC2B0 , 32'h0A591C90 , 32'h091DC7E0 , 32'h022E1090 , 32'hFED54048 , 32'h03DF7B38 , 32'hF6C9F4B0} , 
{32'hF822D2C0 , 32'h0884C4B0 , 32'h004B5715 , 32'hFE8C2568 , 32'hF59C33C0 , 32'hEDB876C0 , 32'h08455620 , 32'h08174900 , 32'hFA26F9E0 , 32'hEBB1F980 , 32'h092804F0 , 32'h033E95CC , 32'hC8944B80 , 32'h4A2FF200 , 32'h110FB980 , 32'h0CBB2930 , 32'hCDBBD480 , 32'h028913D4 , 32'h3645C4C0 , 32'hD79CD980 , 32'hFBB53E80 , 32'hFB447350 , 32'hD434B0C0 , 32'h12650C80 , 32'hF54821E0 , 32'h025A3D44 , 32'hECD64C60 , 32'h00523BC7 , 32'h033DF21C , 32'hFCB5F470 , 32'hF1F31070 , 32'hE429DA20 , 32'hE8E92620 , 32'h015F3B64 , 32'h0C39DB60 , 32'h0C2664D0 , 32'h1456C380} , 
{32'hFFFF61A6 , 32'hFFFFCF3A , 32'hFFFF06AF , 32'hFFFCEFA2 , 32'h0000637C , 32'h0006F7CE , 32'h00030855 , 32'h0002CE93 , 32'h00048734 , 32'h0004556E , 32'h00007EA1 , 32'h0004ADE9 , 32'h00003EB8 , 32'h00002066 , 32'hFFFF0B09 , 32'h0001C8A8 , 32'hFFF8ED5B , 32'hFFFFC022 , 32'h00022EFA , 32'hFFFEE642 , 32'h0000C0BD , 32'h0004829A , 32'hFFFFF02D , 32'hFFFF3046 , 32'hFFFEF1BF , 32'hFFFCA218 , 32'h0005F138 , 32'hFFF8D0CF , 32'hFFFAE114 , 32'hFFFAB9D0 , 32'h00009E0F , 32'hFFFDA720 , 32'h0005EA4D , 32'hFFFD20BB , 32'h0001961E , 32'hFFFF7CF6 , 32'h00033E9B} , 
{32'hFFFECF4F , 32'h0000C08B , 32'h0004D243 , 32'h0000FE1C , 32'hFFFD650E , 32'hFFF8DA89 , 32'hFFFF920E , 32'hFFFF4E0A , 32'h0005FB73 , 32'hFFFB963A , 32'h00043A2D , 32'h0004D830 , 32'hFFFEADE7 , 32'hFFFA25AA , 32'h0003B6C5 , 32'h0000E890 , 32'hFFFD84F9 , 32'h00024DD7 , 32'h000428D4 , 32'h00009874 , 32'hFFFF60F8 , 32'hFFF8FBE8 , 32'h00043928 , 32'h0004B7EC , 32'hFFFF1EC4 , 32'h00044474 , 32'h0001EBAA , 32'hFFFEAAB6 , 32'h0000F889 , 32'h00018E02 , 32'hFFFB319B , 32'h000281B0 , 32'h0000FAE7 , 32'hFFFEE3F5 , 32'hFFFFAD52 , 32'hFFFEF307 , 32'hFFFF137E} , 
{32'h0002918B , 32'hFFFE250D , 32'hFFFF8479 , 32'h0004E4C9 , 32'h0003D526 , 32'hFFFE595C , 32'hFFF77D01 , 32'h0005F8B1 , 32'hFFFAA84C , 32'h0003EF62 , 32'hFFF84AC7 , 32'h0001136F , 32'hFFF895B2 , 32'hFFF776F5 , 32'h0004C2F8 , 32'h0004B6A1 , 32'h000463D2 , 32'hFFFE433E , 32'h00073279 , 32'h00006576 , 32'hFFFD1C51 , 32'h00012173 , 32'h00002575 , 32'h00030461 , 32'h0001DC77 , 32'h0003CD82 , 32'hFFFF236A , 32'hFFFCFE84 , 32'h0004BD1C , 32'h0003CDE6 , 32'hFFF67C7B , 32'hFFFECF27 , 32'h00007482 , 32'hFFFD186B , 32'hFFFF296F , 32'h00056EE6 , 32'hFFFED370} , 
{32'h000242D3 , 32'hFFFFCB7C , 32'hFFFF5891 , 32'h000A4C28 , 32'h000943B5 , 32'hFFFDED2A , 32'hFFF56591 , 32'hFFFE3C3E , 32'hFFFEFE85 , 32'hFFFEE9C2 , 32'h0001ADF3 , 32'hFFFE9F72 , 32'hFFFAD945 , 32'hFFF9D2C2 , 32'hFFFE9EF1 , 32'hFFFCDAB6 , 32'hFFFB6BDD , 32'h00061F5F , 32'h00008C08 , 32'hFFFFDF17 , 32'h0003E915 , 32'h0007269B , 32'hFFFC415A , 32'hFFF56D53 , 32'hFFFDB038 , 32'hFFFD426A , 32'h0000E310 , 32'hFFFED768 , 32'hFFFC4A8F , 32'hFFF9A33D , 32'hFFFB599C , 32'hFFFC9F4F , 32'h000035DC , 32'hFFF72D56 , 32'hFFFA1713 , 32'hFFFE9FD0 , 32'hFFF57B8F} , 
{32'hFFFEBC68 , 32'hFFFF06D4 , 32'hFFF7C1DD , 32'h00015E58 , 32'h0002ADA6 , 32'h000349B4 , 32'h000279EE , 32'hFFF6BCCD , 32'h0006CBE8 , 32'hFFFCDB04 , 32'h0005E3EE , 32'hFFFBE2DB , 32'h00038D6B , 32'h000BE982 , 32'h00003BD6 , 32'h00009F26 , 32'hFFF6CB1B , 32'h000026A5 , 32'hFFF99E5E , 32'hFFFECCCE , 32'hFFFCA358 , 32'hFFF67743 , 32'hFFF62688 , 32'hFFFD3012 , 32'h0003AF1A , 32'hFFFE5DF4 , 32'hFFF5BD06 , 32'h0002D57B , 32'h000683E3 , 32'h000042A1 , 32'hFFF1899B , 32'hFFFE87CB , 32'hFFFBB003 , 32'hFFF6C843 , 32'hFFFFFD66 , 32'h0005F63F , 32'h0005A44A} , 
{32'h0006ED94 , 32'hFFFF5450 , 32'hFFFE3673 , 32'h00032CC7 , 32'hFFFB29A8 , 32'h00059F99 , 32'h0004AD9D , 32'hFFFFD073 , 32'hFFFE81D3 , 32'hFFF9AC3E , 32'h0009F9D6 , 32'hFFFC376F , 32'h0000E4D6 , 32'hFFFBC6DC , 32'h0002E917 , 32'h00043E6C , 32'hFFFE944C , 32'hFFFF0226 , 32'h00002285 , 32'hFFFC3696 , 32'hFFFAF082 , 32'hFFFDD433 , 32'hFFF627F9 , 32'hFFFDBA1E , 32'h00000A03 , 32'h0006331B , 32'h000623CD , 32'hFFFB3A19 , 32'hFFFDFB8E , 32'h0002170C , 32'h0004C6A5 , 32'h00003A43 , 32'hFFFD831E , 32'h0003B2FE , 32'hFFFC136D , 32'hFFF817C5 , 32'hFFFE37FB} , 
{32'h0004F5FB , 32'hFFF7BF62 , 32'hFFFA9B1D , 32'hFFFAEB2B , 32'h00054635 , 32'hFFFC0922 , 32'h000005D2 , 32'hFFF6B409 , 32'h00037141 , 32'h000180B8 , 32'h000366AA , 32'h0004E522 , 32'h00067F93 , 32'hFFFCB4D7 , 32'h000647C4 , 32'h000604CD , 32'hFFFE831D , 32'hFFFCF487 , 32'h00023E23 , 32'h00076EA6 , 32'h0007E7F8 , 32'hFFFC13E8 , 32'h0001548D , 32'hFFFE7B8C , 32'h00061C2E , 32'h00041705 , 32'h0003A642 , 32'h00027DFB , 32'hFFFB3A95 , 32'hFFFB3FE5 , 32'h000093E5 , 32'hFFF73D9B , 32'h000005E3 , 32'hFFFDFB52 , 32'hFFFE475E , 32'h0001028F , 32'h000710E7} , 
{32'h00059E03 , 32'h0000CA3A , 32'h0006FAFA , 32'hFFFF2CFD , 32'h00007D94 , 32'h00045984 , 32'hFFFB2BEE , 32'h000107F2 , 32'h0003500C , 32'hFFFD45C4 , 32'h0008AC86 , 32'hFFFCF948 , 32'hFFFFEA83 , 32'hFFFC8FDF , 32'h00036FB6 , 32'h000486E3 , 32'h00049F94 , 32'hFFFE18EE , 32'hFFFF38FA , 32'hFFFE2DB9 , 32'hFFFC4602 , 32'h000296BF , 32'hFFFDC1E6 , 32'hFFFCBC30 , 32'hFFFF28C4 , 32'h0001E3AE , 32'hFFF75F65 , 32'hFFFDAA2B , 32'h0003B9D4 , 32'hFFFEC061 , 32'h00007334 , 32'h0007B210 , 32'hFFF9AB96 , 32'hFFF7D7EB , 32'hFFFDD340 , 32'h0000532F , 32'hFFFFDD0B} , 
{32'h0065C008 , 32'h012D74E4 , 32'h00914F87 , 32'hFED46FFC , 32'h033A08CC , 32'hFF4343CA , 32'h001372BE , 32'hFF2B1380 , 32'hFE0470B4 , 32'hFF03B148 , 32'h0193E6EC , 32'hFD98EBF4 , 32'h04CEBCE8 , 32'h024FFB3C , 32'hFF2AABE6 , 32'hFEC24644 , 32'hFCF7077C , 32'hFFB0D380 , 32'hFEB1D9DC , 32'h00B54B9E , 32'hF880CC68 , 32'h01A7AC14 , 32'hFF449015 , 32'h03201504 , 32'h00AF838A , 32'hFE7BE840 , 32'h03606DE4 , 32'h00039069 , 32'hFD13CE34 , 32'hFE7353A4 , 32'h00C08525 , 32'h073B4998 , 32'hFE956EF4 , 32'hFE2F6664 , 32'h04C34530 , 32'h07696308 , 32'hFB8C5878} , 
{32'hE81DD380 , 32'h0FD7CD00 , 32'hF767F6C0 , 32'h05E0AED8 , 32'h02231640 , 32'h0C915BA0 , 32'h00209A44 , 32'hFEFCF024 , 32'hF067D5B0 , 32'hF93F7CD8 , 32'h029A8DA4 , 32'hFDAC8308 , 32'hFB6AAAE8 , 32'hE88E3460 , 32'hFB802510 , 32'h036C1440 , 32'hF5BA4620 , 32'h039CA000 , 32'h144BFC80 , 32'hFC7E192C , 32'h0EE3DC50 , 32'hE864A2A0 , 32'hFA5095F0 , 32'hFF2B6502 , 32'hF17A7920 , 32'h01AAB6A0 , 32'h04F82440 , 32'h15F181E0 , 32'hFC505898 , 32'h047AC8A8 , 32'h030C9E40 , 32'h091D0780 , 32'hF6983100 , 32'hF28D3D70 , 32'h040A2E18 , 32'h00A1F54B , 32'hF9B376A8} , 
{32'h1001CFA0 , 32'h209DC700 , 32'h025820BC , 32'hD80AA9C0 , 32'hFF479760 , 32'hE7667FC0 , 32'h0F2F28F0 , 32'hF315AE80 , 32'hF1F71AB0 , 32'h01FBF624 , 32'hF94C2470 , 32'hD65C7940 , 32'hECBCA120 , 32'h2DF08C40 , 32'hFF2FFDAD , 32'h146428C0 , 32'hDC1D8C00 , 32'h06C882E0 , 32'h0CBFC100 , 32'h0E69CE00 , 32'hD32B6240 , 32'hFAAD3510 , 32'hFEFC4C4C , 32'hEBACC560 , 32'h0420D6B8 , 32'hE93268E0 , 32'hE3F11EE0 , 32'h0D6E6570 , 32'h067020B0 , 32'h0F7A58D0 , 32'h186DA2A0 , 32'h1B5E7BE0 , 32'h0C981030 , 32'h04746C60 , 32'h23AAD800 , 32'h01141278 , 32'h1B2CC100} , 
{32'hF81D0FD8 , 32'hF1F18F90 , 32'hEB07DD00 , 32'hE83C0CA0 , 32'h03742974 , 32'h04EF53D0 , 32'h08984740 , 32'h078AE710 , 32'hF66C8370 , 32'hEB96C740 , 32'hFAFB6C88 , 32'hDE417B00 , 32'h18C22520 , 32'h12485020 , 32'hEE74E0C0 , 32'hCCA1BD40 , 32'h00AE3014 , 32'h20A94880 , 32'hFDD6F014 , 32'h1F819480 , 32'hFD42B6F0 , 32'hDE20B800 , 32'hBBD5D780 , 32'hDBDD39C0 , 32'h20CE7600 , 32'h1FBCAD60 , 32'h12D42DE0 , 32'hFCBE8064 , 32'h03CED380 , 32'hD07D8540 , 32'hE8170C20 , 32'h0B641490 , 32'h004065F3 , 32'hFD525DF4 , 32'hDA681740 , 32'h1FA5F400 , 32'hFDA2AD20} , 
{32'hFC8B7518 , 32'hF0BC6CD0 , 32'hCE8B5E80 , 32'hF75EAFB0 , 32'hEC691A00 , 32'hEAA5C4E0 , 32'h0DF55EA0 , 32'h062990D0 , 32'hF68996D0 , 32'h07A83F38 , 32'hFC9480D0 , 32'h06116278 , 32'h1A658980 , 32'h0431F038 , 32'h1E40B400 , 32'hF7425960 , 32'hED12D480 , 32'h1F315020 , 32'hFC99D7AC , 32'hF7F5E5E0 , 32'h052A0458 , 32'hE482D4C0 , 32'hEEDC8D20 , 32'hE7127580 , 32'h02A60E58 , 32'hFE322C34 , 32'hF905C430 , 32'hF00FC510 , 32'h14879060 , 32'hF2E92DA0 , 32'hE916D500 , 32'h145B9A40 , 32'hF9F068F8 , 32'h1FCEDF00 , 32'hFEE240E8 , 32'hE8BE8260 , 32'hFA5BD260} , 
{32'hFE92E470 , 32'h1D60B240 , 32'hCBE55B80 , 32'hF0D507C0 , 32'hF8D24E00 , 32'hDEE895C0 , 32'hEFF5E600 , 32'h276A08C0 , 32'h08E844C0 , 32'hF2099480 , 32'h2C6E1200 , 32'hFD47E8C0 , 32'h01BF5A94 , 32'h015D2414 , 32'hFC5DB44C , 32'hE4468C40 , 32'hDB230100 , 32'h008CB3D5 , 32'hF0109600 , 32'h0A446DF0 , 32'h0C3BAA10 , 32'hEC9CE8A0 , 32'hF74E8D50 , 32'hECBBEB80 , 32'h22C95FC0 , 32'h209E0580 , 32'h00F60FD2 , 32'hDBABACC0 , 32'h09E46720 , 32'h0B30C250 , 32'hFAD4F2F0 , 32'h21D5C3C0 , 32'h2E5DB340 , 32'hF6A864E0 , 32'hF385DF80 , 32'hFDF1DCC8 , 32'h08023F30} , 
{32'hE79752A0 , 32'h02246100 , 32'hEC9F0480 , 32'hEB9D6A80 , 32'h067FA1F8 , 32'hE578C480 , 32'hF9E34E88 , 32'h09E21A10 , 32'h02CCF32C , 32'h0459D440 , 32'h0A677450 , 32'h037DE4FC , 32'h011C8E0C , 32'hFDA83F7C , 32'hE99E04C0 , 32'hEC1B6480 , 32'hF71C7320 , 32'hF56DE7A0 , 32'hF8310858 , 32'hEF4963A0 , 32'h0C597C40 , 32'hFE1FA0CC , 32'hF36BACA0 , 32'hE7DB8B60 , 32'h13DEA140 , 32'h0A162A70 , 32'hF347D5C0 , 32'hFCB2D114 , 32'h00B7E3C8 , 32'hFDF53A80 , 32'h098E1210 , 32'h0632F6C8 , 32'hFE823190 , 32'hF60474B0 , 32'h18B3E4A0 , 32'hF9CC69E8 , 32'h0029EBB9} , 
{32'h08D40240 , 32'h09AAAF00 , 32'hD9C22640 , 32'h0039274B , 32'hED9C2E00 , 32'hC9F68CC0 , 32'hEE526F40 , 32'h04392E40 , 32'h207D7B80 , 32'hE771C760 , 32'h29690EC0 , 32'h1A990F40 , 32'hEEC39D40 , 32'hEB9CD9A0 , 32'hA8C9D100 , 32'h1261EC80 , 32'hCA55DF40 , 32'h07629068 , 32'hF1DAD930 , 32'hFAC29838 , 32'hEF036580 , 32'h154951C0 , 32'h00AB969E , 32'h0911C9C0 , 32'h03CCAC3C , 32'h03CE698C , 32'h277C3140 , 32'hF3F53FA0 , 32'hFFD8D2C7 , 32'hF9EDEC38 , 32'hEF63E3E0 , 32'hFE033EDC , 32'hFBFD18D0 , 32'h0D87F4E0 , 32'hE0E90320 , 32'h02178650 , 32'hD3557440} , 
{32'h03EEF89C , 32'h0E7D27B0 , 32'hE0DD97C0 , 32'hE6F6A700 , 32'h1A608CA0 , 32'hAD9B0980 , 32'hF1826350 , 32'h0F249210 , 32'hFC304100 , 32'hE638BD40 , 32'h2ECCD3C0 , 32'h15AA2D60 , 32'hD2B1F300 , 32'hF33B9A50 , 32'hA6FB9A00 , 32'h3DF44480 , 32'hDFF75AC0 , 32'hF86B6BA0 , 32'hE1B29160 , 32'h08ACCFC0 , 32'h4765D600 , 32'h1CFAFDA0 , 32'h2B8600C0 , 32'hE9C15A00 , 32'hECF0D4C0 , 32'hEEE9DBC0 , 32'h2D4FD080 , 32'hF5FD0730 , 32'h0B5C08C0 , 32'h09D511A0 , 32'h04504908 , 32'hFFF64AED , 32'h0666BD08 , 32'h0D3998D0 , 32'h090D5DE0 , 32'h0D7B4160 , 32'hF8394900} , 
{32'h0590AAD8 , 32'h05BBCA00 , 32'h0CAC5AB0 , 32'h0E1F6D30 , 32'hFAD78330 , 32'hF703DC50 , 32'hF745FB50 , 32'h0DF5D8E0 , 32'h00115CD6 , 32'hDED08DC0 , 32'hFD396BC0 , 32'h1493E040 , 32'hF6789AF0 , 32'h1AF64EE0 , 32'hF5437710 , 32'hFB33DAB8 , 32'hF740B060 , 32'h01345190 , 32'hFC69ABDC , 32'hF0C56BF0 , 32'h04CF6F80 , 32'h0143C940 , 32'hFD8EE4B0 , 32'hF4AF3DD0 , 32'hE28B0A40 , 32'hEBB3E8C0 , 32'h00F7287A , 32'h095DC400 , 32'hF81C3848 , 32'hFBEEC5B8 , 32'hFFABCAF0 , 32'hF33FBDA0 , 32'hF3267730 , 32'h0EE966C0 , 32'h0CEFE4B0 , 32'hF16B4C80 , 32'h00933E26} , 
{32'hF8C77258 , 32'h008E99C8 , 32'hF75369B0 , 32'h27FD0680 , 32'h112AD6A0 , 32'hF3791360 , 32'hEE2F8FE0 , 32'h13A61060 , 32'h01EA881C , 32'hF446C740 , 32'hFDB77448 , 32'h2BCF3B40 , 32'hF56C6270 , 32'h13F9E520 , 32'hB8EB3780 , 32'hFB5BC0B8 , 32'h204AA740 , 32'h24CD80C0 , 32'hE4A633C0 , 32'hF17042E0 , 32'h089C66E0 , 32'hFFD31C8C , 32'hD8A52C40 , 32'h134AB880 , 32'h016E8144 , 32'h029A5578 , 32'h05544C60 , 32'hF8964640 , 32'hD135DA00 , 32'h24C6BD80 , 32'h1FD0AA40 , 32'h0B816B70 , 32'hF61A0B20 , 32'h0BA128D0 , 32'h118A4580 , 32'h02A4BE10 , 32'h1CD56780} , 
{32'hE5B54C00 , 32'h11C5E3C0 , 32'hF47EB570 , 32'h108F4740 , 32'h05564A80 , 32'h1B8524A0 , 32'hE2232A00 , 32'h10A51CE0 , 32'hFF5AE5A9 , 32'h0559C7B8 , 32'h0F8EAED0 , 32'h0F523E40 , 32'hF7A51190 , 32'h1C176D20 , 32'hEE40EA00 , 32'hF96F49B0 , 32'h239C5480 , 32'h0E3B1430 , 32'hEBFB7EA0 , 32'hFF94804D , 32'hE378DEC0 , 32'hE1931780 , 32'hE33622A0 , 32'h25BCCE80 , 32'h02936B14 , 32'h067AB4F0 , 32'h1BC99200 , 32'hF28444F0 , 32'hF49F7530 , 32'hF9FDCDA8 , 32'h1C774080 , 32'hF6625DA0 , 32'h10C502A0 , 32'h1BA6F2A0 , 32'hE7D82DE0 , 32'h01458908 , 32'h0E107770} , 
{32'hFCA70AB8 , 32'h0A350BA0 , 32'hFFB19BDA , 32'h07692520 , 32'h06F2A5F8 , 32'h0152E234 , 32'h00814315 , 32'h0E4AB4C0 , 32'hF9706238 , 32'h079A6EF8 , 32'hFA1A99F8 , 32'h06C3F738 , 32'hF06BE7F0 , 32'h23BC2B00 , 32'hF9D86D90 , 32'h03CE9288 , 32'h14FD7A00 , 32'h09BFF140 , 32'hFBAC39C0 , 32'h1FA3AF80 , 32'hE8D2F820 , 32'hCDC69600 , 32'hE6DEB2A0 , 32'h09DAF020 , 32'hF931F5F0 , 32'h16056240 , 32'hF7285CE0 , 32'hF4B73F50 , 32'hF2D43DA0 , 32'h02413BB8 , 32'h1D620F00 , 32'h0566C350 , 32'h070AA3B8 , 32'h140DAE40 , 32'hEFC51AA0 , 32'hF5775D80 , 32'h00A761EF} , 
{32'h0270C97C , 32'h0E4CEB40 , 32'hF7503440 , 32'hF957E570 , 32'h1319D700 , 32'hFA574B58 , 32'hFA354320 , 32'h0F123C20 , 32'h07B0FB88 , 32'h0BB1AE00 , 32'h1CF73A20 , 32'hFA36DD18 , 32'h0701E998 , 32'h01F1299C , 32'hC91E2640 , 32'hFA4B3A50 , 32'h17D7F760 , 32'hE9F47AC0 , 32'hF9465270 , 32'hEC870B00 , 32'hF16B4DD0 , 32'hF67A0FF0 , 32'hD4E3B3C0 , 32'h129723A0 , 32'hF3981340 , 32'h13A77AA0 , 32'hD65F5780 , 32'hF341B2E0 , 32'h1AD194C0 , 32'h06F24788 , 32'h2A17A1C0 , 32'hF1A16FF0 , 32'h292472C0 , 32'hF3006B80 , 32'hEB7B9060 , 32'h0EB3AD60 , 32'h028A2998} , 
{32'hFE2C4BBC , 32'h16093280 , 32'h0E51D8F0 , 32'hF5ABFD70 , 32'hDF6A21C0 , 32'h04461B50 , 32'h23E77E00 , 32'h36CBB300 , 32'h07ECBA60 , 32'h013D3230 , 32'hFC28DE50 , 32'hDF1D3F40 , 32'hE15C1200 , 32'h22885A80 , 32'hFD2B49E8 , 32'h0DE5BE30 , 32'h3FA17100 , 32'h212F40C0 , 32'hEC84C2C0 , 32'hE88A0AC0 , 32'hE5ED7000 , 32'hDF42CAC0 , 32'h0CC18B80 , 32'hF8384FF8 , 32'hF19EFB80 , 32'h12DD8860 , 32'hCCEF8100 , 32'h27F2A500 , 32'h1131A420 , 32'h394495C0 , 32'hE40005E0 , 32'h08395710 , 32'hD7A81680 , 32'h18286200 , 32'hEB24FF80 , 32'hE7BCB900 , 32'hCC779880} , 
{32'h008E49FF , 32'h193D6240 , 32'hE7A1A020 , 32'hFE779140 , 32'hF02EC320 , 32'h0FB179E0 , 32'h26146C80 , 32'h317A3940 , 32'h1A88D1C0 , 32'hF993BE60 , 32'h2C516E80 , 32'h16FCCD40 , 32'hD3DAB900 , 32'h0D88D620 , 32'h1F8851C0 , 32'h1293F300 , 32'h24547680 , 32'h33215A40 , 32'hF8DE18B0 , 32'h21423300 , 32'h06E6F208 , 32'hE8F00D00 , 32'hF659D0A0 , 32'h08DF45A0 , 32'hF4BB3890 , 32'hDA6A3C80 , 32'h04BDF120 , 32'hF9DBAEE0 , 32'hFF9F404F , 32'hFE38C260 , 32'h099042D0 , 32'h096D64C0 , 32'h13CAC7E0 , 32'hFA27B600 , 32'hE8220DE0 , 32'hECAE53E0 , 32'h1F5B7CA0} , 
{32'h0328F4F0 , 32'h2306A000 , 32'h0238CB6C , 32'h00D2929A , 32'hEA748060 , 32'h13C598C0 , 32'h298F0380 , 32'h34C76780 , 32'h1415A780 , 32'hC5ECBB00 , 32'h1EA2C460 , 32'h018A6128 , 32'hDDD3A940 , 32'h28349100 , 32'h344F7C40 , 32'h1D1E1B60 , 32'h039AB924 , 32'h16816000 , 32'h1E1CBC00 , 32'h03F76A94 , 32'h0968EEF0 , 32'hFE1768FC , 32'h06632DF8 , 32'hE36F0140 , 32'hF1023A50 , 32'hDA38F600 , 32'h0213ABBC , 32'hE9E57A40 , 32'hEEFBA440 , 32'hE5E7D880 , 32'hF71DA2E0 , 32'h08624360 , 32'hF95DE1B8 , 32'h03F99C10 , 32'hFE1620A0 , 32'hEBE05680 , 32'h1A929C60} , 
{32'hE00431C0 , 32'h17BC5C60 , 32'hECF1F840 , 32'h0EDAA8C0 , 32'hF6C18730 , 32'h0C18C170 , 32'h0BABCC00 , 32'h1302B320 , 32'h0369D77C , 32'hEE8782C0 , 32'hF2E4A990 , 32'hEEC3CC00 , 32'hF63F2690 , 32'h1E641D40 , 32'h0E648B10 , 32'h12EF3FE0 , 32'hD1C2F7C0 , 32'h075E39E8 , 32'h167FEEC0 , 32'hE7644FE0 , 32'h0A46B070 , 32'h075BEBC0 , 32'hFF785C4D , 32'h0732A360 , 32'h091849F0 , 32'h0CD4EF20 , 32'hE418E7A0 , 32'hE911B940 , 32'hFC637B78 , 32'h051E6A48 , 32'hFAEE3020 , 32'hEEE79D80 , 32'h05ACF910 , 32'h16592F80 , 32'hF6B945A0 , 32'h1162CBE0 , 32'hFE5961E4} , 
{32'h01C38224 , 32'h0C209ED0 , 32'h0398C844 , 32'h0B403C40 , 32'hFEADF898 , 32'hF86EEAA0 , 32'hFE200E78 , 32'h04E795D0 , 32'h0184534C , 32'hE69D4320 , 32'h096506C0 , 32'hFD20CCE0 , 32'hE0ABDAE0 , 32'h2ECE2F40 , 32'h0A5CA1E0 , 32'hFD56A53C , 32'hF5323BD0 , 32'hFAC7FCE8 , 32'h16292B00 , 32'hF0F0A7A0 , 32'h0FAA6E90 , 32'h067DF338 , 32'hE06FDDA0 , 32'hF991DF40 , 32'hDEEE7580 , 32'hF405A860 , 32'h011F3750 , 32'hFD14C968 , 32'h01FEE634 , 32'hFF12C45D , 32'hF82D76F8 , 32'hF8EE5830 , 32'hFFA68B29 , 32'h00E59051 , 32'hF9DAAC78 , 32'hE2C8AC20 , 32'h083D9120} , 
{32'hED4EE7E0 , 32'h0132F8C4 , 32'h0C8E6FB0 , 32'hF59DCD20 , 32'h02F2C104 , 32'hFDFB85E4 , 32'hEE74F8E0 , 32'h0BE7C500 , 32'h0B05C820 , 32'hEC512460 , 32'h04CC88E0 , 32'h1317D4A0 , 32'hDD71AC00 , 32'h1EFB3700 , 32'h02913018 , 32'hFC5DB3C8 , 32'hF6F74D70 , 32'h06FF82C0 , 32'h07F0ECA0 , 32'hEF7FDDE0 , 32'hF7C571D0 , 32'h00217B73 , 32'hFE3D742C , 32'h006561F1 , 32'hF22783C0 , 32'hF52F3E80 , 32'hF1A55AC0 , 32'h0700D6A0 , 32'h04889AC0 , 32'hF26FE9E0 , 32'hFB22B548 , 32'hFF10CC26 , 32'hF3A29450 , 32'h074141E0 , 32'hFAC86290 , 32'hEC0A55E0 , 32'h0C4BCA40} , 
{32'hE86E29A0 , 32'hF8DFE558 , 32'h06BA2800 , 32'hE8823460 , 32'h0585BE80 , 32'h05AC67B8 , 32'hEEB693E0 , 32'h0992F570 , 32'h0AF1C860 , 32'hFB6583F8 , 32'hFB9C5000 , 32'h0B792A30 , 32'hF7146280 , 32'hFDD15A8C , 32'hF9585588 , 32'h029FF858 , 32'hFD7D2930 , 32'h0ED38010 , 32'hFC015308 , 32'hF5DB25C0 , 32'hF4A57EB0 , 32'h0072E29F , 32'h151191C0 , 32'h1031DD20 , 32'h02689F4C , 32'hFD2D45AC , 32'hF0FA9E60 , 32'h029A6B94 , 32'hFA0BA3F8 , 32'hED44E740 , 32'hF75CCEA0 , 32'h0F2532E0 , 32'hF68F5240 , 32'h02E462C0 , 32'hF815B1A8 , 32'h02B1627C , 32'h061FD390} , 
{32'h00039EF6 , 32'h000278D4 , 32'hFFF796E1 , 32'h00044A49 , 32'hFFFE42E2 , 32'hFFFA1C76 , 32'hFFFD6F53 , 32'h0004124E , 32'h000534ED , 32'h0005FF88 , 32'hFFFC8048 , 32'h00043B8C , 32'h0004513B , 32'h00000D5B , 32'hFFF7FF8D , 32'hFFFC7420 , 32'hFFFCD3CC , 32'h000166F7 , 32'hFFFF02C3 , 32'hFFFE8459 , 32'h00021D5F , 32'h000393CE , 32'h00095D4D , 32'hFFFB567F , 32'hFFFCE077 , 32'hFFFF58FE , 32'hFFFFEE1E , 32'hFFFB0E2D , 32'h0000269E , 32'h00013381 , 32'hFFF7DDB0 , 32'h000414CA , 32'hFFFFFCD9 , 32'h0002BB07 , 32'h0004ACB8 , 32'hFFFE4F5F , 32'hFFF8A644} , 
{32'h00032180 , 32'h0000E3B3 , 32'h00057855 , 32'hFFFCF1DD , 32'hFFFB44DC , 32'hFFFC2812 , 32'hFFFC0031 , 32'hFFFEACD4 , 32'hFFFD9909 , 32'hFFFDD1F3 , 32'h000065B9 , 32'hFFFEFA35 , 32'h00051641 , 32'h0003B9C3 , 32'h00093381 , 32'hFFFA84ED , 32'hFFFC2046 , 32'h00040954 , 32'h00003C8F , 32'h0001FDF5 , 32'h0007F179 , 32'h00031AB6 , 32'h0002AAEC , 32'h00028750 , 32'hFFFAAD13 , 32'hFFFBFF08 , 32'hFFF70CFA , 32'h000A90F1 , 32'hFFFA339E , 32'hFFFE7C8B , 32'h000383F5 , 32'h00026919 , 32'h0005E87F , 32'hFFFF9228 , 32'h0001D71C , 32'hFFFE5EDD , 32'hFFF8D501} , 
{32'hFFFFB0D2 , 32'hFFFA53EB , 32'h00076E50 , 32'hFFFE08BD , 32'h0000F36A , 32'hFFFD7316 , 32'h0009BD81 , 32'hFFFF276B , 32'h00009896 , 32'hFFFC51FD , 32'h0009345B , 32'hFFF9497D , 32'hFFFD3DE6 , 32'h0003EDA2 , 32'h0005C87C , 32'hFFF5DC57 , 32'h00016559 , 32'hFFFED70C , 32'h0006CB0C , 32'h0000FA11 , 32'h00009B9F , 32'hFFFFEC6A , 32'hFFF94B95 , 32'hFFFA8E52 , 32'h0002B00B , 32'h00044630 , 32'h00035833 , 32'h00015F8A , 32'hFFF75FAD , 32'hFFFBF00D , 32'hFFFFCC37 , 32'h000403D8 , 32'hFFFE1115 , 32'hFFF85A7F , 32'h0001880E , 32'hFFFE4D39 , 32'h000210E9} , 
{32'h0001E82D , 32'hFFF5C537 , 32'hFFF6B7F5 , 32'h00030E96 , 32'h00004FBF , 32'hFFFCAC70 , 32'h00040DC0 , 32'hFFFFDAFF , 32'h0003380E , 32'hFFFD98BD , 32'hFFFDAA27 , 32'h0004AF9B , 32'hFFF95562 , 32'hFFFE775A , 32'hFFFF0983 , 32'hFFF6D9BD , 32'h0009DD5C , 32'h0007C67B , 32'hFFFE725A , 32'hFFFB26EE , 32'h0007824C , 32'hFFF5A521 , 32'hFFFBEF90 , 32'hFFFAFD40 , 32'hFFFD6BB7 , 32'h00037D9D , 32'hFFF2C787 , 32'hFFFE598F , 32'hFFFE3747 , 32'hFFFCEB38 , 32'h00019538 , 32'h000868DA , 32'h000611C1 , 32'h00058FB8 , 32'hFFFA6C0C , 32'h00024A28 , 32'hFFFA795D} , 
{32'hFFFE8850 , 32'hFFFF945E , 32'hFFF7C448 , 32'hFFF88167 , 32'h000399AE , 32'hFFF9ED00 , 32'h000532E6 , 32'hFFFEFEAC , 32'h0001DC9B , 32'hFFFB68D3 , 32'hFFFCC47D , 32'h00032C90 , 32'hFFFFDC06 , 32'h00010750 , 32'h00028989 , 32'h00056F29 , 32'hFFF516EC , 32'h0004DDBF , 32'h0004B114 , 32'h00028E2E , 32'h0008C442 , 32'h0000DA02 , 32'hFFF4E414 , 32'hFFFB3446 , 32'hFFFC1C6A , 32'hFFF991FD , 32'hFFF760C9 , 32'hFFF99E6E , 32'hFFFB5B1D , 32'hFFF90E33 , 32'h0002978B , 32'h00042F25 , 32'hFFFED297 , 32'hFFFF9FEC , 32'h00036BAE , 32'h000B076D , 32'hFFFEB491} , 
{32'hFFFD4974 , 32'hFFFA1D83 , 32'hFFFFEC2B , 32'hFFF8D9AE , 32'hFFFE2333 , 32'hFFF98F3B , 32'h00066B44 , 32'h0003CAF7 , 32'hFFF7C660 , 32'h00082FF4 , 32'hFFFF047A , 32'h0003B103 , 32'h000226DD , 32'h00096588 , 32'hFFFD805D , 32'hFFFE614B , 32'h000408C7 , 32'h000A29B6 , 32'h0002C323 , 32'hFFFE3872 , 32'hFFFFDE74 , 32'hFFFF34BF , 32'hFFFE9616 , 32'h00084CD8 , 32'h00028D65 , 32'h00059715 , 32'hFFFEC42B , 32'h00020E9F , 32'h00024C9F , 32'h000177AA , 32'h00008D43 , 32'h00056FCC , 32'hFFFD202A , 32'h0002AE2A , 32'h0003AE29 , 32'hFFFCFDE4 , 32'h000AAF5B} , 
{32'hFFFE08CB , 32'h00025080 , 32'h0002A09D , 32'hFFFD2F25 , 32'hFFFE3B45 , 32'h00028239 , 32'h00048839 , 32'hFFFFEC04 , 32'h0000B1A4 , 32'hFFFB5C68 , 32'h00001942 , 32'hFFF9B604 , 32'hFFFE871A , 32'hFFFFFA47 , 32'h00024C3E , 32'hFFF5A434 , 32'hFFFB7DF7 , 32'h000A1028 , 32'hFFFDCB4B , 32'hFFFAAD19 , 32'h0008B3D3 , 32'h0000F9E7 , 32'h0004C806 , 32'hFFFB3553 , 32'h00036088 , 32'hFFFC0B8C , 32'h00046FDB , 32'h00015465 , 32'hFFFE4A2E , 32'hFFF73496 , 32'hFFF98394 , 32'h00044F5B , 32'h0004CF7E , 32'h00009C32 , 32'hFFFE1E99 , 32'h00031F3A , 32'hFFFF44B6} , 
{32'h05FCECE8 , 32'h01050D1C , 32'hF8A18680 , 32'hFD4CB6AC , 32'hFEC92B2C , 32'h052A6DB8 , 32'hFA9BC5A0 , 32'h02DFDD9C , 32'hF92DC778 , 32'h00614315 , 32'hF7FFA290 , 32'h00B6B277 , 32'h02C4956C , 32'h059800C0 , 32'h0153812C , 32'hFB0AC820 , 32'h0732F2B8 , 32'h0618EAC8 , 32'h01A8577C , 32'hFD7C65C8 , 32'h02CAADF8 , 32'hFCCFF9FC , 32'hF9333580 , 32'hFFD4F981 , 32'h0309767C , 32'h050A5F78 , 32'h0CBA29C0 , 32'h01943D90 , 32'h013E5FF4 , 32'hFE795670 , 32'hFE0FDA84 , 32'h05F9CC50 , 32'h0485BB38 , 32'h0090440F , 32'h01AD7E08 , 32'h03B4DE14 , 32'h0B52ED70} , 
{32'hFFC0D589 , 32'hFFFB96C6 , 32'hFFC84F6F , 32'h0015AB6D , 32'hFFD50ADF , 32'hFFEA9C6C , 32'hFFF4AE3D , 32'h00010573 , 32'hFFE4BE4D , 32'h001162CE , 32'h0022A457 , 32'hFFDEA609 , 32'h000D1F9E , 32'h00102749 , 32'h000A0C61 , 32'hFFE27E17 , 32'h000A1CD4 , 32'hFFE25051 , 32'hFFE629F1 , 32'h00164B97 , 32'hFFEC020A , 32'h002EBC2E , 32'h0005A41A , 32'h001025C9 , 32'hFFAA2D42 , 32'h0007A904 , 32'hFFEE1B8D , 32'h000355AE , 32'hFFCE7DE7 , 32'hFFFA0EC9 , 32'h00085F0F , 32'hFFE57CBB , 32'h000662C1 , 32'hFFFF0605 , 32'h0039D906 , 32'h00048EB3 , 32'h00336FB5} , 
{32'hFF9AB6EF , 32'h099866D0 , 32'h02DF9FB0 , 32'h0B73B9B0 , 32'hE464EC80 , 32'hF1605F50 , 32'hF47CBEA0 , 32'hF94EDAC0 , 32'h07C19CD8 , 32'hFFA2ED16 , 32'h0D12E470 , 32'hE6342660 , 32'h00F9A03E , 32'hF4E34B40 , 32'h0A2FC350 , 32'hE4F8CB80 , 32'hDE50EF00 , 32'h1250ABC0 , 32'hF5F8CB50 , 32'h05C35388 , 32'hFD3DFCFC , 32'hF5723700 , 32'h00F6D6A0 , 32'hFAC44DD8 , 32'h1C56E940 , 32'hFC5D10D4 , 32'h08496180 , 32'hF713DFF0 , 32'hF2A8B3E0 , 32'h0BEC7680 , 32'hEE765860 , 32'h0F2232D0 , 32'h01547454 , 32'h07FB1AA8 , 32'hF9EF9928 , 32'hF00576F0 , 32'h03FBBE4C} , 
{32'hF61E78D0 , 32'hECC13B60 , 32'h09986B30 , 32'hEDCA98C0 , 32'hE2EBBA80 , 32'hFB38EED8 , 32'h280724C0 , 32'h057047E0 , 32'hF8070878 , 32'hF02B25D0 , 32'hF1B713B0 , 32'hE96DE760 , 32'h177A8520 , 32'hFF991A8F , 32'hF8BDF030 , 32'hE14FFBC0 , 32'hF0A06A10 , 32'h27FD4280 , 32'hFC887EE0 , 32'h17C634E0 , 32'h0EFCEAF0 , 32'hF67D8B30 , 32'hD1E2DF00 , 32'hE133F600 , 32'h08FC0010 , 32'hFA5FC2D8 , 32'hEF4235E0 , 32'h0C7055E0 , 32'hF6993270 , 32'hF5C8B140 , 32'hF130A590 , 32'h09DDE640 , 32'hF0B700D0 , 32'h0CF03820 , 32'hCDE75340 , 32'h141B1820 , 32'hE5DEB020} , 
{32'hE6B94DA0 , 32'h1141C4C0 , 32'hE14D58A0 , 32'hEBE831E0 , 32'hDCA782C0 , 32'hDB14FD80 , 32'h089F1590 , 32'hF935BCF0 , 32'hFFB1D41D , 32'h0A204180 , 32'h11C608E0 , 32'h016C55F0 , 32'h0707E2F8 , 32'h006E3999 , 32'hDE0A5E00 , 32'hDF44A800 , 32'hF29417B0 , 32'h18CA5900 , 32'h01A275F4 , 32'h1810D880 , 32'h027EE1C8 , 32'hF15CB180 , 32'hECD1ED00 , 32'hF1BBC340 , 32'h016D66B8 , 32'h1C7D6580 , 32'hFF46C3A0 , 32'hDBD60C40 , 32'hE4F92520 , 32'h1DD0D5E0 , 32'hF40E8590 , 32'h26A4EB00 , 32'hEBF7CE60 , 32'h146C1F00 , 32'h01E5F10C , 32'hF89F1078 , 32'h01D11B84} , 
{32'h0303FB0C , 32'h0CEA5C00 , 32'hF74DED10 , 32'hDC49DA40 , 32'hF87375D0 , 32'hEA256F20 , 32'h18E48D60 , 32'h07586450 , 32'hEDDB41E0 , 32'hFD768F8C , 32'hE82BF920 , 32'hFAEB5640 , 32'h0576F750 , 32'hF39AA900 , 32'hF07DC170 , 32'hF26264F0 , 32'hE366D580 , 32'h1D8BA0E0 , 32'hFD407BC0 , 32'h036C89DC , 32'h1508B420 , 32'hF789E720 , 32'h0E5D1270 , 32'hF986A698 , 32'hF079E4F0 , 32'h10B98BA0 , 32'h16120EE0 , 32'hF6F911F0 , 32'hEF67DBC0 , 32'h0F98C370 , 32'h0764BD50 , 32'h025D05CC , 32'hF2587620 , 32'h21B4F080 , 32'h0D9338D0 , 32'hF009C680 , 32'hF5A9A430} , 
{32'h0B364640 , 32'h24A89800 , 32'h01FD0468 , 32'h05962068 , 32'hEB0D8A40 , 32'hFB4555E0 , 32'hF246F1B0 , 32'h058C7480 , 32'hFC35440C , 32'hF51CD190 , 32'hEF834040 , 32'h0F295310 , 32'hFB619CC0 , 32'hEDDFF080 , 32'hEC778B40 , 32'hFE049940 , 32'hDD793740 , 32'h05E3BC88 , 32'h0CC5D280 , 32'h11D7A140 , 32'h029EC558 , 32'hFD900324 , 32'hF524D2B0 , 32'hFC9C6BE8 , 32'h0F9697F0 , 32'hF8996A70 , 32'h0EB7C870 , 32'h084EB390 , 32'h123CF380 , 32'h02F6C900 , 32'hE8A23220 , 32'h11EE6CA0 , 32'hF3204B10 , 32'hFE120340 , 32'hFCA7E144 , 32'hF06A9070 , 32'hFE07699C} , 
{32'h11724540 , 32'h1AED17A0 , 32'hFE6BC8CC , 32'hFB3B15C0 , 32'h169A26A0 , 32'hE1300820 , 32'hE419B2A0 , 32'h0595D498 , 32'hF23A9930 , 32'hFD9DE4E8 , 32'hDFBF2400 , 32'h1D4B5DA0 , 32'h044E6B00 , 32'h13005A60 , 32'hD6CD8EC0 , 32'hFF0416CD , 32'hD9FAC940 , 32'h0A6BFD90 , 32'hE9FF6E60 , 32'hF8010130 , 32'h11E21400 , 32'h04EEF570 , 32'hEB898560 , 32'hE0257C80 , 32'h08DA1080 , 32'h10186A60 , 32'hF0DEC140 , 32'h09EA6DB0 , 32'h01E0888C , 32'h0C4430E0 , 32'h052A5B28 , 32'h161FFF20 , 32'hE8F08B80 , 32'h23947580 , 32'hF2541BB0 , 32'h03F6220C , 32'hF64D8490} , 
{32'hED33AA00 , 32'h1AA2ABE0 , 32'hFC5423F0 , 32'h05220C40 , 32'hF72B92C0 , 32'hF0750250 , 32'h02B327D8 , 32'h10C73100 , 32'hFE47126C , 32'hF42F2B50 , 32'h0A704BD0 , 32'h0AE5D490 , 32'hFC0307BC , 32'hF0481440 , 32'hC801ED00 , 32'hFD94D9F0 , 32'hEDBA6B00 , 32'h2647A2C0 , 32'hFAAC82C0 , 32'hEB4E4720 , 32'h31810280 , 32'h045D4ED0 , 32'h09468320 , 32'hF0609F00 , 32'hDF81E3C0 , 32'h1CB4AAA0 , 32'h20569E40 , 32'h20A5AB40 , 32'hFEB105F4 , 32'hFB298A60 , 32'h15326F00 , 32'hDF88E400 , 32'hDF1056C0 , 32'h095A3BD0 , 32'hFA22D948 , 32'hF00FFC90 , 32'hFA0D48B0} , 
{32'hF1E4E310 , 32'h199E42E0 , 32'h0D9ACFB0 , 32'hF58201E0 , 32'hF918A7F8 , 32'hE387E600 , 32'hDC4FDA80 , 32'h0488C1F0 , 32'hFA749260 , 32'hFA313378 , 32'h011673D0 , 32'h0021FAC5 , 32'hEC17C6C0 , 32'h278F9C00 , 32'hCEA6F540 , 32'hF660F1A0 , 32'hEDE9D2A0 , 32'hF9DA2738 , 32'h180ABDC0 , 32'hFE2683F8 , 32'h243E9340 , 32'hFB101268 , 32'hF2774470 , 32'hF7BB5CD0 , 32'hC43F4000 , 32'h0D727BB0 , 32'h0DAA1320 , 32'hF21EB6E0 , 32'hE7FDA400 , 32'hF60DBC70 , 32'h0D2C0410 , 32'hD39D4340 , 32'hEB308320 , 32'h03F4D814 , 32'hFA651190 , 32'hD983A500 , 32'hF51B9360} , 
{32'h03212A1C , 32'h4FC3FE80 , 32'hF37BA680 , 32'hDA9B8440 , 32'hEBF0E1E0 , 32'hE42C2220 , 32'h0DD69750 , 32'h1D251EE0 , 32'hF0072050 , 32'hFB952938 , 32'h03D613D0 , 32'hEFAB91E0 , 32'h0C190A50 , 32'hF39446A0 , 32'hAD204280 , 32'h13BE05A0 , 32'h06D21C78 , 32'h0069AEFB , 32'h0677B190 , 32'hFF43D73E , 32'h47476A00 , 32'hF7B53D00 , 32'hFACB7150 , 32'h1CB41380 , 32'hE59E2C20 , 32'hF9284E30 , 32'h1D95DF60 , 32'h0EB2D600 , 32'hE5BCD840 , 32'hFFF62CAD , 32'h028DE21C , 32'hEFDF4B40 , 32'hF02EC940 , 32'hEE1F0960 , 32'h125EEE40 , 32'h0040D4B1 , 32'h03CFA2D0} , 
{32'h1358AAC0 , 32'h205AB940 , 32'h098AF130 , 32'hDF15A700 , 32'h11BAD8C0 , 32'hEA500C20 , 32'h1213A040 , 32'h0C14A1A0 , 32'hF9FA5440 , 32'h008F0103 , 32'hF84ABB48 , 32'h0465CDC8 , 32'hF2754BD0 , 32'h0409F278 , 32'hDBECD440 , 32'hF9895380 , 32'hF90D9608 , 32'h229631C0 , 32'hE6D2B720 , 32'h07BA7800 , 32'h05316AC0 , 32'hF9CB7C78 , 32'hEC427B00 , 32'h093BA750 , 32'h050907E8 , 32'hFD7A87A0 , 32'h0AB05110 , 32'h04878908 , 32'h106BD620 , 32'h19D3E500 , 32'h335F6000 , 32'h0A0C7870 , 32'h0100CAE4 , 32'h097828E0 , 32'h106ADB40 , 32'hF7A810C0 , 32'h0D57E760} , 
{32'hF85605D8 , 32'h0DF90370 , 32'hF0D82A30 , 32'hF4C0F250 , 32'h09573200 , 32'h0233A028 , 32'h048F9EB0 , 32'h0CB97510 , 32'h011270C8 , 32'h0308C37C , 32'h0875F790 , 32'hF9DBD090 , 32'hF8936940 , 32'h05C8A290 , 32'hE9C2D3E0 , 32'hEDAED860 , 32'h16183A60 , 32'h0816B470 , 32'hF842A3E8 , 32'hFAFEBF90 , 32'hEF01A340 , 32'hEA67D6A0 , 32'hEB3E9EC0 , 32'h055BE2E8 , 32'h08E1F6B0 , 32'h20A603C0 , 32'hFED6459C , 32'hE9176060 , 32'hF2D5FED0 , 32'hF97BCAA0 , 32'h08548580 , 32'h05125F78 , 32'h19A8BEC0 , 32'h0DA0C410 , 32'h087F0910 , 32'h0B227520 , 32'h06665CB0} , 
{32'hF1C40A60 , 32'h398AF880 , 32'hF3C99F20 , 32'hF4D46570 , 32'h1963BEC0 , 32'h0E705AA0 , 32'hFE78BF0C , 32'h203E8980 , 32'hF4C64120 , 32'h1F7C87C0 , 32'h201C1400 , 32'hECD57880 , 32'hDEAE2380 , 32'h17C4CC00 , 32'hCBE92280 , 32'hE2219100 , 32'h4755DD80 , 32'h087B05F0 , 32'hE5F70B80 , 32'h0B858F20 , 32'hC1A25300 , 32'hD23E9840 , 32'hD44DE880 , 32'h0E5116F0 , 32'hF793EEC0 , 32'h2150F6C0 , 32'h0DE53440 , 32'h04598228 , 32'h0FCC45D0 , 32'h0B31DCC0 , 32'hEF4033A0 , 32'h089B8FA0 , 32'h0975C790 , 32'h109D85A0 , 32'hFE7E30F4 , 32'h15B80220 , 32'hF5D17040} , 
{32'h0C153810 , 32'h26FF4D80 , 32'h0A03D470 , 32'hFFC9BC3F , 32'h0F9F7650 , 32'h157CA260 , 32'h0290834C , 32'h248B7B80 , 32'h0D048440 , 32'hE146F500 , 32'h16A65B00 , 32'hF19F6FD0 , 32'hDAF25580 , 32'h1D02B840 , 32'h0112A5D0 , 32'h1206F240 , 32'h2A4C1F00 , 32'h067D1168 , 32'h05AB3950 , 32'hF0E380E0 , 32'hF50A85E0 , 32'h150BE540 , 32'hF6D9AA00 , 32'hF16396B0 , 32'hEFFB93C0 , 32'h00DBFC73 , 32'hFB1C09C0 , 32'h0FF71590 , 32'h0010ED6D , 32'h248E2280 , 32'hE4756120 , 32'h05994A40 , 32'hEC3AFFC0 , 32'hF855FEF0 , 32'h0398EAD0 , 32'hF0622F20 , 32'h02BC08BC} , 
{32'h02990E84 , 32'h15F7C240 , 32'hF1C3F0F0 , 32'hECCE5340 , 32'h0135024C , 32'h0FF9DE80 , 32'h1B7E8DC0 , 32'h23BD3040 , 32'h0884E950 , 32'hE38943E0 , 32'h127CD820 , 32'hF2635BB0 , 32'hF330BC00 , 32'h0B3A02D0 , 32'h115B9C40 , 32'h01F1B440 , 32'h11B27D40 , 32'h1A068380 , 32'hF8D5EA10 , 32'h086D5F50 , 32'hEE635D20 , 32'hFF707E1C , 32'h035DC3CC , 32'hEE5DA400 , 32'hFEBC460C , 32'hF90A12F8 , 32'h05C97698 , 32'h0A7811E0 , 32'hFD2D952C , 32'h0C0D51D0 , 32'hDFBD7CC0 , 32'h15755B00 , 32'hEA1773E0 , 32'hF740E1E0 , 32'h01F7BBCC , 32'hFD70EB5C , 32'h1BAB93C0} , 
{32'h03BF5C14 , 32'h19609280 , 32'hF2A53620 , 32'hF3D5B3F0 , 32'hFFEA11C6 , 32'hF946E8E8 , 32'h2E6D5380 , 32'h32A593C0 , 32'h0AF61610 , 32'hD540CB80 , 32'h12B1DBE0 , 32'hFEAB26FC , 32'hB7484D80 , 32'h4A3AF280 , 32'h33C135C0 , 32'hF27C97F0 , 32'hC33EC280 , 32'h01721A90 , 32'h2CDA63C0 , 32'hCB567680 , 32'h130F25A0 , 32'hD0D85200 , 32'hD3949BC0 , 32'hF7396E00 , 32'hC9619440 , 32'hD24F7AC0 , 32'hF1C672A0 , 32'hEAEE5D80 , 32'hFAF1A6F0 , 32'hDDECAB00 , 32'h07EDEC48 , 32'h31D75E40 , 32'hF7A17AB0 , 32'hDD870E40 , 32'hD9DBB600 , 32'h1B3DB140 , 32'h217C0840} , 
{32'hFF23D598 , 32'h032C0284 , 32'hFE5F85D8 , 32'hFD6C1528 , 32'h0209E6A0 , 32'hFB5099E8 , 32'h0CB5D6F0 , 32'h0A0A8420 , 32'h014FF410 , 32'hFFF3E9DB , 32'h03B92DAC , 32'hFF7D03A8 , 32'hF1A7C7E0 , 32'h14DABC60 , 32'h114AE3E0 , 32'hFBD85190 , 32'hE89F68C0 , 32'h0B7E1F30 , 32'h14A27040 , 32'hEEC02F40 , 32'h08491330 , 32'hE977C820 , 32'hF55F2700 , 32'h0969F3E0 , 32'hF1C00E90 , 32'hF4D68630 , 32'hF8DDFB38 , 32'hFB920FA0 , 32'hFA768138 , 32'hFCC6B31C , 32'h05DF1E80 , 32'h0BEB5250 , 32'hF9A63B08 , 32'hF7390860 , 32'hF30F3470 , 32'h0D6C1960 , 32'h0193E588} , 
{32'hF329BEA0 , 32'hFEF3DB50 , 32'hFF9A7DEE , 32'hFAB72CF0 , 32'hFB86DB80 , 32'hF2F10A80 , 32'h0DFF0110 , 32'h07C15530 , 32'hED49ABC0 , 32'hFD28128C , 32'h0D39D900 , 32'h099D3AF0 , 32'hE87C5040 , 32'h27C7FAC0 , 32'h1073CCA0 , 32'h031922D8 , 32'hD8D13B40 , 32'h0BF21FD0 , 32'h2E5F5FC0 , 32'hE59AAB80 , 32'hF68FF0F0 , 32'hE629DEC0 , 32'hF6C68CE0 , 32'h1D7B9DA0 , 32'h24AFA3C0 , 32'h025A0F1C , 32'hF5B589D0 , 32'h06E22728 , 32'h13F226C0 , 32'h076DDA78 , 32'hF5CDE1A0 , 32'hD5111E00 , 32'hE7FF81E0 , 32'h00A375DD , 32'h1BFBC4E0 , 32'h2CA41300 , 32'h07C33AA0} , 
{32'h000E094C , 32'hFFDA4E70 , 32'h0007039F , 32'h00188EAE , 32'hFFFEE457 , 32'hFFEAAC59 , 32'h0000857D , 32'h00025B52 , 32'hFFE597A5 , 32'hFFD82D86 , 32'hFFEF92CD , 32'hFFE845CC , 32'hFFE04943 , 32'hFFF172F2 , 32'h001518C9 , 32'hFFED8DE0 , 32'h001E8B2C , 32'hFFF2060A , 32'h0008CE30 , 32'hFFD9F5C7 , 32'hFFF11B36 , 32'h002300C7 , 32'hFFFC1939 , 32'h001A62EE , 32'h003FC5DC , 32'hFFBFDC7A , 32'hFFED1B70 , 32'h0006D1AC , 32'h002D2A64 , 32'hFFE89538 , 32'h0020C92B , 32'h001B511D , 32'h00228F21 , 32'hFFFD5728 , 32'hFFE8B916 , 32'hFFEE1764 , 32'hFFF0EC56} , 
{32'hFFA2B423 , 32'h015CA494 , 32'h00C525F0 , 32'h00319B14 , 32'h0591C640 , 32'hFF9351A2 , 32'h01923D84 , 32'h0313E8A8 , 32'h008A1449 , 32'h06989720 , 32'h03D6A728 , 32'h02EA2A88 , 32'h00DB837D , 32'h082A10D0 , 32'h0B13EE60 , 32'hF445C500 , 32'hFBA594F0 , 32'h0B1E6A50 , 32'h0C0C3020 , 32'hFEA2C118 , 32'h09D639D0 , 32'hEC788440 , 32'hFAD60C60 , 32'h028DA8EC , 32'hF0BAAE80 , 32'hF72B8560 , 32'h0016FC1B , 32'hFB9B13B8 , 32'h00B55F89 , 32'h062D10E0 , 32'h093F09F0 , 32'h0EED3DF0 , 32'h00DF28A8 , 32'hFFD740C1 , 32'hFC22E3C0 , 32'h02BED32C , 32'hF56582C0} , 
{32'h00069F21 , 32'hFFFBD2E5 , 32'h000319DC , 32'hFFFB0E98 , 32'h00031CBB , 32'h00042A55 , 32'h0001E0AF , 32'hFFFEE3F1 , 32'hFFFF8037 , 32'hFFFCEA57 , 32'h0000246C , 32'h00039AF7 , 32'h0000DC31 , 32'h00032B46 , 32'h0001A777 , 32'h000736EC , 32'h00046BCF , 32'hFFFF1B6F , 32'hFFFDB198 , 32'hFFFC1267 , 32'hFFF94B4A , 32'h0000A2D8 , 32'hFFFE263D , 32'h0007ABDD , 32'hFFFA364D , 32'hFFFB2F8D , 32'h00056CA2 , 32'h0002E736 , 32'h00017498 , 32'h0000EF50 , 32'h0000E875 , 32'h0009E6D7 , 32'hFFFD98C8 , 32'hFFF8699D , 32'hFFFBB65D , 32'h0000B12B , 32'h0001858B} , 
{32'h00035986 , 32'h0003D5A5 , 32'h00035CC3 , 32'hFFFC5CB9 , 32'hFFFA57E1 , 32'h0004AEB2 , 32'h000470E0 , 32'hFFF7AA13 , 32'h000087E7 , 32'h000773A3 , 32'hFFFF71F9 , 32'h0006AA73 , 32'h0005D7B3 , 32'hFFFA74A2 , 32'h0003160D , 32'h0005F1AF , 32'h00038897 , 32'h0001EBE0 , 32'h000076A5 , 32'h000502AA , 32'hFFFDEF7C , 32'h00098679 , 32'hFFF8C4AE , 32'hFFFD28DE , 32'hFFFB834E , 32'hFFFE40EA , 32'hFFF8D023 , 32'h0007C74D , 32'h00031775 , 32'hFFFD6D83 , 32'h0001C524 , 32'h00020E65 , 32'hFFF7FED7 , 32'hFFFAA769 , 32'h0002FDBE , 32'h0001D63A , 32'hFFFC4CFB} , 
{32'hFFFDF7DB , 32'h0000DA21 , 32'hFFFDB442 , 32'h00076567 , 32'h0006167A , 32'h00021C63 , 32'hFFF833D3 , 32'h0006CC2C , 32'h0001D6C8 , 32'hFFFBF5E2 , 32'h000104F9 , 32'h00030242 , 32'hFFF9C061 , 32'hFFFD08EE , 32'hFFFDCAEE , 32'h0001541D , 32'hFFFC4B89 , 32'h00006AB8 , 32'hFFFA483D , 32'hFFFB19CF , 32'h000054A1 , 32'h00016DCB , 32'h000265FA , 32'h00025C08 , 32'h0000D9E0 , 32'h0007B6A1 , 32'hFFF9DFDC , 32'hFFFF4B83 , 32'hFFFE5A1F , 32'hFFF45025 , 32'h000BD24C , 32'h00003C85 , 32'h0004C9D3 , 32'h00082CA7 , 32'hFFFCB7DE , 32'hFFFADE57 , 32'hFFFAEB18} , 
{32'h0005BD83 , 32'h0001923D , 32'h0006E2D3 , 32'h00008674 , 32'hFFFF2354 , 32'hFFFD032A , 32'hFFF997A9 , 32'h00023626 , 32'hFFF4BC0C , 32'hFFFA8C62 , 32'hFFFEA502 , 32'hFFF756BF , 32'h00032493 , 32'h000169C0 , 32'hFFFE729D , 32'hFFFDD2D4 , 32'hFFFE457D , 32'hFFF76A31 , 32'hFFFA667F , 32'h0000DA77 , 32'hFFFC5FF3 , 32'h000ABB23 , 32'h00009426 , 32'h0004D8E9 , 32'hFFF2200E , 32'h000227F3 , 32'h00024E57 , 32'hFFFE36B3 , 32'hFFFCAD5C , 32'h000583C0 , 32'hFFFEC40B , 32'h00010CE8 , 32'h0000D8C3 , 32'h0003C9AC , 32'h0004F13B , 32'h0005F6C5 , 32'hFFFEF2E4} , 
{32'h00077723 , 32'h0000C243 , 32'h0002596B , 32'hFFF7B348 , 32'h0002D3C9 , 32'hFFFC4809 , 32'h00045630 , 32'h0000F7BC , 32'h0006F0EE , 32'h00076E49 , 32'hFFFEDAAF , 32'hFFFBC7A4 , 32'hFFFB6C48 , 32'hFFFCD5D7 , 32'h00016D9F , 32'hFFFA645A , 32'h000803B7 , 32'hFFFBFB5D , 32'h00066E6C , 32'hFFFDE43F , 32'hFFFFD7F7 , 32'hFFFB49FE , 32'h0003BED1 , 32'h000163DC , 32'hFFFBD787 , 32'hFFF02C48 , 32'hFFF9B2FC , 32'hFFFFFAEE , 32'h0001026D , 32'h0006C2B7 , 32'hFFF84889 , 32'h00029048 , 32'hFFFF389B , 32'h000171CF , 32'hFFF91E18 , 32'hFFF960DA , 32'h00029395} , 
{32'h000C3426 , 32'hFFFF01BD , 32'h000343B6 , 32'hFFFE2BD4 , 32'h00089479 , 32'hFFFEA06E , 32'hFFFF5A6C , 32'hFFFBD8AC , 32'hFFFF86C2 , 32'h0002FCD1 , 32'hFFFE49A0 , 32'h0003E5B0 , 32'hFFF8FB04 , 32'h00048BAE , 32'h0000516A , 32'hFFFE65BB , 32'hFFFAC0CE , 32'h00060D8E , 32'hFFFB20F1 , 32'hFFFE08E8 , 32'h0002FC1E , 32'hFFFDBB22 , 32'hFFFF9A07 , 32'hFFFF4A9C , 32'h0003D533 , 32'h00008756 , 32'hFFFA6123 , 32'hFFFF474D , 32'hFFF9F082 , 32'h0005100B , 32'h0002922C , 32'h00025424 , 32'h000555DA , 32'h00083BD1 , 32'h000265C6 , 32'h00001E80 , 32'hFFFE6C5A} , 
{32'hFFF9E53A , 32'hFFFF617C , 32'h00019C74 , 32'hFFF9EB2A , 32'hFFFF83A6 , 32'hFFF73A65 , 32'hFFFAF678 , 32'hFFFBAE89 , 32'hFFFBC2D1 , 32'h00018E7B , 32'hFFFCB5F4 , 32'h0002EFFB , 32'h000350E1 , 32'hFFFC0291 , 32'h00042131 , 32'hFFFE9F1B , 32'hFFFB9368 , 32'h0005B4A7 , 32'hFFFC2CE2 , 32'h000126D5 , 32'h00003A49 , 32'hFFFE2B3D , 32'hFFFBE536 , 32'h000289AB , 32'h0001B08E , 32'h00018D4D , 32'hFFFBDE7B , 32'hFFF9585F , 32'hFFFA4B64 , 32'hFFF6C669 , 32'h00076355 , 32'hFFFD2C1C , 32'h0001E180 , 32'hFFF89A49 , 32'h0008E513 , 32'hFFFFCF3E , 32'hFFF9E35F} , 
{32'h000984C6 , 32'h00063241 , 32'hFFF84D0B , 32'h0003C329 , 32'hFFFCA397 , 32'hFFF59C4A , 32'h00007C1C , 32'hFFFD7234 , 32'hFFF393F8 , 32'hFFF6E215 , 32'h00125E60 , 32'h0003F9A2 , 32'h00002707 , 32'hFFF9F0C3 , 32'h00062710 , 32'h000BB8DC , 32'hFFFE056A , 32'h00071A4A , 32'hFFF8AAD8 , 32'hFFF7D6B1 , 32'h000932FD , 32'h0003A4A1 , 32'hFFFEB454 , 32'hFFF8F250 , 32'hFFFB06D2 , 32'h00100B18 , 32'hFFF75885 , 32'h0008EDC0 , 32'h000036E6 , 32'h000095CC , 32'h00049CEB , 32'h0006EBE9 , 32'hFFFEF126 , 32'hFFF7379D , 32'h000DCDF2 , 32'hFFF8A636 , 32'h00089946} , 
{32'hFFB3D81E , 32'h03B28370 , 32'hF7626040 , 32'hF84FEE48 , 32'hF4E69EC0 , 32'hF89ED830 , 32'h044CE448 , 32'h0AC2A5D0 , 32'h0474EC98 , 32'h10D94320 , 32'h00A00FBD , 32'h0486A158 , 32'hEF8B5AC0 , 32'h09470D70 , 32'hF75CB1E0 , 32'hFEA9A8A4 , 32'h0A5517F0 , 32'h0914CFF0 , 32'hF39013F0 , 32'h0D644790 , 32'hFC198F70 , 32'hE088D040 , 32'hFD82FD4C , 32'h05790870 , 32'h049983A0 , 32'h1AB2FFA0 , 32'hEE90BE20 , 32'hFD341EDC , 32'h0867ACB0 , 32'h056C3E80 , 32'h074C86E8 , 32'h0601C2A0 , 32'h0E52A8E0 , 32'h079780B0 , 32'hFB4529B8 , 32'hF7097F40 , 32'hFC1F4AE0} , 
{32'h04AA4E10 , 32'hFE8AFAB0 , 32'hF8691900 , 32'h046B2378 , 32'hFC937874 , 32'hFC8C18B4 , 32'h055B8E28 , 32'h037FAFA4 , 32'hF7E7B9D0 , 32'h0CD1B6B0 , 32'hE9C2D940 , 32'hFBFDBA00 , 32'hFE6CCA1C , 32'h05429078 , 32'h0B33C600 , 32'hFC386440 , 32'hFDF50670 , 32'h13F452E0 , 32'hF7B6BEB0 , 32'h09416D60 , 32'hFE05DA4C , 32'hDF6BC780 , 32'h02D67F08 , 32'hF51ECA40 , 32'hFDF0C604 , 32'h03953CB0 , 32'h02B5555C , 32'hFDE18530 , 32'h06E807D8 , 32'hF01AC2B0 , 32'hFC084578 , 32'hFF0BB944 , 32'hFCE67EBC , 32'h184B9BE0 , 32'hFD608B20 , 32'hEC9BF0E0 , 32'hF59717C0} , 
{32'hFB9A96D0 , 32'hFF5B805D , 32'h226B43C0 , 32'hF12C8690 , 32'hE70F9100 , 32'h0A935CA0 , 32'h25742E80 , 32'hF638D990 , 32'hDD4E1300 , 32'h173FB800 , 32'hEA625B40 , 32'hF3AF0A40 , 32'h06C23118 , 32'hF707C320 , 32'hFE344A58 , 32'h0D72DB60 , 32'hE57AA9C0 , 32'h1EDD0260 , 32'h0225C708 , 32'h16DE3240 , 32'hF60C19A0 , 32'h021A0640 , 32'hF4BC6860 , 32'hD57E9E00 , 32'h0381DE44 , 32'hE8956B60 , 32'hE9BC1040 , 32'hEBBC7580 , 32'hEAA53E40 , 32'h0DFB51E0 , 32'hF3638660 , 32'h1B88F800 , 32'hFF47279B , 32'h0CD3DCC0 , 32'h0CEE58D0 , 32'hF5624DA0 , 32'h00B66925} , 
{32'h05717770 , 32'h0DA75BE0 , 32'h0B30D540 , 32'hFD0E2B20 , 32'h11E74840 , 32'hFAA74350 , 32'hF9B73290 , 32'hF72CDB40 , 32'hF79D0440 , 32'h049470C0 , 32'hFD1AA220 , 32'h125FE060 , 32'h063ED348 , 32'h050A1590 , 32'hFCBFE7F0 , 32'h0581A088 , 32'hF1AA5800 , 32'h0E071170 , 32'hFCD018E0 , 32'h0D339100 , 32'hFDC84994 , 32'h04F37360 , 32'hF4F24750 , 32'h0F189BA0 , 32'h14A158A0 , 32'hF9683CB8 , 32'h02B9AFA0 , 32'hF36CF130 , 32'h0E1718F0 , 32'hFE498398 , 32'hFEF3E7EC , 32'h10EA92C0 , 32'hF92B42B0 , 32'hF5304B30 , 32'h0404EF20 , 32'h0F6548A0 , 32'hEE13D080} , 
{32'h0A3F5D50 , 32'hFE8E1EC4 , 32'h07CE2348 , 32'h05615698 , 32'hFE0DC484 , 32'hFC4818F0 , 32'h08DCE230 , 32'h0CE27DB0 , 32'h07BA1128 , 32'h020409FC , 32'hF7FE6890 , 32'h003ADE15 , 32'hFE85BD70 , 32'h0165A6B8 , 32'hE186A4E0 , 32'h107FF340 , 32'hF684BDC0 , 32'h17561C40 , 32'h0B5044D0 , 32'h00BB904C , 32'h0967F180 , 32'h007B165E , 32'hFA9D1CC0 , 32'hFE25E114 , 32'h0A378070 , 32'hF5BB45B0 , 32'h06661158 , 32'h0E2449B0 , 32'hF61DF380 , 32'h07E8AAE0 , 32'h09715830 , 32'h00C69869 , 32'hFCDD0E9C , 32'h05DB58C8 , 32'hF60E1250 , 32'h01594770 , 32'hF452B3A0} , 
{32'h07EBA080 , 32'h0D0C1EB0 , 32'h2653A380 , 32'hEEF5D580 , 32'hF86DF408 , 32'hF190FB80 , 32'h0BA50190 , 32'hFD30D024 , 32'hF6BD5E60 , 32'hFA45D3C8 , 32'hF5290B10 , 32'h07C5A838 , 32'h14ED1F00 , 32'hFE47310C , 32'hDA7CEB80 , 32'hFAA61068 , 32'hE779D800 , 32'h3110BF40 , 32'h0FAF3660 , 32'h06BC1CF0 , 32'h1B04F000 , 32'hF44E95B0 , 32'h03ECC558 , 32'hED8F38A0 , 32'hD85257C0 , 32'h2014C2C0 , 32'h0E95FE50 , 32'h021445C8 , 32'h00B5107F , 32'hFF40845B , 32'hFAEBEBC0 , 32'hF35404B0 , 32'hC512E680 , 32'h2484D500 , 32'h012061C8 , 32'hDFEF14C0 , 32'hF5154EF0} , 
{32'h0F1C59E0 , 32'h1776FE60 , 32'h15D24A20 , 32'h0A58AAF0 , 32'hDA493B00 , 32'hFE92E9C8 , 32'hF4743430 , 32'hFC87BB40 , 32'hFF9DF086 , 32'hFC677E88 , 32'hF9CC05E0 , 32'h0CF27820 , 32'h061AAA28 , 32'hFF67B1C8 , 32'hE3FAFC60 , 32'h0BE556D0 , 32'hF7DAA640 , 32'h13B597E0 , 32'hF8C860B8 , 32'hF4ACD0D0 , 32'h019FCC40 , 32'h0DF0F7E0 , 32'hF11C7B60 , 32'hF067B360 , 32'hF5947B60 , 32'hFB3FC470 , 32'h00FFC99E , 32'hFB8D0E70 , 32'h00486398 , 32'hECDA7460 , 32'h01BDC464 , 32'h03B03E7C , 32'hEF21B9A0 , 32'h1F439520 , 32'h08B53E90 , 32'h059E7038 , 32'hF72EC680} , 
{32'h1276A500 , 32'h160FCD80 , 32'h1659EE40 , 32'hF2DF7F10 , 32'hEB878E20 , 32'hEDE05000 , 32'hFB233860 , 32'hFD393BAC , 32'hF86878D0 , 32'hE0DD9B80 , 32'h059CA3F0 , 32'h05E80DA0 , 32'h0CBE0FB0 , 32'hF3E434B0 , 32'hE4805320 , 32'h0AA39A70 , 32'hEFB9EAA0 , 32'h0D008020 , 32'hF4AEE8D0 , 32'hF45C1680 , 32'h11F7C980 , 32'h019925F4 , 32'h150C7DE0 , 32'hEDE9ED60 , 32'hDE591800 , 32'h0F5EA460 , 32'h12EDEEC0 , 32'hFD7C5500 , 32'h1210E3A0 , 32'hE4DBB6C0 , 32'h1AEB2BC0 , 32'hEDF9DDE0 , 32'hE704A160 , 32'h0CC69990 , 32'h0B4F2E90 , 32'hFCE803EC , 32'hF83826F8} , 
{32'h0FD95200 , 32'h1B0439C0 , 32'h011BA988 , 32'hEB1BCE00 , 32'h06A240D8 , 32'hEDCC2780 , 32'h0805C620 , 32'h0B2204A0 , 32'hFA048498 , 32'hEDC5C1E0 , 32'hF8CAF548 , 32'h07D9FB30 , 32'h000FCD9C , 32'hF40F00A0 , 32'hE0EE8A20 , 32'h103E05C0 , 32'hF9984168 , 32'h03B002FC , 32'hF4437670 , 32'h00318199 , 32'h0FADA0A0 , 32'h06D50600 , 32'hFCD81918 , 32'hFE608144 , 32'h02637F34 , 32'h03A31F60 , 32'hFD178488 , 32'h10733E00 , 32'h23E02840 , 32'hF9178318 , 32'h0E86D1F0 , 32'hFC2F2C08 , 32'h0B507B10 , 32'h024CA6A0 , 32'hF988CEA8 , 32'hFCB593A4 , 32'hFCA52AB4} , 
{32'h0BCA2000 , 32'h20B51400 , 32'hFFAA7E46 , 32'hDEBE4C40 , 32'hF4186E30 , 32'hFC9EEB7C , 32'h0E1CAB50 , 32'h0965F200 , 32'hFC4CEBAC , 32'h01A7F768 , 32'h04609F00 , 32'hFD9A2814 , 32'h0AA90F20 , 32'h0F7166C0 , 32'hEDBFA400 , 32'h1D9DB680 , 32'h0CE40C70 , 32'hE3886400 , 32'hF6468BA0 , 32'hFF2637B0 , 32'h084DFAE0 , 32'hFFFF6604 , 32'h02193E38 , 32'h174BF080 , 32'hFE8D53A8 , 32'hED6EF1C0 , 32'hF04CC2E0 , 32'h00F375A6 , 32'hFD95EEFC , 32'hFDF44A8C , 32'h09458810 , 32'h03182EA8 , 32'h011D52D4 , 32'hF73FE930 , 32'h04D76A90 , 32'h00C1D1DA , 32'h09551690} , 
{32'h104E0DA0 , 32'h17A4E100 , 32'h0238A854 , 32'hE87BAC60 , 32'h08C17A90 , 32'h0AA6BB40 , 32'h004B3B36 , 32'hF5EAEB30 , 32'h079AA7D0 , 32'h01AD032C , 32'h163C72A0 , 32'hF986EBC8 , 32'h063B9148 , 32'h02FDF958 , 32'hC53DDB80 , 32'h165B4DE0 , 32'h04D711D0 , 32'hFEB34A2C , 32'hE625EFE0 , 32'hFF908196 , 32'hF41D7FF0 , 32'hE97589C0 , 32'hDF5425C0 , 32'hFE586574 , 32'hEB257780 , 32'hED878B00 , 32'h01D133E4 , 32'hF8449A70 , 32'h04E926C8 , 32'hE6771740 , 32'h0B2FA980 , 32'hF26566B0 , 32'hF6006FF0 , 32'hFD05A984 , 32'h04CE3CD8 , 32'hFA25C648 , 32'h159752E0} , 
{32'hFE38FF18 , 32'h26787C80 , 32'h05DE1FC0 , 32'hCD537C80 , 32'h0A627E80 , 32'hFFF26B90 , 32'h0EB04740 , 32'h08B51DA0 , 32'hF3D94EC0 , 32'h02824924 , 32'h18BB7E80 , 32'hCFE71EC0 , 32'h12611C80 , 32'h08507690 , 32'hEB981340 , 32'hFCAE1E24 , 32'h15436280 , 32'hEC6A67A0 , 32'hFCF74B08 , 32'hFBD43C00 , 32'hFF82CF78 , 32'hF033D0C0 , 32'hFD4C41EC , 32'hE9D679C0 , 32'hF14D1130 , 32'hFF0628FB , 32'hEB3322E0 , 32'h06E3F1F8 , 32'hFFE85E43 , 32'h096206F0 , 32'hF8D3FE90 , 32'hF1ACF8C0 , 32'hFDF865E0 , 32'hFC74E670 , 32'hF9272000 , 32'hEBB6D980 , 32'hFD6BE014} , 
{32'h0ADF5D50 , 32'h149FCD40 , 32'h032F9324 , 32'hDC5890C0 , 32'h08356100 , 32'h0BCC2730 , 32'h1075E800 , 32'h00676714 , 32'h068E69D8 , 32'h060A0140 , 32'h19CBC220 , 32'hEF460260 , 32'hE857FB80 , 32'h01EF1EB4 , 32'h14C1B600 , 32'hFCC771F0 , 32'h1D7A8200 , 32'h19AD1CA0 , 32'hF7BA8AF0 , 32'h23F4F880 , 32'hF46D3DD0 , 32'hFE0518CC , 32'hFCD52F44 , 32'hF55F42D0 , 32'hFF5B7468 , 32'hE2C0AC80 , 32'h01CDA568 , 32'h1B287760 , 32'h051CD678 , 32'hFDC73220 , 32'hF499F3F0 , 32'h06B936D0 , 32'hF3BC0C20 , 32'hF24B2850 , 32'h134B1EC0 , 32'hFECB39F0 , 32'h14720F40} , 
{32'h14072CA0 , 32'h44500680 , 32'hE7793780 , 32'hC9BDD840 , 32'hEBE1D6C0 , 32'h142308A0 , 32'h44905980 , 32'h3C482E80 , 32'h0F818F20 , 32'hE5676520 , 32'h2B5EE800 , 32'hFACFA1C0 , 32'hE1DC4380 , 32'h00C93739 , 32'h05FB3418 , 32'h0DD1E9F0 , 32'h285636C0 , 32'h277F60C0 , 32'h00D22D8B , 32'h2E09F900 , 32'hCA843300 , 32'hFB035C08 , 32'h2884A400 , 32'hE529A440 , 32'hF3B00A40 , 32'h031B0E1C , 32'h132C8EC0 , 32'h224CD180 , 32'hFC6F70BC , 32'h0E0D7D70 , 32'hDE83B040 , 32'hFFACFE2D , 32'hFEB8C288 , 32'h04B3F8D8 , 32'h0C2C7BB0 , 32'hE7B4DFE0 , 32'h092C5F30} , 
{32'hF8884D78 , 32'h2D41FDC0 , 32'h04074AA0 , 32'h01A0BFB8 , 32'h0E22C840 , 32'h077433A8 , 32'hF86DF648 , 32'h13176200 , 32'hF6D2F810 , 32'h01D80068 , 32'hFF863C7E , 32'hFF8896D3 , 32'hFD2ED0F4 , 32'h17DDEFA0 , 32'hF3E2A170 , 32'h0AF8F130 , 32'h115B5E40 , 32'hF9CFE4E8 , 32'h1F490A00 , 32'h1A4BE820 , 32'hF54190B0 , 32'hF6A87FA0 , 32'h17DB2980 , 32'hF367E9A0 , 32'hEDF82CE0 , 32'h10A08C00 , 32'h0B1B8320 , 32'hF01C3A60 , 32'hE2577E40 , 32'h044F0C30 , 32'hEEBD4080 , 32'hFCF54E68 , 32'h07DE4310 , 32'h072D0998 , 32'h0F931980 , 32'hF2DF5B40 , 32'h1DA07140} , 
{32'hFDA129F0 , 32'hFEE1C7AC , 32'hFACB7C78 , 32'h048EF8D8 , 32'h078EC0B8 , 32'hFC97FC6C , 32'h0D9ABA70 , 32'h05734A78 , 32'hFA18F0E8 , 32'hFF6C1073 , 32'h078A9DE0 , 32'hFBD6CE08 , 32'h01718160 , 32'h0F5E9AC0 , 32'h05C9C998 , 32'hF7B8EEE0 , 32'hF5549ED0 , 32'h10FD0420 , 32'h10D5BA60 , 32'hF92E25F0 , 32'h0D93D440 , 32'hEEF83080 , 32'hF5B78680 , 32'h10B6BC60 , 32'hF97AB360 , 32'hEDF8FE20 , 32'h05E8C590 , 32'h0082F8C0 , 32'h07644148 , 32'h0899D590 , 32'hFD1E9340 , 32'h03CB1B78 , 32'h0060883A , 32'hFCCFDB50 , 32'hFE551148 , 32'h02CF958C , 32'hF7EA3700} , 
{32'h0072D1A2 , 32'hFC0699F0 , 32'h0141E1B8 , 32'h01FC0BF4 , 32'hFFCCD6E8 , 32'hFDEBEC80 , 32'h02D3C984 , 32'h0302B8CC , 32'h014CCF84 , 32'hFF771B00 , 32'h02E872B4 , 32'h04877F70 , 32'hFE62CE14 , 32'h033B9C10 , 32'h02586F58 , 32'hFD33F0E8 , 32'hFBEB3530 , 32'h038319E4 , 32'hFAAF4678 , 32'h000E3ECE , 32'h01D8E3A8 , 32'hFDA4C140 , 32'hFB498960 , 32'h03737C08 , 32'hFF6232F4 , 32'hFAF952F0 , 32'hFF225B29 , 32'hFE7CB884 , 32'h02E73808 , 32'h002A49F4 , 32'h00D8F9AB , 32'h040161D8 , 32'hFAE9CAD0 , 32'hFEFC4B24 , 32'h03B52320 , 32'hFE4E15E0 , 32'hFF458CCD} , 
{32'h0183829C , 32'hFC93DF84 , 32'h04BA2E48 , 32'h010484C8 , 32'h06BDAB60 , 32'hFE2E669C , 32'h02685278 , 32'h04EF9940 , 32'h0260C200 , 32'h06D47110 , 32'h076E9E08 , 32'h09012E50 , 32'h0234A988 , 32'h0BB06AC0 , 32'h0CA93450 , 32'hEEA59860 , 32'hFB54D058 , 32'h0DA93730 , 32'h03B50870 , 32'h008D6514 , 32'h0A5740A0 , 32'hEA9122E0 , 32'hF66CF2C0 , 32'h0335CA40 , 32'hEF289AA0 , 32'hF23F59E0 , 32'hFE15B750 , 32'hFC69EA9C , 32'h057C3DF8 , 32'h048F6D30 , 32'h0B152260 , 32'h13D2F280 , 32'hFC6DDAE0 , 32'h00D7AFE7 , 32'h026DF768 , 32'hFD0DE29C , 32'hF2255A70} , 
{32'h00917BA2 , 32'hFF42BE89 , 32'h007CFA2E , 32'h014CC198 , 32'h007A343C , 32'h001EE375 , 32'h00BB97CD , 32'h00262DAF , 32'h0037F9D2 , 32'hFDFD91B8 , 32'h00627483 , 32'h00C80333 , 32'h013A87CC , 32'h007CD889 , 32'hFF98CFDD , 32'h009C47F2 , 32'hFFD20C2D , 32'h007B3749 , 32'hFE8CF124 , 32'hFF0C4A37 , 32'h00036EBD , 32'hFD5089F0 , 32'h014C4C84 , 32'hFEE614E8 , 32'h00006DFE , 32'h006BA2FA , 32'hFFC2AE5D , 32'hFFE49271 , 32'hFF2E90A3 , 32'h004BC1E2 , 32'h00FAE6EE , 32'h00CD8236 , 32'hFF592BD2 , 32'hFF4536B5 , 32'h0038983B , 32'hFFAE609A , 32'h000F7EB0} , 
{32'hFFFF0171 , 32'h0000DEDA , 32'hFFFFEA3D , 32'hFFFDCC2E , 32'hFFFF162A , 32'hFFFD2D11 , 32'hFFFE5B61 , 32'hFFFEF310 , 32'hFFF28BEC , 32'hFFFCF448 , 32'h000476B0 , 32'hFFFB3F5F , 32'hFFFDE8FF , 32'hFFFC3477 , 32'h00012171 , 32'h0001B34F , 32'h00025E2A , 32'h00060DE8 , 32'h00018911 , 32'hFFFF6A33 , 32'hFFFD050F , 32'hFFFD4A80 , 32'h0000EEEE , 32'hFFFEBDF9 , 32'hFFFFE9EA , 32'h000A1374 , 32'hFFFE9EFF , 32'h00009760 , 32'h000075BD , 32'h0004554B , 32'hFFFF3F58 , 32'h0000551C , 32'hFFFD07FF , 32'hFFFC8F43 , 32'h0001B62B , 32'h00031126 , 32'hFFFF8A9C} , 
{32'h00016EC3 , 32'hFFFFF03D , 32'hFFFD62A4 , 32'h0002A265 , 32'hFFFA1628 , 32'h0000CC02 , 32'h0001F86E , 32'hFFFF99D6 , 32'hFFFCCF62 , 32'hFFFE0B0A , 32'hFFFB0088 , 32'h00075F46 , 32'hFFFC9F68 , 32'hFFFD82C0 , 32'h000AA31F , 32'hFFFF8C38 , 32'hFFFB23AF , 32'h00007119 , 32'h00021F92 , 32'hFFF86742 , 32'h00017200 , 32'h0005877D , 32'hFFFB5DA3 , 32'h0000AFCE , 32'h00041D26 , 32'hFFFFD2C7 , 32'hFFFBCCCF , 32'h0006C8B6 , 32'hFFF8D07E , 32'hFFF7DCBE , 32'hFFF92013 , 32'hFFFF0EC9 , 32'h0001BD83 , 32'h00005317 , 32'h00036E39 , 32'hFFFEA16A , 32'h0004E413} , 
{32'h00019AA1 , 32'h0001E1E2 , 32'h0002601E , 32'h00068737 , 32'h00000CD2 , 32'h00010EE4 , 32'hFFF7527A , 32'hFFFDFC4F , 32'hFFF94D4B , 32'hFFFA2AA5 , 32'h0003D90C , 32'hFFFF0CBF , 32'h0002C593 , 32'hFFFDE8A5 , 32'h0001B73E , 32'h0001B0ED , 32'h0003E980 , 32'h00045120 , 32'hFFFDEDEE , 32'hFFFC2581 , 32'h0003C017 , 32'hFFF28309 , 32'hFFFE86BC , 32'h0004CFC7 , 32'h0008859F , 32'h00012913 , 32'h000593E9 , 32'h00062597 , 32'h00047E4F , 32'h00063A57 , 32'h0004BB83 , 32'h00011993 , 32'hFFFB7475 , 32'hFFFE35B0 , 32'hFFFD053D , 32'hFFFA5596 , 32'hFFFEDF6F} , 
{32'hFFF7F927 , 32'h00016372 , 32'h0005354E , 32'hFFFC2A90 , 32'hFFFE296D , 32'hFFFF0865 , 32'h00037394 , 32'hFFFCF11B , 32'hFFFD72B3 , 32'h0002DD8C , 32'h00032BEA , 32'hFFFD90FB , 32'h0000FDC8 , 32'hFFFEA631 , 32'h00031206 , 32'h000058B3 , 32'hFFFFE927 , 32'h00068C58 , 32'h00010AD3 , 32'hFFFCDD3E , 32'hFFF6F404 , 32'hFFFFF23E , 32'h0000FA23 , 32'hFFFEE998 , 32'h0002E6D6 , 32'h0007ECED , 32'hFFFF6FA9 , 32'hFFFE672E , 32'h0001BF32 , 32'hFFFE7909 , 32'hFFFCFCF1 , 32'h00032114 , 32'h0003944C , 32'h00019CA7 , 32'hFFF97032 , 32'h00040ABD , 32'h0005683A} , 
{32'hFFFFE4F8 , 32'hFFFDAC2B , 32'hFFFB7E55 , 32'h000145D3 , 32'hFFFE87FA , 32'h000172ED , 32'hFFFF58F3 , 32'hFFFAB26F , 32'h0003D94D , 32'h0000E3CA , 32'h0001A9D7 , 32'hFFFDF5C2 , 32'hFFFAA03B , 32'hFFFD1EBE , 32'h00033389 , 32'h00063947 , 32'hFFFC228C , 32'h0004C2FA , 32'h0005A58A , 32'h0005A6BC , 32'h00013220 , 32'h000074A7 , 32'h0001E565 , 32'h0005B50A , 32'hFFF944CC , 32'hFFFEC891 , 32'h00076C57 , 32'hFFFD1C7B , 32'h0000CE2E , 32'h0002A088 , 32'h00048A12 , 32'h0007D52B , 32'h00034BC0 , 32'h0003E57B , 32'hFFFC72EF , 32'h00044108 , 32'hFFFF0458} , 
{32'hFFFA0B1B , 32'h0003E3C9 , 32'hFFFED8E7 , 32'hFFFCBBCE , 32'h00014948 , 32'hFFFC9506 , 32'hFFFF02C4 , 32'h000646B6 , 32'h00006A45 , 32'h00022CF2 , 32'h00062D29 , 32'h0001D5BE , 32'h0007CC0C , 32'hFFFAAD0A , 32'hFFFCD911 , 32'hFFFEA99F , 32'h000074A5 , 32'h0001639C , 32'hFFFCF7D5 , 32'hFFFEF286 , 32'hFFF79969 , 32'h0003B358 , 32'hFFFE8387 , 32'hFFFA525A , 32'h000187AE , 32'h0001926E , 32'hFFFABCAA , 32'h00042C96 , 32'h00090E0D , 32'h000381E0 , 32'hFFFC9905 , 32'hFFFCCBCC , 32'hFFFE032F , 32'h00051B1A , 32'h000242C9 , 32'hFFFD8465 , 32'hFFF78856} , 
{32'h000088BA , 32'hFFFF4BCB , 32'h00077193 , 32'h0008A26B , 32'hFFFC6DF5 , 32'hFFFC48C3 , 32'hFFFBEA8D , 32'h00006BDA , 32'hFFFB4384 , 32'h00085C53 , 32'hFFFDCBCE , 32'h00016F26 , 32'h0001D157 , 32'hFFFE6CDC , 32'hFFFBB57B , 32'h000A1B49 , 32'h000860E0 , 32'h0008DE8C , 32'hFFF8D9CC , 32'h0004AB56 , 32'h00063053 , 32'hFFFF021B , 32'hFFFEA126 , 32'h0003A6D0 , 32'h000432AB , 32'hFFF984D3 , 32'h00022D2A , 32'hFFFEBBCE , 32'h0000BAF5 , 32'h0003C280 , 32'h000283F4 , 32'hFFFE280E , 32'h0005C1B3 , 32'h0007D3E1 , 32'h00019175 , 32'hFFF9A561 , 32'h000211D3} , 
{32'hFFFEAFFB , 32'hFFFFD51C , 32'hFFFB1539 , 32'hFFFC3EF2 , 32'hFFFBB1B6 , 32'hFFF9B27F , 32'hFFF9CC7B , 32'hFFFA8142 , 32'hFFFF82AB , 32'hFFFAFBFC , 32'h0006D109 , 32'hFFFD7DBB , 32'h00008041 , 32'hFFFA8CA7 , 32'h00025D12 , 32'h000134EA , 32'hFFF895D0 , 32'h0003F89E , 32'h0002EC0D , 32'hFFFEBBEA , 32'hFFFEBAEC , 32'h0007F6DD , 32'hFFF760EA , 32'h00001BD7 , 32'h0006BAB5 , 32'h000311C5 , 32'h000135AA , 32'h00058202 , 32'h00062FEC , 32'hFFFC5279 , 32'h00070C6A , 32'h00022806 , 32'hFFF965F7 , 32'hFFFF1A8C , 32'hFFFF1333 , 32'hFFFEE5BA , 32'h0009A39F} , 
{32'h00071DFE , 32'h000EE6DE , 32'hFFF8BCD5 , 32'h0009DD6D , 32'h0006C4A7 , 32'hFFF57026 , 32'h000215DF , 32'h00074BCF , 32'hFFED7E0E , 32'hFFF77D43 , 32'h001436F5 , 32'h000DDD01 , 32'hFFFF9DB8 , 32'hFFFB246C , 32'h000D5910 , 32'h000F616B , 32'hFFF9CDC3 , 32'h00067BC8 , 32'hFFF08459 , 32'hFFF6A6F1 , 32'h000B759C , 32'h0000E94F , 32'hFFF9838E , 32'hFFF2DA7F , 32'hFFF57CE1 , 32'h0014CB8C , 32'hFFF55B07 , 32'h000E3A1E , 32'h0000CE91 , 32'h00000D09 , 32'h00040FBF , 32'h000D7402 , 32'hFFFC532D , 32'hFFFC66CF , 32'h000D4FAF , 32'hFFFDEED9 , 32'h0005EF16} , 
{32'hFB8FAE18 , 32'hFD3BC924 , 32'h018C9010 , 32'hF84BA120 , 32'hFC2DDA44 , 32'h029AC0DC , 32'hF587BF30 , 32'h017874FC , 32'hFF83DF0E , 32'hFD659EE0 , 32'hFE7CAC54 , 32'hFFDB0304 , 32'hFF83D49A , 32'h03CEEEC0 , 32'hFD835C50 , 32'h009FC622 , 32'h00F61FA5 , 32'h038CC650 , 32'h00F02B3C , 32'h00736763 , 32'hFEE27194 , 32'hFF117D17 , 32'h01685578 , 32'h00C64200 , 32'h00CB8786 , 32'hFCBF1FA0 , 32'h03052940 , 32'hFF4641BE , 32'hFF3538A2 , 32'hFF253503 , 32'h00E6BC10 , 32'hFDFFDC64 , 32'h03945B0C , 32'hFD792DA8 , 32'hFE4E7734 , 32'hFC397DC8 , 32'hFD409EA0} , 
{32'h01C53494 , 32'hF4EF84F0 , 32'hFD17F60C , 32'hF9692828 , 32'hF6686AD0 , 32'hFA8D19F8 , 32'h02262338 , 32'hF32F8280 , 32'h00E4C2A6 , 32'hFA220AB0 , 32'hF71C55A0 , 32'h0C1ED360 , 32'h057B1840 , 32'hFDCBE644 , 32'h02F3CDD4 , 32'hFBB8CE10 , 32'hE7A59820 , 32'hF5B09310 , 32'h076FC2E8 , 32'h0787E5C0 , 32'h121BE200 , 32'hFF6E1E99 , 32'h064509F8 , 32'hFF083082 , 32'hFDC2A718 , 32'hFB1F0308 , 32'h00DBD91B , 32'h005073F6 , 32'h0045D6A7 , 32'hE3F6A960 , 32'h02CE9854 , 32'h0278E014 , 32'h13CA0F20 , 32'hF2631C70 , 32'h00467CD3 , 32'h0BD54EC0 , 32'h08AC3590} , 
{32'h0C7C3CB0 , 32'h10AEB040 , 32'h09ECAA40 , 32'hF7E2C080 , 32'hEB6A7CE0 , 32'h043D1110 , 32'h0B55EEF0 , 32'h151C86E0 , 32'h11BC1720 , 32'hF5CBC010 , 32'h0FE10590 , 32'h0653C118 , 32'hF9BEFA78 , 32'hE2B5B0C0 , 32'h12AB24C0 , 32'h15FEB840 , 32'h127904E0 , 32'h1C7282C0 , 32'hECF06220 , 32'h1CEAC280 , 32'h0D6FF150 , 32'h0C2E09B0 , 32'h1593CB40 , 32'hF4441430 , 32'hFBC406C8 , 32'h0F03A940 , 32'h111ADCA0 , 32'hEAF18F80 , 32'hEBA5F580 , 32'hDDDDD780 , 32'h2461F900 , 32'hF7AEC990 , 32'h030E7094 , 32'h0316DA54 , 32'h079ACBF0 , 32'hFEACEF90 , 32'hF4D7BA10} , 
{32'h0562E7B8 , 32'hE7BA9860 , 32'h04F9AEA0 , 32'hEA70F260 , 32'hDDBDDEC0 , 32'hDD5BF900 , 32'h0A17AB60 , 32'hF4624F10 , 32'hFF4DB9BF , 32'h11C5EF60 , 32'hF3EBB8A0 , 32'hE92C27A0 , 32'h10EFAEC0 , 32'h0AA9F900 , 32'h1BB23320 , 32'h14360D80 , 32'hF0B00720 , 32'h2622E480 , 32'hEB3CB500 , 32'hF33FE410 , 32'h158CC180 , 32'h12CEBEC0 , 32'h134386A0 , 32'h033979F8 , 32'h0BE165A0 , 32'hE5E2FAC0 , 32'hDA08AEC0 , 32'hE463CFC0 , 32'h1478E700 , 32'h14466A20 , 32'h0062F838 , 32'hFAEB4378 , 32'hFE76D1C4 , 32'hEBC56820 , 32'h03A61B10 , 32'hEA26FB60 , 32'hEE921340} , 
{32'h099FBAC0 , 32'h02B35034 , 32'h00534762 , 32'h01688274 , 32'hFDD2663C , 32'hF147E150 , 32'h04D6AA38 , 32'hFB68D730 , 32'hF4796690 , 32'hF9C76780 , 32'hFC352AE4 , 32'h15AAA280 , 32'hF5C1CFF0 , 32'hFCE3B308 , 32'hE8EA8B40 , 32'h099E7E60 , 32'hED6A3960 , 32'h1C2F4020 , 32'hF7CD1A20 , 32'h0B4F5490 , 32'hFB69A268 , 32'h032F599C , 32'hF58221B0 , 32'hF8E85CF8 , 32'hFFB04F42 , 32'hFEC37640 , 32'h108A5520 , 32'hF1417730 , 32'hF37CB710 , 32'h11013860 , 32'hFDA4F388 , 32'h005D8E01 , 32'hF6C29EE0 , 32'hFED4FA4C , 32'h0941A9B0 , 32'hFFB09241 , 32'hF6084350} , 
{32'h0488C610 , 32'h16F0EAA0 , 32'h101C2560 , 32'h061C14B0 , 32'hE6470100 , 32'hF3582F00 , 32'hF84B4F78 , 32'hFEA37D24 , 32'h0094340A , 32'hF8AF9218 , 32'hFFC176F2 , 32'hFF4A5BF5 , 32'h0286975C , 32'hFF05D1B7 , 32'hF4CB2150 , 32'h01F13974 , 32'hF81136F0 , 32'h0C10C2E0 , 32'hF94576D0 , 32'hF71B2E50 , 32'h093FB450 , 32'h0053B22A , 32'h1196C300 , 32'hEC847700 , 32'hFD48301C , 32'hFFB2793B , 32'h03C25A4C , 32'h08E8A570 , 32'h12F8CD20 , 32'hEF9F6A80 , 32'h0CC810E0 , 32'hF77EA700 , 32'hF6CB8E70 , 32'h016551AC , 32'h062F8B60 , 32'h07861148 , 32'h0290E140} , 
{32'h130D4F00 , 32'h2D161540 , 32'h290CF280 , 32'hEF6FC8A0 , 32'hE65A68C0 , 32'hE8845CE0 , 32'hFF09B4E9 , 32'h0606B800 , 32'hE44319C0 , 32'hF8A85488 , 32'hF888B358 , 32'hE325BD20 , 32'h15FA5100 , 32'h03BF49B4 , 32'hE839BB80 , 32'h077C8F68 , 32'hF8A03388 , 32'h1881CC80 , 32'h18C8D180 , 32'h01933A74 , 32'h047FCF50 , 32'hFE519958 , 32'h0F980400 , 32'hE55DF5C0 , 32'hFC2FB57C , 32'hF214ECB0 , 32'hE53E6800 , 32'hF62836A0 , 32'h0F8E7D70 , 32'hE63E63C0 , 32'h0E3A91A0 , 32'h03F4D07C , 32'h094BA880 , 32'h0C638650 , 32'h08F8FB80 , 32'h0E14FCA0 , 32'h150AFB80} , 
{32'h07946C28 , 32'h0F5FEE50 , 32'h0E5BFBF0 , 32'hF0B2AFF0 , 32'hEA23B2C0 , 32'hE4AC5780 , 32'hFFD1E510 , 32'h10D4A0A0 , 32'hEC189620 , 32'h08E734F0 , 32'h08FE2F50 , 32'hF7F87B50 , 32'h18865820 , 32'h13B1AA80 , 32'hFA133CE0 , 32'h2077F6C0 , 32'hE0CF72E0 , 32'h0D0F1670 , 32'hF3FCFEB0 , 32'h024E1208 , 32'h027D3C7C , 32'h0340FBE4 , 32'h02ECDC28 , 32'hE9A4E380 , 32'hEFBCA980 , 32'h0067D516 , 32'hD2ADC000 , 32'hFEAC3E9C , 32'h18599C40 , 32'hE886F5A0 , 32'hFFF16F44 , 32'hF98ED710 , 32'hFB003378 , 32'hF3829B90 , 32'hFA6DC860 , 32'hEF768B60 , 32'hF5BD6AA0} , 
{32'h0192BE60 , 32'h0E4822E0 , 32'h090E35B0 , 32'hE69616E0 , 32'hF6007CC0 , 32'hEFA045E0 , 32'h05E82608 , 32'hF90E96C8 , 32'hF14B4430 , 32'hF41B15E0 , 32'h00B2E20D , 32'hFE592C08 , 32'h06EE9DA8 , 32'hF0DC1780 , 32'hFE16E2A8 , 32'h030D8978 , 32'h0AAD43A0 , 32'hEF560440 , 32'hE87EFC80 , 32'hFEDAEA38 , 32'h044603A0 , 32'hF5185CC0 , 32'h0BA67700 , 32'hF26AA280 , 32'hEFC58500 , 32'h130BBE00 , 32'h0786EF58 , 32'h06F722F8 , 32'h1D15F680 , 32'hECCDF8E0 , 32'h079D0BC0 , 32'hEF49A7C0 , 32'hF52F12B0 , 32'hFD4D6E04 , 32'h15B7D680 , 32'h056C1B68 , 32'hFD867A60} , 
{32'h0DF61C40 , 32'h177001A0 , 32'h07C19380 , 32'hE95D6840 , 32'hF812AF88 , 32'hFD2FB3D8 , 32'h0EA465A0 , 32'hFB11C2E8 , 32'hE7A67F40 , 32'hEA200100 , 32'hF453B820 , 32'hF0B5EB60 , 32'hFDADA2F4 , 32'h0691C6C0 , 32'hFEE13324 , 32'h2A8D3700 , 32'h0C3E64E0 , 32'hED08F040 , 32'h03C42E3C , 32'h02F795EC , 32'hF23D6EB0 , 32'hEE627580 , 32'h10D3F4E0 , 32'hE7803880 , 32'hEFB4F1E0 , 32'h0380A97C , 32'hD7F4AE00 , 32'hEC34A900 , 32'h090A26D0 , 32'hFC311894 , 32'hFD5E5910 , 32'hFF6F3CA3 , 32'h027745B0 , 32'hE5968740 , 32'h05AF57F0 , 32'h165315E0 , 32'h15096740} , 
{32'h0B457C30 , 32'h1D7BDEC0 , 32'h06F248D0 , 32'hE3132420 , 32'h0B1B1B40 , 32'hFC5489E4 , 32'h0B9704B0 , 32'h005A01E8 , 32'hE4E30740 , 32'hF77C5620 , 32'h019EEECC , 32'hF31BFCF0 , 32'h055696F0 , 32'hFDBDF57C , 32'hE0CF17E0 , 32'h20EB5A40 , 32'h0BEF35B0 , 32'h0288BCCC , 32'h0DA1EB80 , 32'h180A7960 , 32'hE014FAE0 , 32'hEFB51A20 , 32'hEAD8D900 , 32'hDAC5B180 , 32'hFDA23E5C , 32'hFEEE3EB0 , 32'hD1FF2300 , 32'hE6F92B00 , 32'hF68941F0 , 32'hF3FD7FD0 , 32'h023667FC , 32'h0494E1C0 , 32'h0BDBB690 , 32'hF5AA4D70 , 32'hFF6348CC , 32'h04391648 , 32'h1C8FBB00} , 
{32'h13DA6440 , 32'h29A6A240 , 32'hF5D16C20 , 32'hD67D6BC0 , 32'hF23C9720 , 32'h152E9AC0 , 32'h296EC6C0 , 32'h2576E900 , 32'h0D35D670 , 32'hE52A6860 , 32'h21AD54C0 , 32'hE467AB20 , 32'hF9C4E7A8 , 32'h0989DEF0 , 32'hF811C980 , 32'h3266A840 , 32'h37333740 , 32'h00132AC3 , 32'hDC8D1100 , 32'h1AB87400 , 32'hD74728C0 , 32'h1B22BDC0 , 32'hF5ADD2D0 , 32'h193BD620 , 32'h248F8900 , 32'hFEB7E15C , 32'h156060A0 , 32'h1338CD60 , 32'hFA22C550 , 32'hE1895700 , 32'h073F7500 , 32'hD9827480 , 32'hF2569F00 , 32'h00702709 , 32'h22EDD4C0 , 32'hF4C6BBD0 , 32'h32660F00} , 
{32'h230B4540 , 32'h33E881C0 , 32'hFF2AEE45 , 32'hDCBEFF00 , 32'h054CBB90 , 32'hEF1C42A0 , 32'h260A5CC0 , 32'h02161B88 , 32'hDF5E83C0 , 32'h0F08A1D0 , 32'hFBD05170 , 32'hC611C780 , 32'h0791DBD0 , 32'h1CD1FAE0 , 32'hF23C1B90 , 32'h21899900 , 32'h05F49A30 , 32'hE52C37A0 , 32'hFE40C858 , 32'h2A041C80 , 32'hE7DD21E0 , 32'hE69F4C60 , 32'hFD750B88 , 32'hDB702900 , 32'h1375D4A0 , 32'hF8F53ED0 , 32'hE89D9320 , 32'h109CF9E0 , 32'h097CF0F0 , 32'h1BA6E420 , 32'h08110CA0 , 32'h025843D8 , 32'h088147A0 , 32'hFE39D40C , 32'h1B56D200 , 32'hD8A69980 , 32'hF8F17A70} , 
{32'hFE990C84 , 32'h1E962640 , 32'hE8845580 , 32'hE2AA3560 , 32'hE6626FE0 , 32'h0184FBB0 , 32'h0F81F110 , 32'h112A9180 , 32'hFC543914 , 32'hF741D1E0 , 32'hF6246FF0 , 32'hFDF719B4 , 32'hF3D44CA0 , 32'h0751EE80 , 32'hFC743A38 , 32'h0357FCAC , 32'h023DA15C , 32'hEB095800 , 32'hF81E54C8 , 32'hF6F21D40 , 32'h17C46240 , 32'hE56C2860 , 32'hFD6072FC , 32'h02D8C880 , 32'h1E9FF1A0 , 32'h27654D80 , 32'hFB612858 , 32'hED5C4FA0 , 32'hEFF74240 , 32'h08BED4F0 , 32'hFCF82664 , 32'h04DD23B0 , 32'h196D84A0 , 32'h09F61DA0 , 32'h02302820 , 32'h01447470 , 32'hF9946278} , 
{32'hF59080D0 , 32'h058B27E8 , 32'hF9402CE0 , 32'h1302B500 , 32'hFCA8013C , 32'h077F7E60 , 32'hFD270FA0 , 32'h17DB9780 , 32'h0077CD7E , 32'hF2C1BBD0 , 32'hFDF2D9B4 , 32'h09205A40 , 32'hF6FBCD40 , 32'h1063ABA0 , 32'h04FD9E20 , 32'h0B72C920 , 32'h01065A40 , 32'hF97EDE38 , 32'h2527BA00 , 32'hF98057A8 , 32'h0F245670 , 32'hF5BFABF0 , 32'h0D493C10 , 32'hFB222850 , 32'h1780E140 , 32'h15AD7E40 , 32'hF9E36990 , 32'hED236820 , 32'hFB717298 , 32'h0F4C0DA0 , 32'hF5F57B30 , 32'hE2629660 , 32'h095FB260 , 32'h16FDDB20 , 32'hFF08292B , 32'hFAAD1C18 , 32'h0DB993C0} , 
{32'h04F4F200 , 32'h0FD2DA70 , 32'h049F14B8 , 32'hF1ACBEF0 , 32'hFE9CE904 , 32'h01499784 , 32'h05140398 , 32'h004EC0E3 , 32'hF11D5AC0 , 32'h02C4DEB4 , 32'hFB6E9298 , 32'hEF2FC540 , 32'h087F4090 , 32'h05115C18 , 32'hFC6CE320 , 32'h0ED9EBD0 , 32'hFB8EB018 , 32'hF70D9660 , 32'h03127770 , 32'h0C3C2FA0 , 32'hF9FCE888 , 32'hF77A4CE0 , 32'hFC97FEE4 , 32'hF6219BB0 , 32'h00B9503B , 32'hF2727E50 , 32'hF16592E0 , 32'hFA379430 , 32'hF6A50D90 , 32'hFC1C36B4 , 32'hFD9AE5D0 , 32'h0583DF50 , 32'h02C055CC , 32'hF68F1400 , 32'h06097E68 , 32'hF67D19F0 , 32'h0571E4E0} , 
{32'hFA3948E0 , 32'hFB37AE08 , 32'h01D127E8 , 32'hFF701DDA , 32'h02ADFF60 , 32'h0055AFB3 , 32'h08280A70 , 32'h0318FA2C , 32'hF0B5A8E0 , 32'hFB70DAF0 , 32'h0F67C090 , 32'h10A9BA40 , 32'h029A9038 , 32'h1574F7A0 , 32'h026DD3C4 , 32'hF751C770 , 32'hF0A61B30 , 32'h03D0E8AC , 32'h22208C00 , 32'hF9588388 , 32'hFA8D3490 , 32'hEEAB0D60 , 32'hFDCA8CEC , 32'h1976F140 , 32'h20BA2880 , 32'h06C044C8 , 32'h01DAB780 , 32'hFE2D67CC , 32'h12E7C100 , 32'h0B664250 , 32'hF3ED6B20 , 32'hE48A1220 , 32'hE9BFD900 , 32'h00818DC4 , 32'h2BC3D800 , 32'h11284980 , 32'hFE0104E8} , 
{32'h012B68F0 , 32'hFE797EF8 , 32'hFFA2A17B , 32'h00AB2321 , 32'hFFF3F162 , 32'hFFC2AA3C , 32'h007317EF , 32'h0056FF89 , 32'hFEC942FC , 32'hFCFC20D0 , 32'h00ED0BDB , 32'h01ED7750 , 32'h02481240 , 32'h002B16B7 , 32'h011B14C8 , 32'h011960AC , 32'hFFD4062A , 32'h00AB7829 , 32'hFD9B3864 , 32'hFF30A706 , 32'hFFD1B7D7 , 32'hFDA2DA74 , 32'hFFF5748B , 32'hFEA58E70 , 32'hFF4E8A66 , 32'h0158CE9C , 32'hFF4DF360 , 32'hFFAA425B , 32'hFF6CDB96 , 32'h0068628F , 32'hFFDE4FC9 , 32'h00F1F1DB , 32'hFF915748 , 32'hFF576EF7 , 32'hFF4AF017 , 32'hFEFE4194 , 32'h00E621C4} , 
{32'hFB5A1AD0 , 32'hFD4FB4C8 , 32'h027F7BF8 , 32'hFE9F43A0 , 32'h02375A14 , 32'h005DD599 , 32'h053426E8 , 32'h011F8D8C , 32'hF4D7E4E0 , 32'hFE14926C , 32'h0BB26620 , 32'h0B97E470 , 32'h013B5968 , 32'h0FBC6C70 , 32'h0178A4B8 , 32'hF9608D38 , 32'hF5D9E550 , 32'h022079B0 , 32'h1AA859A0 , 32'hFB9B3360 , 32'hFC329AF4 , 32'hF5E975D0 , 32'hFE6023A8 , 32'h1359ECA0 , 32'h19C2DC60 , 32'h04D71488 , 32'h02196D50 , 32'hFF6973AC , 32'h0E556160 , 32'h07CE5138 , 32'hF7183560 , 32'hEB3463C0 , 32'hF096D670 , 32'h010BAAF0 , 32'h204750C0 , 32'h0E0C5400 , 32'hFD3D848C} , 
{32'hFFFF809D , 32'hFFFAD807 , 32'h00013C91 , 32'hFFFCEB68 , 32'hFFFB0196 , 32'hFFFE5EEB , 32'hFFFCA176 , 32'h00018747 , 32'h00047B74 , 32'h0002C850 , 32'h00014745 , 32'h00061829 , 32'hFFF9D2B1 , 32'hFFF9630A , 32'hFFF97929 , 32'hFFFCD3FD , 32'h00014D2F , 32'hFFFFF4CB , 32'h0002F8E5 , 32'h0003AA52 , 32'h0004F379 , 32'hFFFFCBBC , 32'hFFFE2D78 , 32'hFFFC4208 , 32'hFFFBAE05 , 32'hFFF39262 , 32'h00038818 , 32'hFFFA31B9 , 32'hFFFACC55 , 32'hFFFE6490 , 32'hFFF675C0 , 32'h000017E1 , 32'h000028FF , 32'h0002A495 , 32'h0000D58F , 32'h00027CFD , 32'h0006729B} , 
{32'h000919E4 , 32'h00040C37 , 32'hFFFFDBB9 , 32'h00068460 , 32'h00025269 , 32'hFFF8FB65 , 32'hFFFF62EA , 32'h0001E20B , 32'h0004846A , 32'hFFFC29AA , 32'h0000CA60 , 32'h000340C9 , 32'h0002C212 , 32'hFFFEBA41 , 32'h0004B33B , 32'hFFF5D6F4 , 32'hFFFFF1BD , 32'hFFFE27E7 , 32'hFFFD98C1 , 32'hFFFD43E3 , 32'hFFF7B8F9 , 32'h0006D25D , 32'hFFFFFFB5 , 32'h0005A648 , 32'hFFFF16CC , 32'h0005179A , 32'hFFF8CA0A , 32'hFFFD7474 , 32'hFFFB3CBF , 32'h00039A52 , 32'hFFF9F5B6 , 32'hFFFACCC8 , 32'h00002C53 , 32'hFFFE5454 , 32'h00006A57 , 32'h0001C893 , 32'h00028948} , 
{32'h0001972D , 32'h0002BFBA , 32'h0001FE93 , 32'hFFFEB9C4 , 32'h0002D0A5 , 32'h0002FA89 , 32'hFFFD1D47 , 32'hFFFAE04C , 32'h00025D22 , 32'hFFFBCB32 , 32'h00085EBC , 32'h00060711 , 32'h00009399 , 32'h000A831C , 32'hFFFD965F , 32'hFFFA9A8A , 32'hFFF5FC8A , 32'h0006940C , 32'hFFFCA584 , 32'h00001699 , 32'hFFF98465 , 32'h0002729F , 32'hFFFAFF31 , 32'hFFF19E94 , 32'h00053443 , 32'h0002E162 , 32'h000F4262 , 32'h0001838C , 32'h0002AFBC , 32'hFFFDAED0 , 32'h0000061D , 32'h00035DEE , 32'h00065D6B , 32'hFFFE7A6C , 32'hFFFF2A1B , 32'h0005167D , 32'hFFFB9940} , 
{32'h0002918E , 32'h00032A99 , 32'h0003F694 , 32'h0007B75B , 32'hFFFF4397 , 32'h000338EB , 32'hFFFF34FB , 32'hFFF7EDA1 , 32'hFFFCD288 , 32'h00014408 , 32'h0000CF49 , 32'hFFFE9A83 , 32'h00011642 , 32'h000278C1 , 32'hFFFEED37 , 32'hFFFD2E09 , 32'hFFFD0E15 , 32'hFFFBAF63 , 32'h000353DE , 32'h0001CEC9 , 32'hFFFFAA76 , 32'h0000FB60 , 32'h0000163C , 32'hFFFBFF31 , 32'hFFFD5DEE , 32'h00046892 , 32'h00027CEF , 32'h00021028 , 32'h000C846F , 32'hFFFEDA30 , 32'h00057568 , 32'hFFFE1F5D , 32'hFFFD2F55 , 32'hFFFF8621 , 32'h000271D3 , 32'hFFF7601B , 32'hFFF7AD0E} , 
{32'h0004536C , 32'h00000F50 , 32'hFFFF3B76 , 32'h0004604B , 32'hFFF78AAD , 32'hFFFF0721 , 32'hFFF9A32F , 32'h0000BEEC , 32'h0001D9AA , 32'h0003BC92 , 32'h000236FB , 32'h00031B5A , 32'h0002D076 , 32'hFFF80218 , 32'hFFFF5A7F , 32'h0004C63C , 32'hFFFE0DDE , 32'hFFFFB836 , 32'hFFF6AA50 , 32'hFFFF76DC , 32'h0000608B , 32'h0006495A , 32'h000164D7 , 32'h0001F55F , 32'hFFF7FCED , 32'h0000B498 , 32'h0006BB4E , 32'h0002F9BA , 32'h000037A2 , 32'h0002080C , 32'h00026B17 , 32'hFFFE14D9 , 32'hFFFC7F17 , 32'h000AEC15 , 32'hFFFF15AA , 32'h0009C2FC , 32'hFFFBC6BD} , 
{32'h00031F1A , 32'hFFFC74B4 , 32'hFFFBFB28 , 32'hFFF9EAF3 , 32'h0003EAB2 , 32'h0003CC86 , 32'h0006EB9D , 32'h0003FC4E , 32'hFFFD4621 , 32'hFFF85480 , 32'hFFF2EEBF , 32'hFFFFE808 , 32'hFFFC5B86 , 32'hFFFAAC54 , 32'hFFFEBEED , 32'h0002329D , 32'h00034F0E , 32'hFFF65162 , 32'hFFFE09A9 , 32'h000041CB , 32'h00026AD2 , 32'hFFFEB2DE , 32'hFFFE0AB9 , 32'hFFFB579D , 32'hFFFDA5E6 , 32'hFFFFBBCD , 32'h0000E303 , 32'h0000981F , 32'hFFFBFB58 , 32'hFFFDF507 , 32'h0005EBC7 , 32'hFFFD497D , 32'hFFFC48CA , 32'hFFFF6C3C , 32'h0000055D , 32'hFFFEC4A7 , 32'hFFFB0A62} , 
{32'hFFFDFBA9 , 32'hFFFB23B9 , 32'hFFFA4A10 , 32'h0001470B , 32'hFFFDBF5D , 32'h0004CEEE , 32'hFFFFBD25 , 32'h00039D2B , 32'h0000C309 , 32'hFFFA8157 , 32'hFFFF7237 , 32'h0000101D , 32'hFFFA3C65 , 32'hFFFFB3D9 , 32'hFFFC5E5F , 32'hFFFE2DDC , 32'hFFFC9948 , 32'h000CBCEB , 32'h0002EAC0 , 32'hFFFBD3D2 , 32'h00037B00 , 32'hFFFF7B4F , 32'hFFFE185D , 32'hFFFE1E6E , 32'h000306A5 , 32'h000041DE , 32'hFFFA0930 , 32'h0000715D , 32'hFFFF3FC7 , 32'hFFFFA0C7 , 32'hFFF88824 , 32'h0002F2B2 , 32'h00052162 , 32'hFFFD9ADC , 32'hFFFC8FCC , 32'hFFFDFEC1 , 32'h000671D3} , 
{32'hFFF308A9 , 32'hFFFF644C , 32'h00011702 , 32'h00017BDC , 32'h0002B682 , 32'h00020825 , 32'hFFFE967C , 32'hFFFCDCD3 , 32'hFFFB4E9A , 32'h000036D0 , 32'h0004AD86 , 32'hFFFFF391 , 32'hFFFE99F5 , 32'h00038080 , 32'h000263BB , 32'h00018C88 , 32'h00012C1E , 32'hFFFDD50E , 32'hFFFF0035 , 32'h00060393 , 32'h000A0B87 , 32'hFFFC570A , 32'hFFFFC04B , 32'hFFFB4ADA , 32'hFFFF5F56 , 32'hFFFACD3C , 32'hFFFD0370 , 32'hFFFAF613 , 32'hFFFEBCDA , 32'hFFFFF66D , 32'hFFFEA6A5 , 32'h000313FA , 32'h000852A3 , 32'hFFFC2E55 , 32'hFFFE4985 , 32'h0000C56B , 32'hFFFC259E} , 
{32'h025D678C , 32'hFF3A6AC5 , 32'h00FD4393 , 32'hFEE07E78 , 32'hFFA003CE , 32'h015F308C , 32'hFEFD2954 , 32'h0025B7AD , 32'h0269D034 , 32'h02000F10 , 32'hFFA10595 , 32'hFCF051C8 , 32'h045435A0 , 32'h00C00EF9 , 32'hFFCD1049 , 32'hFE9F9858 , 32'h0068DA7B , 32'hFE4FFBFC , 32'hFE2E7244 , 32'h01A86DF0 , 32'h053CF1D8 , 32'h0434B158 , 32'hFBE8A950 , 32'h04BBB2B0 , 32'hFAAAA8D0 , 32'h01E6B408 , 32'hFF769FE5 , 32'hF8398F68 , 32'hFC676350 , 32'hFC0288B4 , 32'hFD090EE8 , 32'h093AF770 , 32'hFD6B7D78 , 32'hFEAAF410 , 32'h05EDBF40 , 32'hFE84A0F0 , 32'hFCC7DCF8} , 
{32'h00A950AB , 32'hFC5FF98C , 32'hFF5AE025 , 32'hFAC2F3F8 , 32'hFB14D100 , 32'hFFDF8E7D , 32'h01AF4A20 , 32'hFBF47E10 , 32'h0125D5B8 , 32'hFA0D8398 , 32'hFBB34F40 , 32'hFF5A4490 , 32'h00E05F28 , 32'hFEA2F750 , 32'hFFF67DB3 , 32'h00F65778 , 32'hFC022134 , 32'hF6E15B90 , 32'h03CF310C , 32'h00A0E7DB , 32'h05538F40 , 32'h016D9204 , 32'h08415370 , 32'hF9F76D98 , 32'h023BC458 , 32'h04BB1A08 , 32'hFE157004 , 32'h05306620 , 32'h02F3CA34 , 32'hF7CA46A0 , 32'hFB3662F8 , 32'hFF9227AB , 32'h033BB8A4 , 32'hFBD1EAE0 , 32'h03DDCDC0 , 32'h045CA8E8 , 32'hFA441E50} , 
{32'h09EA4B30 , 32'hFCCA1DA8 , 32'h0446A690 , 32'hFB27CBC8 , 32'hFE49C9E4 , 32'h05B30540 , 32'hFBC59A00 , 32'h008B7F99 , 32'h0A20A880 , 32'h0817ECB0 , 32'hFE24D3A4 , 32'hF324E6F0 , 32'h12330720 , 32'h031B1814 , 32'hFF4464BA , 32'hFA2BF928 , 32'h017164F8 , 32'hF95A4738 , 32'hF8852D98 , 32'h0706E8C0 , 32'h15E70240 , 32'h11291D20 , 32'hEECA3D40 , 32'h13816FE0 , 32'hEA076DA0 , 32'h08298CC0 , 32'hFDAE81C8 , 32'hDF900300 , 32'hF13BB500 , 32'hEF37C080 , 32'hF3C51A90 , 32'h26508540 , 32'hF56C8FE0 , 32'hFA8F9BC0 , 32'h18945640 , 32'hF9CD3F88 , 32'hF2937F20} , 
{32'h140C3E00 , 32'h1D7BF040 , 32'h2FC9AE40 , 32'hFDE2AFD8 , 32'hC7466440 , 32'h0EA756F0 , 32'h0AAB0EF0 , 32'h0ACBEAE0 , 32'h0048DA38 , 32'h102F04E0 , 32'hEFA60B60 , 32'hE9CD9AC0 , 32'h22E2E440 , 32'h031AF69C , 32'hF9094FC8 , 32'h070E5118 , 32'h10BA9BE0 , 32'h00CC9C65 , 32'hF62152C0 , 32'hF1E68260 , 32'h1C07E080 , 32'h04E06838 , 32'hE8790460 , 32'h238BE000 , 32'hF126A180 , 32'hFCC591B4 , 32'hF1F96D20 , 32'hFD7CC544 , 32'hE910BFA0 , 32'hE797D240 , 32'hF1CF4550 , 32'h18493EA0 , 32'hDF07C880 , 32'h03968E50 , 32'h059FA548 , 32'h0866A390 , 32'hE60F9920} , 
{32'h032AC070 , 32'h2555F680 , 32'h315E0240 , 32'hFDFC54A4 , 32'hEB9BB520 , 32'hF40E2EB0 , 32'h103DE140 , 32'hF64F7650 , 32'h0C7ADD20 , 32'h09101F60 , 32'hD96E0600 , 32'h14995200 , 32'h0FEDBC40 , 32'h040D3F38 , 32'h0AE80890 , 32'h0DD9BDD0 , 32'hF34BABF0 , 32'h1661BDE0 , 32'hFF503112 , 32'hF0526080 , 32'h0FE602B0 , 32'hFAD2E9D0 , 32'hF3A22E60 , 32'h05466798 , 32'h00FF6B98 , 32'hEFD5DDE0 , 32'hF65582A0 , 32'hF9370BB8 , 32'h10FB9CA0 , 32'hE9DF64C0 , 32'hF73D3AD0 , 32'h09DDD4D0 , 32'h0B8AF720 , 32'hFFE31970 , 32'hF7C74940 , 32'h11A5A140 , 32'hFF1682D1} , 
{32'h077C8908 , 32'h12ED89E0 , 32'h231C1A80 , 32'hF3311590 , 32'hED59CD00 , 32'hFF7F1CBB , 32'h16330E60 , 32'h0835EAD0 , 32'hF3C96820 , 32'h083DD6E0 , 32'hDFE51C80 , 32'hF8AF56A8 , 32'h018A6AC8 , 32'h0577E508 , 32'h0EE106B0 , 32'h01C4F298 , 32'hEEF717C0 , 32'h0CE97440 , 32'hF38AF2F0 , 32'hFC0A38D4 , 32'h00117658 , 32'hEF813CC0 , 32'h026F6320 , 32'hFA672BC8 , 32'h0E9ECCD0 , 32'hF8B356F8 , 32'hF476B270 , 32'h06B97DF8 , 32'h12EF6560 , 32'hF3AA9FC0 , 32'hEECD0FE0 , 32'h08B7F800 , 32'hEFD03BA0 , 32'h1944D120 , 32'hEC08DBC0 , 32'h003FC5D2 , 32'hED2E45E0} , 
{32'h113F4300 , 32'h03773F1C , 32'h172F8C20 , 32'hEFD2AC00 , 32'hEAA33AA0 , 32'h1424C8A0 , 32'h2DD1A540 , 32'h09CE7D40 , 32'h0C216930 , 32'hFF4DE4CB , 32'h0EC634D0 , 32'hFC062454 , 32'h1675EAE0 , 32'hE78FF420 , 32'h11D3BC00 , 32'h15820000 , 32'h0D871AF0 , 32'h2FC96940 , 32'h04211D08 , 32'h0B2FB8F0 , 32'hEA7D4E40 , 32'hFE809044 , 32'h0E7FD900 , 32'h1615D220 , 32'h03545000 , 32'hF623F510 , 32'h1041F0E0 , 32'h0E17FB50 , 32'hF730B080 , 32'hF1F4B4B0 , 32'h035CB8A8 , 32'h03A98F10 , 32'hFF0F072E , 32'h0B47C680 , 32'hFE59FA9C , 32'h06E601B0 , 32'hD9EDD680} , 
{32'h0E2C7D30 , 32'h17C74980 , 32'h066A6A88 , 32'h03CBA0C8 , 32'hDD993D00 , 32'hE84BB520 , 32'h0C2FD580 , 32'h14795640 , 32'hF78069D0 , 32'hEF69D840 , 32'h1EE1F800 , 32'h10E78C60 , 32'h01A5D250 , 32'hF6E94760 , 32'hF8EB0C08 , 32'h09D99110 , 32'h039AF294 , 32'h207C36C0 , 32'h0121299C , 32'h0CE682B0 , 32'h035DC4F4 , 32'h1600B220 , 32'h097E7FE0 , 32'h04DB0CF0 , 32'hFAB91630 , 32'h0B40C240 , 32'h15BF04A0 , 32'hF46461E0 , 32'hFE43B854 , 32'hCCEF2900 , 32'h13C34840 , 32'hE8C62200 , 32'hF5CEA4D0 , 32'hFF829E80 , 32'h00EF067D , 32'hFD67FC10 , 32'hE4B077E0} , 
{32'h03382FB4 , 32'h2A9AEB40 , 32'h0C691E60 , 32'hCC31BBC0 , 32'hE9795E60 , 32'h0238A5B8 , 32'h0E407530 , 32'hF9D6BE70 , 32'hE43791C0 , 32'h04706208 , 32'h187F4520 , 32'hECFB7D40 , 32'h244D97C0 , 32'h19679F60 , 32'h0C8D3B10 , 32'h0F160EA0 , 32'h11F66300 , 32'hD3B51F80 , 32'hCAD73DC0 , 32'hE2821580 , 32'h2E162900 , 32'hE742FE40 , 32'hF6774680 , 32'h1B92DB20 , 32'h0C3DCB90 , 32'hEED5C500 , 32'hF5D35D60 , 32'hF4791370 , 32'hF35739D0 , 32'hEA0127E0 , 32'hFBD6B618 , 32'hF50AB050 , 32'hE6769180 , 32'h0165A66C , 32'h0798AD70 , 32'hF525B8F0 , 32'h02923B2C} , 
{32'h0FCF6C40 , 32'h207E2100 , 32'h031F06CC , 32'hCA7204C0 , 32'hF841C590 , 32'h07707658 , 32'h125E3DA0 , 32'hFCC7AAA8 , 32'hE7A7D300 , 32'h3050F880 , 32'h0921D5B0 , 32'hDD7616C0 , 32'h26992D00 , 32'hF1D48C80 , 32'hF1282000 , 32'h46AFC600 , 32'hED987AA0 , 32'hE7E3CC20 , 32'hF702FBD0 , 32'h12999360 , 32'hF09DBE00 , 32'hE2921F40 , 32'h08950900 , 32'hF327CAF0 , 32'h200FF140 , 32'hE82A38A0 , 32'hF1F36030 , 32'hED417840 , 32'h01E4E020 , 32'hE159F940 , 32'h0167FD0C , 32'h0CE99170 , 32'hF9B41708 , 32'hFE716E7C , 32'h09EEBF30 , 32'h01F50B7C , 32'hFD2C3FEC} , 
{32'hFCEE952C , 32'h19997960 , 32'h102CEDE0 , 32'hEE22B220 , 32'hE6CB8400 , 32'hFB395A18 , 32'h273DB7C0 , 32'h0A164A60 , 32'h124FD020 , 32'hF8776660 , 32'h04529980 , 32'hF13E82D0 , 32'h0D5E6120 , 32'h015B9974 , 32'h160B3B00 , 32'h2341EA40 , 32'h05F925C0 , 32'h0BE1C6F0 , 32'h014E009C , 32'h08327100 , 32'hFCE1A914 , 32'hFABB5E48 , 32'h048D9328 , 32'h0439AC20 , 32'h025BABD8 , 32'hE6DFEC60 , 32'h1FF6FB80 , 32'h08595F20 , 32'h1F72A140 , 32'hE0088820 , 32'hF4A278F0 , 32'hECEDEE80 , 32'h115454C0 , 32'h06D0D098 , 32'h0AB90EA0 , 32'hFE8717F4 , 32'hF6A12830} , 
{32'h09186BA0 , 32'h0E472430 , 32'hFB2ED1A0 , 32'hF0B6FBF0 , 32'h0171C564 , 32'h02A5C960 , 32'h0C6A4330 , 32'h0D7225E0 , 32'h0B26E160 , 32'hF02F2700 , 32'h0B978EC0 , 32'hFF76FCA5 , 32'hFB8560F0 , 32'hF9FCA2C8 , 32'hF4160680 , 32'h0EC2CBE0 , 32'h092B92D0 , 32'h08976B60 , 32'hF3C7DE60 , 32'h039E6ED8 , 32'hF069A720 , 32'h055B06F8 , 32'h049EBBC8 , 32'hF1492C70 , 32'h06C105A8 , 32'hE5588680 , 32'h090F48F0 , 32'h08C78B70 , 32'h123825E0 , 32'h074E66E8 , 32'hF02345D0 , 32'hF6E7EAE0 , 32'h012D5CB0 , 32'h0F229AA0 , 32'h09E39A40 , 32'hFB8EA050 , 32'h283AA500} , 
{32'h0F90A130 , 32'h26708D00 , 32'hEC674D60 , 32'hC8AB2280 , 32'h16E5E360 , 32'h19A64220 , 32'hFE002CAC , 32'h2B32EF80 , 32'h161E53E0 , 32'h4234AB00 , 32'h3F36BB40 , 32'hBA8BBF00 , 32'hEB5934E0 , 32'hF6A0FA20 , 32'hDEFE1800 , 32'h00D81AC3 , 32'h35462040 , 32'hFEC0BF74 , 32'h00067401 , 32'hE9329C40 , 32'h006B09A6 , 32'hF8FC0140 , 32'hB81FE280 , 32'h00042610 , 32'h270278C0 , 32'h29F6CB00 , 32'hF7BB30D0 , 32'h0229B21C , 32'h0434F4F0 , 32'h0A616850 , 32'hF0DF5BB0 , 32'hFEFE4C58 , 32'hEBBBA0E0 , 32'h0FE758B0 , 32'hF562C7C0 , 32'hF1DFF230 , 32'hF12F6FF0} , 
{32'h0BEA7640 , 32'h1652A380 , 32'hEA624160 , 32'hF7EF5200 , 32'h194DFD60 , 32'h18F88380 , 32'h0FB2E210 , 32'h1CD15C60 , 32'h072D9168 , 32'hF344C620 , 32'h11C937A0 , 32'hD89917C0 , 32'hF5565120 , 32'h1409D400 , 32'hC657DE80 , 32'hEE15A340 , 32'h2C4E1440 , 32'h26DE4380 , 32'hEB9F7780 , 32'hF2964360 , 32'hF8C24D40 , 32'hE8876720 , 32'hE2036880 , 32'h026ACD80 , 32'h217111C0 , 32'h38761F80 , 32'hF416CD40 , 32'hDD8C5400 , 32'h019ED108 , 32'h1B095520 , 32'hFDA2F5C8 , 32'hFEC12648 , 32'h0C843910 , 32'h133D1120 , 32'h02B754A0 , 32'h0C73B8E0 , 32'h026B8EE4} , 
{32'h065DAD88 , 32'h0ABD3570 , 32'hF9528110 , 32'h09287680 , 32'h0A6F5F50 , 32'h0296DD20 , 32'h147E5560 , 32'h0CEC64C0 , 32'h02EAF45C , 32'hFF537908 , 32'h07B12B88 , 32'hED654C00 , 32'hFA5DF540 , 32'hFC7012B4 , 32'h01BB3C64 , 32'h00809F1D , 32'h108B77C0 , 32'hFD7DEA98 , 32'hFD2A9A58 , 32'hF62FFE80 , 32'hF730A280 , 32'hFF682BD1 , 32'hFC308FB0 , 32'hF86E4F10 , 32'h019DFC84 , 32'h0A2F61B0 , 32'hF9053720 , 32'h053DDC40 , 32'h0A09EB00 , 32'h13DE1FE0 , 32'hF45C4230 , 32'h077285C8 , 32'hEE306F20 , 32'h06A84AB8 , 32'h006737EE , 32'hFD480754 , 32'hF4584710} , 
{32'hFFACBD06 , 32'h05BF08B8 , 32'h00D43E57 , 32'hF805F8A0 , 32'h06163438 , 32'h01F6EAB4 , 32'h09389AA0 , 32'h0E71CA50 , 32'hF375AA00 , 32'hF6137500 , 32'h06AAAD58 , 32'hF9058158 , 32'hFD38ED28 , 32'h10BF7CE0 , 32'h02196004 , 32'h03E00828 , 32'h019EFD60 , 32'hFA7116A8 , 32'h13371320 , 32'hF81F1F48 , 32'hEBBD51A0 , 32'hF2ABCC40 , 32'hFDCBA004 , 32'h0FCBBE30 , 32'h1F8381C0 , 32'h0CB32100 , 32'hFF4C8EB6 , 32'h0E3F55B0 , 32'h20C25C80 , 32'h118EC4C0 , 32'hEC138DE0 , 32'hEA4F6FE0 , 32'hE93E9B40 , 32'h083A13B0 , 32'h239E8040 , 32'h05860610 , 32'hEDC240A0} , 
{32'hFF087D0A , 32'h00ABEC5F , 32'hFE68A64C , 32'h0172EE0C , 32'hFF77F5D1 , 32'h001566C5 , 32'h00EB0DE0 , 32'h01316774 , 32'h008864D0 , 32'hFF8C2B61 , 32'hFE6BDFBC , 32'hFF18EB58 , 32'hFEA6055C , 32'h00B71698 , 32'h00DD1F10 , 32'h00C1C514 , 32'hFDA54468 , 32'h0198BDCC , 32'h000C2CEF , 32'hFE768098 , 32'hFEA64E4C , 32'hFE24E0F4 , 32'hFF5D665B , 32'h000BCC2E , 32'hFE2F1664 , 32'hFE9A69B4 , 32'hFEBE34CC , 32'hFF3A0017 , 32'h00DADF83 , 32'h00946776 , 32'h000F5412 , 32'h00A83790 , 32'h0017EBA5 , 32'h007DBC1A , 32'hFF41DFC8 , 32'hFE5BA8EC , 32'h00503134} , 
{32'hFACCF580 , 32'hFC3CBC18 , 32'h01D00328 , 32'hFD5452C8 , 32'hFFEEEE7C , 32'hFBBACE30 , 32'h04159E00 , 32'h069AB340 , 32'hF4219EA0 , 32'hF9306550 , 32'h069EDAB8 , 32'h0FB55CD0 , 32'hFFC05196 , 32'h0D95F170 , 32'h04D96040 , 32'hF63FF8E0 , 32'hF29AB520 , 32'h0261B6B0 , 32'h1C89B720 , 32'hFAD222C0 , 32'hFB15A968 , 32'hF6E6DF20 , 32'hF804D2D0 , 32'h108EC340 , 32'h197AF3E0 , 32'h0070B29B , 32'hFECF8C98 , 32'h0356D65C , 32'h149D6F20 , 32'h069C47C8 , 32'hED80F640 , 32'hE8F56400 , 32'hEA734940 , 32'h03C994BC , 32'h2312F500 , 32'h0D5721C0 , 32'hFA81A800} , 
{32'hFD5B880C , 32'hFDAE7C54 , 32'hFF7D992E , 32'hFE860364 , 32'hFF1CA8F9 , 32'hFFCB5DDE , 32'h0298D700 , 32'h00E96EA3 , 32'hF747E6C0 , 32'hFD6D3038 , 32'h05910BF8 , 32'h06BF6BF0 , 32'h00A5CB27 , 32'h080C3830 , 32'h04101B10 , 32'hFD269E2C , 32'hFA4DE450 , 32'h0168D178 , 32'h0D2FE440 , 32'hFDB25FC0 , 32'hFDB37310 , 32'hFBD12EB8 , 32'hFBFA5DD8 , 32'h0AF42360 , 32'h0CF45960 , 32'h02990404 , 32'hFF811522 , 32'hFEBD2DE8 , 32'h08C0AF90 , 32'h047BD7D0 , 32'hF92C7228 , 32'hF58EA7B0 , 32'hF8E977E0 , 32'h01438A4C , 32'h0FC40030 , 32'h064DB6B0 , 32'hFEDE1618} , 
{32'h0094D214 , 32'hFE76E7B8 , 32'hFEC7BD5C , 32'hFE8D0650 , 32'hFDFF8654 , 32'hFF1AD336 , 32'hFF3A1406 , 32'hFFB11C49 , 32'hFCB491F8 , 32'hFE08F1C4 , 32'h0043BE79 , 32'h0103D230 , 32'h00FC65A6 , 32'hFFDB1958 , 32'h0344D144 , 32'h00C68F49 , 32'h009E598E , 32'h003A63DC , 32'hFF478FB0 , 32'h008225A1 , 32'h000F6CA0 , 32'h018DA054 , 32'hFCEDBC58 , 32'h00823D2A , 32'h00149B6E , 32'h00B3015A , 32'hFEACB7CC , 32'hFF773097 , 32'h00E7D386 , 32'hFFF2623B , 32'hFDA99EFC , 32'h00C47FBD , 32'h010290AC , 32'h00A167E1 , 32'hFE7BAC0C , 32'hFF958F11 , 32'h000BBEAE} , 
{32'h00025768 , 32'h0005FA2E , 32'h00019F21 , 32'h000720E3 , 32'hFFFCA180 , 32'hFFFE43EA , 32'hFFF99C50 , 32'hFFF86F1C , 32'h00002FF2 , 32'hFFFD0557 , 32'h00090AB5 , 32'h00042F6B , 32'h00025F82 , 32'h00029BEA , 32'h0008850C , 32'hFFFE3B62 , 32'h0002D77F , 32'hFFFFCDEE , 32'hFFFCCDB1 , 32'h0003B8FC , 32'hFFF9B003 , 32'hFFFEA74F , 32'hFFFB9BC0 , 32'h0005DCCA , 32'h000051C3 , 32'h0005C384 , 32'h000A1D91 , 32'h00055220 , 32'hFFFF1C3C , 32'h00035AD1 , 32'h000087C2 , 32'h00024235 , 32'h0002F816 , 32'hFFFB341D , 32'h0002405B , 32'hFFFD7366 , 32'hFFFEFE55} , 
{32'h00045896 , 32'h000061B2 , 32'hFFFC4880 , 32'hFFFD96F2 , 32'hFFF32D72 , 32'h0004AD77 , 32'hFFF7EBF4 , 32'h0003DDDB , 32'h000DA9B4 , 32'h00048D3B , 32'hFFFCD152 , 32'h00001161 , 32'h000360A4 , 32'hFFF738CA , 32'hFFFFC9F3 , 32'h0007226F , 32'h00056051 , 32'h00029370 , 32'hFFFC1F01 , 32'hFFF6F8B4 , 32'h0000BDDE , 32'hFFFDBCC1 , 32'hFFFB81BA , 32'h0004D49B , 32'hFFFB73A8 , 32'h00030BA7 , 32'h00013970 , 32'h0005400F , 32'h0000CDC9 , 32'h00055BE2 , 32'h0001FF14 , 32'h0002C465 , 32'h0004B562 , 32'hFFFF1AAA , 32'hFFFFC3BF , 32'hFFFDB3C6 , 32'h00045035} , 
{32'hFFFE66A3 , 32'h0001FA78 , 32'h00004099 , 32'hFFF9D3D4 , 32'hFFF9204B , 32'h000022BF , 32'hFFFBB30C , 32'hFFFF25C0 , 32'h000C25C0 , 32'h0006C5B0 , 32'h0000A73E , 32'h00082263 , 32'hFFFB34DA , 32'h0007E37D , 32'hFFFBDEFE , 32'h00033072 , 32'h00024718 , 32'h0000B5AB , 32'h0000A4BB , 32'hFFFCEACC , 32'hFFFC509F , 32'hFFFA8B3C , 32'hFFFABF7A , 32'hFFFFD6A7 , 32'h0004A580 , 32'h000246F2 , 32'hFFFC3439 , 32'h00106ADE , 32'h00042A32 , 32'hFFFE7F14 , 32'hFFFD66CA , 32'hFFF157C6 , 32'h0001EBA4 , 32'hFFFEDC27 , 32'h0003B987 , 32'hFFFDB4CD , 32'h00041EFA} , 
{32'hFFFDB423 , 32'hFFF7C76B , 32'hFFFE7B83 , 32'hFFFC3A61 , 32'h00065710 , 32'h0002279F , 32'hFFFEDDC4 , 32'hFFFD191D , 32'h000B1181 , 32'hFFFF5C53 , 32'hFFFEBBB3 , 32'h00027964 , 32'h0008BEF8 , 32'hFFFD35DE , 32'hFFFCBCD2 , 32'h0005178D , 32'hFFFC157F , 32'h000569FC , 32'h00015D3D , 32'h00013897 , 32'hFFF8C3B3 , 32'hFFFAA9EA , 32'h0004FB2B , 32'h0007592B , 32'h0003092C , 32'h00007078 , 32'hFFFE66F6 , 32'hFFFF5942 , 32'h0002674C , 32'h0003AF0A , 32'hFFFA9E50 , 32'hFFFAAB16 , 32'hFFFF6A7A , 32'h0000AA26 , 32'hFFFDC7F6 , 32'hFFF7B670 , 32'h00085993} , 
{32'h0004E0F2 , 32'h00030C96 , 32'h0003AC5D , 32'h000465B1 , 32'h00008B5A , 32'hFFFE8B9E , 32'hFFF8AE2F , 32'hFFFDA4E8 , 32'hFFF7DD2E , 32'h000693DD , 32'hFFF67D7D , 32'hFFFAF826 , 32'hFFFBA591 , 32'h000364ED , 32'hFFFC9277 , 32'h00020C10 , 32'hFFFCA9D8 , 32'h0000E6FE , 32'h0003DCF5 , 32'h00000F5D , 32'hFFFACA4E , 32'h00035EB7 , 32'hFFFA210A , 32'h0002752E , 32'hFFF3001F , 32'hFFFB24DB , 32'hFFF68F55 , 32'hFFF8BD12 , 32'hFFFD738E , 32'h0008E626 , 32'hFFF432BA , 32'h0001D15D , 32'hFFFF4B83 , 32'hFFF96BFF , 32'h0002D711 , 32'hFFFF6A08 , 32'hFFFDB1AB} , 
{32'hFFFE7A1E , 32'hFFFFEC4A , 32'hFFF9B30E , 32'hFFFEE660 , 32'hFFFE0B1A , 32'hFFFEE562 , 32'h00000A6D , 32'h0000872C , 32'hFFFF4E29 , 32'hFFFFD30D , 32'h000245B8 , 32'h0004F3FD , 32'h00007148 , 32'hFFFF889E , 32'h00010BB0 , 32'h0002FDB9 , 32'h000357D6 , 32'h00017C1C , 32'h0003338C , 32'hFFFA508B , 32'h0007AF66 , 32'hFFFDE2C5 , 32'hFFFDF985 , 32'hFFFE2CAD , 32'h000329D0 , 32'h0007102C , 32'hFFFCE63D , 32'hFFF6AF6C , 32'h0000DE20 , 32'hFFFC6B34 , 32'hFFFBB2C6 , 32'h000667C9 , 32'hFFFCA022 , 32'h0000E717 , 32'h000212AB , 32'hFFFD4479 , 32'h0002252C} , 
{32'h0003AD62 , 32'h0000FF97 , 32'hFFF75E82 , 32'hFFFCDA5A , 32'hFFFA2FD3 , 32'h000901F0 , 32'hFFF7DAF6 , 32'h00030F30 , 32'h0000ED69 , 32'h00002322 , 32'h0002ED1B , 32'hFFFF10D1 , 32'h000A9401 , 32'hFFF521A2 , 32'hFFFD4FC2 , 32'hFFF8FA7B , 32'hFFF7AAA0 , 32'h00005053 , 32'h000ABAE9 , 32'hFFFD3260 , 32'h000558A0 , 32'hFFFED967 , 32'h0002EBAB , 32'hFFFC702C , 32'hFFFCC888 , 32'h0005EB7C , 32'hFFFA7AFA , 32'h000331D1 , 32'hFFFBF085 , 32'h0006A82E , 32'h00050154 , 32'h0006CDC9 , 32'h00024395 , 32'h0006DD52 , 32'h000091EF , 32'hFFF9415D , 32'hFFFF3B62} , 
{32'h000084F0 , 32'h0002CB7B , 32'hFFFBFE9D , 32'hFFFDF6E1 , 32'h0007E95D , 32'hFFFF309D , 32'h0001B44E , 32'hFFFBE0EF , 32'hFFFA91C9 , 32'h00014FF1 , 32'hFFFDA5B0 , 32'hFFFDB9EB , 32'h00002959 , 32'h00017EC7 , 32'h0004AE31 , 32'h00024BC4 , 32'h0003DCDE , 32'h000884E4 , 32'h0005B91C , 32'hFFFFFE1A , 32'h000BABDB , 32'hFFFCCA98 , 32'h000709C0 , 32'h00003F00 , 32'h000A1CCA , 32'h0001FB75 , 32'h00030CDC , 32'hFFFAC3BC , 32'h00055CD1 , 32'hFFFDFA94 , 32'h00076116 , 32'h00010D67 , 32'h00076550 , 32'hFFFCFF77 , 32'hFFF9B444 , 32'hFFFBCA76 , 32'h00016F59} , 
{32'hFFFFBFFA , 32'h000680CD , 32'hFFFE31C8 , 32'hFFFE6B34 , 32'hFFFF4FA6 , 32'h00045FA6 , 32'h0001BE96 , 32'h0001B662 , 32'h00042686 , 32'hFFFB37EC , 32'hFFFDE5D8 , 32'h0006AF5B , 32'hFFFFF5B2 , 32'hFFFD15D4 , 32'h0009D875 , 32'h0003B502 , 32'h0002ABA6 , 32'h00025052 , 32'h0008B33C , 32'hFFFAC55B , 32'hFFFE30AD , 32'hFFF67CCC , 32'h0000AB46 , 32'hFFFD743D , 32'h00041E02 , 32'hFFFF669C , 32'hFFF96E50 , 32'hFFFB0608 , 32'h00044217 , 32'h00051AE5 , 32'h00028776 , 32'h0007A632 , 32'hFFF9D763 , 32'hFFFEA89B , 32'h0005A2B5 , 32'hFFFF357E , 32'hFFFC3C4F} , 
{32'hFBAE7498 , 32'hFEC4BB38 , 32'h0388BEC8 , 32'h0120F838 , 32'h040613B8 , 32'h0418F850 , 32'hFBFD0700 , 32'h019DDDF4 , 32'h01FEA0D4 , 32'h01997DF8 , 32'hF9D80A18 , 32'hF7BAFE50 , 32'hFF79F32E , 32'h013376D0 , 32'h03A593F4 , 32'h030C1BA4 , 32'h05B99BF0 , 32'hFBF2E488 , 32'h015B8F90 , 32'hFD624AF8 , 32'h0C89E390 , 32'hFFE887A9 , 32'h025CEAB4 , 32'h01AC5E08 , 32'h0447C6B0 , 32'hFEE668C0 , 32'hF8C62618 , 32'h0175D3D8 , 32'hFDD248A4 , 32'hFBC650D8 , 32'h03FEDE54 , 32'h04D60490 , 32'h00EDE7EE , 32'h0AAE3B40 , 32'h0249797C , 32'hFFCEFBD3 , 32'h07B1F5F0} , 
{32'h05EFDC70 , 32'hFE06F7DC , 32'h02728CA8 , 32'hFD19BC7C , 32'hFF0EDFA2 , 32'h03698268 , 32'hFD73CF40 , 32'h007451A9 , 32'h06184AD0 , 32'h0503F588 , 32'hFF10C8FC , 32'hF8532148 , 32'h0AEA1900 , 32'h01E71B6C , 32'hFF8328BC , 32'hFC9915E8 , 32'h00FB995E , 32'hFBD76E48 , 32'hFB701550 , 32'h042EE6B0 , 32'h0D2E2AB0 , 32'h0A95B5E0 , 32'hF5A72840 , 32'h0BD35170 , 32'hF2AC8560 , 32'h04BAD0D0 , 32'hFEB241CC , 32'hEC824F40 , 32'hF70FACC0 , 32'hF5FCDD90 , 32'hF89596B0 , 32'h17202A80 , 32'hF98312B8 , 32'hFCAE7850 , 32'h0EDEC2D0 , 32'hFC610910 , 32'hF7E2BD40} , 
{32'h04727070 , 32'h018EE394 , 32'h0113401C , 32'hFDDC8574 , 32'hFF45324E , 32'h0F09F510 , 32'hFFF0D8D0 , 32'hFD02998C , 32'h0FCDF080 , 32'hFD087958 , 32'hF93D5D58 , 32'hF5B44140 , 32'h0E828A60 , 32'h05457D88 , 32'hFD65C4F8 , 32'hF7B4E9D0 , 32'hFC9C85BC , 32'hFF6FD569 , 32'hFAFDBC30 , 32'h08001A80 , 32'h0F298D40 , 32'h106F1000 , 32'hF27170F0 , 32'h12622920 , 32'hF4194B70 , 32'h09B0CFC0 , 32'hF8FA5CB8 , 32'hEFF449A0 , 32'hFB2E2B78 , 32'hF8CA1568 , 32'hFC4934AC , 32'h1504CB40 , 32'hFCF676F8 , 32'hFADE7A00 , 32'h0D9F43C0 , 32'hF95311A8 , 32'hF7EA0D80} , 
{32'h09DFAE60 , 32'h129865A0 , 32'h083E7030 , 32'hE9085160 , 32'hFA608FD8 , 32'h0B214690 , 32'hFF188ADB , 32'h12A0A320 , 32'h020E0E68 , 32'h0ECEB4C0 , 32'hF412D2A0 , 32'hD9B70800 , 32'h1F23FDE0 , 32'h0CB84EE0 , 32'hF8A5E068 , 32'h0F04CC20 , 32'h0E8628F0 , 32'hD4C49080 , 32'hE4F35920 , 32'hFF984FBC , 32'h39C69AC0 , 32'hF4D9F430 , 32'hEA174DE0 , 32'h2D621140 , 32'h088C2EE0 , 32'hF15202E0 , 32'hF5BA1E30 , 32'hF04C0050 , 32'hDFE39BC0 , 32'hE5CFE820 , 32'hF9A11A00 , 32'h13F03360 , 32'hE257E400 , 32'hFE515840 , 32'h0F1F92A0 , 32'hEA71CF60 , 32'h0182AE8C} , 
{32'h0F4A3530 , 32'h065CCF78 , 32'h05D8A428 , 32'hE28C7BA0 , 32'hFB0BCEE0 , 32'hFC34E67C , 32'h0819C210 , 32'hF696C7F0 , 32'hF7A13BB0 , 32'h18014AC0 , 32'hFD5916E0 , 32'hF3A0B6B0 , 32'h1167C4E0 , 32'hF45B5640 , 32'hEE5D24C0 , 32'h00E99326 , 32'h0DA084E0 , 32'hECE8AB60 , 32'hD3A7CEC0 , 32'h0B1B1AF0 , 32'hFFF81C24 , 32'hE6B4F680 , 32'hEF36AC20 , 32'h251B9FC0 , 32'h0A9F9960 , 32'hE732C280 , 32'h08635CD0 , 32'h1BA747A0 , 32'h0660FDA0 , 32'hEEBB5640 , 32'h040A3010 , 32'hFE5E2C04 , 32'hEAB25E80 , 32'hE87857C0 , 32'h081540F0 , 32'hFE6205D4 , 32'hFCB73EC0} , 
{32'h10B062A0 , 32'h15398100 , 32'h14C87E00 , 32'h0704C440 , 32'hDA043740 , 32'hFD558978 , 32'hF23A9240 , 32'h02460A08 , 32'h0461E7D0 , 32'h00BD4FE8 , 32'hFA533AF0 , 32'hEF804D80 , 32'h15CCFCE0 , 32'hFA994450 , 32'h01DDF6DC , 32'hF5EFCDC0 , 32'h00C78BF1 , 32'h09EF8B30 , 32'hFB3B2750 , 32'hFD66632C , 32'h1373B820 , 32'h0FBEEA10 , 32'hF79819B0 , 32'h0F2D3540 , 32'hF46CC440 , 32'h14FCF280 , 32'hFCFAA50C , 32'hE6878A60 , 32'hF8F85618 , 32'hDD2D90C0 , 32'hF9C6E8B8 , 32'h208C2A40 , 32'hF2487C50 , 32'hF7F0F160 , 32'h1BB42020 , 32'h0D98B450 , 32'hF1167830} , 
{32'h11FBEAC0 , 32'hFB41BB78 , 32'hFDBE7F40 , 32'hFC8486CC , 32'hF7596DC0 , 32'h02856AF8 , 32'hFA26D580 , 32'h0ABDB770 , 32'hEF3CA480 , 32'hF72C7590 , 32'h0079AC84 , 32'hFE9E315C , 32'hFA13C3F8 , 32'hEDD7AFE0 , 32'h123FF4C0 , 32'h03AD05C0 , 32'hFCD5FDA4 , 32'hF94A1FD0 , 32'h063368E8 , 32'h07235AE8 , 32'hFFA8D948 , 32'h0A56E900 , 32'hF84A99B8 , 32'h2438C380 , 32'hF17771F0 , 32'h115F03A0 , 32'h0038A1D5 , 32'hEAD5FF20 , 32'hFA299E78 , 32'hF5F77120 , 32'hEAFCD900 , 32'h0953FB10 , 32'hFF566603 , 32'h0A6387D0 , 32'hFCDAD56C , 32'h04B17E78 , 32'hEA771920} , 
{32'h12EE3E20 , 32'hFAD39800 , 32'h0AE57B10 , 32'hF0C80940 , 32'hECA26080 , 32'h0B4B9D70 , 32'h00F775B1 , 32'hDE716200 , 32'hF5237330 , 32'h23386000 , 32'hEF5E9400 , 32'h0D24C210 , 32'h08A92C60 , 32'hE5A062C0 , 32'h0C8B8800 , 32'hF9158568 , 32'h18B86020 , 32'h0D9B4520 , 32'hDF28DB40 , 32'h0B388320 , 32'hE702B280 , 32'hE90CD0A0 , 32'hEAA28480 , 32'h15050200 , 32'h082E2350 , 32'h04F5DC60 , 32'h0AC1C2F0 , 32'h326150C0 , 32'h0659B6C0 , 32'h06DEABC8 , 32'h0890B6D0 , 32'h08CB6330 , 32'hF7B5A800 , 32'hECEA8160 , 32'h00C0AA8E , 32'h16EC21A0 , 32'h164017C0} , 
{32'h098EDB10 , 32'h020FDC48 , 32'h173CFD40 , 32'h03784BAC , 32'hF4635100 , 32'h117386E0 , 32'hFE2AC558 , 32'h0CB250A0 , 32'hFA098660 , 32'h0E03BD50 , 32'hF8A59448 , 32'hFD91DC68 , 32'h214C0E40 , 32'h01222AE0 , 32'h0FFD1EB0 , 32'hF66374E0 , 32'h085496A0 , 32'h08D6A0D0 , 32'h16269C00 , 32'hF86DD7E0 , 32'hF7BD13A0 , 32'hF381CBD0 , 32'hFE2D5B40 , 32'h07C11A30 , 32'hF946E888 , 32'h008AE7AD , 32'hF2087BE0 , 32'h1885FB80 , 32'h03016B78 , 32'h04AB8040 , 32'hFD717A90 , 32'h0553CE60 , 32'h00C9BAAF , 32'h06162030 , 32'h04137EF0 , 32'h00AA6D3A , 32'h14FF4020} , 
{32'h0DE74050 , 32'h075FE218 , 32'hFF7DE896 , 32'h015700C4 , 32'hF9413E30 , 32'h08179DC0 , 32'h0849EA20 , 32'hFF49FF73 , 32'hF8786478 , 32'h026EE8A4 , 32'hF7236630 , 32'hF2D6F940 , 32'h0D8DACB0 , 32'h0ECD9460 , 32'hF79F88E0 , 32'h0DF3E0B0 , 32'h023E9540 , 32'hEF56CA00 , 32'hF3BBFC90 , 32'hFF6B18D3 , 32'h1524DCC0 , 32'hF9A26828 , 32'h087255B0 , 32'h15F548C0 , 32'h012C7B2C , 32'hE64E1100 , 32'h043BE0B8 , 32'h04CCC028 , 32'hF0E1F640 , 32'hF34B1730 , 32'hF18A5050 , 32'hF570B260 , 32'hEFFE4FC0 , 32'hFAD53BF8 , 32'hFE0E3828 , 32'hF51553A0 , 32'hFEA9CBFC} , 
{32'h0CC90D50 , 32'h16DA1EA0 , 32'hFF0F52E0 , 32'hF35B7710 , 32'h03AF67F4 , 32'hFD7261E8 , 32'h033EEDB8 , 32'h0BBE9CD0 , 32'hFF9107BD , 32'h015D197C , 32'hFECC922C , 32'hFCA58A24 , 32'h083E68C0 , 32'h009AFC7A , 32'hF4CFA620 , 32'h0C228BE0 , 32'h028DA994 , 32'hEA940180 , 32'hF0310CE0 , 32'h0324FC14 , 32'h177FA600 , 32'hF6DE1440 , 32'hFAD39FF8 , 32'h1567DB20 , 32'h0C91C200 , 32'hF781F380 , 32'hFD9F6CF4 , 32'h0A0B1D20 , 32'hF8499578 , 32'hF43B4720 , 32'hF66F9B70 , 32'h000F1CB0 , 32'hF6C76660 , 32'hFA331058 , 32'h00559FAC , 32'hECBF9B00 , 32'hFAE49810} , 
{32'hF91BCA10 , 32'h008FA4BE , 32'hF3805D10 , 32'hE1B3E9C0 , 32'hFE2DB810 , 32'h1198BD20 , 32'hDF07BCC0 , 32'h0DE8D9C0 , 32'hECC08EE0 , 32'h1302D120 , 32'h00796888 , 32'hF11ED270 , 32'hE7DB89A0 , 32'hEA7F9740 , 32'hFA2BD230 , 32'hFFB5B377 , 32'hFE4BCD00 , 32'h0488A908 , 32'h0EDFC5E0 , 32'h083BED40 , 32'hF4E1A7E0 , 32'h00F6D031 , 32'hDB240480 , 32'h0AE16BE0 , 32'hEF9E3A20 , 32'hE2CED260 , 32'h04547EB8 , 32'hF7B5A870 , 32'h020F6FFC , 32'h23CE3A80 , 32'hD7705AC0 , 32'hE9E1D140 , 32'h3B6DD100 , 32'h206FD900 , 32'h0C0F89C0 , 32'h15432CC0 , 32'hE0DBB740} , 
{32'hF747FCF0 , 32'h0E23C150 , 32'hEFE56CE0 , 32'h0060F378 , 32'h05FFD0D8 , 32'h038DD14C , 32'hFE0E1948 , 32'h0B46FB70 , 32'hF52C2A90 , 32'hFD244548 , 32'h0BB15C60 , 32'hF9F94460 , 32'h0479A6B0 , 32'hF8BA2AB8 , 32'h01AE3834 , 32'hFB7E44C0 , 32'hFE7BF7CC , 32'hF9EF87E0 , 32'hFA2616B0 , 32'hFD0CCC94 , 32'hFB3CB6C0 , 32'hFF316052 , 32'h01C1ACB8 , 32'h08171A00 , 32'h05BCCC50 , 32'hF8FE8AE0 , 32'hFDA27758 , 32'h089782D0 , 32'h0873E660 , 32'hFC6D106C , 32'h06D52B38 , 32'hF65D0810 , 32'h144D5520 , 32'h01131B10 , 32'hFB717A08 , 32'hFFBA20F2 , 32'h02E8931C} , 
{32'h00840C22 , 32'hFFA34899 , 32'hFF26E4E1 , 32'hFFB5A0F2 , 32'hFF73C168 , 32'hFEE25624 , 32'h003DA347 , 32'h028FA0C0 , 32'hFCFBA838 , 32'h00B14ACE , 32'hFECF40A0 , 32'hFFE3C61A , 32'h00ECA22F , 32'h0024C414 , 32'h00BA3FF5 , 32'hFF976437 , 32'hFF7C0A7A , 32'hFE599334 , 32'hFF6D0764 , 32'h00AF1062 , 32'hFEAEB5C8 , 32'h02B95BCC , 32'hFEDAF978 , 32'h035F30EC , 32'hFF5A390C , 32'hFE0DFE8C , 32'h0166730C , 32'h00379619 , 32'h01C62F00 , 32'h003F61C6 , 32'hFF4B146E , 32'hFF18B762 , 32'h0143AC78 , 32'h0110FAAC , 32'hFED6670C , 32'hFF1E2AD2 , 32'h005C9641} , 
{32'h134219A0 , 32'hFADE78C0 , 32'hFD58D0C0 , 32'hEC63A640 , 32'h0050B08A , 32'h01684698 , 32'hF9B9D6D0 , 32'h086EACA0 , 32'hE8516FA0 , 32'hEE70FC20 , 32'hF8F59F30 , 32'hFD30B048 , 32'hF906C148 , 32'hDA000B00 , 32'h0DDFCE20 , 32'hFD8F6E64 , 32'hFB9D00A8 , 32'hEE0DEA80 , 32'h07509CD0 , 32'h10C33F20 , 32'hF23E5B80 , 32'h06C7F9F0 , 32'hEEB2A8A0 , 32'h293D0980 , 32'hE2E87A60 , 32'h02995F20 , 32'hF65FE560 , 32'hE71DF200 , 32'h13871540 , 32'hFD95FE44 , 32'hD5A1B840 , 32'hFE4EA744 , 32'h03B939DC , 32'h16294A20 , 32'h06D263F8 , 32'hF7B04290 , 32'hFCCF6B3C} , 
{32'h1199B280 , 32'hFAEA5730 , 32'h0403BB70 , 32'hFD01A500 , 32'hFDBBE88C , 32'hE85AF880 , 32'hFC809D0C , 32'h110FA0C0 , 32'hD4275B80 , 32'hED8F4980 , 32'hFCF02138 , 32'hF4E7CD70 , 32'hF45ECE50 , 32'hE85DBC20 , 32'h0B1E7D60 , 32'hEFBAE6A0 , 32'h0F5EDFA0 , 32'hF712BE00 , 32'h15294080 , 32'h04728260 , 32'hF59F2C30 , 32'h19984020 , 32'hF712AE50 , 32'h282C52C0 , 32'hFB8641A0 , 32'hFD0A85DC , 32'hFFBDED56 , 32'hF2939290 , 32'h07563E30 , 32'hF95FA0D0 , 32'hEEAE2960 , 32'h01C7E2EC , 32'h0DDB3C80 , 32'h1762F2E0 , 32'hE8109FA0 , 32'hFA8C3B68 , 32'hF35D36F0} , 
{32'h0010F7BF , 32'hFFE28169 , 32'h0010347F , 32'h0004EF3C , 32'h00074980 , 32'hFFE85E6A , 32'h0000661D , 32'hFFF1BD20 , 32'hFFDA07E2 , 32'hFFDDD483 , 32'h0023FB94 , 32'hFFFE995B , 32'hFFFD5616 , 32'hFFF9C2F6 , 32'h002B4C32 , 32'hFFF31452 , 32'h00141B43 , 32'hFFEE09EC , 32'hFFFCA79B , 32'hFFC01A92 , 32'hFFFE54AD , 32'h00283ABE , 32'hFFFFA6A1 , 32'h0012B737 , 32'h0041E8C4 , 32'hFFC67FF6 , 32'hFFDF9887 , 32'h0006E35E , 32'h002CE277 , 32'hFFE94781 , 32'h00144404 , 32'h00181417 , 32'h0028C83B , 32'h000D7D0F , 32'hFFED2838 , 32'hFFEB92AB , 32'hFFF5608B} , 
{32'h004498F9 , 32'hFF85F435 , 32'h004E7593 , 32'hFFC60DA7 , 32'hFFDA9633 , 32'hFFAD04F3 , 32'hFFAA6575 , 32'h001A4CC7 , 32'hFF066186 , 32'hFF107DBF , 32'h008EEDD6 , 32'h00350241 , 32'h00619D33 , 32'h00160928 , 32'h00C7205C , 32'hFFF04D7C , 32'h006EC129 , 32'hFFF22EB8 , 32'hFFBA3CB9 , 32'hFFEF2C41 , 32'h001FFF81 , 32'h00C3919B , 32'hFF458CFB , 32'hFFD1AAEA , 32'h008EA855 , 32'hFFD9C8C9 , 32'hFF68D771 , 32'h00615B2E , 32'h006F500B , 32'hFF8B5212 , 32'h002199BD , 32'h0030A2F7 , 32'h008D17C5 , 32'h002CBEF7 , 32'hFF30700F , 32'h008373D6 , 32'hFF73F4AC} , 
{32'h003F0A62 , 32'hFF812D13 , 32'h004CE872 , 32'hFFBE38BD , 32'hFFC25A71 , 32'hFF95F467 , 32'hFF9D3E76 , 32'h0014EDE0 , 32'hFEE0E3C4 , 32'hFEF9CAD8 , 32'h00A0024B , 32'h00580601 , 32'h007D508F , 32'h003973AE , 32'h00E999FB , 32'hFFF924F3 , 32'h00730DA3 , 32'h00041C0A , 32'hFFA34589 , 32'hFFF6633B , 32'h0031C35A , 32'h00E3EA09 , 32'hFF2BDAAB , 32'hFFA9CD13 , 32'h009EC5FA , 32'hFFE10A1A , 32'hFF5C270F , 32'h007F6217 , 32'h006BFD85 , 32'hFF892AC7 , 32'h001D84EE , 32'h0046156F , 32'h00899A48 , 32'h003BFDB4 , 32'hFF29353A , 32'h0089DC6B , 32'hFF6C45C6} , 
{32'hFFFE3B53 , 32'hFFFCA5FD , 32'hFFF81413 , 32'hFFFF5233 , 32'h00019986 , 32'h0002D01D , 32'hFFFF71E1 , 32'h00003557 , 32'hFFFFB972 , 32'h0000AEB6 , 32'hFFFECAED , 32'h000012F4 , 32'hFFFB9009 , 32'h00026357 , 32'h000068C6 , 32'hFFFD0173 , 32'h00032A64 , 32'hFFFE90E7 , 32'h00072489 , 32'h000193FD , 32'hFFFF74AA , 32'hFFFA1F03 , 32'h000765A2 , 32'h000C6C80 , 32'hFFFE62EA , 32'h000659E6 , 32'hFFFF5410 , 32'hFFFB4353 , 32'h0003EA8D , 32'hFFFDF9E7 , 32'h00042950 , 32'hFFF9CEE3 , 32'hFFFA9341 , 32'hFFFF34DB , 32'hFFFCE362 , 32'hFFFD464E , 32'hFFF6F8D0} , 
{32'hFFFF650A , 32'h0002EE53 , 32'hFFFCDBFE , 32'h00049238 , 32'h00016591 , 32'hFFFEF408 , 32'hFFF9ED0C , 32'hFFFDA11F , 32'h000497F7 , 32'h00072F7E , 32'hFFF6C087 , 32'hFFFB15C8 , 32'hFFFB5238 , 32'h0000C23E , 32'h0005D90B , 32'h0000071E , 32'hFFFA6449 , 32'h000A4B22 , 32'h0000B756 , 32'h0008994F , 32'hFFFEAB3A , 32'h0003A78C , 32'hFFF7910A , 32'hFFFEDEE2 , 32'h0000DE60 , 32'h00003858 , 32'hFFF5D318 , 32'hFFFE4150 , 32'hFFFC0D4D , 32'hFFFBC3EB , 32'h000202A6 , 32'hFFFB30CF , 32'hFFFF5A57 , 32'h0001C548 , 32'hFFF3A615 , 32'hFFFCC7EC , 32'hFFFA55C8} , 
{32'h00072433 , 32'h0002DCB3 , 32'hFFFD2F47 , 32'h00010DD5 , 32'hFFFE4DCB , 32'hFFFF24D1 , 32'h0007BDCE , 32'h0002B262 , 32'hFFFD4F6B , 32'hFFFFEAF4 , 32'hFFFF305A , 32'h00079D26 , 32'hFFFF29CD , 32'hFFFFD3F8 , 32'hFFFD9C88 , 32'hFFFB935D , 32'h00035B4C , 32'hFFF8771D , 32'hFFF9D325 , 32'h000278C9 , 32'h00018750 , 32'h0000B74B , 32'h0001C652 , 32'h000051CD , 32'h00022B64 , 32'h0004829D , 32'h0005A980 , 32'hFFFF3AEF , 32'hFFFE4C36 , 32'hFFFE926A , 32'h00094404 , 32'hFFFAD9AE , 32'h0001D2EB , 32'h0001204D , 32'hFFFE8D14 , 32'h000BB55A , 32'h000A1814} , 
{32'h00002443 , 32'hFFFD6433 , 32'h00020D7E , 32'hFFFF2FC9 , 32'h0001046C , 32'hFFFF8930 , 32'hFFFDF42A , 32'hFFFB2F46 , 32'hFFFA3519 , 32'h0006BFB7 , 32'hFFF9A4ED , 32'h000687DD , 32'hFFFD22C3 , 32'hFFFB41C8 , 32'h000028A9 , 32'h0007EE7D , 32'h00068FF3 , 32'hFFFA3859 , 32'h0003E005 , 32'hFFFE6783 , 32'hFFFAC2DF , 32'h000D4124 , 32'hFFF3C8A7 , 32'hFFFF5B8A , 32'hFFFD7070 , 32'h00007341 , 32'hFFFBD04A , 32'h0000298B , 32'h000191D3 , 32'h0001F487 , 32'h00077661 , 32'hFFFDB02D , 32'hFFF95354 , 32'h0002357A , 32'hFFFB12D0 , 32'h000653F8 , 32'h00029E8E} , 
{32'h0004FCF6 , 32'h00035E10 , 32'hFFFC4D7B , 32'hFFF99AE7 , 32'hFFFFFB8C , 32'hFFFE3189 , 32'hFFF9D191 , 32'hFFF88841 , 32'hFFF0ACEE , 32'h0002FBFF , 32'h00086C06 , 32'h0003E903 , 32'h000270A0 , 32'h000278EB , 32'hFFFD5C9C , 32'hFFFE38EC , 32'h0000CFD7 , 32'hFFFD161A , 32'h0003D794 , 32'h00065458 , 32'hFFFCBF6D , 32'hFFFD1EE2 , 32'h0002F195 , 32'hFFFF1515 , 32'hFFFE917A , 32'hFFF9A077 , 32'h0012D48D , 32'hFFFBC5EE , 32'h0001B019 , 32'hFFFFB66B , 32'hFFFB5C9B , 32'hFFFB7473 , 32'h0001933F , 32'hFFFCA41E , 32'h0004591D , 32'h0001528C , 32'hFFF8067C} , 
{32'h0000A796 , 32'h00004DF2 , 32'h0001B0D5 , 32'hFFFD17E7 , 32'hFFFFAE38 , 32'h00061C20 , 32'hFFF76B65 , 32'h0001347E , 32'h000E5866 , 32'hFFFC6AEB , 32'hFFF7B00C , 32'h0000B619 , 32'h000425FE , 32'h0003CB1E , 32'h000124CB , 32'h00028F71 , 32'h0001A34C , 32'hFFFF165B , 32'h0001F85B , 32'hFFFCBC53 , 32'h0005FB8C , 32'h0000D637 , 32'hFFFEB785 , 32'h0009A708 , 32'h00036054 , 32'hFFFA43FF , 32'hFFFD4314 , 32'h00005CFC , 32'h0003E7DC , 32'h0006E135 , 32'h000B47DF , 32'hFFFF41AB , 32'h000136C1 , 32'h0007A001 , 32'h0004235F , 32'h00086C0A , 32'h00034E91} , 
{32'h00054381 , 32'h000981AF , 32'hFFFF4C18 , 32'h00069AB9 , 32'h00020B0F , 32'h000155FB , 32'h0001037D , 32'h00063A18 , 32'hFFFB67A4 , 32'h000B6D04 , 32'h00059FE1 , 32'hFFFEFB7C , 32'hFFFD3423 , 32'h0001D219 , 32'hFFFCB818 , 32'hFFFBCEBA , 32'h00044452 , 32'hFFFE5B4E , 32'hFFFEA72E , 32'h0004F571 , 32'h00048528 , 32'hFFF9B301 , 32'h0001C8C6 , 32'h000217FA , 32'h000926F0 , 32'hFFFFB449 , 32'hFFFFA964 , 32'h0000C003 , 32'hFFFA99C9 , 32'hFFFDB33D , 32'h0002EFDA , 32'h00032485 , 32'h0002B3DB , 32'hFFFE9626 , 32'hFFFD9130 , 32'hFFFD8ED8 , 32'h00053EB8} , 
{32'h0001474F , 32'hFFFD95E9 , 32'hFFFB6AC9 , 32'hFFFCA263 , 32'h000218E1 , 32'hFFF9F1D6 , 32'hFFFBEAB3 , 32'h0002FE21 , 32'hFFFFDCB2 , 32'hFFFF36CA , 32'h0004264F , 32'hFFFCDBC7 , 32'hFFF9C55E , 32'h0007DAF4 , 32'hFFF8F628 , 32'h00017071 , 32'hFFFAF8FF , 32'hFFF694F2 , 32'h0000D067 , 32'hFFFF3FD2 , 32'hFFF8A403 , 32'hFFF6C9E8 , 32'h00069A09 , 32'hFFF73044 , 32'hFFFF3C7E , 32'h00049AC3 , 32'hFFF63E9E , 32'hFFF9DEF6 , 32'h0001E885 , 32'hFFFAB2AF , 32'h0002E310 , 32'h000BCCAC , 32'hFFFC7D31 , 32'h00084B77 , 32'h00002761 , 32'hFFFBB8FB , 32'h00043AB3} , 
{32'h00085F36 , 32'hFFFB08E7 , 32'h0004B4FE , 32'h0002421C , 32'hFFFA1804 , 32'h0001D9C7 , 32'hFFFFC67B , 32'hFFFD5C66 , 32'h00040270 , 32'h00010D67 , 32'h000465B1 , 32'hFFFD6B76 , 32'h00043407 , 32'h00000198 , 32'h0001D1F3 , 32'h0001968E , 32'h0000CD35 , 32'h00005B73 , 32'h0004E3E7 , 32'h000387DF , 32'h0001427E , 32'h00037396 , 32'hFFFDD548 , 32'hFFF65D41 , 32'h00053D15 , 32'hFFFDD616 , 32'h0004F86E , 32'hFFFF75B5 , 32'h0000FCDD , 32'h00049573 , 32'h00067642 , 32'hFFFD84D6 , 32'hFFFD1093 , 32'h00014740 , 32'hFFFE7F91 , 32'hFFFDB25B , 32'hFFFFDE7C} , 
{32'h0016BCD5 , 32'hFFE28315 , 32'hFFD6A730 , 32'h00452EEB , 32'hFFEC48D5 , 32'hFFE3D022 , 32'h00010D03 , 32'h0077B9F5 , 32'h00485D55 , 32'h0020A17C , 32'hFF7B2A4B , 32'hFFC6A17B , 32'hFFC1C866 , 32'hFFD05EA7 , 32'hFFD29C1F , 32'hFFF85FA4 , 32'hFFEBD2CF , 32'hFFFDA8CF , 32'h002C269F , 32'h00361BB5 , 32'hFFE253FB , 32'hFFE39B52 , 32'hFFFB0CED , 32'h000B191B , 32'hFFF4F635 , 32'hFFFAC449 , 32'h000AE344 , 32'hFFF82526 , 32'h001EE36A , 32'hFFF982CA , 32'h0015F9C2 , 32'h00038017 , 32'hFFF4881B , 32'hFFDF463F , 32'h001C47F1 , 32'h0008617A , 32'h00171F22} , 
{32'h001325B3 , 32'hFFE2375F , 32'hFFDC333E , 32'h0049797A , 32'hFFE37D3A , 32'hFFE7B3E5 , 32'h000B3984 , 32'h00753940 , 32'h004E2793 , 32'h0028689B , 32'hFF7FCB85 , 32'hFFCF4B55 , 32'hFFC76F98 , 32'hFFCFAF1A , 32'hFFD4744B , 32'h00013585 , 32'hFFE9A099 , 32'hFFFDD107 , 32'h00272F60 , 32'h002FED8D , 32'hFFDD9153 , 32'hFFEA2869 , 32'hFFF2DEEB , 32'h001561E5 , 32'hFFF7BB43 , 32'hFFFCA5C7 , 32'h0002AD30 , 32'hFFF9C730 , 32'h0019305D , 32'hFFFD586F , 32'h0018E5A0 , 32'h00031867 , 32'hFFF2E205 , 32'hFFDDF9A6 , 32'h0017F755 , 32'h0009F51F , 32'h0020B4E5} , 
{32'hFFFC14C9 , 32'hFFFC574E , 32'h00064991 , 32'hFFFEB52C , 32'h000243FB , 32'hFFFB81B5 , 32'hFFFEA4FF , 32'hFFFA441B , 32'h000690C3 , 32'hFFFE36C6 , 32'h0002338D , 32'h000389D6 , 32'hFFFEB2BF , 32'hFFFC33C6 , 32'h0000013A , 32'hFFFFA78A , 32'h0002759B , 32'h0007FA63 , 32'h0003089A , 32'hFFFC8037 , 32'hFFFBE56F , 32'hFFF90A66 , 32'h0004508D , 32'hFFFFD9B6 , 32'hFFFD5C26 , 32'hFFF3FE40 , 32'hFFFE0BA4 , 32'hFFFB6A9F , 32'hFFFA2F0A , 32'h00036E75 , 32'hFFF97C3A , 32'h0008436C , 32'h0008E2B8 , 32'h00027793 , 32'hFFFEEBA0 , 32'h000413CD , 32'hFFFC8B2A} , 
{32'hFFF6FD82 , 32'hFFFB0386 , 32'hFFFD5DBD , 32'hFFF732C9 , 32'hFFFE100B , 32'hFFFFBDCF , 32'h000D6846 , 32'hFFFE11C6 , 32'hFFF75C15 , 32'hFFFC9112 , 32'h0003A052 , 32'h0006121D , 32'hFFFB72DF , 32'hFFF9EDC4 , 32'h000111E0 , 32'h0004845B , 32'h00040DB9 , 32'h0003DD1C , 32'hFFF6B2F8 , 32'h000788F8 , 32'hFFFB0FB6 , 32'h0009515C , 32'hFFF49485 , 32'hFFF4E36E , 32'h0004C5AC , 32'hFFF42D3D , 32'h000A0DC5 , 32'hFFFA29FC , 32'hFFF965CE , 32'hFFF9336A , 32'h00020B79 , 32'h00024841 , 32'h00034329 , 32'h00014F76 , 32'hFFFDD483 , 32'h000370D9 , 32'h000187E3} , 
{32'h000A16A8 , 32'h000DE13D , 32'h000E5CA6 , 32'hFFF7B751 , 32'h000F11F2 , 32'hFFED200C , 32'h000C09A9 , 32'h0006B002 , 32'hFFF9D365 , 32'h000AF081 , 32'hFFFDA587 , 32'h0004B9F5 , 32'hFFF23ED3 , 32'h0005A42D , 32'h000B9F97 , 32'h0011CC12 , 32'hFFF426AD , 32'h001B2FDB , 32'h0005CB21 , 32'hFFF6D3FB , 32'h000D48B2 , 32'hFFF5FED0 , 32'hFFF4B29B , 32'h0003B001 , 32'h000B5FF5 , 32'hFFFDE161 , 32'hFFF4B514 , 32'h0009AE6F , 32'hFFF0FF17 , 32'hFFF9FA29 , 32'hFFFE1A48 , 32'hFFF836EF , 32'hFFFCB57B , 32'hFFF9D2A6 , 32'hFFEF65B8 , 32'h000EE298 , 32'h00024B53} , 
{32'h141E05E0 , 32'hF9A590E0 , 32'hFC7D0A70 , 32'hF801F6A8 , 32'hFE838510 , 32'h0665DDB8 , 32'hF7E4A890 , 32'h07381760 , 32'hF0C09880 , 32'hF2E638B0 , 32'h02846E0C , 32'hF7705310 , 32'hF6130770 , 32'hE8D2B8A0 , 32'h0A657C70 , 32'h02AB39A4 , 32'hFC931ABC , 32'hF5426110 , 32'h08732790 , 32'h05658EA8 , 32'hF5538FB0 , 32'h05075380 , 32'hF34CE500 , 32'h243FE2C0 , 32'hEB584840 , 32'h044042D8 , 32'h0010E433 , 32'hE6F584C0 , 32'h0729BD48 , 32'hFF3E90F9 , 32'hE7907C60 , 32'h012C1CDC , 32'h08223F90 , 32'h15C76740 , 32'hF8CB7EE0 , 32'h0076A1B6 , 32'hF30D7BD0} , 
{32'hFF251FE0 , 32'hFFD6AFFD , 32'hFE99DE64 , 32'h0024664A , 32'hFE9D4488 , 32'hFEF0EE9C , 32'h0008BBE2 , 32'hFF1D8915 , 32'h0046D58E , 32'hFED29388 , 32'h000340C0 , 32'hFF36643A , 32'h00194E49 , 32'h0065BB52 , 32'h00E22FB6 , 32'hFF7BCB13 , 32'h00A23192 , 32'h00121A00 , 32'h009D1E04 , 32'h00792C82 , 32'hFF9E599C , 32'h005B8938 , 32'hFF68F5F8 , 32'h0160325C , 32'h004FAACB , 32'hFFD5EF27 , 32'hFE241584 , 32'h000EBD39 , 32'h00AE1768 , 32'hFFFF51F6 , 32'h01375CD8 , 32'h005E71D6 , 32'hFFBDA5E3 , 32'h0080DDBD , 32'hFF170571 , 32'hFF5DAFE6 , 32'h0036C2B2} , 
{32'hFFB00EF8 , 32'hFFA51D72 , 32'hFFACE80C , 32'h0008A1E7 , 32'hFF8FBFCE , 32'hFFEB5902 , 32'h00640CE1 , 32'hFFE42FF7 , 32'h00050FAE , 32'hFFA441AF , 32'hFFE565B5 , 32'hFFDCAD2C , 32'h003E136A , 32'h0021DC5E , 32'hFFDB5AB1 , 32'hFFA61BDF , 32'h0020A146 , 32'hFFF001FB , 32'h003ED48D , 32'h000D3944 , 32'hFFF7A1F3 , 32'h007C485E , 32'hFFC7164B , 32'h004AE21C , 32'h003C5AB4 , 32'h00046CFE , 32'hFFAB7208 , 32'h0011C3B7 , 32'h006A3B42 , 32'h000758DF , 32'h00375A3E , 32'h000DAB30 , 32'h001AEBB8 , 32'h0026D6F6 , 32'hFFC8806A , 32'hFFDC8411 , 32'h001A1CD4} , 
{32'h100FD940 , 32'hFBC0AA30 , 32'hFED436FC , 32'hFAD27908 , 32'hFF2FE5D5 , 32'h06CFD4B8 , 32'hF9FFB070 , 32'h05E52E80 , 32'hF4CFA560 , 32'hF779BB60 , 32'h02EBCC80 , 32'hFA743670 , 32'hF8F92AF8 , 32'hEE6F6280 , 32'h0814D550 , 32'h01B41818 , 32'hFE7D0070 , 32'hF7C1DE40 , 32'h0637AC68 , 32'h045A3AB8 , 32'hF7956120 , 32'h023ED978 , 32'hF6F24090 , 32'h19C4E600 , 32'hEF373DA0 , 32'h02F11940 , 32'h01287FBC , 32'hECB30D20 , 32'h04C8BC40 , 32'hFE03342C , 32'hECFEE8A0 , 32'h0156D088 , 32'h06AAEE88 , 32'h0FE71D90 , 32'hFA229E08 , 32'h00B4AC3B , 32'hF7423560} , 
{32'h04EA5E50 , 32'hFEA5FA14 , 32'h00BFBBCF , 32'h0331A0D8 , 32'h04117E18 , 32'h0B3C9540 , 32'hF931F158 , 32'hFB7B0F90 , 32'hFFE60374 , 32'hFDF1EDB8 , 32'hFE80DE48 , 32'h08443B60 , 32'h11A24800 , 32'hE7DC2300 , 32'hF7F3BA80 , 32'hF5897EE0 , 32'h16E902C0 , 32'hF7738030 , 32'hF745B740 , 32'h162E83A0 , 32'hFFB96871 , 32'h078E31B8 , 32'h079B1FF8 , 32'hFD89A9FC , 32'hFAB5D6E8 , 32'h031D426C , 32'h08B69C50 , 32'hFBDD2600 , 32'h01DF5EC0 , 32'h06051AE8 , 32'hFD3D9808 , 32'h0AD459B0 , 32'h05C655C8 , 32'hFF6B127F , 32'h05855C68 , 32'hE767B640 , 32'hFF1108C7} , 
{32'h007E5C3E , 32'h00015AE8 , 32'h00575911 , 32'h004A9A1F , 32'h0227D1C0 , 32'h02034258 , 32'hFEEB2BB4 , 32'hFDCF4458 , 32'h0095B0F6 , 32'h00893929 , 32'h01097ED4 , 32'h013E9134 , 32'h018F9FA0 , 32'hFDCC13A8 , 32'hFF2E832A , 32'h0051DB3A , 32'hFF8464ED , 32'hFF59C61E , 32'h00AD1F6C , 32'h00F53DFC , 32'h016D5E24 , 32'h0000649F , 32'h003D4807 , 32'hFE554FE0 , 32'hFF4029F8 , 32'hFF4A584C , 32'h02571648 , 32'hFDA96508 , 32'hFFD02678 , 32'hFF738786 , 32'hFE464C28 , 32'h0065D2AB , 32'h022FB95C , 32'hFF9F593B , 32'h02D6DD90 , 32'hFE39C930 , 32'h01BE35F4} , 
{32'hFEFD0B98 , 32'h01126BA4 , 32'hFFF10606 , 32'hFB1FFE28 , 32'hFFB77A81 , 32'h00BEAAF8 , 32'hFE100888 , 32'hFE6EFEF0 , 32'hF90C2FB8 , 32'hFD5599D4 , 32'h00349AAE , 32'h003E4EDA , 32'hFFCDFCB5 , 32'hF1F0CBE0 , 32'h02D35848 , 32'hFAA89100 , 32'h00311737 , 32'hF9FC7BB8 , 32'h034EDB64 , 32'h0C79B2F0 , 32'hFDFEB280 , 32'h001C7042 , 32'hFE664720 , 32'h0C144B80 , 32'hF03E4CA0 , 32'h033DED44 , 32'hF8723F40 , 32'hF36007C0 , 32'h03775728 , 32'h01DEA9C4 , 32'hF4FDF550 , 32'h00537513 , 32'hFE2E63A8 , 32'hFFC1BD50 , 32'h082F2BD0 , 32'hFDF9FF48 , 32'h0A466410} , 
{32'h104CB360 , 32'hFB19C9E8 , 32'hFE0FFDCC , 32'hF99FB140 , 32'hFF77461C , 32'h05B080B0 , 32'hF9A25B08 , 32'h06221D38 , 32'hF3D38E00 , 32'hF6720460 , 32'h0223C024 , 32'hF9BFB980 , 32'hF7B7F2E0 , 32'hED7F8F00 , 32'h08107E20 , 32'h028ED908 , 32'hFCDD17F0 , 32'hF78E3060 , 32'h0642E6F0 , 32'h04285418 , 32'hF7C53510 , 32'h03724434 , 32'hF63062A0 , 32'h1C13D1E0 , 32'hEF402AE0 , 32'h0386EC10 , 32'h00E07B90 , 32'hEC0FD620 , 32'h0548D890 , 32'hFF89246D , 32'hEC305E20 , 32'h00EAA19D , 32'h06930EA8 , 32'h10F52AE0 , 32'hFAD0F1F8 , 32'h006EE059 , 32'hF5C71020} , 
{32'h16B36260 , 32'hF9250E10 , 32'hFD4C7E64 , 32'hF700BAA0 , 32'hFF2FAE32 , 32'h06FEE938 , 32'hF7448DE0 , 32'h08920990 , 32'hEEA99360 , 32'hF3E648A0 , 32'h02832208 , 32'hF79766A0 , 32'hF4F01C90 , 32'hE70E29C0 , 32'h0B5FAA20 , 32'h0238DDCC , 32'hFBFA1150 , 32'hF4D2E4A0 , 32'h0809FF30 , 32'h05CD4FE8 , 32'hF45FD4D0 , 32'h05E2FAD8 , 32'hF1F327B0 , 32'h26F08B00 , 32'hEA3014E0 , 32'h02BDBEA4 , 32'h026C8944 , 32'hE682B520 , 32'h08D0BA30 , 32'hFFD2563D , 32'hE5E11FC0 , 32'h01917094 , 32'h0933FF80 , 32'h164AB160 , 32'hF7BB3060 , 32'hFF871331 , 32'hF34DEB50} , 
{32'h021C3138 , 32'h00123CF6 , 32'hFFBADB54 , 32'hFF6FC5A9 , 32'h00572061 , 32'hFF5019C6 , 32'hFF866854 , 32'h00512552 , 32'hFE337CF8 , 32'h0056744A , 32'hFF2F581F , 32'h00327A8B , 32'hFF95BAA3 , 32'hFEBFE118 , 32'h00D25CA9 , 32'hFE7A8E4C , 32'h0082D730 , 32'h00478450 , 32'h000203B4 , 32'h007389A1 , 32'hFEF71F2C , 32'h01DAC4D0 , 32'hFE6B7D34 , 32'h02BCD660 , 32'h003B286F , 32'hFDF002F8 , 32'h0107E250 , 32'h0041BB33 , 32'h021F9B8C , 32'h00077932 , 32'hFF1F43AF , 32'h0108C1A4 , 32'h00FCDA99 , 32'hFFA2A009 , 32'hFE0133B0 , 32'hFE6EFF40 , 32'h0078D047} , 
{32'h01074EF0 , 32'h002537F6 , 32'h00259C25 , 32'hFF916015 , 32'h00370FB9 , 32'hFFA01DAA , 32'hFFBF6725 , 32'h0027FA7B , 32'hFF374385 , 32'h003F4F8B , 32'hFFD4AFD1 , 32'h0042D43E , 32'hFF88A11F , 32'hFF6BC2D4 , 32'h00909DF9 , 32'hFF3675E8 , 32'hFFF43AAE , 32'h0004AB71 , 32'h003C23E8 , 32'h0002700E , 32'hFF81DC55 , 32'h008FCD1F , 32'hFF344B21 , 32'h017608AC , 32'h003A6AB8 , 32'hFF31EDF6 , 32'h004ADB68 , 32'h00072110 , 32'h0171B264 , 32'hFFCF4F94 , 32'hFF663604 , 32'h003FA8B1 , 32'h001B3036 , 32'hFFF1B995 , 32'hFF5DCAE9 , 32'hFF9DD982 , 32'hFFE6C1C7} , 
{32'hFFFFA6DF , 32'h0000E3ED , 32'hFFF91128 , 32'h0001F179 , 32'hFFFFE639 , 32'hFFFD7991 , 32'h000207E9 , 32'h0000EE39 , 32'h00012691 , 32'h00055DA0 , 32'hFFF86654 , 32'h0001CEB5 , 32'h0000475A , 32'hFFFF6810 , 32'hFFFAC697 , 32'h0004DE46 , 32'hFFFB8BE3 , 32'h0003C5EB , 32'h00042526 , 32'hFFFEA5B7 , 32'hFFF7FA50 , 32'hFFFCCD82 , 32'h0005092D , 32'hFFFF5593 , 32'h0004D86B , 32'hFFFF5620 , 32'hFFFC1251 , 32'h00032D6D , 32'h00015E8E , 32'h0000490F , 32'hFFFC549B , 32'h0004C414 , 32'hFFFDEB57 , 32'h0001B04A , 32'hFFFF98BD , 32'h0007CC17 , 32'h00035F16} , 
{32'h00031A4D , 32'hFFFF2BC5 , 32'h0004C1A2 , 32'hFFF64844 , 32'h000209B6 , 32'hFFFF7873 , 32'hFFFE7AC6 , 32'hFFF8EA4D , 32'h000701B8 , 32'hFFFC399C , 32'hFFFC99B3 , 32'hFFFBB7BD , 32'h00002DDC , 32'h00006F75 , 32'h00044A0E , 32'h00036908 , 32'hFFFC3661 , 32'hFFFDDAD3 , 32'h0004B1B9 , 32'h0004760B , 32'hFFF9A0E3 , 32'h00086325 , 32'h0002940F , 32'h000501DA , 32'h00050592 , 32'hFFFC012A , 32'h0005E849 , 32'hFFF3F115 , 32'h00086C30 , 32'h0002E79D , 32'h000174AE , 32'h000698C5 , 32'hFFF8B640 , 32'h0006E7A2 , 32'hFFFFA0ED , 32'hFFF59744 , 32'h0002F65E} , 
{32'h00049450 , 32'hFFFD61B4 , 32'hFFFF3769 , 32'hFFFF9AD6 , 32'h0009CA9B , 32'h00026EF4 , 32'h0001E8EC , 32'h0001CCB5 , 32'hFFFD2074 , 32'h000DBD52 , 32'h0000DF47 , 32'h0001475E , 32'h000250F3 , 32'hFFFF87C6 , 32'h00015AAA , 32'hFFFD2A30 , 32'h00088883 , 32'hFFFC8DCE , 32'h00032435 , 32'hFFFCF356 , 32'hFFFF5F48 , 32'hFFFE8765 , 32'h0008C9A3 , 32'h00001AF6 , 32'hFFFE5825 , 32'h00004F91 , 32'hFFFDA7F2 , 32'h000069BD , 32'hFFFFCE1F , 32'h00054FE5 , 32'h0001B31D , 32'hFFFCA869 , 32'h00027E39 , 32'h0005405F , 32'h00088A44 , 32'hFFFDC111 , 32'h00003A78} , 
{32'h0004245C , 32'h00000E3E , 32'h00019F37 , 32'h000034ED , 32'hFFFCF00E , 32'hFFFFC2F4 , 32'hFFF86E2B , 32'hFFF4F011 , 32'h000477E9 , 32'hFFF8CE23 , 32'hFFFEF54E , 32'h0002D241 , 32'h000D803F , 32'h0000BA86 , 32'h0001342C , 32'h000508FD , 32'hFFFDE797 , 32'hFFFB8C6E , 32'h000494F8 , 32'h0000BE22 , 32'hFFFF1B6F , 32'h00059CD6 , 32'h00032A26 , 32'hFFFBB585 , 32'h00019E0A , 32'hFFFB3C1B , 32'hFFFB112F , 32'h00028955 , 32'hFFFEF5A5 , 32'h0003B486 , 32'h00034259 , 32'h00031CA7 , 32'hFFF8F431 , 32'h00050654 , 32'h000CAF5D , 32'h00067651 , 32'h00016CF2} , 
{32'hFFFE9E55 , 32'hFFFE4D10 , 32'h0001BE45 , 32'hFFF646EB , 32'hFFF2442B , 32'h0000D1D4 , 32'h0001E73D , 32'hFFFFE90D , 32'h0009008E , 32'hFFFEA3FD , 32'h0003A3DE , 32'h00041620 , 32'h0003F8B6 , 32'h0003B2A8 , 32'h0003637C , 32'h0005E368 , 32'h000A1E81 , 32'h00051AA9 , 32'hFFFEBAAD , 32'h0005EF14 , 32'hFFFCC967 , 32'h000382DC , 32'hFFFEF1D9 , 32'h0009AC16 , 32'h00014D84 , 32'h000871DA , 32'hFFFAFD4C , 32'h0000E1BC , 32'h000492D8 , 32'h0000E52C , 32'hFFFDFA34 , 32'hFFF9F9D6 , 32'hFFFB8B0C , 32'hFFF8026D , 32'h00047552 , 32'h0004CC65 , 32'hFFFE3434} , 
{32'hFFF67844 , 32'h00032B58 , 32'hFFFF98EF , 32'hFFF515AE , 32'hFFFFFF4B , 32'hFFFE565E , 32'hFFFE47C7 , 32'hFFFCE858 , 32'h000132E9 , 32'h0002946C , 32'h00080268 , 32'hFFFC5370 , 32'hFFFEDA03 , 32'hFFF76840 , 32'hFFFA2DAF , 32'h00021FD4 , 32'hFFFE5217 , 32'h00020F2F , 32'h00006061 , 32'hFFFFB66C , 32'hFFFF9B55 , 32'hFFF92161 , 32'h0009487A , 32'hFFF9722C , 32'h0002BD65 , 32'hFFFEBC2A , 32'h0003058D , 32'h0002E790 , 32'hFFFA365D , 32'hFFFCD1B2 , 32'h0001B767 , 32'h0002374B , 32'hFFFA3036 , 32'h0005F64D , 32'hFFF94266 , 32'h000435E6 , 32'h0004F648} , 
{32'hFFFB8D7E , 32'hFFF73489 , 32'hFFF972AC , 32'hFFFB7F9A , 32'h00013949 , 32'h0009F09E , 32'hFFFEB886 , 32'hFFFD0DCB , 32'h00050330 , 32'hFFFE1DE0 , 32'hFFFE151E , 32'h0001CF72 , 32'hFFF853D1 , 32'h00028B94 , 32'h0002143B , 32'hFFFA680D , 32'hFFFE5E2F , 32'h000293DA , 32'h00002343 , 32'h00038267 , 32'h0007A3F4 , 32'hFFFF5336 , 32'hFFF99A8E , 32'h000192A6 , 32'hFFF76394 , 32'h000F4B1C , 32'hFFFC2A0E , 32'hFFFE6C79 , 32'hFFFC76DE , 32'hFFF690AD , 32'hFFF7163C , 32'h0001AA18 , 32'h0003EC03 , 32'hFFFF0580 , 32'h0002C384 , 32'hFFFAF8B1 , 32'hFFF60C5B} , 
{32'hFFFB84BF , 32'hFFF82E4A , 32'h00028139 , 32'hFFFFAAAB , 32'h00062A65 , 32'hFFFB6F52 , 32'hFFFABC7D , 32'hFFFCC269 , 32'h000523A3 , 32'h00061953 , 32'h000081F2 , 32'hFFF76BEE , 32'hFFFC732C , 32'h0000D3C7 , 32'h0002BEC5 , 32'hFFFB199D , 32'h0003CDDC , 32'h0000CF3D , 32'h00028D7A , 32'h00049510 , 32'h0003F942 , 32'h000540B0 , 32'hFFFABCEF , 32'hFFFF0BB0 , 32'hFFFFB3DA , 32'hFFFE7458 , 32'hFFFFBB9E , 32'h00063F26 , 32'h0004165B , 32'hFFFD8480 , 32'h000804EB , 32'h0007E8AF , 32'h00025569 , 32'h00058A4D , 32'hFFF7A590 , 32'hFFFD1695 , 32'h000CD827} , 
{32'hFFFED7CE , 32'hFFF90E70 , 32'h00061C89 , 32'h0006E69A , 32'hFFFF83E0 , 32'hFFFFEEA9 , 32'h00092A09 , 32'h000B919D , 32'hFFFE59FE , 32'hFFFD400A , 32'h0005F116 , 32'hFFFA31B6 , 32'h00028F11 , 32'h0003CF62 , 32'h00104AF6 , 32'hFFFBBE78 , 32'h00000CFB , 32'hFFF98E4A , 32'hFFF379CE , 32'h0003B309 , 32'hFFFDB167 , 32'h0001DC6E , 32'h0006465A , 32'h000172EB , 32'hFFF95593 , 32'h000201B2 , 32'h00000933 , 32'hFFFD1307 , 32'hFFF96B1F , 32'h0001198D , 32'hFFFD07B8 , 32'h000945AD , 32'h0003C54C , 32'h0003A988 , 32'hFFF5284B , 32'hFFF3A284 , 32'h0001F798} , 
{32'h0006C31E , 32'h0010565B , 32'hFFFD7070 , 32'hFFFE623E , 32'hFFFF0EF7 , 32'hFFFE180A , 32'hFFFC3D8B , 32'hFFF5EFCA , 32'hFFFF32ED , 32'hFFFFCAB6 , 32'hFFF9F259 , 32'hFFFACD53 , 32'hFFF78FA2 , 32'h000540F2 , 32'hFFFDF2E6 , 32'h0002BFF1 , 32'hFFF6E005 , 32'hFFF44B85 , 32'h0000FF76 , 32'hFFFB29A6 , 32'h00001FCB , 32'h0002F8A8 , 32'hFFF783A4 , 32'hFFFF73CA , 32'h000268E2 , 32'h0004CFFF , 32'hFFFADE6A , 32'hFFF9FC84 , 32'h00007D61 , 32'h00071543 , 32'hFFFF1F21 , 32'hFFFC4F7C , 32'hFFF8FBF1 , 32'hFFFC0DC4 , 32'hFFFE4007 , 32'h00006BF5 , 32'hFFF8862A} , 
{32'h000659A8 , 32'h00014912 , 32'hFFFE6064 , 32'hFFFA0C2E , 32'h00048BAA , 32'h000005C4 , 32'h00039374 , 32'hFFFE4153 , 32'h0008021B , 32'h00005016 , 32'h0001BB60 , 32'hFFFA63D1 , 32'hFFF99346 , 32'h0003F11B , 32'hFFFCC2A2 , 32'h0001868E , 32'h0006B96F , 32'hFFF9E3D4 , 32'h0000D186 , 32'h00041F62 , 32'h00017756 , 32'hFFFFDAFA , 32'hFFF236E6 , 32'hFFF9CEC5 , 32'h00016664 , 32'h0002DD46 , 32'h0004AB57 , 32'h0000F722 , 32'h00045304 , 32'hFFFD6FDA , 32'h00020053 , 32'hFFF85BD8 , 32'h00026778 , 32'hFFFBF244 , 32'hFFFA1F38 , 32'hFFFA63DA , 32'h000ACDE5} , 
{32'h00004305 , 32'h0000014F , 32'hFFFD62BC , 32'h0002983C , 32'h0004505E , 32'hFFFBEDC1 , 32'hFFFF23D6 , 32'h00010170 , 32'hFFFF6EE5 , 32'hFFFC4518 , 32'h0006EC8B , 32'hFFF8BE73 , 32'hFFFD58C5 , 32'h000D7465 , 32'hFFFCC607 , 32'hFFFFEF5B , 32'hFFF57231 , 32'hFFFD2A42 , 32'hFFF79AB1 , 32'h0007B296 , 32'h00018BA9 , 32'hFFF8298A , 32'h00027AE4 , 32'h0004AC1A , 32'hFFFF8B5D , 32'hFFFD3DB0 , 32'hFFFF57CD , 32'h0003D62B , 32'h00034D10 , 32'hFFF673A4 , 32'h0007C5C5 , 32'hFFFFD1BC , 32'h00023407 , 32'hFFFE31CC , 32'hFFFA3086 , 32'h000D7177 , 32'h000B4308} , 
{32'h0005744F , 32'h0001C993 , 32'h0002373F , 32'hFFF9187C , 32'hFFFE7EB7 , 32'hFFF84FEC , 32'hFFFF2F95 , 32'hFFF80A28 , 32'hFFF9031F , 32'hFFFF185C , 32'hFFFB89EC , 32'hFFF8EA5A , 32'h00016BED , 32'hFFFEEF58 , 32'hFFF6CC1C , 32'hFFFD24C8 , 32'h00058A38 , 32'h00031718 , 32'hFFFD57F3 , 32'hFFFC2BF5 , 32'h000798D4 , 32'h00040E01 , 32'h00061070 , 32'h00049C1B , 32'h0005E18A , 32'h0008CCA8 , 32'h000F252C , 32'hFFFC467F , 32'hFFFB9386 , 32'h00025074 , 32'hFFF928A1 , 32'h0000B083 , 32'hFFFAFF0E , 32'hFFFB2359 , 32'hFFFFA7E4 , 32'hFFFDA8B0 , 32'hFFFC6ADF} , 
{32'h000AA204 , 32'h0000FB82 , 32'h0009148B , 32'hFFFDBD46 , 32'h000E0053 , 32'hFFFE76B5 , 32'h00085F35 , 32'hFFF63BCA , 32'h0006C90F , 32'hFFFEF79A , 32'hFFFC0BFA , 32'h00056523 , 32'hFFF6AD64 , 32'h0001417F , 32'hFFFD8DF6 , 32'hFFFF8199 , 32'h00041A78 , 32'hFFFD237D , 32'h00021A11 , 32'h000BCCBC , 32'hFFFF6828 , 32'h0000EA20 , 32'hFFFDD0F3 , 32'hFFFB310F , 32'hFFF7EEF7 , 32'h000096B7 , 32'hFFFEE641 , 32'hFFF9BB1B , 32'hFFFCCA8D , 32'h00014A32 , 32'hFFFFBD7C , 32'h00011A62 , 32'h000283B1 , 32'h0004C9F8 , 32'hFFFA1AED , 32'hFFFC8F1D , 32'hFFFCEE97} , 
{32'h00068DEF , 32'hFFF775D8 , 32'hFFF83513 , 32'h0000F8F3 , 32'h0005A830 , 32'hFFFB3EF5 , 32'hFFF65EBB , 32'h000112EC , 32'hFFFE3BC2 , 32'h0001E223 , 32'hFFFF4B6B , 32'hFFF862A0 , 32'hFFF8CC73 , 32'h00041602 , 32'h000430E4 , 32'h000B1A73 , 32'h0000330B , 32'hFFFF409F , 32'hFFF9CCB3 , 32'h000258FB , 32'h00049451 , 32'h00025778 , 32'hFFFAAE87 , 32'h0006EC64 , 32'h000436AA , 32'hFFF8439F , 32'h00031075 , 32'hFFFFB6C6 , 32'h00054E67 , 32'h00036D6F , 32'h00009C90 , 32'hFFFC9F9B , 32'hFFFD5BB8 , 32'h0004C3FD , 32'hFFF5D03C , 32'h0000F8DE , 32'hFFFBAA4D} , 
{32'h0003AE78 , 32'hFFFE52C8 , 32'h00069C74 , 32'hFFFD5950 , 32'h0008EFB6 , 32'h0002314B , 32'h0005BC6E , 32'h000016DC , 32'hFFFDABE0 , 32'h000BBF94 , 32'hFFFBBEBB , 32'hFFFBEC78 , 32'h000705F4 , 32'hFFF9817C , 32'hFFF636F8 , 32'h000031C3 , 32'h0001017C , 32'h00036277 , 32'h000A6BB7 , 32'hFFFC5DE7 , 32'hFFFF72D0 , 32'h0001362F , 32'hFFFE9C7C , 32'h00027099 , 32'hFFFFAEFD , 32'h00004AA7 , 32'hFFFBFDCF , 32'h00003AC8 , 32'h0008E1C8 , 32'hFFFBD3FA , 32'h00078982 , 32'hFFFA0900 , 32'hFFFC5D09 , 32'h00045676 , 32'hFFFE1A01 , 32'h00008184 , 32'h00022C01} , 
{32'h0001463B , 32'h0006DCCC , 32'h0001CEA7 , 32'h00051BBC , 32'h0009C299 , 32'h000CEAFE , 32'h0003E853 , 32'hFFFF5E58 , 32'hFFFD3D70 , 32'h00022249 , 32'hFFFD3243 , 32'hFFFCB146 , 32'hFFFFC1E1 , 32'h0001C9BE , 32'hFFFDAEDA , 32'hFFFA35EF , 32'h000475FB , 32'h0005449B , 32'hFFFC681E , 32'hFFFE36FD , 32'hFFFB39A5 , 32'h0006BE0B , 32'hFFFF804D , 32'h0005AF23 , 32'h000110EE , 32'hFFF99638 , 32'hFFFF2BCA , 32'hFFFDF149 , 32'hFFFF5BA3 , 32'h00029E37 , 32'hFFFD885B , 32'hFFFB0B9F , 32'h00021886 , 32'h000774EB , 32'hFFF6C894 , 32'h00032934 , 32'h000532DB} , 
{32'h00004341 , 32'h00018083 , 32'hFFF9A7AF , 32'h0004D4CF , 32'hFFFE67C9 , 32'h00034E0E , 32'h0008D2A6 , 32'h0004BC60 , 32'hFFF82CFF , 32'hFFFE065D , 32'h00015974 , 32'hFFFF236C , 32'hFFFD4508 , 32'h00044869 , 32'h00075B6E , 32'h00089DFC , 32'hFFFFEA17 , 32'h0004830E , 32'hFFFC53FD , 32'h00048898 , 32'hFFFF6EC7 , 32'hFFFC1128 , 32'hFFF44A10 , 32'hFFF7D430 , 32'h0007D1FF , 32'h000C00ED , 32'hFFFA28C8 , 32'h0007C815 , 32'h00012F80 , 32'hFFFFB8CF , 32'h0005E7F6 , 32'hFFF648FC , 32'h0002D60C , 32'hFFFA7D5E , 32'hFFFC5412 , 32'hFFFA41C0 , 32'hFFFD58DA} , 
{32'h0003C47B , 32'h0000920B , 32'h0000B6FD , 32'hFFFEB779 , 32'hFFFE121F , 32'hFFFE801B , 32'hFFF84708 , 32'h0007A3D1 , 32'h00057492 , 32'h0000DBE0 , 32'hFFFDB0B0 , 32'hFFF5EA42 , 32'hFFFE8906 , 32'h0008C4E2 , 32'hFFFA8930 , 32'hFFFF35EE , 32'hFFFF0F8D , 32'hFFFCB57B , 32'hFFFBC204 , 32'hFFFBE732 , 32'hFFFB5A98 , 32'h0001C446 , 32'hFFFE2880 , 32'h00017270 , 32'hFFFE8BF8 , 32'hFFFCD6F9 , 32'h0002B5F1 , 32'h0002B3D4 , 32'hFFFB2EBC , 32'hFFF2873D , 32'h000B5CC8 , 32'hFFFF28F4 , 32'h0004CD4D , 32'hFFFE0CDF , 32'h0005113D , 32'h0007E607 , 32'hFFFD7A18} , 
{32'h00070CD3 , 32'hFFFD0A8F , 32'h00068626 , 32'h000366C5 , 32'h0003C167 , 32'hFFF9A04A , 32'hFFFDB060 , 32'hFFFC4CB3 , 32'hFFFA8F27 , 32'hFFFFDC0E , 32'h00087F5F , 32'h0004D72C , 32'h00048B0A , 32'h0005B960 , 32'hFFF648C1 , 32'h00033750 , 32'hFFFA3CB2 , 32'hFFFE13B9 , 32'hFFFED9E3 , 32'hFFFF0926 , 32'h00046F4C , 32'h0005387F , 32'hFFFE85DC , 32'hFFFDCAE1 , 32'hFFFB0EFA , 32'h00024AB8 , 32'h0004BF45 , 32'hFFFC824B , 32'hFFFC571C , 32'h0005F5E1 , 32'h000056B1 , 32'h0006A8BE , 32'hFFFE04EF , 32'h000385A1 , 32'hFFFF37E4 , 32'hFFFC316E , 32'h0004BCDC} , 
{32'hFFFE1499 , 32'h00037143 , 32'hFFF891D1 , 32'hFFFC3185 , 32'h0000F709 , 32'hFFFA9256 , 32'h0004E550 , 32'h0004762E , 32'h0006430E , 32'h00010827 , 32'h000737EC , 32'hFFFFCFB4 , 32'hFFFEC9C5 , 32'hFFF72C50 , 32'hFFFABFEE , 32'h0009273F , 32'h0005FE22 , 32'h0002E097 , 32'hFFFEC958 , 32'hFFFEED0E , 32'hFFFF8FB9 , 32'h00003FB0 , 32'h00007C92 , 32'hFFFD9E5B , 32'h00009B4F , 32'h0002FA45 , 32'h000072E2 , 32'hFFF3DA14 , 32'hFFFB47D5 , 32'h0004A25F , 32'hFFFE023A , 32'hFFF9C823 , 32'h0007A679 , 32'hFFFE492F , 32'h000174F7 , 32'hFFFA0A14 , 32'hFFFC02AB} , 
{32'hFFFB2553 , 32'hFFF2AA3E , 32'h0007550B , 32'h000DF46D , 32'hFFF96E70 , 32'h000180FF , 32'h0003867A , 32'hFFFDBD0F , 32'hFFFF7100 , 32'h0005788A , 32'hFFFA220E , 32'hFFF54999 , 32'hFFFD9AA2 , 32'hFFFE4E7A , 32'h0004DFC8 , 32'h000C4AC1 , 32'h0004FED7 , 32'h0000EA3E , 32'h0000A820 , 32'h0001B335 , 32'h0007E925 , 32'hFFFECC63 , 32'h0002CDE7 , 32'hFFF6ECF0 , 32'h000776F0 , 32'h00029969 , 32'h00067034 , 32'hFFF2A06D , 32'h000611DB , 32'h00022BD0 , 32'hFFFCA0EF , 32'hFFF7731C , 32'hFFF6A257 , 32'hFFFD1177 , 32'hFFF1C812 , 32'hFFF6F7C8 , 32'h0005C39B} , 
{32'h000438E5 , 32'h0008E4CC , 32'hFFFD5F31 , 32'hFFFCC5AA , 32'hFFF94632 , 32'h0002BC9A , 32'hFFFE5CC6 , 32'hFFFE0D11 , 32'h0000AEC6 , 32'h0009EDFE , 32'h0000B12C , 32'hFFFA2219 , 32'hFFFED541 , 32'hFFFC68B3 , 32'hFFFEF469 , 32'hFFFAE80C , 32'hFFFBBC29 , 32'hFFFF0119 , 32'h00012FA9 , 32'h0000915D , 32'hFFF59E65 , 32'hFFFDC11A , 32'hFFFD03B6 , 32'hFFFA5CF5 , 32'hFFFE1C9B , 32'hFFFE6234 , 32'hFFFE6D2F , 32'h000261EB , 32'h00026A73 , 32'h0001E8F8 , 32'hFFFD28BB , 32'hFFFD19C2 , 32'h00009A3C , 32'h0001C6AB , 32'hFFFAFE3F , 32'hFFF9108B , 32'hFFFBBDB5} , 
{32'h000100DC , 32'hFFF7A997 , 32'h0002ABC9 , 32'h0003BEF7 , 32'hFFFC21BE , 32'hFFFBA756 , 32'hFFFB6EBC , 32'hFFFD5FD0 , 32'hFFFE0728 , 32'h0005883E , 32'hFFFF73D3 , 32'h0004A110 , 32'hFFFE2E46 , 32'hFFFF8689 , 32'hFFFEB54F , 32'hFFFE67A6 , 32'h000163C3 , 32'h000204FF , 32'hFFFE5B30 , 32'hFFFAE5B8 , 32'h0005F8BD , 32'h0001B969 , 32'hFFFB2932 , 32'h00049E9F , 32'h0000D9F5 , 32'hFFFBE510 , 32'hFFFC0C69 , 32'hFFFFE076 , 32'h0002ED90 , 32'h0004F86C , 32'hFFFCDF65 , 32'h00007D5D , 32'h0000CD60 , 32'hFFF63434 , 32'hFFFB8579 , 32'hFFFAD959 , 32'h000322BB} , 
{32'h00061797 , 32'hFFF9F88A , 32'h0001A043 , 32'h00080094 , 32'h0005D1F4 , 32'h0000B704 , 32'h0000C75B , 32'h00051A20 , 32'h00048532 , 32'hFFFFADD5 , 32'h0004907B , 32'hFFFE2DEB , 32'h00040090 , 32'hFFFD7F25 , 32'hFFFEC6FB , 32'hFFFF8EA9 , 32'hFFFF02D6 , 32'h0000AEEA , 32'h0001EECC , 32'hFFFF0F1A , 32'h00042635 , 32'h00006664 , 32'hFFFF9796 , 32'h00096C23 , 32'hFFF7F7E4 , 32'h00014CEF , 32'hFFF6CFEC , 32'h0008A91D , 32'h00017B5D , 32'h00058A68 , 32'h000366B6 , 32'h0009A4EE , 32'hFFF9EDE4 , 32'h00022858 , 32'hFFF616EE , 32'h00061452 , 32'h0003ED48} , 
{32'h0002D158 , 32'hFFFF365E , 32'h000020B1 , 32'h0001674B , 32'h00012790 , 32'hFFFF1A82 , 32'hFFFD3EBD , 32'hFFF90200 , 32'hFFFD90B2 , 32'hFFF8C2DD , 32'hFFF4D401 , 32'h000417BD , 32'hFFFAB236 , 32'h0006C1B3 , 32'hFFFF191E , 32'h0004FD69 , 32'h00021A27 , 32'hFFFF3070 , 32'h00048E83 , 32'h0000E3A5 , 32'h0001914E , 32'hFFF55D36 , 32'h0003CE9E , 32'hFFFF1173 , 32'hFFFC87E2 , 32'h0002B0B8 , 32'hFFF61113 , 32'hFFFDE874 , 32'hFFFAEA0F , 32'h00030EB2 , 32'hFFFFDAB0 , 32'h0003E009 , 32'h0003B572 , 32'hFFF919C7 , 32'hFFFC3AFE , 32'hFFFDEBB5 , 32'hFFFE2DC6} , 
{32'h000E4624 , 32'hFFFCE670 , 32'h0001658C , 32'hFFFCF631 , 32'h000163CC , 32'hFFF5750D , 32'h000595A5 , 32'h000344D3 , 32'h00058C0A , 32'h00066537 , 32'h0003AB6D , 32'hFFFFB3A4 , 32'h00049D85 , 32'h0007E5F3 , 32'h00009A48 , 32'hFFFE73DE , 32'h00006CAE , 32'hFFFF6029 , 32'hFFFB834D , 32'h00090DCF , 32'hFFFF8F08 , 32'h00037C0A , 32'hFFFE39D9 , 32'h0004CE3D , 32'hFFFFB10B , 32'hFFFDCD4B , 32'h00030DFC , 32'hFFFDA08E , 32'hFFFF83A7 , 32'hFFFC6513 , 32'hFFFBE1F9 , 32'h0001C91C , 32'hFFF79100 , 32'hFFFCF314 , 32'h00072030 , 32'hFFFDCF75 , 32'hFFFC9C6E} , 
{32'hFFFA8BC6 , 32'h000448DE , 32'h00027CAA , 32'h000926DB , 32'hFFFE2E62 , 32'hFFFAD8EB , 32'hFFF86A67 , 32'h000139B2 , 32'hFFFEEA49 , 32'h00055996 , 32'hFFFC7432 , 32'hFFFC2B25 , 32'h00015A34 , 32'hFFF5DA16 , 32'h000240DF , 32'hFFFB17FF , 32'h000293FC , 32'hFFFA3090 , 32'hFFFEF636 , 32'hFFFA1EA4 , 32'hFFFEB70C , 32'hFFFA9247 , 32'h00054ED6 , 32'hFFFE9434 , 32'hFFF8A4A1 , 32'hFFFDA995 , 32'hFFFF2914 , 32'hFFFCD3F3 , 32'h0005462B , 32'hFFFE5E62 , 32'hFFFC6EF7 , 32'h00057F9B , 32'hFFFD3B43 , 32'h00048D17 , 32'h0005B7C5 , 32'hFFFE09CE , 32'hFFFFC587} , 
{32'hFFFA856C , 32'h00018E4F , 32'h0009E45E , 32'hFFFC5D0A , 32'h000255BE , 32'hFFFFE618 , 32'hFFFD2F74 , 32'hFFFFD3B6 , 32'hFFF86466 , 32'hFFFC2023 , 32'hFFFD3C90 , 32'hFFFDB50B , 32'h00025921 , 32'h000016FD , 32'h000757D2 , 32'hFFF3CDA8 , 32'hFFFEB773 , 32'hFFF5BC66 , 32'h0002A087 , 32'h00083CA1 , 32'hFFFD63F0 , 32'h00030977 , 32'h0005CC7F , 32'hFFFA466B , 32'h00058BE2 , 32'h0003078C , 32'hFFF82F9B , 32'h000737FF , 32'hFFFCC2BC , 32'h00005FA4 , 32'hFFFBAD88 , 32'hFFFE178A , 32'h00058602 , 32'h00069CE7 , 32'hFFFB49FD , 32'h0003D782 , 32'hFFFD4FA1} , 
{32'h0006D1D5 , 32'h0007CD4D , 32'hFFFA28D4 , 32'h000319A2 , 32'h0003A822 , 32'h00038C64 , 32'hFFFBD46B , 32'h00027133 , 32'h0009B0F2 , 32'hFFFD87C6 , 32'hFFFF4E59 , 32'h0005E6FA , 32'hFFF8F441 , 32'hFFFA631C , 32'h0001232C , 32'hFFF94ADD , 32'hFFFE9605 , 32'hFFFF53B1 , 32'h00026EE2 , 32'hFFFE2F30 , 32'hFFFF2CBE , 32'h0002E293 , 32'h00042647 , 32'h0005121E , 32'h000764EE , 32'h00024832 , 32'hFFFA9301 , 32'hFFFC68EA , 32'hFFF8AF45 , 32'hFFFDB2EF , 32'hFFFC19B2 , 32'h0008827D , 32'hFFFEE179 , 32'hFFFCF22A , 32'hFFFD04A9 , 32'h00029E0C , 32'h0002516B} , 
{32'hFFF9EB7E , 32'h0000EECA , 32'h0008C0A4 , 32'h0003A264 , 32'hFFF9EAC5 , 32'hFFFE861C , 32'hFFFB9C44 , 32'h000066AD , 32'h00021483 , 32'hFFF8F5EA , 32'h00017014 , 32'h0005BEBB , 32'hFFFFE5AC , 32'hFFF7D191 , 32'hFFFD7956 , 32'hFFFE751A , 32'hFFFE73F0 , 32'hFFFBB035 , 32'hFFFF4085 , 32'hFFFA4820 , 32'h0002390E , 32'hFFF50281 , 32'h000DDFA1 , 32'hFFF916BA , 32'hFFFA0647 , 32'hFFF73BE7 , 32'hFFFAB599 , 32'h0002DA2F , 32'hFFFF8957 , 32'hFFFAFE3B , 32'hFFFB5C69 , 32'hFFFDA868 , 32'h0005B035 , 32'h00027F50 , 32'h00087FB4 , 32'hFFFFEC1B , 32'h0003E0D8} , 
{32'hFFFAC8AD , 32'h00002152 , 32'h0008DFD2 , 32'hFFFFE39F , 32'hFFFF85F4 , 32'hFFFEAB1D , 32'h00031A3B , 32'hFFFF960A , 32'h0002ABF3 , 32'h0002074A , 32'hFFFD7FEF , 32'hFFFFCC46 , 32'h00025056 , 32'h00000CF9 , 32'h0002C3A6 , 32'h0000DA10 , 32'h0008201B , 32'hFFF35EB8 , 32'h000620FB , 32'h0006D13E , 32'h00018E2C , 32'hFFFCEB94 , 32'hFFF6DA44 , 32'hFFFAF1B1 , 32'hFFFBF99B , 32'hFFFDB312 , 32'h0004EE97 , 32'h00034A65 , 32'hFFFE0FB5 , 32'h000594BE , 32'h0001441D , 32'h00036490 , 32'hFFFE15E7 , 32'hFFFE216F , 32'hFFFF119A , 32'hFFFB26EA , 32'hFFFEA10C} , 
{32'hFFFF556D , 32'h0006DB03 , 32'hFFFD42EE , 32'h000A75FF , 32'h0003298D , 32'hFFFD3616 , 32'h0000BACD , 32'h0000DBFA , 32'hFFFFC267 , 32'h000275A0 , 32'hFFFC3094 , 32'h0003A485 , 32'h000026E5 , 32'h00050CB3 , 32'hFFF9083E , 32'h0009C78B , 32'hFFF726B8 , 32'h0003EB1B , 32'h00065223 , 32'hFFFC7DEF , 32'h000105AC , 32'h00011A61 , 32'h00034340 , 32'h00043988 , 32'h00079DA3 , 32'hFFFDC5DF , 32'hFFFFFDB4 , 32'h000010AD , 32'hFFFE96BF , 32'h00037BDC , 32'h00011084 , 32'hFFFD0C9E , 32'h0001C127 , 32'h00066D3A , 32'h0005982B , 32'h00037B08 , 32'hFFFFEA27} , 
{32'h000184AF , 32'h0002FD1C , 32'hFFF9B1CB , 32'h0008566F , 32'hFFF3C878 , 32'hFFFDEE4D , 32'h0008E4EB , 32'h0000CC29 , 32'h00025B3E , 32'hFFFE22D7 , 32'h00014C53 , 32'hFFFDF18C , 32'h0007B47A , 32'hFFFE4F16 , 32'h000125D6 , 32'h0001565E , 32'h000A05AB , 32'h0002BE90 , 32'hFFFA1FEE , 32'hFFF9E315 , 32'hFFF58B2B , 32'h00022451 , 32'h000976FD , 32'hFFFB603A , 32'h00003CB2 , 32'hFFFDDFD6 , 32'hFFF8F663 , 32'hFFFF6073 , 32'hFFF5C679 , 32'hFFFBC326 , 32'h00007B11 , 32'hFFF8BDC1 , 32'h0002E7E6 , 32'h00004D3C , 32'hFFFD2241 , 32'h0006F9FD , 32'hFFFB51B8} , 
{32'hFFFE147E , 32'hFFFD3558 , 32'h0005931C , 32'hFFFD2A11 , 32'hFFFBC4B3 , 32'h00045A36 , 32'hFFFEB513 , 32'h000558AE , 32'h0000238E , 32'hFFF8CBD4 , 32'hFFFDB50B , 32'hFFFC3094 , 32'h0006C43D , 32'hFFF2AF62 , 32'h000B27BD , 32'hFFF8AA63 , 32'hFFFC11CF , 32'h00074265 , 32'h00068B22 , 32'hFFFC7D3C , 32'h0005278D , 32'h0005EE8E , 32'hFFFCC184 , 32'hFFF3698D , 32'h0000BD08 , 32'h0001FDF0 , 32'hFFFFB4FA , 32'hFFF5187D , 32'hFFFB6AC4 , 32'h00020E76 , 32'hFFFB0B21 , 32'hFFFD68F1 , 32'h00075896 , 32'h00012AD6 , 32'hFFF90331 , 32'h00026E00 , 32'hFFFC8090}
};

logic signed [31:0] US_1 [37][37] ='{
{32'hF24FAF50 , 32'h087A4890 , 32'hE8309380 , 32'h0AE123A0 , 32'hF6CAD420 , 32'hD6541940 , 32'h0B6E5990 , 32'h090CE7D0 , 32'h0BF11770 , 32'hD8383400 , 32'h0B3B3FF0 , 32'h0AE1B0A0 , 32'h028B8F14 , 32'h11577280 , 32'hE6F93860 , 32'hEA5726E0 , 32'h17EFE440 , 32'h07B11818 , 32'h156D0600 , 32'h11F2AEE0 , 32'hD55E71C0 , 32'hF16F5440 , 32'h09FC94F0 , 32'h028D4E0C , 32'h01322A28 , 32'h05F65F88 , 32'h1F344140 , 32'hEC949A20 , 32'h1D4F7760 , 32'h08ACA090 , 32'hEF7BFD00 , 32'hFFCC44A7 , 32'hFAE41048 , 32'h0A727F70 , 32'hDFF3F140 , 32'h021C1270 , 32'hCBD2A180} , 
{32'hF1928B10 , 32'h081A3C90 , 32'hD29B2780 , 32'hF6CCCBB0 , 32'h14EC59A0 , 32'h12E0AD40 , 32'h190DB920 , 32'hF3BE4010 , 32'hFC6F2164 , 32'hF73C5000 , 32'hFBB6C398 , 32'h1454FE80 , 32'hF4ED6CC0 , 32'hF2DF7780 , 32'hE68C23C0 , 32'h071CD468 , 32'hFDAB10A0 , 32'hC968C540 , 32'h0D3B4C60 , 32'h01B1F560 , 32'hE2193520 , 32'h094C3B20 , 32'h03634CB4 , 32'h1D7E49C0 , 32'hF308C630 , 32'hECE27BC0 , 32'hD9E5B140 , 32'h1B541D20 , 32'h064FD2E0 , 32'hDB0D3780 , 32'h10EA2020 , 32'hF59F05D0 , 32'h16BEBFA0 , 32'h071C9128 , 32'hECE34940 , 32'hEEDD2C00 , 32'h09BEE0D0} , 
{32'hDE607AC0 , 32'hDAFBBA40 , 32'hECE44820 , 32'hEC616AC0 , 32'h1B356F00 , 32'h04479B28 , 32'h1B099A20 , 32'hFC97EA68 , 32'h1ACA2620 , 32'h09AFC360 , 32'h167E8F60 , 32'hE1CDD400 , 32'hE5EBFBE0 , 32'h0891D570 , 32'h10288CE0 , 32'h21E82980 , 32'h02A10794 , 32'h22DB1300 , 32'h217FDC40 , 32'hF645EED0 , 32'h1E3C9D00 , 32'h06D29CB8 , 32'h104AF280 , 32'h03C7FF7C , 32'hFE42B768 , 32'h0CA71460 , 32'hEC365960 , 32'h07656FB0 , 32'hEA090B60 , 32'hFBAA0F10 , 32'hEF6B6A40 , 32'h12F210E0 , 32'h0A22C210 , 32'hFAD41328 , 32'hEBF68B00 , 32'h043F7708 , 32'hDC6C84C0} , 
{32'hFBC75D58 , 32'h0B492690 , 32'h0C080210 , 32'hD7525F00 , 32'h0C662650 , 32'hE2779F20 , 32'h0126152C , 32'hFC09BEE0 , 32'hFA437F08 , 32'hF5F2F8F0 , 32'h3094AD00 , 32'h00D0FE9E , 32'hDFC7EF00 , 32'h0853AE10 , 32'hED898960 , 32'hF711D240 , 32'hF34F4850 , 32'hFEE6ADFC , 32'h04F34B10 , 32'hFACAF2D8 , 32'hFDFDB8E4 , 32'hEDE78500 , 32'h1651E980 , 32'h0C42D180 , 32'h08623A10 , 32'hE234AF40 , 32'h0B004F40 , 32'h05AF0848 , 32'h01FD4C4C , 32'h0C103F90 , 32'h13A34CA0 , 32'h274B39C0 , 32'hF49A84D0 , 32'h100A01E0 , 32'h01F0E9F8 , 32'h2E57E0C0 , 32'h31815CC0} , 
{32'h1F1BF1A0 , 32'h03FAAF40 , 32'h13D0F1E0 , 32'h1E0889A0 , 32'hF669FBD0 , 32'hE325D540 , 32'hF6FE1820 , 32'h03C7620C , 32'hF913EDC8 , 32'hD57CF980 , 32'hE082B3A0 , 32'hF634ACD0 , 32'h0E07B1E0 , 32'h120CF000 , 32'hF1057A70 , 32'h16CC2E20 , 32'hFC55CBC0 , 32'h19C14E60 , 32'h15CB14E0 , 32'hFB6AF598 , 32'h0ECFDB50 , 32'hEF588B00 , 32'h172EDB00 , 32'h09125F40 , 32'hF5B1F930 , 32'hEC4F10A0 , 32'hCFEFBBC0 , 32'h12E54F20 , 32'h0BC5BDB0 , 32'hF6E3C3F0 , 32'hE3A61B40 , 32'h015786AC , 32'h210743C0 , 32'hEADC83C0 , 32'hF5CACE40 , 32'h10DEE080 , 32'h15BCCB80} , 
{32'hFDC58474 , 32'h0F258DD0 , 32'h1C179460 , 32'hF8E13690 , 32'hF7E48920 , 32'hF413B5E0 , 32'h00836DAC , 32'hE684CA00 , 32'hF5C03B90 , 32'h065AD018 , 32'hE981BC20 , 32'h235839C0 , 32'h02C10FE4 , 32'hFE6A3958 , 32'h00510B10 , 32'h07B7CF08 , 32'hFC4862DC , 32'hE94EA9A0 , 32'hF71A0A80 , 32'h0B689070 , 32'h3356DD00 , 32'h16EA1AE0 , 32'hF4A18DC0 , 32'h06691830 , 32'hFB9B0348 , 32'h0829F9D0 , 32'h0086D39D , 32'hEF35BBC0 , 32'hFF00951F , 32'hEA66CA80 , 32'hFAD29920 , 32'h0DFA58B0 , 32'h123B3A20 , 32'h379C4A00 , 32'hE12FF080 , 32'h2B609DC0 , 32'hDED9A7C0} , 
{32'hF7D3C2C0 , 32'h251E27C0 , 32'hF4EB07F0 , 32'hF6AA6CA0 , 32'h1242D640 , 32'hF3290AB0 , 32'hE8B03F60 , 32'hF3B41870 , 32'hFA9DEDF0 , 32'h11C793C0 , 32'h2C551EC0 , 32'h0AA79290 , 32'h0E842C10 , 32'h22E5D400 , 32'hE4E5DDC0 , 32'hF98CC2E0 , 32'hF753EF80 , 32'h05CC53D0 , 32'h0627B550 , 32'hE7D4BD60 , 32'h0DBD0C20 , 32'h10BE0940 , 32'hFA13C6C8 , 32'hEA77ED20 , 32'h1E0050E0 , 32'h1E9D34C0 , 32'hE19C9DC0 , 32'hEF12BF80 , 32'h06D849C0 , 32'hFC5C1790 , 32'h02E36FCC , 32'hC7146200 , 32'h0E843CB0 , 32'hE9FDAD60 , 32'hFDF12AB4 , 32'h0C6BD1E0 , 32'hFFD7127C} , 
{32'h088E0930 , 32'h10AAD1E0 , 32'hF752D9F0 , 32'hF40E0010 , 32'h20B9C240 , 32'hF643BE90 , 32'hF03C2210 , 32'hF3C4C3A0 , 32'hF2CCD150 , 32'hFC888428 , 32'hE6134860 , 32'hFDA0D860 , 32'hECE9F460 , 32'h00E173E2 , 32'hF432AB30 , 32'h01FF5AC0 , 32'hCF989140 , 32'hF1A5C430 , 32'h16B35EA0 , 32'h15D6E000 , 32'h1C293CC0 , 32'hE0587420 , 32'h05F849F8 , 32'hF47BD740 , 32'hE05D0340 , 32'h2DB93640 , 32'h1E34D6C0 , 32'h0188E414 , 32'h0DC26EE0 , 32'h16B6AAE0 , 32'h16F71F00 , 32'h0FA00190 , 32'h11EEE100 , 32'hE8E6AFC0 , 32'hF8EDCFE8 , 32'hE0AB6A40 , 32'hFDE16290} , 
{32'hDD36CC00 , 32'hDC41C2C0 , 32'h18299AC0 , 32'hE3947620 , 32'hE7A4B380 , 32'hF118A800 , 32'hFE18BCFC , 32'hF7872820 , 32'hE77C64E0 , 32'h0D2AAA40 , 32'hE7E9CFC0 , 32'h235C8640 , 32'hFD4700C4 , 32'h12C18E40 , 32'hFAF26708 , 32'hE814D5C0 , 32'hF3C5B870 , 32'hF33042F0 , 32'h16E75540 , 32'hE9F6CDC0 , 32'hF83F7A10 , 32'hE0D6BFA0 , 32'hFAB0EE70 , 32'hFF050408 , 32'h05B61090 , 32'hF422C3C0 , 32'hE0F53B20 , 32'hD4F29280 , 32'hEFF37380 , 32'hF16BF9F0 , 32'hF4E5E6F0 , 32'h10CC2A80 , 32'hED8B4D00 , 32'hE4AE5BC0 , 32'h04451958 , 32'hE6192280 , 32'hFAE1E1A0} , 
{32'h0B330FD0 , 32'h03E104BC , 32'hF80076A8 , 32'hFB3AE4B8 , 32'h0792F558 , 32'h2F77FC00 , 32'h17044180 , 32'hF3976800 , 32'h0FCE4A20 , 32'h02460E40 , 32'hF1E19D10 , 32'h09C1CD10 , 32'hFDF56E34 , 32'h1F83F6E0 , 32'hD226DFC0 , 32'h00146B99 , 32'h05A66EE0 , 32'h1DBED080 , 32'h0525D3E8 , 32'hF50FC730 , 32'h13710EC0 , 32'hDADF5740 , 32'hD32A5C80 , 32'hD6FDB580 , 32'hF944A458 , 32'hD0F1CF00 , 32'h0B8DA980 , 32'h0893B150 , 32'h07DCF498 , 32'h05556620 , 32'h06B79848 , 32'hFBBC7498 , 32'hFAC07798 , 32'h1157C4A0 , 32'hFA793A60 , 32'hFFDE7FBC , 32'hFB2D9E08} , 
{32'hE36BB920 , 32'hCE2A1500 , 32'h040820C0 , 32'h00A1BE47 , 32'hFEEBCB58 , 32'hF5774210 , 32'h09BBA860 , 32'h139242C0 , 32'h04511BA0 , 32'hEF2497A0 , 32'hE536C080 , 32'hFB6E7988 , 32'h03057F1C , 32'hF87A4148 , 32'h02998698 , 32'h0354F17C , 32'hE99C1A60 , 32'h0D39E9D0 , 32'hEC81C480 , 32'h15C87860 , 32'hF5190AD0 , 32'hF4E11380 , 32'hEFDCD040 , 32'hE8157300 , 32'h1CCB81E0 , 32'h1853A520 , 32'hFBDC66F8 , 32'h0BEAE370 , 32'h0DCED5A0 , 32'hEE70D2E0 , 32'h33158740 , 32'hE39ABE60 , 32'hF9631CF8 , 32'hFB491EC0 , 32'hDB191C00 , 32'h24958FC0 , 32'h160937A0} , 
{32'h1050E900 , 32'hE9757BC0 , 32'hFAA93D58 , 32'h131E9BC0 , 32'hFCA4BC0C , 32'hD533FC80 , 32'hEC5027C0 , 32'h032458B8 , 32'hF9B41548 , 32'h14858A00 , 32'h1054B040 , 32'hFB20A688 , 32'hEF7A9E00 , 32'h02653F18 , 32'hFA33EC18 , 32'h1D269800 , 32'h0D1ECEB0 , 32'hF3477750 , 32'hF6153100 , 32'h15743B20 , 32'h16746EC0 , 32'hDF9FE9C0 , 32'h08EF2930 , 32'h0F004170 , 32'hFCD015C0 , 32'hDC50D5C0 , 32'hEB7622C0 , 32'hFCA9A3CC , 32'hF3453D50 , 32'h112200E0 , 32'h30207D00 , 32'hDAD209C0 , 32'hF5242AC0 , 32'h161C76C0 , 32'h1089DDE0 , 32'hEBBB06A0 , 32'hDE14DEC0} , 
{32'hFDA9743C , 32'hF5843900 , 32'h12C5AC00 , 32'h129145A0 , 32'hF7461360 , 32'hFFF06C81 , 32'h13E681A0 , 32'hFF7858D0 , 32'h0B1EAEA0 , 32'h1B9E6160 , 32'h27109740 , 32'h2C27AD80 , 32'h0E196A20 , 32'hF1809AE0 , 32'h01B4CBA8 , 32'hE9249820 , 32'hF28756A0 , 32'h29486900 , 32'h02ECC5E0 , 32'h2648A7C0 , 32'hF69EA1A0 , 32'h11DB8040 , 32'hECE869C0 , 32'h0950A330 , 32'hDF4C9400 , 32'hFD0744B4 , 32'hE2C41AC0 , 32'hFFD1E6C8 , 32'h154FE2E0 , 32'h18FFA760 , 32'h1693D1E0 , 32'h157491A0 , 32'h24EAB5C0 , 32'hF4215B70 , 32'hFE18D200 , 32'hF69FA610 , 32'h02AA0E38} , 
{32'hD8888100 , 32'h173E48A0 , 32'hC97E9700 , 32'h2EF032C0 , 32'hE7FA1060 , 32'hDBC67F80 , 32'h14F06200 , 32'h01A5A0E4 , 32'hE20EF900 , 32'h14F22CA0 , 32'hF93F8BB0 , 32'hF17489B0 , 32'h06F8B7B0 , 32'h1086A400 , 32'h08354FE0 , 32'h0AECB260 , 32'hF1D9D3E0 , 32'hFEA2464C , 32'hF75A1520 , 32'hF757C500 , 32'h0D9517D0 , 32'h0F3FA010 , 32'hE91384E0 , 32'hF283D330 , 32'hEDD040C0 , 32'hE8A41540 , 32'h1269EF20 , 32'hF8246E80 , 32'hEA8779C0 , 32'hFF082C01 , 32'h05E02268 , 32'h16AD7560 , 32'h019C2F18 , 32'hEC5F8FC0 , 32'hFD645CDC , 32'h0E0ABBC0 , 32'h12069900} , 
{32'h039B9BF8 , 32'h04883340 , 32'h0226A708 , 32'hE7B46920 , 32'hD9C34700 , 32'h00E125B9 , 32'hFED36324 , 32'hDAB53B40 , 32'h1458D100 , 32'h02923378 , 32'h04C0E528 , 32'hED519D00 , 32'hE23FE0C0 , 32'h14AC9AC0 , 32'hFD538F14 , 32'hFEB67EB0 , 32'h1903D4C0 , 32'hF5A0EEB0 , 32'hBF72AE00 , 32'h1287B9E0 , 32'hEDD6D1A0 , 32'hF2445AF0 , 32'h156C7420 , 32'hDE781EC0 , 32'hE1C5DD60 , 32'h096E0E80 , 32'hF5AD9600 , 32'hFE25596C , 32'hF07AB520 , 32'hF5FDA8D0 , 32'hFDD5413C , 32'h03BC8C2C , 32'h20977500 , 32'hE53631E0 , 32'hF36D6760 , 32'h0372E04C , 32'hFB90C910} , 
{32'h0C705450 , 32'hF60027C0 , 32'h07B6B6D0 , 32'hEA51AC40 , 32'h09886E70 , 32'hEB1DD3A0 , 32'h1C141700 , 32'h06E61DE8 , 32'hEA134380 , 32'hFCD02AE0 , 32'hFDD552BC , 32'h025B47A0 , 32'h0E6F8AC0 , 32'h1E6B5A00 , 32'hF3B83F40 , 32'hF9930B60 , 32'hD0592C80 , 32'hFA633270 , 32'hE8A7EEE0 , 32'h1D8BFF20 , 32'hF7333F50 , 32'h22415C80 , 32'h0A9F9F50 , 32'hE7F794A0 , 32'h1DD755E0 , 32'hEE1C4240 , 32'h006E6E68 , 32'h33524E40 , 32'hF35528D0 , 32'h0175EF48 , 32'hEB4F4080 , 32'h08390260 , 32'hFC1E5E50 , 32'hFEB390BC , 32'h1BA98340 , 32'hF1885D70 , 32'hDC95D640} , 
{32'h05436000 , 32'hFCF25978 , 32'hF15FCBC0 , 32'h0B4867B0 , 32'h07141840 , 32'hFFEEAD66 , 32'hDB1A6480 , 32'hE8280020 , 32'hFD84203C , 32'hF363DDC0 , 32'hF778E0C0 , 32'h099C6800 , 32'hDE39BAC0 , 32'hF9E48780 , 32'hDBEDB500 , 32'hFFE7E029 , 32'h149DF360 , 32'h23D11780 , 32'hFC06CEEC , 32'h2D3808C0 , 32'h09808030 , 32'h1AA624A0 , 32'hEB244C60 , 32'h17FC4520 , 32'h2F00A400 , 32'hFFE201F4 , 32'h0BADC8D0 , 32'hF51D6DF0 , 32'hE48235E0 , 32'hE24D3940 , 32'hFF5F8E34 , 32'h166922A0 , 32'hFDB25B18 , 32'hEEF88400 , 32'h00863D6E , 32'hE925D540 , 32'h0EA72EB0} , 
{32'h0C0807F0 , 32'h1B763F40 , 32'h06090BF0 , 32'hFC4E8314 , 32'h21F5AA00 , 32'hE9E5F720 , 32'h0AA74400 , 32'h26D22700 , 32'h13393080 , 32'h104B5A80 , 32'h05DE6F08 , 32'h1C7D8B60 , 32'hF6C94890 , 32'hF3ECD2A0 , 32'h22738D80 , 32'hF406D2D0 , 32'h099861A0 , 32'hFA872D28 , 32'h0BCDCCC0 , 32'h259F5E40 , 32'h001442C2 , 32'hDBF1D2C0 , 32'hF00E01D0 , 32'hEABE1D40 , 32'hF8BD7800 , 32'hF626FED0 , 32'h04EBEB80 , 32'h05D233C8 , 32'hD2671080 , 32'hDFCE3180 , 32'hDEA93380 , 32'hE99E6180 , 32'h00C2816E , 32'hF4747A20 , 32'hF4141730 , 32'h07909238 , 32'h0D5D7670} , 
{32'hDD31AB40 , 32'h1CCEFE20 , 32'hF6A43A20 , 32'hF2ECE160 , 32'hE646DDA0 , 32'h11B21E00 , 32'h093675C0 , 32'hFFD670E5 , 32'h10D835C0 , 32'h236EBDC0 , 32'hD925A440 , 32'hFC2201F8 , 32'h07AB3188 , 32'hE3B8CB60 , 32'hE548BDA0 , 32'hFAB4A5E0 , 32'hFB726398 , 32'h0B194DA0 , 32'h1266AB00 , 32'h28363AC0 , 32'h087BF320 , 32'hFDA18DAC , 32'h38972BC0 , 32'h02A5B454 , 32'h12A34C40 , 32'hF1DB2CB0 , 32'hFAE0D9D8 , 32'hF9F153F8 , 32'hFC0D2AE4 , 32'h21BDA780 , 32'hF5159F50 , 32'hE768E360 , 32'hFB188038 , 32'hFFA5F2C9 , 32'h09250030 , 32'h11EEA720 , 32'h077FFC40} , 
{32'h04A1DFC8 , 32'h16CC3100 , 32'hEF12CEC0 , 32'hF4EB1C20 , 32'h1AEFC960 , 32'h12366E60 , 32'hF981D028 , 32'h1B109BC0 , 32'hF4301DB0 , 32'h014F7980 , 32'hFC9466B0 , 32'h0B751800 , 32'h277A6480 , 32'hF71A1A80 , 32'h02DB93E0 , 32'hF3868210 , 32'h0E78A770 , 32'h0AAEF9A0 , 32'hD04E0940 , 32'hF3ED5480 , 32'h15D4BD60 , 32'hE656E360 , 32'h150E65A0 , 32'h1A3A7900 , 32'h0EEC6A60 , 32'hF4F97E60 , 32'hF2FEFD80 , 32'h02AA3F74 , 32'h0289A2C8 , 32'hFCB2248C , 32'h1888E400 , 32'h24ACE040 , 32'hF209E110 , 32'hD5FC9480 , 32'hE5BAC3C0 , 32'h0A8AA7E0 , 32'hDC83C9C0} , 
{32'hFE361B28 , 32'h091413B0 , 32'h065CEA18 , 32'h20A85D00 , 32'h0AAA8E10 , 32'h0D746340 , 32'hEE9676C0 , 32'hFEB65B2C , 32'h01325D5C , 32'hFA7933F0 , 32'hFE72D374 , 32'hF4FD0040 , 32'hCC7F6040 , 32'hEF2A5A00 , 32'hF1F83170 , 32'hEBF76840 , 32'hEB3021C0 , 32'hF0B8A240 , 32'hFC832F50 , 32'h066894E0 , 32'hF7614860 , 32'h09596000 , 32'hE7A6FAC0 , 32'hFA9564F0 , 32'hE94BCB20 , 32'h044A60E0 , 32'hD3F620C0 , 32'h08D0B880 , 32'h04860318 , 32'h134C53A0 , 32'hEDC752C0 , 32'h03F6B2E4 , 32'hC88F2B80 , 32'hEB8BC440 , 32'h020B162C , 32'h2967F380 , 32'hE210E4C0} , 
{32'h3590E940 , 32'hF3746E40 , 32'hE7D02D00 , 32'h06F67350 , 32'hEFBC2CC0 , 32'h013025B8 , 32'h0FA82A40 , 32'hE40FC720 , 32'h26997100 , 32'h092D5CA0 , 32'h03EF402C , 32'hF17386E0 , 32'h1ABC8DE0 , 32'h12294D00 , 32'hFDE341C8 , 32'hE03995C0 , 32'hCF3B8140 , 32'h05C77908 , 32'h06D18210 , 32'h00328BF8 , 32'hFEBD91A8 , 32'hFDFB35F4 , 32'h0C7EF970 , 32'h21A1FEC0 , 32'hF4AA8530 , 32'h088885A0 , 32'h021452DC , 32'hEA870B40 , 32'hDDCFA800 , 32'hEB0327C0 , 32'h08CF6C90 , 32'hF803DB20 , 32'hE1F49F20 , 32'h05E82B10 , 32'hED546E80 , 32'h094F7470 , 32'h058A27E8} , 
{32'h29DB7740 , 32'h0D81BCB0 , 32'hEC83F880 , 32'hD9FCAE80 , 32'hD17388C0 , 32'hF21D9680 , 32'h2FA65100 , 32'h1F937AC0 , 32'hE545F3C0 , 32'hFD616AD8 , 32'hFC66D3D4 , 32'h10E78720 , 32'hE14E1140 , 32'hE2ADBE60 , 32'hECA391E0 , 32'h1533D580 , 32'h07450D10 , 32'h15EBA560 , 32'hFD754028 , 32'hEC4BCFA0 , 32'h08319EF0 , 32'h01D2E2F8 , 32'hEA90DE00 , 32'h0D1C0B70 , 32'h005002FE , 32'h233BED80 , 32'hF8472150 , 32'h01949F08 , 32'hF9B19110 , 32'h098F31C0 , 32'h007C18A9 , 32'hF4D1F210 , 32'hF6E73600 , 32'hF8283588 , 32'h0349C088 , 32'h001D7684 , 32'hFD6BA268} , 
{32'h0556CFB8 , 32'hF29291A0 , 32'hE21278E0 , 32'hE3A6C5E0 , 32'h0A48EAA0 , 32'h0B1B7A80 , 32'hFA96C778 , 32'hE1D55D00 , 32'hDF5AAF80 , 32'hE7A616C0 , 32'hF86E4F88 , 32'h02B5875C , 32'h17D51400 , 32'h189DEEA0 , 32'h23057080 , 32'hFE238A24 , 32'h17AD89A0 , 32'hF963D7C8 , 32'h05AC9D18 , 32'h203B0300 , 32'hF98A8568 , 32'hF9D98870 , 32'hE19197A0 , 32'h117C0B60 , 32'h0228186C , 32'h05050300 , 32'hECF40880 , 32'h0196ACC4 , 32'hE7ECB560 , 32'h41541B80 , 32'hF2E9E560 , 32'hF5E83820 , 32'h00688E90 , 32'h043A29D8 , 32'hF5EC94F0 , 32'h134513C0 , 32'h0DABD040} , 
{32'h013A1DEC , 32'hFE55F9E0 , 32'hEDDBE0E0 , 32'h04F7B558 , 32'hE0AB1460 , 32'h100D3AA0 , 32'hEF4E3B60 , 32'h1271EEE0 , 32'h37F58FC0 , 32'hDB71DA00 , 32'h09A55F60 , 32'h2AF97D40 , 32'hEF41BBA0 , 32'h04429B30 , 32'h16966DC0 , 32'h19F774E0 , 32'hDCB38AC0 , 32'hE0CBF700 , 32'hFE099888 , 32'hF6041A50 , 32'h0F1906D0 , 32'h035FB0EC , 32'hFA55CFC0 , 32'hFEEEE970 , 32'h214E79C0 , 32'hEC1D37A0 , 32'h08D72BE0 , 32'hF55C4070 , 32'hFC04C0E4 , 32'h1C8791C0 , 32'hFF791740 , 32'h04723A90 , 32'h16184CC0 , 32'hE8744FA0 , 32'h04F5D060 , 32'h042B8D40 , 32'hF8DDACB8} , 
{32'hE338E7E0 , 32'hF818B650 , 32'h0360B81C , 32'h0A28A510 , 32'h1BFA53E0 , 32'hFEE053A8 , 32'hFC40736C , 32'h001F1F15 , 32'h00470169 , 32'hE36E4B40 , 32'hED97FAA0 , 32'h2DDF7700 , 32'hF443B280 , 32'h06677028 , 32'hF1D117A0 , 32'hF9881BC0 , 32'hF902A190 , 32'h22FD61C0 , 32'hE0240F20 , 32'hDE0E31C0 , 32'hF7742340 , 32'h09147EE0 , 32'h18C4F5E0 , 32'h15205360 , 32'hD70FDA80 , 32'h07C08C30 , 32'h1350C640 , 32'h081885A0 , 32'hD0E8E6C0 , 32'h0D6E9080 , 32'h0339EA4C , 32'hE00B6040 , 32'h04F72AF8 , 32'h0AEA59E0 , 32'h152DB860 , 32'h06E10E90 , 32'h003FD6C6} , 
{32'h0DE28830 , 32'h08953C50 , 32'hF7ACBB80 , 32'hFF6DA6FA , 32'h22CCE0C0 , 32'hD134A040 , 32'h1E1361C0 , 32'hC68EC900 , 32'h1F402020 , 32'hF4D5DA50 , 32'hE7B9F500 , 32'h0CA8A250 , 32'h05790440 , 32'hD304A940 , 32'h11F0AE00 , 32'hFE531570 , 32'h0C8C7D50 , 32'h06CDBE48 , 32'hF7C65280 , 32'hE734FE80 , 32'hFE91A204 , 32'h0A63F650 , 32'h01C314CC , 32'hDCFE3480 , 32'h137C31C0 , 32'hF57D7140 , 32'hEEF8A6C0 , 32'hF34D90B0 , 32'h0B740940 , 32'h0FE2EB80 , 32'h099D65D0 , 32'h07A1D720 , 32'hF1468C10 , 32'hFA80DC20 , 32'h0AE2B490 , 32'hF4ADE3C0 , 32'h04828D30} , 
{32'h08134EC0 , 32'h02C1DA48 , 32'h02DF1A4C , 32'hDC91E400 , 32'hFD2A3FE8 , 32'hFBA8A968 , 32'hF4CFD960 , 32'hFF96EE6A , 32'h028E8860 , 32'h010290D0 , 32'hF0CF9310 , 32'h0FC1D480 , 32'hF459B510 , 32'h1BA05480 , 32'h1D6C64A0 , 32'h0AD2DB80 , 32'h0DBC9110 , 32'h0BB8DBF0 , 32'h105E58E0 , 32'h0B42BCF0 , 32'h0C3C5F30 , 32'h3415A6C0 , 32'h0A58C440 , 32'h04B02858 , 32'hDA86DE80 , 32'hDCC12F00 , 32'h149EC6A0 , 32'h0250568C , 32'h25543C80 , 32'hF0FD0E30 , 32'h10B802A0 , 32'hE4F62500 , 32'hD9A63940 , 32'hDAE59A80 , 32'hF029EAB0 , 32'hFF69F346 , 32'h031D2BE0} , 
{32'h0839BA70 , 32'h10DE51C0 , 32'h20547D00 , 32'h0F9B0400 , 32'hF2697EF0 , 32'h086CBCC0 , 32'h04625A80 , 32'h0889F830 , 32'h01A6FD58 , 32'hF3312150 , 32'h00F4978A , 32'h0410FCE8 , 32'h0A7A30A0 , 32'h08E32110 , 32'hF2F33240 , 32'hFDA34BE8 , 32'h1F170540 , 32'hECFB9B20 , 32'h2AF4EF80 , 32'hF842D9F8 , 32'hF950FA18 , 32'h1B3F3B80 , 32'h0FEADFC0 , 32'hDE86BBC0 , 32'h027FB294 , 32'h0B87D360 , 32'hFB42DC00 , 32'h145223C0 , 32'hC57F0700 , 32'h12BD27C0 , 32'h33E92140 , 32'h136336E0 , 32'hF4819540 , 32'hF87BF070 , 32'hE44C2EC0 , 32'hF844FED0 , 32'hFBD7B470} , 
{32'hFC304D80 , 32'hF0E1ACB0 , 32'hFA48C3D0 , 32'hE06AB380 , 32'h01398A70 , 32'h01BAC9F8 , 32'hF487A5E0 , 32'h0B3186B0 , 32'hF8399CE0 , 32'hD255DE00 , 32'h13C35620 , 32'hE268A6E0 , 32'h232B5E80 , 32'hCEAD32C0 , 32'hE5F248A0 , 32'hF8DAC3F8 , 32'hF8F295D8 , 32'hF9A177A0 , 32'h0A51D1C0 , 32'h0E0BCB50 , 32'h0F710340 , 32'h109503C0 , 32'hF28268F0 , 32'hE8F78360 , 32'hDEC65C80 , 32'hE75B7A60 , 32'h036CA380 , 32'hDB09ABC0 , 32'hEBE91AA0 , 32'hF06812B0 , 32'h05B1EF40 , 32'hF7217910 , 32'h1072FD20 , 32'hF2033350 , 32'h19A37140 , 32'h0F3074F0 , 32'hF1477780} , 
{32'h0F372680 , 32'hF2E997A0 , 32'h101BEDC0 , 32'h0594BEC8 , 32'h0DFDC8A0 , 32'h02FE279C , 32'h022D9E24 , 32'h075EC178 , 32'hE47FBDA0 , 32'h0B189210 , 32'h052773F0 , 32'hEE38C5A0 , 32'hE8570A00 , 32'hE84A5920 , 32'hF968EEA8 , 32'hF26AED10 , 32'hEB8FE1C0 , 32'hFEAA5250 , 32'hEF2627C0 , 32'hEC4FD940 , 32'hFC1CF35C , 32'h13C23A60 , 32'h07131F00 , 32'hFDD5CEC4 , 32'h0BB41F90 , 32'hDA28A200 , 32'h0D890520 , 32'hE8FBC740 , 32'hF7395750 , 32'h20DAF100 , 32'hE983E500 , 32'hE9274280 , 32'h15E7D220 , 32'hFD646D44 , 32'hB42CFD80 , 32'hE832FB60 , 32'h05EE77A8} , 
{32'h0C36A4C0 , 32'hE39C73C0 , 32'hF0E38F20 , 32'hF5C15DE0 , 32'h15B722E0 , 32'hE6B128C0 , 32'hFDAE1838 , 32'h310CBC80 , 32'h26989CC0 , 32'h16C8DD00 , 32'hDE680580 , 32'hF3835F30 , 32'hFB0FAC58 , 32'h1A12E560 , 32'hE2F6F100 , 32'hD94D7FC0 , 32'h1EE78900 , 32'hE47A9D40 , 32'hF6AEC210 , 32'hF83B7148 , 32'h135324C0 , 32'h1D0A8340 , 32'hF47DD730 , 32'h05DDF530 , 32'hF86C4A88 , 32'h08525BB0 , 32'hF55DC350 , 32'hF5A751D0 , 32'h06D97508 , 32'h15B67CE0 , 32'hFD56F490 , 32'h0EA94E20 , 32'h14386840 , 32'h04C24730 , 32'h0BF47E80 , 32'h04C3F5B0 , 32'h11829DA0} , 
{32'hE9F94580 , 32'h05A1D288 , 32'hFBA71A28 , 32'hFE6B16D4 , 32'hFBBF7DA8 , 32'hFD5F8F10 , 32'hFF27DFAF , 32'h11E60740 , 32'h0ECE34F0 , 32'hE64A0900 , 32'h161FE580 , 32'h090D1210 , 32'h15A193A0 , 32'h04389750 , 32'hEFB52A20 , 32'h18124080 , 32'hFAC94CF0 , 32'hFCB81EE4 , 32'hE193A4E0 , 32'h12CE8AE0 , 32'h1C886840 , 32'h04F8CFE8 , 32'h08F893F0 , 32'hEEF89C40 , 32'hEBF6F0A0 , 32'h10056EE0 , 32'hE4404420 , 32'hF6B5DFC0 , 32'h049911A8 , 32'h0744B420 , 32'hE6F76360 , 32'h093B2F20 , 32'hCC47C500 , 32'h1E0B2B20 , 32'hE642ACC0 , 32'hCF999DC0 , 32'h242A9780} , 
{32'hFCEC4234 , 32'hFAEEBAB0 , 32'hE6090300 , 32'h0CB45620 , 32'hEA3CFC20 , 32'h0BA31B90 , 32'h06B618C8 , 32'hFFAE585C , 32'hEAAEEB60 , 32'hE0DE88C0 , 32'h0B092A30 , 32'h02309930 , 32'hE42541A0 , 32'hFD4C0D50 , 32'h20909C40 , 32'hB2EE2E80 , 32'h094ECB50 , 32'h072571D0 , 32'h07333248 , 32'hFE708F70 , 32'h339249C0 , 32'hFC11E01C , 32'h19EC59E0 , 32'hED78C5C0 , 32'h08EE8BD0 , 32'hFEA66D8C , 32'hF4E24DE0 , 32'h13185700 , 32'h0AA9E800 , 32'hF3EC87C0 , 32'h0761CD78 , 32'hF4458100 , 32'h06FB7C18 , 32'h11004460 , 32'h0729EDE0 , 32'hF0FBDBE0 , 32'h02B50934} , 
{32'hDC99D480 , 32'h20EA7C80 , 32'h1730E880 , 32'hE42DEF20 , 32'hE7E3F0A0 , 32'hE3938920 , 32'hEED354E0 , 32'hF74EFE60 , 32'h21937F00 , 32'hF8024580 , 32'hF8DE27E0 , 32'hDF41ABC0 , 32'h094058F0 , 32'hF48F7100 , 32'h038068E8 , 32'hE768FAC0 , 32'hF6E5C700 , 32'h089761E0 , 32'hFDF9A240 , 32'hF00DC900 , 32'h08EFE0E0 , 32'hF9CF22B0 , 32'hD0432AC0 , 32'h2592A040 , 32'hFF3905F2 , 32'hF6A34BD0 , 32'hFF24F62F , 32'h2FC93800 , 32'hF6DD8260 , 32'h06469728 , 32'h04986A68 , 32'hF430C750 , 32'h03C1BA0C , 32'h01560B9C , 32'hF15113B0 , 32'hE6A05640 , 32'hF7704A30} , 
{32'h017D7CBC , 32'hD0E0F180 , 32'hFC71286C , 32'h0C4875D0 , 32'hF33BC7F0 , 32'hF51FB940 , 32'hFAA851B0 , 32'hE3708CE0 , 32'h00AE8A43 , 32'h126369A0 , 32'h188C5240 , 32'h1A52E0C0 , 32'h16C78580 , 32'hE5FB99C0 , 32'hE094FAC0 , 32'hFEC0B790 , 32'h1638E6E0 , 32'hE49A7420 , 32'h04E34AC0 , 32'hF712BEB0 , 32'h1D9A9BE0 , 32'hF4C1D460 , 32'h038E0CB8 , 32'h0129D38C , 32'hFA5B5BF8 , 32'h09031550 , 32'h2253EF40 , 32'h32A96A00 , 32'h044D4808 , 32'h04A0BBD8 , 32'hE0E04FC0 , 32'hF7103810 , 32'hF36B7B50 , 32'hDD8AA580 , 32'hF4D87A10 , 32'h0E5FF370 , 32'h081B1EB0} , 
{32'hF131DA70 , 32'h08E808B0 , 32'h2D19E5C0 , 32'h16811000 , 32'h0EE38580 , 32'h0A642F90 , 32'h47416880 , 32'hF65F0880 , 32'h018EF334 , 32'hE66E4C00 , 32'h09CDC970 , 32'hEE2E9560 , 32'hF9B638F8 , 32'h141CE580 , 32'hF9988950 , 32'hFEE88FD0 , 32'h0CE63B30 , 32'hE55DA5C0 , 32'hF4EA1E00 , 32'h12A98C40 , 32'h1C4172A0 , 32'hFC341E90 , 32'hF95C6188 , 32'h252B6C80 , 32'h0B2FCEE0 , 32'h03FE991C , 32'h0D18AB60 , 32'hE63D6AE0 , 32'h04DB4CB0 , 32'h0396D820 , 32'h0469ED28 , 32'hEB69AB80 , 32'hFD3329DC , 32'hDE9A6100 , 32'h1051EFE0 , 32'hFC0D0530 , 32'h06873300}
};

logic signed [31:0] US_2 [300][100] ='{
{32'hF34311C0 , 32'h7FFFFFFF , 32'h48BF6080 , 32'h3338DA80 , 32'h147EE6E0 , 32'hE87B4B60 , 32'h26B10C40 , 32'h01F31E14 , 32'hCE49DB00 , 32'hD1750200 , 32'hDA2A3AC0 , 32'h19F424C0 , 32'h0DE8D470 , 32'hDA4D5100 , 32'h16FAC2E0 , 32'hF5103AB0 , 32'hE187CA00 , 32'h1068B680 , 32'h087D1000 , 32'hF1E6E4C0 , 32'h03FA18C0 , 32'hE0F3A4C0 , 32'h27DE35C0 , 32'hEE27A360 , 32'hD45C5C40 , 32'hE8F33DC0 , 32'hF081F770 , 32'hEC97CE40 , 32'h0915C190 , 32'hF571C2E0 , 32'hFF596CE6 , 32'hFF716B3D , 32'hE1386C20 , 32'hFF7983D2 , 32'h05D25118 , 32'h04D88FF0 , 32'hFD43BE64 , 32'hE7123FC0 , 32'hF98058E8 , 32'hFFEAA9BB , 32'hF5E41AA0 , 32'hF952B3E8 , 32'h029E22D4 , 32'h25E63300 , 32'hE51CDFA0 , 32'hEEA79D00 , 32'hFD4B3690 , 32'hF83E8630 , 32'h0674D2C8 , 32'h0BD94320 , 32'hFFF5C64D , 32'h047E9808 , 32'hFE6E82F8 , 32'h02680AB8 , 32'hF272EF10 , 32'h03E79034 , 32'hF5A2F190 , 32'h07DAFC08 , 32'h0D35B980 , 32'h11D5D980 , 32'hFE31DB50 , 32'h05B353A8 , 32'h051BA0F8 , 32'h052AA2C0 , 32'h04595D68 , 32'hFFF6FB5E , 32'hFA414A58 , 32'hF6E99D40 , 32'h068200E0 , 32'h0085501A , 32'h06ED3D20 , 32'h02ACD400 , 32'h0085E8F3 , 32'h0E15CF50 , 32'hFC2280D8 , 32'h0496E120 , 32'hF7DEB020 , 32'h02683B9C , 32'h0B2D1860 , 32'hFACBFBA0 , 32'h057B33D8 , 32'h023FE984 , 32'hFBBD0298 , 32'hF76F7F00 , 32'hF6D37990 , 32'hFE1B348C , 32'h0453DB50 , 32'hFD6FCF7C , 32'hFAEF7B98 , 32'h005B1F9B , 32'h00014F2F , 32'h00019D0F , 32'hFFFF79AB , 32'hFFFCC74B , 32'h00035193 , 32'h00002D75 , 32'hFFFF7665 , 32'hFFFE4899 , 32'h000009F5 , 32'hFFFE41A3} , 
{32'h3D39CF00 , 32'h7FFFFFFF , 32'h3695EF80 , 32'h6EA88400 , 32'hFFD5C48C , 32'hA6ECD080 , 32'hECB5AA00 , 32'h60C98F80 , 32'h2CB0F400 , 32'h538C0880 , 32'h07E3C5D8 , 32'h08BF25D0 , 32'h18096360 , 32'hE67B6E80 , 32'hE31AA860 , 32'hE6A709C0 , 32'h08BDFF40 , 32'h30F7D180 , 32'h50E5E300 , 32'h0E2B0C90 , 32'hF16545C0 , 32'hE2198980 , 32'hC197D040 , 32'hEE737040 , 32'h06BBBBD8 , 32'h043A7998 , 32'hD4F1A680 , 32'h02B708E0 , 32'h00EC6370 , 32'h20733C00 , 32'h1E6C1880 , 32'h03E23A2C , 32'h03756284 , 32'h0EEF6270 , 32'h07BFCA38 , 32'h0E490380 , 32'hFC67F164 , 32'hEC0BC340 , 32'h1E837800 , 32'hE7E28FC0 , 32'h0B7E2F90 , 32'hF5203DA0 , 32'h2008C980 , 32'hF7F75F60 , 32'hFF88E832 , 32'h089E2D10 , 32'h136B5180 , 32'h0318CEFC , 32'hF5FFA0B0 , 32'hFD20DA60 , 32'h042E91F8 , 32'h12E32B00 , 32'hEEDA4640 , 32'hF4DA80F0 , 32'hF87DEFD0 , 32'h01E4642C , 32'hF50809E0 , 32'hFFFF9A79 , 32'h06E75480 , 32'h0BAFE200 , 32'h01C62940 , 32'hFA2BD2A8 , 32'h139D5B80 , 32'hFD087468 , 32'h044BDBE8 , 32'h0385C240 , 32'h033D81C8 , 32'hFA6A3CD8 , 32'hFB100638 , 32'hF743E1C0 , 32'hF41AC420 , 32'hFD1AFFBC , 32'h07CCCF90 , 32'h00D8BBA9 , 32'hFE75A494 , 32'hF60931D0 , 32'h049D7590 , 32'hFC27C978 , 32'h04DF45E8 , 32'h03F8F394 , 32'h081F6010 , 32'h042137B0 , 32'h03147D20 , 32'h0271D930 , 32'h00BAD040 , 32'h05CC2E98 , 32'h01B7D3A8 , 32'hFF1F3D15 , 32'hFC3D1640 , 32'h00CB9AF2 , 32'hFFFFB465 , 32'h00003339 , 32'hFFFE7EA1 , 32'hFFFBFA69 , 32'hFFFE1DB4 , 32'h0001702D , 32'hFFFF98D7 , 32'h00038A39 , 32'hFFFF7F4F , 32'hFFFEE7DA} , 
{32'h0005DF8F , 32'hFFF633CF , 32'h00023CDA , 32'hFFFBF484 , 32'h000089B1 , 32'hFFFDC6BE , 32'h00018C65 , 32'h00059BA2 , 32'h00070BF9 , 32'hFFFB6FE6 , 32'hFFF6891D , 32'h00011FAB , 32'h00024FAB , 32'hFFF96ED8 , 32'h0006BE61 , 32'hFFFC3BA6 , 32'hFFF51EBA , 32'h0002380C , 32'hFFFE9DDF , 32'hFFFAE902 , 32'hFFFBB820 , 32'h00021ABE , 32'hFFFAC2F4 , 32'h0009C01A , 32'h000446B7 , 32'hFFFE322E , 32'h000649D4 , 32'hFFFFBD30 , 32'hFFFE5ACC , 32'h000310A5 , 32'h00007D4D , 32'h0001AEC1 , 32'h00011A2B , 32'h00011165 , 32'h00040560 , 32'h00044FD7 , 32'hFFFB2003 , 32'h00073262 , 32'hFFFCFB39 , 32'h0007036B , 32'hFFF70FBE , 32'hFFF8C3A4 , 32'hFFFE6129 , 32'h00031D79 , 32'h0003F34C , 32'h0005C4F5 , 32'hFFFFDC54 , 32'hFFFAA24F , 32'hFFFA42F8 , 32'h00031D3D , 32'h00037DDA , 32'h000581AB , 32'h0003F19B , 32'h0005CEEA , 32'hFFFC161E , 32'hFFFF5503 , 32'h0006E98D , 32'h00073944 , 32'hFFFF08CD , 32'hFFF903B4 , 32'hFFF93398 , 32'hFFFF1CC7 , 32'hFFFDA6D6 , 32'h0005CE19 , 32'h0002DE29 , 32'hFFFFD7D8 , 32'h0003E58B , 32'h0003D403 , 32'hFFFCECB9 , 32'hFFFA0913 , 32'hFFFCA5FB , 32'hFFFFB8F7 , 32'hFFFC062A , 32'h00082C65 , 32'hFFF9CBAF , 32'hFFF9C222 , 32'h0001B538 , 32'h000048A5 , 32'h0000B75C , 32'hFFFD3FD4 , 32'hFFFC62E8 , 32'hFFF23989 , 32'h00014F3B , 32'hFFFB2BEC , 32'h00014A8E , 32'hFFFE2FC5 , 32'h0007C357 , 32'h000110C0 , 32'h0007C041 , 32'hFFFF7944 , 32'h0000C822 , 32'hFFF7108B , 32'hFFFA309E , 32'h0002A62F , 32'hFFFEB3C6 , 32'hFFFAD6C0 , 32'h00024F72 , 32'hFFFEE9B0 , 32'hFFF9B9F7 , 32'hFFFC3DF0} , 
{32'hD0AA1500 , 32'h11CCE6A0 , 32'hFAFC7118 , 32'h48183180 , 32'h05D2CC10 , 32'h022641B4 , 32'hDC1FA380 , 32'hD8A56540 , 32'hE0A23440 , 32'h2C53F980 , 32'hF6F6BF10 , 32'hEC42A6E0 , 32'hC4C94700 , 32'h20FFC740 , 32'h0093173F , 32'h07DBDD90 , 32'h0A42D6F0 , 32'h33F47C40 , 32'hF97C4F70 , 32'hE4BEEEE0 , 32'hEE2F99A0 , 32'h2B544400 , 32'hCB8BBCC0 , 32'hFC848DF4 , 32'hF6404730 , 32'h169D48E0 , 32'h0BCC7820 , 32'hF0B4E3D0 , 32'hE2EE5960 , 32'hDD5EE8C0 , 32'hFE6BFC04 , 32'hEF7F56A0 , 32'h2D0DED00 , 32'h12018FE0 , 32'hF3F46E30 , 32'h11392740 , 32'h06BDD638 , 32'hF3CAFCD0 , 32'h1D827C80 , 32'hFB92CB70 , 32'hEE223500 , 32'hED377CE0 , 32'hDDA52580 , 32'hFF2C3372 , 32'hFB15FF68 , 32'h18ECF840 , 32'hF756F2C0 , 32'hEE5C69E0 , 32'hFDA62CA8 , 32'hFEAA8770 , 32'hF7E5C630 , 32'hFA60FE30 , 32'h0E2DB0D0 , 32'hF5CD7360 , 32'h0B5492A0 , 32'h0058049A , 32'hFBE13AA8 , 32'hFBA9BE00 , 32'h05E08398 , 32'h01EC10DC , 32'hFB959E10 , 32'h023B7304 , 32'h0122F92C , 32'h0159B0AC , 32'h06FAB9C8 , 32'hED5FF220 , 32'hF52DDF90 , 32'hFDC07030 , 32'hFAA145C0 , 32'hFF017280 , 32'h0043D7C7 , 32'h0ECCD940 , 32'h00008CD6 , 32'h01D6E2AC , 32'h0F40BC80 , 32'hFFD36FAD , 32'hF67ED6F0 , 32'h0198414C , 32'h0ACCBA40 , 32'h04720780 , 32'hFF3D9D18 , 32'hFEF52594 , 32'hFF44EE70 , 32'hFCF7C1EC , 32'h04D598F8 , 32'hF824A6B8 , 32'h02466884 , 32'h01C5DA30 , 32'hFDC10D98 , 32'hFF4AC428 , 32'h00010ED5 , 32'hFFFF007D , 32'h000137EB , 32'hFFFCC77F , 32'h0003363A , 32'h0002549A , 32'h0001981B , 32'h00018F80 , 32'hFFFBDCF9 , 32'hFFFEF2CA} , 
{32'h0004E9AD , 32'hFFFB65B5 , 32'hFFFE059F , 32'hFFFFCAD5 , 32'hFFFD96B1 , 32'hFFFD07CE , 32'h00027E3E , 32'hFFFE9B55 , 32'h00028544 , 32'h0001E84B , 32'h00025AF7 , 32'hFFFE1F00 , 32'hFFFEB15B , 32'h00053F29 , 32'h00012968 , 32'h00043794 , 32'hFFF8A476 , 32'h00075AF3 , 32'hFFFAD20E , 32'h0004FDD7 , 32'h0000A8C3 , 32'h0003430A , 32'hFFFEDD38 , 32'h0001FDDE , 32'h00002F17 , 32'h00057D88 , 32'hFFFE9E2F , 32'h0001EE5D , 32'hFFF67963 , 32'h000342E1 , 32'hFFF773CA , 32'hFFFD91B9 , 32'h0009C57C , 32'h0005734F , 32'hFFFC5B97 , 32'hFFFF7DF9 , 32'h0002742A , 32'h00026F52 , 32'hFFFEFF75 , 32'h0004729E , 32'hFFFCE6D4 , 32'h0004A9F4 , 32'hFFFB029E , 32'h00023230 , 32'h0006DBB3 , 32'h0005B9B6 , 32'hFFF507F1 , 32'h00085941 , 32'hFFFC52A8 , 32'hFFF6E376 , 32'h0003F08C , 32'hFFFD6245 , 32'hFFFDFE13 , 32'hFFFE8B80 , 32'hFFFB3AFF , 32'h00025B8F , 32'h0008B84D , 32'hFFFB24E0 , 32'h0003C5B3 , 32'hFFF9BC50 , 32'h0003B365 , 32'h0000A07D , 32'hFFF8E788 , 32'hFFF99A3F , 32'hFFFAA5B5 , 32'hFFF4C739 , 32'h000101D0 , 32'h0000D640 , 32'h00020011 , 32'hFFFE7819 , 32'hFFFAD8CD , 32'hFFFB15FA , 32'hFFFAD443 , 32'hFFF84CD1 , 32'hFFFF0D92 , 32'hFFF97A98 , 32'hFFFEFDB0 , 32'hFFFA50E3 , 32'h000097C8 , 32'hFFFAD316 , 32'h00011461 , 32'hFFF7B8D6 , 32'hFFFB8CEC , 32'hFFFEBB98 , 32'hFFFB92DB , 32'hFFFCECA0 , 32'hFFFD7257 , 32'hFFFCCC02 , 32'h00026CBE , 32'hFFF78A16 , 32'hFFF7C844 , 32'h000044C5 , 32'h0002651A , 32'h0000B097 , 32'hFFFD6F63 , 32'hFFF7425D , 32'hFFFFB299 , 32'hFFFB0FC8 , 32'hFFFD2D59 , 32'hFFFDE571} , 
{32'hF8D9B120 , 32'hECD3D1A0 , 32'h087E6630 , 32'hF075FA40 , 32'hE4119020 , 32'h004C9302 , 32'h0FFA41B0 , 32'hDA286280 , 32'hF9183788 , 32'hF4880080 , 32'h0CAF6080 , 32'hFEFE5D94 , 32'hFB3CA430 , 32'h001F2D64 , 32'hF9CF71B0 , 32'hF80999D8 , 32'hFFC3E224 , 32'h05170FF0 , 32'hF9085270 , 32'h20FDDC40 , 32'h20A2EFC0 , 32'h08CB6910 , 32'hFBBCBC38 , 32'hD74A8600 , 32'hFD038688 , 32'h1268A100 , 32'h12F97760 , 32'h0A853240 , 32'hFE8A7974 , 32'hEB694BE0 , 32'hFE8C67C8 , 32'h0D028290 , 32'h052D3710 , 32'hF75B5570 , 32'h1ECB5900 , 32'h0D84A9A0 , 32'h007835A7 , 32'hF8896BE0 , 32'hFB28C2C8 , 32'hEAC8B9C0 , 32'h05B88F30 , 32'hFAFB3008 , 32'hF6F38E60 , 32'hF6C865D0 , 32'h051DA5E8 , 32'h1948E600 , 32'h14EC6000 , 32'hF02B4FB0 , 32'h07C38A38 , 32'hFEE20BA8 , 32'hF4F0CBC0 , 32'hF9347C90 , 32'h10D7F3E0 , 32'hFA54FFB8 , 32'hFC3B0534 , 32'h0367B65C , 32'hF3627820 , 32'h0409E8F0 , 32'h021F2BA0 , 32'hFD3D1F48 , 32'h0C70BBC0 , 32'hFCBFC448 , 32'h093FA4A0 , 32'h05FE86B0 , 32'hF96392A0 , 32'hF75C8D80 , 32'hFF80F4B1 , 32'hFE3769F4 , 32'hFADA0E88 , 32'hF40F31B0 , 32'h00E35D75 , 32'hF4A99530 , 32'hFD53BF64 , 32'h06339660 , 32'hFD53CF10 , 32'h040A0BA0 , 32'h031FF368 , 32'h05285A20 , 32'hFF3C243A , 32'hFBADE9F8 , 32'h01024348 , 32'hF9FDAE88 , 32'hF80B3230 , 32'h00F2A505 , 32'hFF8A91E5 , 32'hFCB51468 , 32'hFE90A268 , 32'hFA43A838 , 32'h059818F8 , 32'h017E8E20 , 32'h0002ED39 , 32'h000279E3 , 32'hFFFF8319 , 32'h00010A2C , 32'hFFFF73A1 , 32'h0000FB9D , 32'h0002A37E , 32'hFFFC80C9 , 32'hFFFD3E13 , 32'hFFFCF2E7} , 
{32'h000901D8 , 32'h0001004A , 32'hFFFFC5C7 , 32'h00050ED1 , 32'h0001EC1F , 32'hFFFCDC74 , 32'h0000E2D6 , 32'h0000E9ED , 32'h000B70FA , 32'h0000F8F4 , 32'hFFFF1347 , 32'hFFF9DB8D , 32'h0005CAC8 , 32'h00043377 , 32'hFFF82377 , 32'h00012679 , 32'hFFF64110 , 32'h0002B6A7 , 32'hFFFE2243 , 32'hFFF6CB02 , 32'h00010D75 , 32'h0000A5E4 , 32'hFFFFF023 , 32'h00024366 , 32'h00005D84 , 32'h0000007C , 32'hFFFF716B , 32'hFFFB60D5 , 32'hFFF23309 , 32'h000D99E2 , 32'hFFFAC765 , 32'h00015EDE , 32'hFFFD7C37 , 32'hFFFC4E4F , 32'hFFF8C82F , 32'hFFFD75A4 , 32'h000418DC , 32'h0006EF0B , 32'hFFF810A8 , 32'h0000E75B , 32'hFFF7B38A , 32'hFFFE584D , 32'hFFF925D6 , 32'h00026EE3 , 32'hFFFFF6B9 , 32'hFFFCA602 , 32'hFFFEECED , 32'h0002F1FA , 32'h0000D626 , 32'h00019F97 , 32'hFFFD461E , 32'hFFFF7BA3 , 32'h000B1750 , 32'hFFF4E014 , 32'h0000EBFA , 32'hFFF7C52A , 32'h00032C2E , 32'h0001DFA1 , 32'h0001C217 , 32'hFFFEDFBA , 32'hFFFED08B , 32'hFFFBA88C , 32'hFFFE147E , 32'hFFFA590C , 32'hFFFF19D0 , 32'h000BC2A7 , 32'hFFFFEEC0 , 32'h0004BDA9 , 32'h0002C143 , 32'hFFFE60D2 , 32'h00012232 , 32'hFFFB3527 , 32'hFFFF6A06 , 32'hFFFF2340 , 32'hFFFD94D4 , 32'hFFFF9594 , 32'h00040BB9 , 32'h00082AAF , 32'h0004C992 , 32'hFFFDBA3E , 32'hFFF9CB70 , 32'h000016CD , 32'h00017C58 , 32'hFFFE306B , 32'h0003EFFA , 32'h00045BD7 , 32'h00027C0E , 32'h0001D16E , 32'hFFFF19F5 , 32'h000172E7 , 32'hFFFFBDDC , 32'hFFF4E6BE , 32'hFFFDC5AA , 32'hFFF27259 , 32'hFFF9630D , 32'h000338F7 , 32'h0000A15A , 32'hFFF777BB , 32'h000CF677 , 32'hFFFAF0FE} , 
{32'hFFFFD112 , 32'hFFFC70BD , 32'h00058AF8 , 32'h0008128B , 32'hFFFEB644 , 32'hFFFB7C08 , 32'h0005197F , 32'h00028DA4 , 32'hFFFFE9D4 , 32'h0004EA61 , 32'h0005FC78 , 32'h000528DC , 32'h00046130 , 32'hFFFCB439 , 32'hFFFFE2A7 , 32'hFFFEC970 , 32'h00020BA2 , 32'h000531B6 , 32'hFFFBE5E7 , 32'hFFFCAB46 , 32'h00016D23 , 32'hFFFEDB31 , 32'h0006420B , 32'hFFFB3831 , 32'hFFFFD472 , 32'h0004AC23 , 32'h00064F9C , 32'hFFFFB5FA , 32'hFFF95AA3 , 32'h0003959F , 32'h0004505D , 32'hFFFBF653 , 32'h000049C1 , 32'hFFFE10CB , 32'h00007026 , 32'h0003F18A , 32'h00034CF1 , 32'h00047274 , 32'h000184DD , 32'h0004AD31 , 32'h00060460 , 32'h0003F353 , 32'h0002B834 , 32'h0002DE95 , 32'h00015A76 , 32'hFFF83CE3 , 32'hFFFFE257 , 32'h0001DCCA , 32'hFFFC4673 , 32'hFFFE68DB , 32'h0007E1E5 , 32'hFFFFEB3C , 32'hFFFAE5A1 , 32'hFFFA297F , 32'h000268C0 , 32'hFFF7D9A2 , 32'hFFFEEFF9 , 32'h0000AB9B , 32'hFFF82F61 , 32'hFFFF129D , 32'h00034825 , 32'hFFFF9AAA , 32'hFFFCCF25 , 32'h00068703 , 32'hFFFCCBFB , 32'hFFFF4A20 , 32'hFFFF6C94 , 32'h000112C7 , 32'hFFFDF673 , 32'hFFFD6F4B , 32'hFFFF2124 , 32'hFFFF0193 , 32'h0006136C , 32'h0003B247 , 32'h00028A4B , 32'hFFFCCD2C , 32'h00023E4A , 32'hFFFC5C35 , 32'hFFFB900E , 32'hFFFF2E02 , 32'h000426EF , 32'h0002591F , 32'hFFFA659C , 32'hFFFE9637 , 32'hFFFE3929 , 32'hFFF6276A , 32'h0005061D , 32'h0004312D , 32'h00011920 , 32'hFFFDE662 , 32'h0001B7FE , 32'hFFF9E259 , 32'hFFFB73EA , 32'hFFFF6D8F , 32'h0005FBD5 , 32'hFFFDD391 , 32'hFFF72089 , 32'hFFFD1601 , 32'h00053961 , 32'hFFFE0CFE} , 
{32'h0004732E , 32'hFFFA094D , 32'h000287D8 , 32'h00027FBF , 32'hFFFDFF12 , 32'h00060946 , 32'h0005A5FB , 32'h0002494C , 32'hFFF87234 , 32'h000514CA , 32'h000730DC , 32'h00073B30 , 32'h0009DEBB , 32'h0000C5FA , 32'h00072463 , 32'hFFFC6E41 , 32'h00000391 , 32'hFFF9579D , 32'h0001FA28 , 32'hFFF6895A , 32'hFFFD2EE4 , 32'h0009340D , 32'hFFFFB48C , 32'hFFFC1ECD , 32'h00024FC7 , 32'hFFFD989B , 32'hFFFEA24F , 32'hFFFD97BE , 32'hFFF6E042 , 32'hFFFCF21E , 32'hFFF91B71 , 32'hFFFF12F1 , 32'h00001E22 , 32'hFFFA2717 , 32'h0005F578 , 32'h00010CCB , 32'h0001B033 , 32'hFFF70976 , 32'h0002C43B , 32'hFFFD0501 , 32'hFFFECBDF , 32'h0000FF21 , 32'hFFFA1EF1 , 32'h00093EF6 , 32'hFFFC85AF , 32'hFFFF37C2 , 32'h0003FEC0 , 32'h00076C45 , 32'hFFFF4F8A , 32'hFFF60522 , 32'h00091CCE , 32'hFFFF9FA5 , 32'hFFFF20E2 , 32'hFFF87B39 , 32'hFFFC564A , 32'h000404A5 , 32'h0003CF4A , 32'h0000873D , 32'hFFFCD172 , 32'h00027501 , 32'h00049339 , 32'h00096E3A , 32'h0002555F , 32'hFFFBA1B4 , 32'hFFFE729E , 32'hFFF865A0 , 32'h0006D805 , 32'h00003EA4 , 32'hFFF64B8C , 32'h0004C465 , 32'hFFFF88C2 , 32'hFFFBECC3 , 32'h000496EB , 32'h00052B84 , 32'h00085AC7 , 32'h0002BC26 , 32'hFFF8FCD2 , 32'hFFFE329B , 32'h0005B554 , 32'hFFFED2E3 , 32'h000B92CE , 32'h0001DF71 , 32'h000464D7 , 32'hFFFAE585 , 32'hFFFC9FA6 , 32'hFFFB9F4A , 32'h00056B87 , 32'h00082C5A , 32'hFFFF86A4 , 32'h0001F224 , 32'hFFFBC0C1 , 32'h0000EDCF , 32'h0001BB78 , 32'hFFFA0AE9 , 32'h000A3D2B , 32'hFFFD7CFE , 32'hFFFF84EB , 32'hFFFA73F0 , 32'h00022C7A , 32'h00014D15} , 
{32'h00057F49 , 32'hFFFB12EC , 32'h0005BCF3 , 32'h000788EB , 32'hFFFB8403 , 32'hFFFDA0FF , 32'hFFF76AC5 , 32'hFFFE22F8 , 32'h0000A20D , 32'hFFFC094E , 32'hFFFB4735 , 32'h000324FE , 32'hFFFEAE22 , 32'hFFFD2D11 , 32'hFFFB6C4F , 32'h000E37A6 , 32'hFFFBF9FB , 32'hFFFDA0E6 , 32'h0004B066 , 32'hFFFBB8A2 , 32'h0005ECB6 , 32'hFFFC285C , 32'h0003A314 , 32'h00008E82 , 32'hFFFC7CF7 , 32'hFFFF6811 , 32'h000505DC , 32'h00056EDD , 32'h000382AA , 32'hFFF7FF8E , 32'hFFFFB249 , 32'hFFFD21CC , 32'h00068D79 , 32'h00074A6D , 32'h00026705 , 32'h000169B9 , 32'h0009E6AD , 32'h000016DE , 32'h0004175D , 32'h0007CF4F , 32'h000440A1 , 32'hFFFB07DD , 32'hFFFDDFB2 , 32'h00087D8A , 32'hFFFF68D9 , 32'hFFF46FAB , 32'hFFF8F2CD , 32'hFFFB2AED , 32'h0000933C , 32'hFFFCDC56 , 32'h000161F6 , 32'h00082B20 , 32'hFFFB1CDD , 32'hFFFFD3AE , 32'hFFFBA913 , 32'h00060372 , 32'hFFF651C8 , 32'h0003BEC9 , 32'h00074784 , 32'hFFFC31F7 , 32'hFFF7E3FA , 32'h000469A6 , 32'hFFFCF11D , 32'h00059ACF , 32'hFFF6042B , 32'h00039485 , 32'hFFFE4C46 , 32'h0003D523 , 32'h00029452 , 32'hFFF737F2 , 32'h00031218 , 32'hFFFC7240 , 32'h0005D769 , 32'hFFFD11BD , 32'h00082C08 , 32'h000714AC , 32'hFFF92E75 , 32'h000AA26D , 32'h0000FF4B , 32'hFFF7ADF5 , 32'h0007CA54 , 32'h00063698 , 32'h0005BBD1 , 32'hFFFBC7B1 , 32'hFFF4DE33 , 32'hFFFA9699 , 32'h00051AC1 , 32'h0004EAC0 , 32'h0007CFB8 , 32'h0007917B , 32'h00073936 , 32'hFFFFCC97 , 32'h00053689 , 32'hFFFA2392 , 32'hFFF8831C , 32'h0002C1C5 , 32'h0004EC30 , 32'hFFFCF4D2 , 32'h000238F6 , 32'h0000FC03} , 
{32'h3D398740 , 32'hDF8AFDC0 , 32'h0F66ADA0 , 32'hF63B4DB0 , 32'hEC78C580 , 32'h1CE668A0 , 32'h3F699F40 , 32'h107953E0 , 32'hD47E6000 , 32'h1B8575E0 , 32'h1352E3C0 , 32'hEEDB8F00 , 32'hFA6A77F8 , 32'hF9418598 , 32'hFB63B110 , 32'h2BA33080 , 32'hEFD7CC00 , 32'h1F22C180 , 32'hEC57B3E0 , 32'h0FC91380 , 32'hE41E8E00 , 32'hF6425F00 , 32'h10D8EE60 , 32'h16A80180 , 32'hF4C57030 , 32'h119FB780 , 32'h0C26E420 , 32'h057A3060 , 32'h0F50A6C0 , 32'hFB698B60 , 32'h141B9E20 , 32'h0B7DC530 , 32'hE25FE9A0 , 32'hD61DC380 , 32'h093B98A0 , 32'h0ADB5BF0 , 32'hEDA53A20 , 32'h12386360 , 32'h0C6D0270 , 32'hF4AF6BE0 , 32'hF3896060 , 32'h03044418 , 32'hD91A6400 , 32'h124CEC00 , 32'h02E743D0 , 32'h11EA2700 , 32'hFD469CE0 , 32'hFB6187D0 , 32'hFB3371B8 , 32'hFF711BBD , 32'hF434FA00 , 32'h0B38E300 , 32'hE5F4D7C0 , 32'h14794C80 , 32'h0AD36EE0 , 32'h08F733D0 , 32'h08856090 , 32'hFF293DD0 , 32'hEF2653E0 , 32'h00574DB3 , 32'hFE26E92C , 32'hFE63FA50 , 32'hFC63E6F0 , 32'h025C6E78 , 32'h06F7C6A0 , 32'hFE827630 , 32'h07FF22B0 , 32'hF7CD0D60 , 32'hF69B8490 , 32'h029DFA0C , 32'hFB3C1098 , 32'hFDC185B8 , 32'h0FAC8FB0 , 32'h017A3954 , 32'h06359658 , 32'h0278D854 , 32'hFC9B7618 , 32'h10702980 , 32'h01A5FEB4 , 32'h044E5570 , 32'h016119EC , 32'h01A46964 , 32'hF73558C0 , 32'hFA91F308 , 32'h0364ED1C , 32'hFDABFD38 , 32'hFCF85A24 , 32'hFE5B9060 , 32'h0266C860 , 32'h00E96A9A , 32'h0000BD7F , 32'h000272EC , 32'h0000A1B8 , 32'hFFFB043F , 32'hFFFE1976 , 32'hFFFE584B , 32'hFFF74205 , 32'hFFFF4EC7 , 32'hFFFD10CF , 32'hFFFDEE46} , 
{32'h46B3C400 , 32'hEB63A680 , 32'h969A5980 , 32'hD7BBB680 , 32'h45D8DA80 , 32'hF6560E40 , 32'hC9966C00 , 32'h0BDD8A80 , 32'hEEB8D840 , 32'hFB572DD0 , 32'h883A7180 , 32'h193C65E0 , 32'hEE31AFA0 , 32'h0D9C7D20 , 32'h20F70240 , 32'hEACD7DE0 , 32'h064E6270 , 32'h097AF2E0 , 32'h14C1EFE0 , 32'h0A556E70 , 32'h07273F90 , 32'h34FD9F00 , 32'h266B5780 , 32'h23C7CDC0 , 32'hE6A61780 , 32'hEF39FC80 , 32'hF1DDF020 , 32'hE1D8E440 , 32'h0E30EE20 , 32'hFE97F808 , 32'h018A54CC , 32'h12A68E60 , 32'h09A28D60 , 32'hF3E1A5A0 , 32'h04C8B050 , 32'h11DE0360 , 32'hE9B78240 , 32'hEC57A760 , 32'h05D74310 , 32'hE0028EC0 , 32'hFCE89F74 , 32'h0DCB9AE0 , 32'hE3A19280 , 32'hF62100F0 , 32'hFE59A944 , 32'hED7EDC40 , 32'h166AD940 , 32'h009CA73F , 32'h04033D88 , 32'hFCDB4D04 , 32'h1033EDE0 , 32'h0194A864 , 32'hF9E1EE88 , 32'hFE2F03BC , 32'hFA96E838 , 32'hFAF8AA78 , 32'h058677B8 , 32'h04360260 , 32'hFEF1D678 , 32'hF352CE90 , 32'hF2406BD0 , 32'h0480E200 , 32'hFAABE1B0 , 32'hF8DB34F8 , 32'hFCDDABB8 , 32'h07500170 , 32'h0584D490 , 32'h033D4454 , 32'h07B22640 , 32'hFE5CF4EC , 32'hFDD18150 , 32'h0362E448 , 32'hFFC930B2 , 32'h02BA4970 , 32'h03303B0C , 32'hFE676DFC , 32'h05E14CE8 , 32'hF39AB8F0 , 32'hFE45AF1C , 32'h05E98918 , 32'h098D5140 , 32'h09F628A0 , 32'h04C332C8 , 32'hFB567AE0 , 32'h019F96C0 , 32'hFF9EA024 , 32'hFD84E468 , 32'hFFFD1ED1 , 32'h0399636C , 32'hFE060C0C , 32'hFFFDC0A3 , 32'h0002B8B9 , 32'hFFFA42E9 , 32'h0000AABC , 32'hFFFC4E57 , 32'hFFFE2A35 , 32'hFFFFE161 , 32'hFFFECE94 , 32'h0000A994 , 32'hFFFC89B9} , 
{32'h148AD920 , 32'h42CA8E00 , 32'hEE07F8C0 , 32'h0A5B6090 , 32'hED75A120 , 32'h0E193F00 , 32'hCC963B40 , 32'h0DF59030 , 32'hEB88F960 , 32'h191B1DA0 , 32'h034C5F48 , 32'h03C30500 , 32'hF0A34E60 , 32'hE1304BA0 , 32'hE0FB1B60 , 32'h020C6C90 , 32'h0A15CCB0 , 32'hFFB4276F , 32'h1DCA9FE0 , 32'hFF287F57 , 32'hFE17D35C , 32'hE75776E0 , 32'hF6A988E0 , 32'hF6E04350 , 32'h029C1670 , 32'h09A1C170 , 32'h06F0E0A8 , 32'hFBAE2E08 , 32'h12F68B20 , 32'h0E8EB2B0 , 32'hFB94BD38 , 32'hF1DFE1D0 , 32'h178519A0 , 32'hF5DB1CC0 , 32'h1A4F3220 , 32'h0D65B6D0 , 32'h0268B688 , 32'h0BA52050 , 32'hFDF075FC , 32'hE874FAC0 , 32'hFE6247F4 , 32'h14905AE0 , 32'h1F360280 , 32'h055C0740 , 32'hF6A576B0 , 32'hD93C5000 , 32'hEDCD3AC0 , 32'hECC08B80 , 32'h06BF34C0 , 32'h0EF00CB0 , 32'hEE570DA0 , 32'h01821634 , 32'hFAEED950 , 32'h1F5AE980 , 32'hEE1568C0 , 32'h0A128440 , 32'hFF311A82 , 32'hFACD9AF8 , 32'h08571390 , 32'hFBFAC520 , 32'hF6A52280 , 32'h03770134 , 32'hED5374A0 , 32'hF0101480 , 32'h0F6475F0 , 32'hFEAD8F18 , 32'hF6217E10 , 32'h01A0EAE8 , 32'hFB8ECA38 , 32'h06112BD0 , 32'h04577290 , 32'hFB4CBA40 , 32'hF57A8130 , 32'h0B9F4290 , 32'h051F4970 , 32'h052D6450 , 32'hF20A11D0 , 32'hFAA463F0 , 32'hFE41293C , 32'hFBEBF678 , 32'hFD23B7CC , 32'hFD554C58 , 32'hFD6B8A28 , 32'hFED76C00 , 32'h062C2FE8 , 32'h0190FA08 , 32'h0340BDBC , 32'h0299A374 , 32'h02778448 , 32'hFFD94820 , 32'hFFF995C7 , 32'h0000831C , 32'h00025EB2 , 32'hFFFBBC49 , 32'hFFFB98B5 , 32'h0001C73D , 32'h00020584 , 32'hFFFEC180 , 32'h0000B28B , 32'h0000163B} , 
{32'h000139E7 , 32'h00001015 , 32'h0003186D , 32'hFFF9E163 , 32'hFFFA2786 , 32'hFFFF40F1 , 32'h00055272 , 32'hFFF8F711 , 32'hFFFEBA34 , 32'hFFF95901 , 32'h0007A54F , 32'h0000B975 , 32'h0000A8F9 , 32'h0003F1D1 , 32'h00078E50 , 32'h0004594B , 32'h0002E825 , 32'h0000DF09 , 32'h0006F7EE , 32'h00022ABD , 32'h00015371 , 32'hFFFE2EEF , 32'hFFFB1EA3 , 32'h00040C7E , 32'hFFFB282B , 32'hFFF8C0D3 , 32'hFFFF123F , 32'h00005668 , 32'h00045177 , 32'hFFFEEC87 , 32'h00018A29 , 32'h0004DB29 , 32'hFFF9AB5F , 32'h000189B1 , 32'hFFFD1C87 , 32'hFFFD4B56 , 32'h00003DC4 , 32'h0005998F , 32'hFFF9DBCE , 32'h000345ED , 32'hFFFA7D93 , 32'hFFF8468D , 32'hFFFF49B1 , 32'h00007C7C , 32'hFFFE1141 , 32'hFFF78014 , 32'hFFF8C179 , 32'h0000E6B2 , 32'h0005199C , 32'hFFFC48F7 , 32'hFFFB2BD0 , 32'hFFFD8FD8 , 32'h0009CB17 , 32'hFFFC33DD , 32'h0000BB5A , 32'h0000EF87 , 32'hFFFCDCB6 , 32'h00015113 , 32'hFFFDB149 , 32'h00014493 , 32'h00030C23 , 32'hFFF9B65B , 32'h00003AA1 , 32'h00018C03 , 32'hFFFCE72A , 32'h0002F296 , 32'h00031B52 , 32'hFFFC8E7A , 32'hFFFE3AB9 , 32'h0006FCA0 , 32'h0005205C , 32'hFFFD78C6 , 32'hFFFACB3E , 32'hFFFF5DA5 , 32'h000459AA , 32'h000080BC , 32'h0000EEDF , 32'hFFFB919D , 32'h00007F8A , 32'h0002714B , 32'h00027AF5 , 32'hFFFF5EE2 , 32'h0001D081 , 32'hFFFEE637 , 32'h0005A5BC , 32'hFFFE437B , 32'hFFFE039C , 32'hFFFC8290 , 32'hFFFFC03B , 32'h0002A3F9 , 32'h0003806C , 32'hFFFB883D , 32'hFFFE5CA0 , 32'h0008637A , 32'h0003D8FE , 32'h000443AF , 32'h00034CF1 , 32'hFFFBBD79 , 32'h00007A27 , 32'hFFFBBE60} , 
{32'h000717B4 , 32'hFFFD9021 , 32'h0008857C , 32'hFFFFF335 , 32'h00023E2B , 32'hFFFCABE6 , 32'h00014A13 , 32'h00005140 , 32'hFFFEE087 , 32'hFFFE43EF , 32'hFFF90051 , 32'hFFFBD9EB , 32'hFFFE9E2C , 32'hFFFCD955 , 32'h0000DC71 , 32'hFFFA93A3 , 32'h0002E7ED , 32'hFFFF9AEF , 32'hFFF9BE26 , 32'h000375B1 , 32'hFFFCCA6C , 32'h00011814 , 32'h000290C1 , 32'hFFFCB346 , 32'h0000CB0B , 32'h0004F343 , 32'hFFFA405F , 32'hFFF63E40 , 32'h00013D11 , 32'h000086BC , 32'hFFFED2D4 , 32'h0002632F , 32'hFFFB906E , 32'hFFFDD20B , 32'hFFFB5063 , 32'h00005ED6 , 32'h00014432 , 32'h000CA2AE , 32'hFFFE1313 , 32'hFFFDFEC8 , 32'h0001196C , 32'h00087317 , 32'h0001936A , 32'h0007E760 , 32'h0003F8F9 , 32'h00021967 , 32'hFFF996D1 , 32'h0002CA80 , 32'h0007A7BF , 32'h00015959 , 32'hFFFAEF00 , 32'h0000AF17 , 32'h00027EE1 , 32'hFFFAB561 , 32'hFFFF7E6D , 32'h0003BF2D , 32'hFFF93D92 , 32'hFFF83B00 , 32'h00011A58 , 32'hFFFFCF72 , 32'hFFFD7C61 , 32'hFFFEFFA7 , 32'h0005AE7A , 32'hFFFD9ED8 , 32'hFFFD596A , 32'hFFFCA3B3 , 32'h00015C02 , 32'h0000D20A , 32'h00006DF6 , 32'hFFFEE239 , 32'hFFFD6CE0 , 32'h000875BC , 32'hFFF1B3FA , 32'h000742DC , 32'hFFFF8990 , 32'hFFFBCB92 , 32'h00040642 , 32'hFFFC0E48 , 32'h0004CBA1 , 32'hFFFBBDE5 , 32'hFFFED21D , 32'h000BF763 , 32'hFFF84BC2 , 32'hFFFB63D8 , 32'h00000129 , 32'h00027F9A , 32'h000429B3 , 32'hFFFCC799 , 32'hFFFC6A6B , 32'hFFFF6664 , 32'h0004A8C8 , 32'hFFFFABF7 , 32'h0003CFB8 , 32'hFFFBB699 , 32'hFFF9CBC7 , 32'hFFFFCD94 , 32'hFFFD1A97 , 32'h0000AA49 , 32'h0001C582 , 32'hFFFAE593} , 
{32'h7FFFFFFF , 32'h29291F80 , 32'h55EBD980 , 32'hE003F3E0 , 32'hDA6A2140 , 32'h05270480 , 32'h0A532E10 , 32'h06DC6FE8 , 32'hD0C21D40 , 32'hE3F34EA0 , 32'hB6257880 , 32'h1C765BC0 , 32'h02F7BE6C , 32'h044D6E90 , 32'hEB853660 , 32'hE7C2A180 , 32'h24F5D7C0 , 32'hED69C9E0 , 32'h21A5FE80 , 32'h1C164F60 , 32'hEDC7E2C0 , 32'hF550CB80 , 32'hDF6D64C0 , 32'hF91B0568 , 32'hFDD91244 , 32'h12FB3960 , 32'h00DABD74 , 32'h0BE5F280 , 32'h207BFD00 , 32'h1157FDA0 , 32'hF8AABA10 , 32'h0BB31480 , 32'h069A4B20 , 32'h07743420 , 32'h0ABDE620 , 32'hE5DA1820 , 32'h11778180 , 32'hFE7D3D68 , 32'h07782060 , 32'hFE7834E4 , 32'h0BFDCD80 , 32'hFBAA2CC0 , 32'h054C13D0 , 32'hF6900F00 , 32'hEB5154A0 , 32'hEA6A8020 , 32'hFBA14BB8 , 32'hFF21ADED , 32'hF879DD48 , 32'h0229A1A0 , 32'hF2AF6D70 , 32'hF9603EA0 , 32'h1C996EC0 , 32'hFE9F74B4 , 32'h062A4C48 , 32'h09C75B80 , 32'hED12CAA0 , 32'h0951A2D0 , 32'hF6B88180 , 32'h012938F4 , 32'h09D8BC00 , 32'hF93ABC68 , 32'hF76FCE70 , 32'h0BD086F0 , 32'hF8E3F1B0 , 32'hF7394080 , 32'h037C240C , 32'h0013CAFD , 32'h1ABCC520 , 32'hFF906CBB , 32'hFC2C3048 , 32'hFCEE39B8 , 32'hFEED9610 , 32'h0C774A70 , 32'h095AD4F0 , 32'hFD985740 , 32'h03C92264 , 32'h0C7D1FF0 , 32'h03DC287C , 32'hFF25C0E0 , 32'hEDF10320 , 32'h01B7B024 , 32'h0A1ECAD0 , 32'hFFFEC650 , 32'h0346FFB0 , 32'h04EF96D0 , 32'h01574E50 , 32'hFA5951C0 , 32'h06384BD0 , 32'h0132F8F0 , 32'hFFFE26DC , 32'h00011123 , 32'hFFF911C8 , 32'h00033F07 , 32'hFFFF660C , 32'hFFFE1852 , 32'hFFFD39D8 , 32'h0000EA58 , 32'hFFFF1928 , 32'h0001AE43} , 
{32'h0005CB38 , 32'hFFFFB384 , 32'hFFF5987D , 32'h000AC69A , 32'hFFFF9ECF , 32'h000139E9 , 32'hFFF750AF , 32'h0001CB99 , 32'hFFFB0C5A , 32'hFFFE2039 , 32'hFFF7938D , 32'h00038425 , 32'h0001268C , 32'hFFFB5422 , 32'hFFFAD2F6 , 32'h0000C075 , 32'hFFFA1824 , 32'hFFF9CD14 , 32'h0004614C , 32'h0001B483 , 32'hFFFF03D7 , 32'hFFF9BF09 , 32'h000223EE , 32'h00034853 , 32'h0002D008 , 32'hFFFBBCE1 , 32'hFFFF4725 , 32'h00037041 , 32'hFFFFC4A0 , 32'hFFFB5573 , 32'h00010292 , 32'hFFFF0614 , 32'hFFFFEF92 , 32'hFFFA4CA3 , 32'hFFFAC177 , 32'h000259AE , 32'h00018B87 , 32'hFFFDDD48 , 32'h0003D205 , 32'hFFFF4CD2 , 32'hFFFD953C , 32'h0002A66F , 32'h000414F7 , 32'hFFFD9903 , 32'hFFFBEA28 , 32'hFFFC62BE , 32'h00043067 , 32'hFFF8D769 , 32'h0001323A , 32'h00023428 , 32'hFFFF08C6 , 32'hFFFA57E4 , 32'h0008EFE3 , 32'hFFFB7452 , 32'hFFFD4FB6 , 32'h000659B0 , 32'h000561F3 , 32'h000412F6 , 32'h000386C0 , 32'h000101FA , 32'h0000891A , 32'h0002F8E2 , 32'hFFFF2698 , 32'hFFF80C3E , 32'h00087B84 , 32'h00014D4C , 32'hFFFF9D74 , 32'hFFFA4AF2 , 32'hFFFE4079 , 32'hFFFE5DA7 , 32'hFFFD1757 , 32'h000241F3 , 32'hFFFC767B , 32'hFFFFEC0D , 32'h00035B85 , 32'h00087A4F , 32'hFFF55AF7 , 32'hFFFA141D , 32'h0002B7C7 , 32'hFFFFB079 , 32'h00011933 , 32'hFFF67B60 , 32'hFFFD4B5A , 32'h0000F9A9 , 32'hFFFA3F76 , 32'hFFFABC7F , 32'h0000F38C , 32'hFFFA3FC5 , 32'hFFFF5D20 , 32'hFFFBF16D , 32'h0008E405 , 32'hFFFB4678 , 32'hFFF8A2D1 , 32'h0004EC82 , 32'hFFFADDAE , 32'hFFFE4102 , 32'h0005FBD3 , 32'hFFFEDCE0 , 32'h0000BEC9 , 32'hFFF8CC38} , 
{32'hB9319300 , 32'h3549A340 , 32'h1DD608A0 , 32'h571C1600 , 32'hF97AE280 , 32'hC3C16180 , 32'h3E9C3300 , 32'hF6BDA9B0 , 32'hB020A680 , 32'h07D8F5D8 , 32'hF1E6EEA0 , 32'h0206BE60 , 32'h25C07C80 , 32'hE4CF5DE0 , 32'hFD722DE0 , 32'h22F48700 , 32'h02AB8330 , 32'hEB6A3A00 , 32'h07DA3608 , 32'h152C1480 , 32'h2B870980 , 32'h0152A6A4 , 32'h08F48C10 , 32'h0913C170 , 32'hFE9C7BF0 , 32'h143898C0 , 32'h0C0C7880 , 32'hF30D7A00 , 32'hFE3A7360 , 32'hD9DF8E80 , 32'h1DA58E40 , 32'h084859B0 , 32'h112E1FA0 , 32'h02F3BFB0 , 32'hF25BAD30 , 32'h158ED760 , 32'h1061C1A0 , 32'hFCDCF054 , 32'h0A3EC6F0 , 32'hF3AFDEF0 , 32'hFFACA0DF , 32'h04EA8618 , 32'h0A03E0B0 , 32'h0EC48510 , 32'h068F1120 , 32'h071E7B08 , 32'h04854CE0 , 32'hFDA375A0 , 32'h2328B140 , 32'h0B8B55A0 , 32'h0C9BDA80 , 32'hFC605214 , 32'hE7F67660 , 32'hE9B580A0 , 32'hF36B3960 , 32'h0E9CC7B0 , 32'hF9FD8910 , 32'hED6052C0 , 32'hF2CBE5D0 , 32'hFDE90244 , 32'h0282EDF8 , 32'hFBC9B5A8 , 32'h0E4A2D80 , 32'hFB714F80 , 32'hF884D2A8 , 32'hF841C280 , 32'hF742EA20 , 32'hF42F1C90 , 32'h08122B00 , 32'hFECA2124 , 32'h035819BC , 32'h0B487370 , 32'hF8EDB460 , 32'h01B6BC78 , 32'h068F2EC8 , 32'h06335C58 , 32'hFD7B5E44 , 32'h02ABB744 , 32'hF7937FF0 , 32'hFD51D1B4 , 32'hF9D44760 , 32'h02DB2A98 , 32'hFE901EA0 , 32'h01A2A660 , 32'h0492A240 , 32'h033C3C20 , 32'hF66CF940 , 32'h036D64BC , 32'hFFBF9038 , 32'h011E2C58 , 32'hFFFFC506 , 32'hFFFA7B95 , 32'hFFFEBE5F , 32'h0002E4F3 , 32'hFFFDE357 , 32'h00009C07 , 32'h00018291 , 32'h00014CF5 , 32'h0002AD6A , 32'hFFFEB68A} , 
{32'h0833F8B0 , 32'h11B56320 , 32'hE7C871C0 , 32'h07419410 , 32'h08FE2B60 , 32'h33E16E00 , 32'h062747E8 , 32'hFD6B9E3C , 32'hF9039F98 , 32'hF2571130 , 32'h11D61840 , 32'hEFE0EF80 , 32'h0D0297E0 , 32'h08138DA0 , 32'hFBFB8BB8 , 32'h0222C358 , 32'h0C0BEE10 , 32'h0BDEBDF0 , 32'h04109B40 , 32'h16C1D200 , 32'hF162B5D0 , 32'hFE673F90 , 32'h25983EC0 , 32'hEED307C0 , 32'hF35607B0 , 32'hFB289518 , 32'h152AEA00 , 32'h11DAC7A0 , 32'hF2A3AAB0 , 32'hFC5EC1A8 , 32'h11FE19E0 , 32'hF2304030 , 32'h1D0F28E0 , 32'hDB84D840 , 32'hE3A41AE0 , 32'hE019C040 , 32'h007B1569 , 32'hFDBBC574 , 32'h1154D300 , 32'h0D3E4020 , 32'hE52E9FA0 , 32'h1534A3A0 , 32'hF7314000 , 32'hF6FC2420 , 32'h016C900C , 32'hE64207A0 , 32'h1A123640 , 32'h08AF4DF0 , 32'h0EFFAEA0 , 32'h03C8DDAC , 32'hEABE6FE0 , 32'hFF5C0339 , 32'hF7D5AD50 , 32'h050CE140 , 32'hFA4CFDC0 , 32'hFB81C7E8 , 32'hFB737048 , 32'h00E6AAE1 , 32'h05F6CBA0 , 32'h00D51257 , 32'hFADB7B10 , 32'h0E8DCBF0 , 32'h0087B145 , 32'h0274DAE8 , 32'h0DFD7860 , 32'h036F1618 , 32'hFD8C70D4 , 32'h082EF350 , 32'hFA7FD8E0 , 32'hFC204888 , 32'h0CC5DF20 , 32'hF67AD640 , 32'hFA095020 , 32'h051E9590 , 32'hFCB58D18 , 32'hF74FC5B0 , 32'h18784060 , 32'h0218B868 , 32'h06C77460 , 32'h08BB7460 , 32'hFCE3A5EC , 32'h07CA5398 , 32'hFD0AA62C , 32'hF46DBA40 , 32'h00F5F1D4 , 32'h053FD290 , 32'h050447F0 , 32'hFE5B12AC , 32'hFFCAA9F2 , 32'h00946E69 , 32'hFFFDDCBF , 32'hFFFE8B1B , 32'h00028C17 , 32'h00004C45 , 32'hFFF9E026 , 32'hFFFE6E2D , 32'h00002F4C , 32'h0000E327 , 32'hFFFC8C0A , 32'hFFFF4072} , 
{32'hFFFE6A44 , 32'hFFFFF1F2 , 32'h0006F1DC , 32'h00017A7D , 32'h0007225B , 32'h00055734 , 32'hFFFB40F8 , 32'h00025B3D , 32'h00016567 , 32'hFFFDC94A , 32'h0009495A , 32'hFFFF9CCB , 32'h0000CA26 , 32'h0000DE76 , 32'h000902BE , 32'hFFF6DE98 , 32'hFFFD23E7 , 32'hFFFDD491 , 32'h000341ED , 32'hFFFC04EB , 32'hFFFF45A0 , 32'hFFFDA4CD , 32'hFFFA7D76 , 32'h0005E51C , 32'hFFFB040E , 32'h0004EBCE , 32'h00020017 , 32'h0000C6F0 , 32'h0001524D , 32'h00044807 , 32'h0003A90C , 32'hFFFCD946 , 32'hFFFDD3FF , 32'hFFF7FD82 , 32'hFFFFC0D3 , 32'hFFFABD5A , 32'h0002B3C2 , 32'h000279F3 , 32'h0003EAED , 32'hFFFA43AA , 32'h0003F00B , 32'hFFF57381 , 32'hFFFA71DB , 32'hFFFF02E4 , 32'hFFF6A0E3 , 32'hFFF6382C , 32'hFFF9B17D , 32'h0003A468 , 32'hFFF9EFBC , 32'hFFFB3AE2 , 32'h0001DC6F , 32'h00003B2E , 32'h0003D10A , 32'hFFFE36EE , 32'h0002EE66 , 32'h000479EC , 32'hFFFED3C5 , 32'h00031FE8 , 32'h00065984 , 32'h00048702 , 32'h0001829C , 32'hFFFD4CA9 , 32'h00038449 , 32'hFFFE6E43 , 32'h00027300 , 32'h00043674 , 32'hFFFA6171 , 32'hFFF6F1DE , 32'hFFFD6E3A , 32'h0006F24F , 32'hFFFE5674 , 32'h00067EC1 , 32'h00022EB2 , 32'hFFFB1539 , 32'h0007D7A4 , 32'hFFFF81DA , 32'h000697DE , 32'hFFFE5F57 , 32'hFFF7C8B3 , 32'h0003D613 , 32'hFFFECF70 , 32'hFFFE25B7 , 32'h00054584 , 32'hFFFCBABA , 32'h000831A0 , 32'hFFFE1261 , 32'hFFFD61FA , 32'hFFFC7F44 , 32'hFFFCCCC4 , 32'hFFF9C741 , 32'hFFFD47A5 , 32'hFFFC2C91 , 32'h0004F14B , 32'h0002B8D8 , 32'h000127BA , 32'hFFF809C7 , 32'hFFFFADF0 , 32'h0000984B , 32'hFFFF8E6F , 32'h0008007D} , 
{32'h00031ADA , 32'h0002EA68 , 32'hFFF7F849 , 32'hFFF92CC3 , 32'hFFFF38B8 , 32'hFFFF6BC2 , 32'hFFFE0248 , 32'h00009209 , 32'hFFFA5AF6 , 32'h0008B8D8 , 32'hFFFC5B1B , 32'hFFFC06F4 , 32'hFFFA5E03 , 32'h000096BD , 32'hFFFEABBB , 32'hFFF8C482 , 32'hFFFA414E , 32'h0006384E , 32'hFFFC7A88 , 32'hFFFEC9F3 , 32'hFFFFBA5B , 32'h00049979 , 32'h0000B538 , 32'hFFFC38B0 , 32'h0002AEBF , 32'hFFFE657D , 32'h000997A0 , 32'h0003FE28 , 32'h0001F8D7 , 32'hFFFE5EE2 , 32'hFFF9F8EE , 32'h00069B67 , 32'hFFFF1E23 , 32'h0004331A , 32'hFFFEE1F2 , 32'h00007B4A , 32'hFFFFBB0A , 32'hFFFC5B1A , 32'hFFFAE2A6 , 32'hFFFFB063 , 32'h0000F39B , 32'hFFFB47C9 , 32'h00030D65 , 32'h0008815B , 32'h00033A05 , 32'hFFFE6E07 , 32'hFFF973A0 , 32'h00069212 , 32'h000909EA , 32'hFFF84DB2 , 32'hFFFDB5F9 , 32'hFFFE45DC , 32'hFFFED6B7 , 32'h0008B700 , 32'hFFFD5A57 , 32'h000C1CC4 , 32'h0004E0B6 , 32'h00021A55 , 32'h00010298 , 32'h0002108E , 32'hFFFAF047 , 32'h00013FAB , 32'h000F6AF4 , 32'hFFFE7392 , 32'h00003C6B , 32'h000040D3 , 32'h00032F78 , 32'hFFFB9773 , 32'h00051968 , 32'hFFFFD572 , 32'h0008C74F , 32'hFFFEC3B9 , 32'hFFFF792D , 32'h00008F49 , 32'h00057199 , 32'hFFFF3A7B , 32'h00060CBA , 32'h000723E0 , 32'h0000063B , 32'h0002EF9B , 32'hFFFF3C38 , 32'hFFF68356 , 32'hFFFA76CF , 32'h00087B01 , 32'hFFFC94FF , 32'hFFFF6122 , 32'hFFFE2FDB , 32'h000A28BB , 32'hFFF94946 , 32'hFFFD1F57 , 32'h0002EE52 , 32'hFFF7E785 , 32'hFFFD01D3 , 32'hFFFFA8BF , 32'hFFFC94EE , 32'h0000CDB4 , 32'h000121A6 , 32'hFFF9EAFE , 32'hFFFD5C97 , 32'hFFFF6C60} , 
{32'hF9FCDA20 , 32'h012FCABC , 32'h0DB2DA20 , 32'h0C13E710 , 32'hFFA22C99 , 32'hF19CB650 , 32'hF4AAA220 , 32'hFC36FE04 , 32'hFF76B771 , 32'h00EAC183 , 32'h0CC4D830 , 32'hFB7C78C0 , 32'h0CFA0BD0 , 32'h0237AB4C , 32'h0B4A3410 , 32'h01E89500 , 32'h0B6C71E0 , 32'hF74E9310 , 32'h0B951DD0 , 32'h029D5A90 , 32'hF79E8F70 , 32'hF8793B10 , 32'hFB5BE5A8 , 32'hFE0E7F94 , 32'h05FA9670 , 32'h0E59F020 , 32'hFD621020 , 32'hEF1141C0 , 32'hFA94DD98 , 32'hF08D9CA0 , 32'hF6E840B0 , 32'h0E62F600 , 32'h046AE8F8 , 32'h00B900BA , 32'hFF528BC3 , 32'hF3AF0310 , 32'hFF66663D , 32'h02B08BBC , 32'h0029F297 , 32'hF8FB05F8 , 32'hFF00131E , 32'hFF8DCED4 , 32'h02ECB73C , 32'hFC8B21F8 , 32'hFC88AA34 , 32'hF9D46480 , 32'hF51F17C0 , 32'hF14242B0 , 32'hF81AC530 , 32'h03F24924 , 32'hFA878848 , 32'h0351BA38 , 32'h01C0B45C , 32'h059D71F0 , 32'h051CFE48 , 32'h0244650C , 32'hFEE5C538 , 32'hFFE8F54D , 32'h022C39F8 , 32'h0232DBF8 , 32'hFDD432E0 , 32'h084039E0 , 32'h002F0098 , 32'hF8212BC8 , 32'h05986518 , 32'hEF47C600 , 32'hFFB33336 , 32'h0317B328 , 32'hFBBD78B8 , 32'hFD9D0DA8 , 32'h072A2430 , 32'hFC690F24 , 32'hFBFF97E0 , 32'hFCD38264 , 32'h00EAF50A , 32'h0049951F , 32'hFADA4C58 , 32'hFD99B958 , 32'h0227D588 , 32'h03919D2C , 32'h025E3774 , 32'hFF37741F , 32'hFFDEE871 , 32'h0050943F , 32'h00ED2603 , 32'h04DA8D48 , 32'h024A8098 , 32'h02FD5560 , 32'h04B62678 , 32'hFF40D16F , 32'h0003ED87 , 32'hFFFCD551 , 32'hFFFC9579 , 32'hFFFC48AB , 32'h00018F70 , 32'h00008EC1 , 32'h00022011 , 32'hFFFD54C4 , 32'h0006E8EA , 32'h00002E5C} , 
{32'h11E9CCA0 , 32'hF790EE60 , 32'h460F2580 , 32'hEBF852E0 , 32'hDADBB180 , 32'h0EFB93B0 , 32'hF38BD540 , 32'hCECDDB80 , 32'h14A94B80 , 32'hF7DB6900 , 32'hF5A5DE80 , 32'hF85F77D8 , 32'hFC209E8C , 32'hEB1E7980 , 32'h00ACF885 , 32'hED086800 , 32'hEF8BD800 , 32'hF3803380 , 32'h171FB8E0 , 32'h07806680 , 32'hF2D4CD30 , 32'hF9DB2908 , 32'hE9AFD480 , 32'hF7D04030 , 32'hEBB8FD60 , 32'h03BB0ACC , 32'hE8BD64A0 , 32'h040E1780 , 32'hF564CAE0 , 32'hF3953AC0 , 32'hDA5CB840 , 32'h03403668 , 32'h0F1FA4F0 , 32'hEBEA7220 , 32'hFDC0D4A4 , 32'hF4669060 , 32'h1A850D20 , 32'hF5367760 , 32'hF81880B0 , 32'h15292840 , 32'h08C83BA0 , 32'h10BCC680 , 32'hEF5B4040 , 32'hFC158808 , 32'hEB91C4E0 , 32'hEE84A3E0 , 32'hFC38E214 , 32'hFAE8CC68 , 32'h10D1B400 , 32'hFAD58110 , 32'h0D719130 , 32'hF057ED30 , 32'hFBA3C620 , 32'hEF2EADA0 , 32'hEE878B00 , 32'hF24A6500 , 32'hEF82DE80 , 32'hF11976B0 , 32'hF6DD3800 , 32'h0E5B9F40 , 32'hFAB92C70 , 32'hFF3FEFAB , 32'h00631A41 , 32'hFD3048F8 , 32'hED2CFDC0 , 32'h04A479D8 , 32'h0B12C4A0 , 32'h02DE319C , 32'hFF3638D6 , 32'h0A808470 , 32'h04BEBF60 , 32'h0E523260 , 32'hFBC7F338 , 32'hF566B890 , 32'h055ADAE8 , 32'h0900FE20 , 32'hFD1BE384 , 32'h05931DC0 , 32'h0D191750 , 32'h08959550 , 32'h077C99F8 , 32'hFE543ACC , 32'hFC7A5200 , 32'h04BCCE28 , 32'h00E42F4E , 32'h077E5298 , 32'hFD320360 , 32'h019B099C , 32'hFF96CC1F , 32'hFFF8534C , 32'hFFFDC143 , 32'hFFFB2AB5 , 32'hFFFEE858 , 32'hFFFDAE78 , 32'h00015F00 , 32'h00014F33 , 32'hFFFA4171 , 32'hFFFF3726 , 32'h0005D961 , 32'hFFFE79D1} , 
{32'hD07ABA40 , 32'h08E9DD00 , 32'h24A44240 , 32'hCA5A4740 , 32'hE970B120 , 32'hE2E3A780 , 32'h0B456EB0 , 32'hE2EB24C0 , 32'h10E1D460 , 32'hD0192D80 , 32'hF7DDE800 , 32'h23F9D680 , 32'h1847DE80 , 32'hFD302BC0 , 32'hF4212410 , 32'hE33513C0 , 32'hED782000 , 32'hED0E03C0 , 32'hE4C6C8C0 , 32'h25D29700 , 32'hEAE1B7C0 , 32'hEE787F00 , 32'hF8E58680 , 32'hECA0B100 , 32'hEC9448A0 , 32'h279F8E40 , 32'h06288120 , 32'h10CC2940 , 32'hF1B4C520 , 32'hD8310180 , 32'h15D137C0 , 32'h0154BF90 , 32'hDE077C80 , 32'hE687E5A0 , 32'hF7F51580 , 32'h0356775C , 32'hEE28FC20 , 32'h019912D0 , 32'h0068E76A , 32'h08EE3880 , 32'h08990AD0 , 32'h11F37F20 , 32'h08DF8130 , 32'h056338C8 , 32'hFB5003C8 , 32'hFB391598 , 32'h09978970 , 32'h04626E18 , 32'h04DB3380 , 32'h0179F250 , 32'hF88CFEF0 , 32'h03C547D4 , 32'hFC34F5C0 , 32'hF86E6580 , 32'hF6717630 , 32'h0B5FABA0 , 32'h13E6D700 , 32'h01A27738 , 32'h0EFC1470 , 32'hED43E720 , 32'h0E76C9C0 , 32'hFCC49FCC , 32'h0F96BB20 , 32'hE8F7D840 , 32'h09B9F120 , 32'h04F00E28 , 32'hF7CEB950 , 32'h0321E98C , 32'h00EBC733 , 32'hFDC24D10 , 32'h05FC1610 , 32'h0BC4AA50 , 32'h058517C8 , 32'h093BC150 , 32'h01243AC0 , 32'hF47E7950 , 32'hFEE2572C , 32'h027B0688 , 32'hFC5E864C , 32'hFD7A60A4 , 32'hFD615D70 , 32'hFF89EE0E , 32'h0772E3B8 , 32'h03241930 , 32'h013052C8 , 32'hF9A7EE48 , 32'hFFDC6205 , 32'h011E4384 , 32'hFBEEA290 , 32'hFFACB1B5 , 32'hFFFEAA24 , 32'hFFFC8FEB , 32'h0000CB25 , 32'h00026DCD , 32'h00004D2A , 32'h00045702 , 32'hFFF8FB08 , 32'h0001AB74 , 32'h0004F718 , 32'hFFFF4450} , 
{32'hB1A73F80 , 32'h273F09C0 , 32'h3DB22180 , 32'hFCD63CE0 , 32'hFEB6B694 , 32'h14C18520 , 32'h1A0E10A0 , 32'hED481BA0 , 32'hE81A8E20 , 32'h278C77C0 , 32'hDAE2D000 , 32'h0FB078B0 , 32'hFB733AE8 , 32'hFA43FEE0 , 32'hDF037480 , 32'hD28D0B00 , 32'h22737500 , 32'h03B44C28 , 32'h0FC57B20 , 32'hEA1FD1A0 , 32'h00E1FFDD , 32'hE8303040 , 32'h00E9E694 , 32'h024633C0 , 32'h236A9400 , 32'hE64ED6E0 , 32'hFC8B6794 , 32'hEEDCBBC0 , 32'hF9D0F6B8 , 32'hD89DC180 , 32'h0AE40F80 , 32'h16BE8EE0 , 32'hFEF6A5BC , 32'h0981C3F0 , 32'hF1964C20 , 32'h04963018 , 32'hF6A60C70 , 32'hF5947BC0 , 32'hF803FB18 , 32'h14A24560 , 32'h0355CD44 , 32'h09946360 , 32'hEBB91680 , 32'hFAD87898 , 32'hFF3919C5 , 32'hF76A5D40 , 32'hE89B43A0 , 32'h03ECC258 , 32'hE6752880 , 32'hFE621A44 , 32'h0501D430 , 32'hF27FE0F0 , 32'hFE98332C , 32'h13998F40 , 32'h11883380 , 32'h0CD0F710 , 32'h06E52F48 , 32'hE3B75B20 , 32'h0E84EBE0 , 32'hFF10A7E2 , 32'hFE48A9A4 , 32'hF12707E0 , 32'h1579A7C0 , 32'hEBD03F00 , 32'h17C0E360 , 32'h04148610 , 32'h06B85488 , 32'hFD18A604 , 32'hFDABEED8 , 32'hFAADB598 , 32'hFCE63420 , 32'h007DC9FE , 32'h0B2BBA30 , 32'hF1B71CE0 , 32'hF4B68CB0 , 32'h0DE471E0 , 32'h003026C7 , 32'hFF8383A9 , 32'hFFB8D974 , 32'hF75BAB70 , 32'h00F9AFBB , 32'h049EF5A0 , 32'h022FCF20 , 32'hF725D440 , 32'h0389CA44 , 32'hFF08BB46 , 32'h01480E8C , 32'hFDC50578 , 32'hFD099D74 , 32'hFF262372 , 32'h00028C69 , 32'h0003000B , 32'hFFFBE9FE , 32'h00017CDE , 32'hFFFD6CF7 , 32'hFFFBE7E1 , 32'h00010C59 , 32'h000095DB , 32'hFFFECE9E , 32'h00025C9F} , 
{32'h0001FB00 , 32'hFFFBFD89 , 32'h00054AC2 , 32'hFFFC5C36 , 32'h00031A1C , 32'h000B0749 , 32'hFFF766E5 , 32'h00020110 , 32'h0005FE08 , 32'h00006C9C , 32'hFFF6010C , 32'hFFFF050E , 32'hFFFE076A , 32'h000A4A8F , 32'h0005DE1E , 32'hFFFE25F1 , 32'h00058FBA , 32'hFFFE90E7 , 32'h0004739A , 32'h00039437 , 32'h0003C502 , 32'h00005406 , 32'h00024392 , 32'h00013617 , 32'hFFF78EB5 , 32'h00016CCB , 32'hFFFB67F9 , 32'h000B9716 , 32'hFFFCAFF8 , 32'h000281E7 , 32'hFFFC7272 , 32'h0003F408 , 32'h0005744A , 32'hFFFD065B , 32'h0002B03E , 32'h0003F1A9 , 32'hFFFEB0B1 , 32'hFFFFA7A5 , 32'hFFF8E186 , 32'h0001C54A , 32'hFFFDA93D , 32'h00040134 , 32'h00040656 , 32'h00056550 , 32'hFFFE6FDA , 32'h0007BF94 , 32'hFFF7241D , 32'h00047C25 , 32'hFFFC9A06 , 32'hFFFEA257 , 32'h00018C65 , 32'hFFFF8B14 , 32'hFFFDC02E , 32'h0003C07E , 32'hFFFC0149 , 32'h0001B899 , 32'hFFFFE916 , 32'h00020080 , 32'h000898EB , 32'h00096F2C , 32'h0005DF9C , 32'h000340C6 , 32'h0006BA6E , 32'hFFF7C58F , 32'h0001B2B0 , 32'hFFFBD70D , 32'hFFFD2C33 , 32'h00061F92 , 32'h0003BD85 , 32'h0009D29E , 32'hFFFD37D6 , 32'h0000D61E , 32'h0000111D , 32'hFFFDB3A1 , 32'h0002CA0B , 32'h00013FC6 , 32'hFFFDA972 , 32'h000501F7 , 32'h0003B19B , 32'h00089A08 , 32'h0000488E , 32'h0002B701 , 32'h00043271 , 32'hFFFA56D3 , 32'h000AAD94 , 32'h0002CB77 , 32'hFFFED6D0 , 32'hFFF8984D , 32'h000063A5 , 32'hFFFEAB4F , 32'hFFF8561F , 32'h00049A06 , 32'hFFFA923D , 32'hFFFA7709 , 32'h00043478 , 32'hFFFFDF10 , 32'h000400A7 , 32'h00009BFF , 32'hFFF8BB1A , 32'h000072BA} , 
{32'h000EEF35 , 32'hFFB7D63C , 32'h016C93F4 , 32'hFC316890 , 32'hE9DD16A0 , 32'h03B594DC , 32'h057054B8 , 32'hFFAC6BB0 , 32'h084DDCD0 , 32'h0EBCBC60 , 32'h02483CA0 , 32'h052DAC78 , 32'hF71FF500 , 32'h0D657B70 , 32'h072B7E48 , 32'hF6B6EB10 , 32'h0C780E20 , 32'hFDBCE88C , 32'hFEF90208 , 32'h0515C218 , 32'h019C6BE4 , 32'h0F292DD0 , 32'h0A0A7330 , 32'hF28EF000 , 32'h00BBC9AA , 32'h1771AD40 , 32'hEF294380 , 32'hF6A67690 , 32'h0E5BC7A0 , 32'hFE523A4C , 32'h01AA1080 , 32'hFB4FC910 , 32'h0BF27DB0 , 32'hF4750830 , 32'h0A4F5F00 , 32'hFC5F5440 , 32'hF1A972B0 , 32'hF723AAD0 , 32'h118E3BE0 , 32'hFE0BFFF4 , 32'h02342140 , 32'hFA8150D8 , 32'h0ECF19B0 , 32'hEAE3E380 , 32'h0C72C0B0 , 32'hFF0680C8 , 32'hFC112980 , 32'hF02ABC00 , 32'hF78DCF40 , 32'hF50F9CA0 , 32'h013E1FC8 , 32'hFE1F367C , 32'hFFB7CFFB , 32'hF76F19C0 , 32'hFB118CA8 , 32'hFEC4080C , 32'h07C25BE8 , 32'h0A4886A0 , 32'h045141F8 , 32'h03FE4BDC , 32'h00A03320 , 32'hFA6174B8 , 32'hF8C662A0 , 32'hF8C88D30 , 32'h05AAA160 , 32'hFC1427CC , 32'hF7C88950 , 32'hF7AAD760 , 32'h0103A85C , 32'h04483F88 , 32'h0B753890 , 32'h026FEB3C , 32'h077DF470 , 32'hFD0C6154 , 32'hFFB3370A , 32'hFB79D578 , 32'h007F69B5 , 32'hFF501F5B , 32'h082362A0 , 32'hF7893A20 , 32'hFB262AD0 , 32'hFE8A4994 , 32'hFD954D54 , 32'hFE0F5B70 , 32'h031AA094 , 32'hF79C02A0 , 32'hFBBBC3D0 , 32'hFBC29C10 , 32'hFB6B11E8 , 32'hFFB186ED , 32'h0000A4E2 , 32'hFFFE0967 , 32'hFFFA4490 , 32'hFFFCEDB2 , 32'hFFFE5C5F , 32'hFFFE6ED0 , 32'hFFFC12CA , 32'hFFFE7681 , 32'h00017DFB , 32'h00007913} , 
{32'hF27836E0 , 32'h0D96C850 , 32'h01514218 , 32'h0AF5D9D0 , 32'h04114CD0 , 32'h0332691C , 32'hF9307D48 , 32'h00083815 , 32'h0C68BAF0 , 32'hEE69DFA0 , 32'hFEE9EEAC , 32'h01ED1CD8 , 32'h038911D0 , 32'h15DD1F40 , 32'h035491EC , 32'hEFAEDDA0 , 32'hFBB03C00 , 32'hF7D6E020 , 32'h0F42FE00 , 32'hFB1211D0 , 32'h13D67620 , 32'hFFB6DF27 , 32'h03F83150 , 32'hF99CA3D8 , 32'hFFC8EE79 , 32'hFB6BA7E8 , 32'h03496F20 , 32'h00DE9CF3 , 32'h08891F30 , 32'hF91EC960 , 32'h0145B238 , 32'hFC51F62C , 32'h05F6F080 , 32'h0615C6B0 , 32'hFC1C93C8 , 32'hFEA06EE8 , 32'hFF8ACC4E , 32'h0256E520 , 32'hFE8464AC , 32'h02F777D0 , 32'h01893E8C , 32'h07DDFEF0 , 32'h02066648 , 32'hFD95A504 , 32'h09AB2390 , 32'hFC7A1C78 , 32'hFB4AFD68 , 32'hFF567B0C , 32'h01D9C6A4 , 32'hF5D8B4E0 , 32'h01828254 , 32'hF775FC50 , 32'hFC85A3AC , 32'h01ACE41C , 32'h08AD2AB0 , 32'hFC97D788 , 32'hFAA62680 , 32'hF47A3370 , 32'h030AC7F0 , 32'hF7F18930 , 32'h0A1ABCC0 , 32'h01424BA8 , 32'hFFCC1A03 , 32'hFF31701E , 32'hF94CD6E0 , 32'h0618EB00 , 32'hFBDBBD68 , 32'hFEAD6B50 , 32'hF8EC8420 , 32'h093F92F0 , 32'h07F04600 , 32'h04ECEFE0 , 32'hFDA6CBF0 , 32'h03D09DC8 , 32'h0178D294 , 32'h07D2EF48 , 32'h02202B34 , 32'h016002EC , 32'hFF6BD87D , 32'hF6E5CD80 , 32'h00A35037 , 32'h050AD8D0 , 32'hFD12C9FC , 32'h023D0644 , 32'h02E1CE68 , 32'h011FD434 , 32'hFABBCEA0 , 32'hFC2490C4 , 32'h0021828F , 32'h0079AA41 , 32'h0002F1AA , 32'hFFF9BF87 , 32'hFFFDF17F , 32'hFFFFA909 , 32'h00077E56 , 32'h0002B425 , 32'h0004662A , 32'hFFFA9F51 , 32'hFFFE261C , 32'h0001DCF8} , 
{32'hFFFF6204 , 32'hFFF9B925 , 32'hFFFFEE9A , 32'hFFFA39FA , 32'hFFFD7188 , 32'hFFF8E09E , 32'hFFFCFE0F , 32'h000482CD , 32'hFFF99673 , 32'hFFFFBD87 , 32'hFFFBF264 , 32'hFFFF0EF8 , 32'hFFFE10E5 , 32'h00078B05 , 32'hFFF9883A , 32'h0002C015 , 32'hFFFB967E , 32'hFFFDE33D , 32'hFFFF4383 , 32'hFFFD562A , 32'hFFF70DEA , 32'h00002192 , 32'hFFFA9575 , 32'h00016C68 , 32'h0006B6A7 , 32'h0009A3AC , 32'h00040C31 , 32'hFFFEF84C , 32'hFFFD9321 , 32'h000140C7 , 32'h00065B9D , 32'hFFF95576 , 32'hFFF5DB6A , 32'h00009B40 , 32'hFFFF65FE , 32'h00022A54 , 32'hFFFE2A2C , 32'hFFFF12B1 , 32'h0006D529 , 32'h0001930A , 32'h00025018 , 32'h0004A0EE , 32'hFFFDD131 , 32'hFFFCF62B , 32'hFFF6BEAE , 32'hFFFE7643 , 32'hFFFFC3B0 , 32'hFFFA15C5 , 32'hFFF0D2B3 , 32'hFFF8B68E , 32'hFFFFD92A , 32'h0004E5EB , 32'h00010EDC , 32'hFFFE556B , 32'hFFFE9139 , 32'hFFFCC4F6 , 32'h00089071 , 32'h0003BDFA , 32'h00053DCE , 32'h00020017 , 32'h0001329B , 32'hFFFCC520 , 32'hFFFFDE70 , 32'h00036E8B , 32'hFFFBF59D , 32'h00066B59 , 32'hFFFD3023 , 32'h0002BDE2 , 32'h0000EF1F , 32'hFFFE6E15 , 32'hFFFE07B7 , 32'h0003EC98 , 32'hFFF95327 , 32'h0002E8D9 , 32'h00005801 , 32'hFFFF8BD8 , 32'hFFFAAFE7 , 32'hFFFDAF13 , 32'hFFFF400A , 32'h0003A28F , 32'h00021C3D , 32'h00023FD2 , 32'h00008C43 , 32'h000367EB , 32'h00069E4D , 32'hFFF85C68 , 32'h00008DB9 , 32'hFFF88231 , 32'h0003B607 , 32'hFFFFE6DE , 32'h0003AD15 , 32'hFFFB9061 , 32'h00070713 , 32'h00005CBF , 32'h0004721D , 32'hFFF8A287 , 32'h0002C86F , 32'hFFF69812 , 32'hFFFFFD22 , 32'hFFF941F1} , 
{32'hC3D4C3C0 , 32'hEA658440 , 32'h5B36E980 , 32'hBFEB2380 , 32'h1C02F1C0 , 32'h2267E640 , 32'hB9E55280 , 32'hB95F8200 , 32'hDDA24A80 , 32'h0452ADF8 , 32'h11F21680 , 32'h30F8ACC0 , 32'hF474DE50 , 32'hDD9856C0 , 32'hF812E3A8 , 32'h1202FC80 , 32'h3A942000 , 32'h06DA4D98 , 32'h093645D0 , 32'hB919AC80 , 32'h2FC7FF40 , 32'hF4717F20 , 32'hC1284C80 , 32'hEACF1700 , 32'h071DA2D0 , 32'hFC2A55F8 , 32'h04030DB0 , 32'hF8DA3E78 , 32'hE4184620 , 32'h101CB400 , 32'hFC291CDC , 32'h00A98ED9 , 32'h1A1BDEE0 , 32'hE27BE7C0 , 32'hEC6F0500 , 32'h20312340 , 32'h03E5CF04 , 32'h28F77240 , 32'h1F721200 , 32'h0D10EAF0 , 32'hEB89BE80 , 32'h02ECAFF8 , 32'hF424E790 , 32'h15D1B400 , 32'h082D1390 , 32'h01FC9DAC , 32'h139000C0 , 32'hF08A2170 , 32'h0C978E50 , 32'h15CAF440 , 32'hF34BBCB0 , 32'hF986CA30 , 32'hF7163690 , 32'h05551560 , 32'hFBE794F0 , 32'h0273880C , 32'h2002DE80 , 32'h01BDF818 , 32'hF82D08F8 , 32'h0006DE3B , 32'hE93E7C40 , 32'h07F581A0 , 32'h060C4420 , 32'h06608150 , 32'hF7BD1B10 , 32'h0AAB0CC0 , 32'h10D8AA00 , 32'hFD57A078 , 32'h041580C8 , 32'hFC06E03C , 32'h07006BF0 , 32'h01DE910C , 32'hFC645078 , 32'hF6B8C240 , 32'hF9FAA860 , 32'h03075104 , 32'hFFD6706E , 32'h036234B0 , 32'h04FA5A48 , 32'hFD6DE114 , 32'hFD995C7C , 32'hFD91606C , 32'h035B1FFC , 32'hFFC804CB , 32'hF8985F60 , 32'hFFF6BDD4 , 32'hFB859820 , 32'h00961DB0 , 32'h00DDE342 , 32'h001D9005 , 32'hFFFF85B3 , 32'h000271E6 , 32'h0000DEF5 , 32'hFFFA3B43 , 32'hFFFB7742 , 32'hFFFF36F3 , 32'h0001EE9D , 32'hFFFF02D5 , 32'hFFFFFA77 , 32'h00010071} , 
{32'hFFFA0A94 , 32'h0008594D , 32'hFFFD1D57 , 32'hFFFEBF21 , 32'hFFFF55CE , 32'hFFFCBB4B , 32'hFFFB8DDB , 32'h00088E7B , 32'h000337A0 , 32'h000E18DC , 32'h00044C11 , 32'h0001781A , 32'h0003D0DA , 32'hFFFF1958 , 32'hFFFE4590 , 32'hFFFC79C6 , 32'h000178BA , 32'hFFFC4DCD , 32'h0001E2FA , 32'hFFFF6D77 , 32'hFFFFDF42 , 32'hFFFD038D , 32'hFFF74AAC , 32'h0007B6DD , 32'h00022B32 , 32'hFFFCC8E5 , 32'hFFF7D018 , 32'h0000E8E4 , 32'h00003BE6 , 32'hFFFD8BCD , 32'h00039080 , 32'hFFFC941E , 32'h00015CD7 , 32'hFFFEB540 , 32'h00056872 , 32'h000E2C5A , 32'hFFFCBB1B , 32'hFFFBB52D , 32'h000559E4 , 32'hFFF69B3C , 32'hFFFCBC9D , 32'h000A0343 , 32'hFFFC7A83 , 32'hFFFE2132 , 32'h0004A041 , 32'hFFFCA210 , 32'hFFFA9041 , 32'h00003B76 , 32'hFFF9A022 , 32'hFFF6D0E2 , 32'hFFFB2238 , 32'h000985AD , 32'hFFFF8F34 , 32'h0004D369 , 32'hFFF9D3BC , 32'h0004E6B5 , 32'hFFFD8363 , 32'hFFFA21A1 , 32'hFFFDBB72 , 32'hFFFEE3E0 , 32'hFFFD81E4 , 32'h000233A9 , 32'h000216F1 , 32'hFFFCFBE5 , 32'h00005BAE , 32'hFFFE029C , 32'h00087D46 , 32'hFFFE06C6 , 32'hFFFB7C82 , 32'h0000AB77 , 32'h00035E30 , 32'hFFFFE48D , 32'h00022889 , 32'h000B3E01 , 32'hFFFDCC35 , 32'h00095E26 , 32'h0005123F , 32'hFFFB6E1C , 32'h0002F7DC , 32'h00009210 , 32'h00021CB0 , 32'hFFFCE7B4 , 32'h00065AA8 , 32'hFFF744F8 , 32'h000077AD , 32'h00027B09 , 32'hFFFE02A8 , 32'h00013F46 , 32'hFFFED210 , 32'h00005819 , 32'h00041F91 , 32'h0002EDF7 , 32'h00040479 , 32'h000471A3 , 32'hFFF82E22 , 32'hFFF642FB , 32'h00001AAF , 32'h00060615 , 32'h0006428C , 32'h0000021E} , 
{32'h18541C60 , 32'h3D842B00 , 32'hF3815570 , 32'h06241DE0 , 32'h043BDDE8 , 32'h21E7DE40 , 32'hE8990E80 , 32'hFABC4428 , 32'h16A7BE60 , 32'hF87916B0 , 32'hFD7B1C60 , 32'hE922CCA0 , 32'hF10501F0 , 32'hE4AFCEC0 , 32'hED469420 , 32'h2844CF40 , 32'h0334CC40 , 32'hFDBDF4E4 , 32'h17666A80 , 32'h302A9C00 , 32'h1262A460 , 32'hFED15AE0 , 32'hEECE01E0 , 32'hF564B0E0 , 32'h127C3DC0 , 32'h08619450 , 32'h1259BCC0 , 32'hF2E9C1B0 , 32'hFCB26AA4 , 32'h0479E1C0 , 32'hFE112D20 , 32'hFF22365E , 32'h050E49D0 , 32'hE44BE2A0 , 32'h134076E0 , 32'hFDE55B24 , 32'h0B656230 , 32'h0A002DE0 , 32'hF0D43BA0 , 32'hEA15B8A0 , 32'hFD5CB070 , 32'hF2765770 , 32'h05F984D0 , 32'h03AB9BC0 , 32'h02E3DEEC , 32'hFDD33E20 , 32'hFB00ECE8 , 32'hFB520200 , 32'h0B98FC70 , 32'hFB5F3C70 , 32'h10619DC0 , 32'h16F20D80 , 32'h0211FFAC , 32'hF79ECDF0 , 32'h09A69AB0 , 32'h054CE3B8 , 32'h0B9D97E0 , 32'h013FEC94 , 32'h0006771D , 32'hFB2CB478 , 32'hF3438D10 , 32'hE93BCB60 , 32'h04AB9CE0 , 32'hFCE266A4 , 32'hF2B5BDE0 , 32'hFCABFED0 , 32'hFE79C80C , 32'h00D46692 , 32'hFD017E8C , 32'h04AD44B8 , 32'h0DC16520 , 32'hF767F5E0 , 32'h062E7170 , 32'h046783F8 , 32'hF6CB84D0 , 32'h01B9E838 , 32'h0A8A1F90 , 32'h0182349C , 32'h0185CAAC , 32'hFA457600 , 32'h035F5564 , 32'h05A59A28 , 32'hFD4C7500 , 32'h0096A51C , 32'h01BDDF20 , 32'hFA2751C0 , 32'h002C80BD , 32'hFF8CD0A1 , 32'h0344101C , 32'h0050AD9F , 32'hFFFCDCB9 , 32'h0000198C , 32'h00016993 , 32'h0005B266 , 32'h0005DC76 , 32'hFFFD7736 , 32'h000261B3 , 32'h000AF03F , 32'h0003B886 , 32'hFFFDD8A0} , 
{32'hFFFF904B , 32'hFFFF7617 , 32'h0004E783 , 32'h00022EEC , 32'hFFFD5AD3 , 32'h0003979D , 32'hFFFE0EF1 , 32'h00006151 , 32'hFFFB3E98 , 32'hFFF6ACC3 , 32'h000162AA , 32'hFFFB14B9 , 32'hFFFD38AD , 32'h000693FB , 32'hFFFF1BB3 , 32'h00061DD9 , 32'h0001A0D0 , 32'hFFFCB50C , 32'h0004FB8D , 32'h00036934 , 32'h00034AAD , 32'hFFF98892 , 32'hFFFE48AC , 32'h00019A62 , 32'h0001AE88 , 32'h00009D32 , 32'h000047B9 , 32'hFFFDF9FA , 32'hFFFED7ED , 32'h0002B922 , 32'hFFFA1DFF , 32'hFFFA672E , 32'hFFF96007 , 32'hFFFB36C6 , 32'hFFFB5964 , 32'hFFF7E84B , 32'hFFFEE29E , 32'hFFFD804B , 32'hFFFFBE6C , 32'hFFFABE97 , 32'hFFFF3033 , 32'hFFFFC2B0 , 32'hFFF5F66B , 32'hFFFED36D , 32'hFFFDDEB7 , 32'hFFFBD31D , 32'hFFF9DACF , 32'h0003A8F8 , 32'h000658D1 , 32'hFFFB2056 , 32'hFFFD43E2 , 32'hFFFF6B77 , 32'h00054D44 , 32'hFFFB2192 , 32'hFFF87B2D , 32'h000511EB , 32'hFFFEA6C2 , 32'h00032BD3 , 32'hFFFF4118 , 32'h00095C13 , 32'h00016FF4 , 32'hFFFE6EA9 , 32'h000721F8 , 32'h00021598 , 32'h0003DF3D , 32'h0001DA06 , 32'hFFFB38F1 , 32'hFFFCF6EF , 32'hFFFD5E1D , 32'h000C11AB , 32'h000B56C9 , 32'hFFFEA179 , 32'hFFF958A3 , 32'h000150CE , 32'hFFFA59C4 , 32'hFFFBA032 , 32'h00034A47 , 32'hFFFD02DA , 32'h0003BA5E , 32'h00054012 , 32'h0006CC87 , 32'hFFFD348F , 32'hFFFE98BB , 32'hFFF9C8E5 , 32'hFFFBECE6 , 32'hFFFE8370 , 32'h0001533B , 32'hFFFB76C2 , 32'hFFFD8341 , 32'h000548E5 , 32'h0007DBFB , 32'hFFFEAD44 , 32'h0009E799 , 32'h000C5B02 , 32'hFFFEAA0B , 32'hFFFD1FF5 , 32'h00014BE3 , 32'hFFFCF49C , 32'hFFFD05E1 , 32'h000070F3} , 
{32'hFFFEC1F1 , 32'hFFF6C3D3 , 32'h00029A78 , 32'h00027FFD , 32'h00033A0D , 32'hFFFBB632 , 32'h00062864 , 32'h0002DA1A , 32'hFFFDBA7C , 32'hFFFC322A , 32'hFFFE16C6 , 32'hFFFFD5CF , 32'hFFFE5C3B , 32'h0004092B , 32'hFFFC544D , 32'h00059701 , 32'h00015C64 , 32'hFFFBC430 , 32'h00090264 , 32'hFFFAE628 , 32'h000318D5 , 32'hFFFF64DF , 32'h0005D25A , 32'hFFFE323A , 32'hFFFF075D , 32'hFFFA9674 , 32'h0000C203 , 32'hFFFE55C9 , 32'h0006E7C4 , 32'h0000D721 , 32'hFFF9C408 , 32'hFFFF01CB , 32'h0003601D , 32'h0006D774 , 32'h0005F67E , 32'hFFFF3E79 , 32'h0000D05A , 32'hFFF75487 , 32'hFFFE7B1E , 32'h0003847D , 32'h0001D480 , 32'h0003C578 , 32'h00019743 , 32'h0002C34D , 32'hFFFF5EF0 , 32'h00047186 , 32'h000072BC , 32'h00052324 , 32'h00010B4F , 32'hFFFB1902 , 32'hFFFCA0E7 , 32'h000006BE , 32'hFFFFB64F , 32'hFFF82D69 , 32'h0007993F , 32'h00047A8D , 32'h00017EE3 , 32'h00074507 , 32'h0002F471 , 32'hFFF8B4AD , 32'hFFF9E740 , 32'h00040AF7 , 32'hFFFCD8A4 , 32'hFFFF0677 , 32'h0001A324 , 32'hFFFF7D51 , 32'h0006F12D , 32'hFFFCA7B7 , 32'hFFF6BCE1 , 32'hFFFF2ADC , 32'hFFFDEB27 , 32'hFFFB4A57 , 32'hFFF95364 , 32'h000617C3 , 32'hFFFB40AA , 32'h00007FBB , 32'hFFFD5A57 , 32'h0000E80D , 32'h00013997 , 32'hFFFA2804 , 32'h0007EB9F , 32'h0002FA0E , 32'h0007751B , 32'h000197BC , 32'h00016281 , 32'h00049274 , 32'hFFFC1417 , 32'h000556E3 , 32'hFFFFA900 , 32'hFFFC5C97 , 32'hFFF0A28E , 32'hFFF8F12E , 32'hFFFAB8E7 , 32'h0001BC98 , 32'hFFFF94F0 , 32'h000440BF , 32'h0006C778 , 32'h0005B5B0 , 32'h0003C9A4 , 32'h00067BFD} , 
{32'hFFFF94AD , 32'hFFFEA081 , 32'hFFF82D27 , 32'h0001D6B0 , 32'hFFF11686 , 32'hFFFE7224 , 32'h0001CA13 , 32'h00025539 , 32'h0000CCBA , 32'h0009A8B8 , 32'hFFF58FD0 , 32'h00036788 , 32'hFFF70DB1 , 32'h00027A1C , 32'h0005DEF0 , 32'hFFFC487C , 32'h000AE4D3 , 32'h0006A062 , 32'h000DB70A , 32'h0008B780 , 32'hFFFC0002 , 32'hFFFD2A3B , 32'h00037C40 , 32'hFFFDCE46 , 32'h0008A069 , 32'hFFFDB9CA , 32'hFFFEFE12 , 32'hFFFACDAC , 32'h000A84F3 , 32'hFFFF554A , 32'hFFFE565C , 32'h00004A01 , 32'h000331D6 , 32'h0002B8AB , 32'hFFFFE92F , 32'hFFFCA6BB , 32'hFFF721D1 , 32'hFFF9E5FB , 32'h0006856C , 32'h000465D9 , 32'hFFFE7BE9 , 32'hFFFDCF61 , 32'hFFFF534F , 32'hFFF9C7A0 , 32'hFFF7FF60 , 32'hFFFBEDF0 , 32'h00073656 , 32'hFFFE75A4 , 32'hFFFE42C5 , 32'h0000E8E9 , 32'h0005A6F7 , 32'hFFFFCAE2 , 32'h00039A60 , 32'h0002B1A2 , 32'h00009134 , 32'hFFFEC187 , 32'hFFFDD350 , 32'hFFFFCBE8 , 32'hFFFEC79A , 32'h0002205C , 32'hFFFFE0E3 , 32'hFFFE9523 , 32'hFFF05D18 , 32'h00079D9F , 32'hFFF9F4DC , 32'hFFFFAA48 , 32'hFFF1E74A , 32'hFFFC6C46 , 32'hFFF4E239 , 32'h00013588 , 32'h0001910E , 32'h0001AD43 , 32'hFFF566D5 , 32'hFFFD7374 , 32'hFFFC66A6 , 32'hFFF5E640 , 32'hFFF7CFA0 , 32'h0003B781 , 32'h0004A323 , 32'h00099ACE , 32'h00012FDA , 32'h00055F9C , 32'h0000752F , 32'h000BB88A , 32'h0005D53D , 32'hFFFE325E , 32'h0001C82E , 32'hFFFF575D , 32'h00030567 , 32'h00072FC3 , 32'hFFF9985D , 32'h0000F6E2 , 32'hFFFBE8FA , 32'h00011E40 , 32'hFFFE40A9 , 32'h0002667E , 32'h0008235B , 32'h00008443 , 32'hFFFF3335 , 32'h0003D536} , 
{32'hAA089C00 , 32'hCA72A500 , 32'h86130180 , 32'h2947B440 , 32'h5AAD9980 , 32'hBEEC2200 , 32'hFA55A320 , 32'h06E0F518 , 32'hFB100FA8 , 32'hC4925C40 , 32'h0A70D220 , 32'hDB524E40 , 32'h1FD47E40 , 32'h0A8008A0 , 32'hC96BD600 , 32'h0FCACD80 , 32'hD95634C0 , 32'hD4F06C40 , 32'hF518D330 , 32'h1C52A000 , 32'h27F68D80 , 32'hF163C7B0 , 32'hE3245320 , 32'h0B1D2890 , 32'h06026F88 , 32'h21B59840 , 32'hC764A880 , 32'h03BD60E4 , 32'hFA201440 , 32'h1BE95FC0 , 32'hF90AB7E0 , 32'hF34354E0 , 32'hFB4623F0 , 32'h25099800 , 32'hEBB4B3A0 , 32'hE80BFA20 , 32'hE98A2D00 , 32'h130C2AE0 , 32'hFF7F4F6D , 32'h069E6B88 , 32'hE459CDC0 , 32'h1890AB00 , 32'hE301BD60 , 32'hFE24E168 , 32'h0681CF90 , 32'hF50E2520 , 32'hFB6512F8 , 32'h1AD7F580 , 32'h0CF08CA0 , 32'h0B3BCAD0 , 32'h05726830 , 32'hF2EADD80 , 32'hEDA1A360 , 32'hF24CDF90 , 32'hFB4A6B50 , 32'h101C77C0 , 32'hFBC5FA00 , 32'hF36A62C0 , 32'h07F4EB88 , 32'h08E8E240 , 32'h038956CC , 32'hF0119560 , 32'hF9CA1E28 , 32'h09D7A9A0 , 32'h10DE5C40 , 32'hFAFD8B78 , 32'h07B10FF8 , 32'hEFA28940 , 32'h05BBD940 , 32'h10001580 , 32'h0A67A750 , 32'h01680B94 , 32'hFDD44754 , 32'hFBE67528 , 32'hFF58EDDE , 32'h01D550A4 , 32'hF2AFE0C0 , 32'hFDFF12C8 , 32'hFDE9D3F0 , 32'h0965E890 , 32'h01A00150 , 32'hFAF0C748 , 32'h02DDC548 , 32'hFB8E1728 , 32'h056ADC00 , 32'hFE225C9C , 32'hFD803A6C , 32'hFFB05299 , 32'h0218C874 , 32'hFFB5E188 , 32'hFFFF3C71 , 32'h0000B8FE , 32'h00033C1D , 32'hFFFE31CD , 32'hFFFFACE5 , 32'h00000B84 , 32'hFFFF3E55 , 32'hFFFF297C , 32'hFFFE0429 , 32'h00026ADC} , 
{32'h18D32BC0 , 32'h22B13300 , 32'h4884FD00 , 32'hB636A480 , 32'h5795FA00 , 32'hDFA0EE00 , 32'hD4964000 , 32'h02CEE7F0 , 32'h459A5E80 , 32'hFC96E850 , 32'hC9A70F40 , 32'h096D0030 , 32'h051316A8 , 32'h22A85900 , 32'h05722990 , 32'hF893D1C0 , 32'hF2E3A070 , 32'h1B24CFA0 , 32'hE9214200 , 32'hE5BA3200 , 32'hF6E110A0 , 32'h1034C2C0 , 32'hDFA58EC0 , 32'h181B30C0 , 32'h061FCCF0 , 32'h0F6E98B0 , 32'hD4B12700 , 32'h1C3EC900 , 32'h290C7500 , 32'hCF8E2C00 , 32'hFBE618E0 , 32'hE0603140 , 32'hEC732000 , 32'h10ADD460 , 32'hF4621190 , 32'h1260F540 , 32'hFA8DFAB8 , 32'h18F00840 , 32'hFD91FB28 , 32'h144879C0 , 32'hF6023180 , 32'h031E0FAC , 32'h09080FD0 , 32'hF56E8100 , 32'hF5E09190 , 32'hF0EFA010 , 32'hEF6A0040 , 32'hF8E158C8 , 32'hF4CBFA60 , 32'hED39D8E0 , 32'hFB5A9118 , 32'hF6A33340 , 32'hEF8D3CA0 , 32'h0AA4ADF0 , 32'hE39D85C0 , 32'h06B59D28 , 32'h028A4E80 , 32'h05390DF0 , 32'hF5B3B5D0 , 32'hFC5E5130 , 32'h0204E59C , 32'h0B988520 , 32'hFD0C22CC , 32'h0C300A10 , 32'h01BE2D00 , 32'hE58D0680 , 32'hF68F8CB0 , 32'h039D0FB4 , 32'hF84F3338 , 32'h006CA8B1 , 32'hF6BDFBD0 , 32'hFE356928 , 32'hFEFCF7B4 , 32'h0339D46C , 32'hF6C1AB60 , 32'hF7B76430 , 32'h0274A2BC , 32'h018ED244 , 32'h023F72B0 , 32'hFC158D6C , 32'hFDF20D08 , 32'h011CED6C , 32'hFC602F2C , 32'h03175C98 , 32'hFB60D780 , 32'h01BDD308 , 32'h0212E44C , 32'hFD074DF4 , 32'h00A48E27 , 32'h00F754B6 , 32'hFFFF20EC , 32'h00022F56 , 32'h00022C42 , 32'hFFFF933B , 32'h00001B4B , 32'h0003FE5C , 32'h00029C7A , 32'hFFFD4188 , 32'h0000DEBE , 32'hFFFC141E} , 
{32'h1F92D760 , 32'hCAF94580 , 32'hB0CCD080 , 32'h3FFCEB00 , 32'h17423AC0 , 32'hA8F72D80 , 32'hDF2B7640 , 32'h2D882880 , 32'hEEAB9280 , 32'h1B3CA4A0 , 32'hC9FB0300 , 32'h2CF6C3C0 , 32'h10560CE0 , 32'h358E0F80 , 32'hE780E880 , 32'h12E1EA00 , 32'hFE8C9214 , 32'hFE52DD44 , 32'hDCC03E80 , 32'h01DE3CEC , 32'h39993180 , 32'hF7BB3720 , 32'hF918CAE0 , 32'h0EE42600 , 32'h0ECD3050 , 32'h0E940970 , 32'hF779DCA0 , 32'h06BD1D98 , 32'hF8CB3300 , 32'h12721460 , 32'hDB03F740 , 32'h07F90288 , 32'hEF634800 , 32'hC6AEF380 , 32'h11BB4D20 , 32'hF2F45440 , 32'h20789900 , 32'hF8C881C0 , 32'hF940C1E8 , 32'h0FCBDA40 , 32'h06339858 , 32'h040094E8 , 32'hEDC5AFC0 , 32'hFC805AB0 , 32'h052D3DC0 , 32'h0BC0FAC0 , 32'hFCACA75C , 32'hFD97F670 , 32'hEA73FE60 , 32'hE06E7060 , 32'h0243E46C , 32'hF8F1D238 , 32'h0926C1B0 , 32'h00DD8C0B , 32'h12EE5FC0 , 32'hF6838A90 , 32'hFDF3D7AC , 32'h095E83D0 , 32'hF88F0398 , 32'h19D4E540 , 32'h1063C580 , 32'h0E2048F0 , 32'hFA7B2168 , 32'hEBFD7CC0 , 32'h0C696DD0 , 32'h042B4BB0 , 32'hF8F0FC58 , 32'hFFAED917 , 32'hF3D3A170 , 32'h037F37D4 , 32'h0984D1D0 , 32'h010B6C80 , 32'h056B1D68 , 32'h08E60C00 , 32'h040A9218 , 32'h01871D8C , 32'hFAE2E600 , 32'hFD993BA4 , 32'h01C5A320 , 32'h01CA1070 , 32'h0060FF02 , 32'h01291CA8 , 32'hFA8F7CB0 , 32'hF84C17B8 , 32'hFC1F0714 , 32'h067DC6E0 , 32'h00945A55 , 32'h043DC720 , 32'hFFC2ED5D , 32'h01626D34 , 32'h00044FF4 , 32'hFFFF9A52 , 32'hFFFDBBFD , 32'hFFFD2404 , 32'hFFFE9F4B , 32'h00016AE7 , 32'h0001321A , 32'hFFFFF078 , 32'h00011F04 , 32'h0002083A} , 
{32'hFFFC87FA , 32'hFFFBAC72 , 32'hFFFDA67A , 32'hFFFD82F6 , 32'hFFFCC599 , 32'h0004A9B2 , 32'hFFFF6478 , 32'hFFFA35FF , 32'hFFFEC983 , 32'h000DDF3B , 32'h0000E434 , 32'hFFFE88AC , 32'hFFF56484 , 32'hFFFFE5A2 , 32'hFFFD225F , 32'hFFFDAD54 , 32'hFFFF78A3 , 32'hFFFC9FFF , 32'hFFFCDFFF , 32'hFFFA47DA , 32'h0002A9FF , 32'h0006F25F , 32'h000BF9C5 , 32'hFFFFBB45 , 32'h0001F9A0 , 32'h00076A73 , 32'hFFFBF152 , 32'h0002713A , 32'hFFFEAAFD , 32'hFFFF3B93 , 32'hFFF8ED44 , 32'hFFFDCAF8 , 32'hFFFCE8A2 , 32'hFFF5DB59 , 32'hFFFFB24D , 32'hFFFC5DDA , 32'hFFFC600F , 32'hFFF67FA5 , 32'h0000B201 , 32'h000427BC , 32'h00015AE4 , 32'hFFFE5B4C , 32'h0003876C , 32'hFFFCB3B7 , 32'hFFFC0643 , 32'h00046049 , 32'hFFFCD313 , 32'hFFFF6CBC , 32'hFFFA54BF , 32'hFFFC92FA , 32'h0004B232 , 32'hFFFA726E , 32'h00014BCE , 32'hFFF5C57B , 32'hFFFF9F38 , 32'hFFF84688 , 32'h000146CC , 32'h0000680B , 32'hFFFD27A7 , 32'h0005B0A4 , 32'h00049627 , 32'hFFFBBFA5 , 32'hFFFA8285 , 32'hFFF3A05E , 32'hFFF83110 , 32'hFFFBED89 , 32'hFFF5DDE7 , 32'h00025E18 , 32'hFFFF9F57 , 32'hFFFECC32 , 32'h0001B23D , 32'h000780A5 , 32'h000210A5 , 32'hFFFEBC4F , 32'hFFFE3F29 , 32'hFFFCA7D2 , 32'h0001F1E9 , 32'h0002037F , 32'hFFFCE2AC , 32'h0002B3C7 , 32'h0001BFD7 , 32'h0005EED3 , 32'h0002A593 , 32'h0003759B , 32'h00003519 , 32'h00040AE4 , 32'hFFF8AA80 , 32'hFFFDD9D1 , 32'hFFFFD057 , 32'hFFFFEBFD , 32'hFFFB4F69 , 32'hFFFBFB11 , 32'h00027420 , 32'hFFFCCF98 , 32'h0000F5B7 , 32'h0002867A , 32'h0007CCE8 , 32'hFFFF42D6 , 32'h00052544 , 32'h00016E49} , 
{32'h3BC19940 , 32'h39EE3080 , 32'h0C7C9F10 , 32'h13B195E0 , 32'hFA538788 , 32'hC63BBB00 , 32'hDDDC3B00 , 32'hF9DA9C00 , 32'h7C82CC80 , 32'h37CC67C0 , 32'h00CA7155 , 32'hFA95CA78 , 32'h13E785A0 , 32'h0F198300 , 32'hC59EA080 , 32'hE50D04A0 , 32'hF7ABF070 , 32'hD6EA7940 , 32'hF1847060 , 32'hD66E4780 , 32'h10307260 , 32'h02F67A50 , 32'h2EA560C0 , 32'h038BB438 , 32'h0C115EC0 , 32'hF52EB570 , 32'hEA609E60 , 32'h06BE2020 , 32'hE99F9CA0 , 32'h1E7AC500 , 32'h0062C0E8 , 32'h04B54690 , 32'h0267E91C , 32'hF29C5950 , 32'hF017F5F0 , 32'hF3E6E0A0 , 32'h0A2A9EC0 , 32'h0C99C360 , 32'hE7625760 , 32'hF8AF3DD0 , 32'h0BA138F0 , 32'h05C62C68 , 32'hE808A760 , 32'h11BF9380 , 32'h0666BB20 , 32'h06F102E8 , 32'hFBD2D788 , 32'hE788C5C0 , 32'hFB5572C0 , 32'hFB51B708 , 32'hEC9A5160 , 32'hFB048A30 , 32'hF8AB2148 , 32'hF7D0C9B0 , 32'hF82F11D0 , 32'h100BEB40 , 32'hF3794000 , 32'hF5DA2850 , 32'hF74C4440 , 32'hEFF07A00 , 32'hFB170328 , 32'hF4A76820 , 32'hFCE55FFC , 32'h0D330420 , 32'hEFE89920 , 32'hE41072E0 , 32'h040BE438 , 32'hFCEBCB4C , 32'h0DD6D830 , 32'hFD90FBCC , 32'h0238DABC , 32'h05F9ED80 , 32'hFF351985 , 32'h12DA54E0 , 32'hF9DBD8E0 , 32'h02A43214 , 32'h071C09D8 , 32'hFCE75128 , 32'h0033D1DA , 32'hFF33A134 , 32'h053D5948 , 32'h068D2790 , 32'hFFBEA180 , 32'hFB54D668 , 32'h0351154C , 32'hF7C9A770 , 32'hFEC2E1E8 , 32'hFAD0D7B0 , 32'hF9C5BA40 , 32'h018EE318 , 32'h0005B308 , 32'hFFFF57CC , 32'hFFFD0AAF , 32'hFFFF1CE5 , 32'hFFFF834B , 32'hFFFDC538 , 32'hFFFEEA84 , 32'h0003AEE2 , 32'hFFFE29FB , 32'h00001515} , 
{32'h21FE10C0 , 32'hFAD012F0 , 32'h5C1E3F00 , 32'h25CC3640 , 32'h20D6E780 , 32'h2C100240 , 32'h0F2644A0 , 32'hFDFA8224 , 32'h2E53D980 , 32'h0C977E00 , 32'hDEF89200 , 32'hE6AE9C40 , 32'hC9445CC0 , 32'hBE8E3B80 , 32'hF18E9670 , 32'h05712DF8 , 32'hCD711140 , 32'h097CC080 , 32'h1F8F0160 , 32'h147F9C80 , 32'h27FED8C0 , 32'hD77A1900 , 32'h1DF44D00 , 32'hFD8FC7A4 , 32'hFC358234 , 32'h11552A20 , 32'h1EDF60A0 , 32'hF34B6C60 , 32'h03D35490 , 32'h04A76170 , 32'hE96AC600 , 32'hFA987408 , 32'h179E2A80 , 32'h14C95B80 , 32'hE7DAD480 , 32'h012B2500 , 32'hED51C1E0 , 32'h03278C38 , 32'hF2F98B10 , 32'hF7C7C020 , 32'h00DDDB8E , 32'hFD6D42F4 , 32'hEB8AA240 , 32'h094D2FC0 , 32'h05D526E0 , 32'h076A0148 , 32'hE871DE00 , 32'hE9CE8300 , 32'h0F582070 , 32'hF505D5E0 , 32'hF49CBBB0 , 32'hED9AE480 , 32'hF8BEA030 , 32'h050C58A0 , 32'hFC8D8794 , 32'h010476B4 , 32'hF474A7C0 , 32'h1AA27500 , 32'hF53DA410 , 32'hF6D603D0 , 32'h14DB0F20 , 32'h0414EC80 , 32'h04C99B58 , 32'h0439B820 , 32'hFB739178 , 32'hFBA53D48 , 32'hEB6EA820 , 32'h07B6C488 , 32'hEE3C9120 , 32'hF76C2510 , 32'hFE69913C , 32'h051FC6C8 , 32'hFC621B8C , 32'hEA7C9B20 , 32'hFDE84010 , 32'hFCF46840 , 32'hFBC8B178 , 32'hF8185CD8 , 32'h061CCF00 , 32'h0023744D , 32'hFFB2C2CF , 32'h0147C1A0 , 32'hFB673850 , 32'h013EFD00 , 32'h0267E38C , 32'h00509EED , 32'h0078ABCF , 32'hFDBA2424 , 32'h00A79A1E , 32'hFFF6AFBC , 32'h00013D07 , 32'h0000A77D , 32'hFFFBAD5D , 32'h0003CB3F , 32'hFFFB2AFA , 32'hFFFE1278 , 32'h0001605B , 32'h0003777D , 32'hFFFF8C38 , 32'h00016CD6} , 
{32'h00009CC0 , 32'h0009D889 , 32'h000206BB , 32'h00044165 , 32'hFFFE4B55 , 32'h000173D4 , 32'hFFFF3DAD , 32'h0006984E , 32'h000192F5 , 32'h00067882 , 32'h0001F862 , 32'hFFFABCC6 , 32'h0006C65A , 32'hFFF3536B , 32'hFFFAC16F , 32'h00046E82 , 32'h0001EBF5 , 32'h0004F4D9 , 32'hFFFC4837 , 32'hFFFD692C , 32'h00021D52 , 32'hFFFCF10C , 32'h00045287 , 32'hFFFF4CC3 , 32'h0001FA0A , 32'h0002B83D , 32'h0004FAAF , 32'hFFFC0B4D , 32'h0001051E , 32'hFFF9B9BC , 32'hFFF9D458 , 32'hFFFEB57C , 32'h00004DAD , 32'h000544D5 , 32'h000606B2 , 32'hFFF8BCE1 , 32'hFFFC066B , 32'hFFFDC15E , 32'hFFFA082C , 32'hFFF9CA62 , 32'h00021DC0 , 32'hFFFD1DC1 , 32'h00032B1B , 32'hFFFA901F , 32'h0005E1A6 , 32'hFFFB2AA7 , 32'h00044501 , 32'hFFF7A5C6 , 32'h0000E0E3 , 32'hFFFCE048 , 32'h000402D7 , 32'h00054956 , 32'hFFFF2E62 , 32'h000154FE , 32'h0001DE1B , 32'hFFFF7BE6 , 32'hFFF84AF3 , 32'h0000AD1E , 32'h00057D30 , 32'h00041154 , 32'hFFFF40C7 , 32'h0002748F , 32'h00059D86 , 32'h0002C616 , 32'hFFFD7F04 , 32'hFFF902AA , 32'h0000168B , 32'h0003D5EC , 32'h0004EF81 , 32'h00021C97 , 32'h000329DA , 32'h0007C426 , 32'h00021457 , 32'h00099400 , 32'h0005DEDF , 32'h00019D5D , 32'hFFFBF4DB , 32'hFFF66DAC , 32'h000021B2 , 32'hFFF37B81 , 32'h00004BBD , 32'hFFFF2D2E , 32'hFFFDE9C4 , 32'h0000CD68 , 32'hFFFE3062 , 32'h0005C169 , 32'hFFFEF399 , 32'hFFFD3446 , 32'h0001D007 , 32'hFFFF9E40 , 32'h0007C34D , 32'hFFFC6532 , 32'hFFFF9ACD , 32'hFFFDFAA6 , 32'h0004813F , 32'hFFF8D839 , 32'hFFFFEC83 , 32'h0005FF44 , 32'hFFFCDD07 , 32'hFFFD1EFB} , 
{32'h00014924 , 32'h00013075 , 32'h000707EE , 32'h0001F27B , 32'h00094BDB , 32'hFFFD2DEB , 32'hFFFFAFBC , 32'h0000831F , 32'h00008E59 , 32'h0004453F , 32'h0005C0C1 , 32'hFFFA56F6 , 32'hFFFFC326 , 32'hFFFAD0C4 , 32'h00015656 , 32'h00059BFB , 32'h00047156 , 32'hFFFF5F55 , 32'h0002B59C , 32'hFFFCB27F , 32'hFFFD8B24 , 32'h0009759A , 32'hFFF8309C , 32'h00003D28 , 32'h00019A5B , 32'h00014AD4 , 32'hFFF87366 , 32'h00020643 , 32'h000182A5 , 32'h0005AC8A , 32'h00008E07 , 32'hFFFD47BB , 32'h00032F7F , 32'hFFFEE5EA , 32'hFFFFA8E5 , 32'hFFF710E4 , 32'hFFFC1C53 , 32'h0008D28B , 32'h0000636E , 32'hFFFDC376 , 32'h00052117 , 32'h00019866 , 32'hFFFCD908 , 32'h00033138 , 32'hFFF6B559 , 32'hFFFC7E39 , 32'h00057708 , 32'h00026580 , 32'h00041564 , 32'h000610C8 , 32'hFFFCC97B , 32'h0001651B , 32'hFFF7074F , 32'h000445EC , 32'hFFFF0B8E , 32'hFFFF914B , 32'h0003EE20 , 32'h00003B7C , 32'h0004788A , 32'h00039A93 , 32'hFFFA0EA0 , 32'hFFFD857A , 32'hFFFFAF03 , 32'h00033197 , 32'hFFFDB8E6 , 32'h0000D5A5 , 32'h0003255A , 32'h0005F50F , 32'h0001C5B2 , 32'h00089D88 , 32'h00033A99 , 32'h00038A21 , 32'hFFFE1717 , 32'h00018CCD , 32'hFFF96E5E , 32'hFFFFBC69 , 32'h0003A715 , 32'hFFFCB602 , 32'h000255A2 , 32'h0002F071 , 32'h0000675D , 32'hFFFF4100 , 32'h0006DB7E , 32'hFFFC69DA , 32'hFFFD146D , 32'h0002CAED , 32'hFFFFB565 , 32'h0005ED8B , 32'hFFFB99BF , 32'hFFFF1FCA , 32'hFFFCA985 , 32'h00018B07 , 32'h0003B47C , 32'h00009049 , 32'h00055402 , 32'hFFFAA7FA , 32'h00048459 , 32'hFFFAA3DF , 32'hFFFDD795 , 32'h000776F5} , 
{32'h0811F4F0 , 32'h015CFA8C , 32'h0BA5FC80 , 32'hF4056CD0 , 32'hE47FCDA0 , 32'hE1AAB580 , 32'hE568A720 , 32'hFC96A67C , 32'hEB7C4460 , 32'hFA115E10 , 32'h0E1FBE30 , 32'hEBB70EA0 , 32'hD61CF880 , 32'h0D445DE0 , 32'hF5999980 , 32'hEFF2BF00 , 32'h05BF7258 , 32'hF62ED8C0 , 32'h05D1D2F0 , 32'hFEA73DE4 , 32'h07C38810 , 32'h0DF8B400 , 32'h00DC02A8 , 32'h03E684D8 , 32'h07B775D8 , 32'h0D52F480 , 32'hF954B480 , 32'h03D5E0E4 , 32'hFAEB9480 , 32'hFABF6400 , 32'hF7E94AF0 , 32'h0AF85C30 , 32'h088DE630 , 32'hFBC45A70 , 32'hE3536B80 , 32'hF6527DF0 , 32'hFB6B3B48 , 32'hF7BA4830 , 32'hEE5D2A00 , 32'h057B3110 , 32'h03210D3C , 32'h0B35BA60 , 32'h1C363B20 , 32'h08D3D5D0 , 32'hEE49DB00 , 32'h0632C230 , 32'hEEA42B20 , 32'hFF3E17FD , 32'hFB3D7DD0 , 32'hF82FB2C8 , 32'h02BD9364 , 32'hFD96CDE8 , 32'hFDF9D7E8 , 32'h0B01A020 , 32'hF9100240 , 32'hF531A370 , 32'hFFFB5740 , 32'h02675EA4 , 32'hEF8289E0 , 32'h0B129690 , 32'hF27A8DA0 , 32'h0753CCB8 , 32'h119A8280 , 32'h137B6300 , 32'h0DAC16C0 , 32'h064A14D0 , 32'h02740518 , 32'hFFCD989D , 32'h02B55F28 , 32'h08635520 , 32'h03D9BC6C , 32'hF4DC29B0 , 32'hF656A410 , 32'h011F21E8 , 32'h04F49EF8 , 32'h05327248 , 32'hF543D8A0 , 32'hFA936590 , 32'hFE8BB2EC , 32'hFFF50B80 , 32'h02F2F628 , 32'hFCBEC77C , 32'hF79159B0 , 32'h04E95668 , 32'hF7E71920 , 32'hFE8F64CC , 32'hFEC20390 , 32'h044DFC60 , 32'h01B7DAB4 , 32'hFFF9669A , 32'h0003ED28 , 32'h0002F30F , 32'hFFFF42E0 , 32'hFFFEAE23 , 32'h00012D8D , 32'hFFFFEC0E , 32'hFFFEB5D7 , 32'h0007375E , 32'h0002450A , 32'hFFFECF22} , 
{32'h7FFFFFFF , 32'hC215E480 , 32'hCED86D40 , 32'hE57B5780 , 32'h71E0FB00 , 32'h0EA08170 , 32'hA1186880 , 32'h02E93EF4 , 32'h084823A0 , 32'hDD7A4900 , 32'h0710EAF0 , 32'h2EDECC80 , 32'hEB7CD1C0 , 32'h2C739080 , 32'h15EE7BA0 , 32'h0F3FE850 , 32'h3309ACC0 , 32'h19CC2480 , 32'hFDFBF8C8 , 32'hFF47E50F , 32'h20F24380 , 32'hE7C7A600 , 32'hEAC2BB20 , 32'h0A734D00 , 32'h06839298 , 32'h1901ABC0 , 32'h0C51E4E0 , 32'h0F1AD4D0 , 32'h0F87A520 , 32'hF9A6CD38 , 32'h2A814C40 , 32'h0279DCD0 , 32'hF23D31E0 , 32'hEDFC1A00 , 32'h142085E0 , 32'h0C002930 , 32'hFB712B40 , 32'hF5BA2940 , 32'hED2904A0 , 32'hED982580 , 32'hFF3828F2 , 32'hED8C7740 , 32'h0ECB5340 , 32'h14B61DC0 , 32'hF3FB7920 , 32'hF49871F0 , 32'hFEE66AD4 , 32'h080A4B20 , 32'h04350040 , 32'hE6AC0CE0 , 32'hFD8EE9D0 , 32'hFC933F04 , 32'hEABF5A20 , 32'hFFF3112E , 32'h01C0A34C , 32'h0702B728 , 32'h01C0AC24 , 32'hFA8B43B0 , 32'hFCCB7B7C , 32'h07649040 , 32'hF4B6A3A0 , 32'hF7FFE230 , 32'h030FEDEC , 32'h01596F70 , 32'hFC279374 , 32'h008AA884 , 32'hFA92F3B8 , 32'hFB3BC2D8 , 32'h05B1E0D8 , 32'h0658D920 , 32'hF8057E00 , 32'h0725CC70 , 32'hFEEA5F24 , 32'hFFDF3FB1 , 32'h025C0AA0 , 32'h0599FB58 , 32'h02E0AB80 , 32'hEBC7FC80 , 32'hFD7D7C70 , 32'h03DD3234 , 32'h0287E6CC , 32'hFABAD148 , 32'hF6A2C310 , 32'hFB2A2D98 , 32'h02355A54 , 32'hFD8B3A1C , 32'h00954C9F , 32'hF643FF20 , 32'hFF48716D , 32'hFF6BCD3B , 32'hFFFB1D71 , 32'hFFFE6BB0 , 32'hFFFFD451 , 32'h000413F0 , 32'hFFFD8177 , 32'hFFFE94B9 , 32'hFFFBD729 , 32'hFFFF1D24 , 32'hFFFE6E14 , 32'hFFFFF1B5} , 
{32'hBD545C80 , 32'h7FFFFFFF , 32'h70ECEC00 , 32'h44A0C300 , 32'hF8E185B8 , 32'hF559B8C0 , 32'hFBF55E30 , 32'hF8266FB8 , 32'hFDB5B538 , 32'h02044800 , 32'h0D1EC9C0 , 32'h3C36AB00 , 32'h12D28E20 , 32'hE07BC620 , 32'hFD0F099C , 32'hEFE64CC0 , 32'hE9594BE0 , 32'hDA139D00 , 32'hE6D351A0 , 32'hEC34D700 , 32'h18AFC100 , 32'h26539700 , 32'hE4830240 , 32'h361F5A80 , 32'hEE1E9600 , 32'hF25B5CD0 , 32'h0BEFC150 , 32'h0FB01450 , 32'hEC0526A0 , 32'h17F3C2E0 , 32'h23DC6040 , 32'hEFC55D80 , 32'h1A1015E0 , 32'hD323B500 , 32'h04E12988 , 32'hE7C478C0 , 32'h0A78E770 , 32'hEEDACCA0 , 32'h066979E0 , 32'hE495D520 , 32'h10B84160 , 32'h08510340 , 32'hFCF59B14 , 32'hEAE5D460 , 32'h01E5B67C , 32'h0048F8A5 , 32'h024308E4 , 32'h101A0F80 , 32'hFED140F0 , 32'h1BC23DC0 , 32'hFD8809BC , 32'hFBB395F8 , 32'hFC627100 , 32'h0D1703E0 , 32'h0596FB40 , 32'hF9A00448 , 32'hFCC1EFCC , 32'h076DB630 , 32'h0D2D2760 , 32'hF86752C8 , 32'hFED7D664 , 32'hFD6D1B30 , 32'h046BEBA8 , 32'hF63B6DD0 , 32'h082343D0 , 32'hEED28FA0 , 32'hFD225228 , 32'h01B26FA4 , 32'hF4FAF630 , 32'hFD683430 , 32'h001A327E , 32'hFE45DB28 , 32'hFB7E3F08 , 32'hFDB93028 , 32'h09EBE7E0 , 32'hFEBE0468 , 32'hFE70E714 , 32'hF72C0B70 , 32'h0077FF24 , 32'hF9D2D1F8 , 32'hFEACEFA0 , 32'hFE8825D8 , 32'hFEDF6D40 , 32'h06C627F0 , 32'hFDDE2DC8 , 32'hFE691854 , 32'hFF1746C5 , 32'hFEAEB94C , 32'h03435388 , 32'h0174BCD8 , 32'h00002B82 , 32'hFFF8EC2D , 32'hFFFEB39B , 32'h00038B8A , 32'h0000CC7B , 32'h0002247D , 32'h00015CFB , 32'hFFFF7910 , 32'h00012213 , 32'h0002F5C5} , 
{32'hD2F2BC80 , 32'h3B4AACC0 , 32'h3D1A1200 , 32'h4909F480 , 32'h0026E810 , 32'hD7EC8480 , 32'h0E9234A0 , 32'hF5C364C0 , 32'h08DAF3A0 , 32'h1FA7A7A0 , 32'h36952F40 , 32'hFFE02127 , 32'hFEE7F1C0 , 32'hEB8A7160 , 32'h25A01BC0 , 32'h0C010FC0 , 32'h049C59B0 , 32'hEA30D540 , 32'hF82CE510 , 32'hFF8762BA , 32'hF70ECF70 , 32'h195C63C0 , 32'h0856A640 , 32'h0390881C , 32'h2430E7C0 , 32'h26732D40 , 32'hD89BAD00 , 32'h032574AC , 32'h167ED000 , 32'h02C59A4C , 32'hF923D4E8 , 32'hF565EC70 , 32'hEDBCA8A0 , 32'h128DFB00 , 32'h17515280 , 32'hFF1F1A30 , 32'h065BC840 , 32'hF300FD50 , 32'h0BC51A90 , 32'hE68EA9E0 , 32'hF9FE4E88 , 32'hEF570D40 , 32'hF6AD6650 , 32'hF0FC87E0 , 32'hE2778940 , 32'hFD0D80D0 , 32'h1BAA9160 , 32'hF41F4690 , 32'h07466048 , 32'hE79D6540 , 32'hFE5A9654 , 32'hF955AD50 , 32'hF3A4AE90 , 32'hF22C1A60 , 32'h0215DCB8 , 32'h0B4EAD90 , 32'h143E2FE0 , 32'hFCC2936C , 32'h112BF8A0 , 32'hFB4583C8 , 32'hF8AA4128 , 32'h15CB7000 , 32'hF3FD7B40 , 32'h0485FE58 , 32'h00959DA7 , 32'h03C7A484 , 32'hFD12FB64 , 32'hFB691010 , 32'h0C204480 , 32'h04120BC0 , 32'h0106A144 , 32'hFD28FE90 , 32'h028C2750 , 32'hF0A93230 , 32'h0D5DEB30 , 32'hFBA70550 , 32'hFCF41668 , 32'h01549F28 , 32'hFB9ACDE8 , 32'hF049EEA0 , 32'hFD6E2528 , 32'h03301AB8 , 32'hFC5E8700 , 32'hFD9C4278 , 32'hFEBCE000 , 32'hFE86B524 , 32'hFFC91322 , 32'hFF814B1F , 32'hFE265EFC , 32'hFF519E60 , 32'h0003559C , 32'h0001B9BC , 32'hFFFF3DCE , 32'h00015FD6 , 32'h00008155 , 32'hFFFBF492 , 32'h0002C64C , 32'h00002879 , 32'h00029F9B , 32'hFFFEADE3} , 
{32'hFFFB75B9 , 32'h0002B493 , 32'hFFFE219F , 32'h0003CBDB , 32'hFFF7A22E , 32'h0000A901 , 32'hFFF6F90C , 32'h0000628D , 32'hFFFDB321 , 32'hFFF49CC9 , 32'hFFF81D67 , 32'hFFF426BC , 32'h000597D8 , 32'h000A3D13 , 32'hFFFB1629 , 32'h0006828C , 32'h00030420 , 32'h000440B3 , 32'h0000EE78 , 32'h0008426B , 32'h00078184 , 32'hFFFE2EA2 , 32'hFFF56A2F , 32'hFFFB752B , 32'h00081566 , 32'hFFFCC167 , 32'hFFFEFB70 , 32'hFFFFA827 , 32'h0004D171 , 32'h000D0C58 , 32'h000032A9 , 32'hFFFCB30F , 32'hFFFF3864 , 32'h0009DE34 , 32'h0001036C , 32'h0001D9FE , 32'h0004B26D , 32'h0004BFFC , 32'h00096674 , 32'hFFF3A320 , 32'hFFF8FA96 , 32'hFFFF0E6C , 32'h0008C5C1 , 32'hFFFEA502 , 32'h000AB7F9 , 32'hFFFA119B , 32'h0001B957 , 32'hFFFD95BF , 32'hFFFAE91B , 32'h000C317D , 32'h0003B006 , 32'h00080E6A , 32'hFFFB4A16 , 32'h000627E0 , 32'h0000EFA0 , 32'h0005FFC0 , 32'hFFFFC4E3 , 32'hFFFB44F2 , 32'h0000C0A4 , 32'hFFFBB519 , 32'h0002996F , 32'h0000A12F , 32'h00012768 , 32'h0002B0B6 , 32'h0001F1A0 , 32'h00013E3A , 32'hFFFDE56B , 32'h000AA1B7 , 32'hFFFDA0A3 , 32'h00025DA6 , 32'hFFF500E5 , 32'h0003219F , 32'hFFFE13EF , 32'hFFFDFB36 , 32'hFFFAA6CE , 32'hFFF7C059 , 32'hFFF7221B , 32'h00019304 , 32'hFFFBD5D3 , 32'hFFFB66CE , 32'h0000139F , 32'h000A5DD1 , 32'h0003FA87 , 32'hFFFC5FD8 , 32'hFFF9E936 , 32'hFFFFB409 , 32'hFFFAE2CD , 32'hFFFE3623 , 32'h0007D13E , 32'h00018644 , 32'h0008BB44 , 32'h0003B0B4 , 32'hFFFBCD0C , 32'hFFFFC209 , 32'h00016693 , 32'h00003D0A , 32'hFFFE89DE , 32'h0005C91D , 32'hFFFCCCC5 , 32'hFFFFF80A} , 
{32'h3726A540 , 32'hDE0EF6C0 , 32'h0872E660 , 32'h1551F7C0 , 32'hE8E5C940 , 32'h3E421900 , 32'hEAA433A0 , 32'hDB335BC0 , 32'hF736B230 , 32'hD9196840 , 32'h13E55760 , 32'h0BACA850 , 32'h0AEF6D60 , 32'h09B6F500 , 32'h056BC9D0 , 32'h08E8E370 , 32'h1193D820 , 32'h08543840 , 32'hF7A22830 , 32'h210850C0 , 32'h0E932F70 , 32'hF805A6C0 , 32'hFF85E697 , 32'h0A13A4C0 , 32'h2896FD00 , 32'hEE2B62C0 , 32'hDDFAD2C0 , 32'hF57F5690 , 32'h131270A0 , 32'h11EAB7C0 , 32'hF0BF67A0 , 32'hFC75F71C , 32'h0D041D80 , 32'h06DE24C0 , 32'h0F86E630 , 32'h174D35C0 , 32'hF4006480 , 32'hED60C740 , 32'hFABBED38 , 32'hF3FB0AE0 , 32'h0E708770 , 32'h0C3F0A70 , 32'hECCC2840 , 32'hF365DF70 , 32'h20EFC7C0 , 32'hF7DA3DD0 , 32'hF84DD908 , 32'h0977AC70 , 32'h04D9FD78 , 32'h042D5C40 , 32'hF1667680 , 32'hF984C738 , 32'h013C0604 , 32'hDCDA2B80 , 32'h06626810 , 32'h0B124310 , 32'hF9730C88 , 32'hE2A0C520 , 32'hF6F14580 , 32'h15AC2000 , 32'hFE6D9E60 , 32'h01BE2048 , 32'h0E3E6A80 , 32'h089D9DE0 , 32'h082B6BD0 , 32'hFA14D6E0 , 32'hF4898EA0 , 32'h136F2DA0 , 32'h0D06C1B0 , 32'hFF0FBB28 , 32'hF747BCC0 , 32'hF42EA510 , 32'hF8639868 , 32'hFC8F8520 , 32'h091D5BF0 , 32'hF88F74B8 , 32'h023A8554 , 32'h02D64030 , 32'h0BEB70F0 , 32'hFDE83D28 , 32'h066623D0 , 32'hFFB95903 , 32'hFB7C7EF0 , 32'hFF3DB526 , 32'hFF1639DB , 32'hFC0C3B84 , 32'h022A73CC , 32'h00A15364 , 32'h00D6934B , 32'h0050915C , 32'hFFFCFFE5 , 32'h0000747E , 32'h00024853 , 32'h0002B780 , 32'h00041258 , 32'h00016CAB , 32'hFFFD9083 , 32'h00000C40 , 32'hFFFF102C , 32'hFFFEA178} , 
{32'hD937D640 , 32'h2CAEF300 , 32'h6517E300 , 32'hE92725E0 , 32'h27DAE840 , 32'hC37AB300 , 32'hDB577740 , 32'h0AAFD8F0 , 32'h01B25180 , 32'hDEBF6700 , 32'h239AAF80 , 32'hF454D710 , 32'h0AB92DA0 , 32'hE1022020 , 32'h025E3CF4 , 32'hC3B59480 , 32'hF8B73E00 , 32'hE1C23A00 , 32'h06E135D0 , 32'hF1D48E30 , 32'h05F1A630 , 32'hD9997C40 , 32'h05559A70 , 32'hEDABABA0 , 32'h101B74A0 , 32'hF4AF36D0 , 32'hF86D5EA0 , 32'hD3C6CBC0 , 32'h005EEC59 , 32'hC8FD5BC0 , 32'hE795C820 , 32'h0B6A6CB0 , 32'h056AF610 , 32'h0384D6B4 , 32'h1AD06AA0 , 32'hDB87BA00 , 32'h077A4F50 , 32'h1A3B2400 , 32'hFAC9AC90 , 32'h04EF3588 , 32'h00783360 , 32'hEDB84640 , 32'hF7C95F40 , 32'hFF75B48B , 32'h06A69518 , 32'h020C68E8 , 32'h1436E700 , 32'h096BE100 , 32'hEEA470A0 , 32'hF722BDD0 , 32'hFEC98B54 , 32'h154922A0 , 32'hF5C953B0 , 32'hEF045F00 , 32'h14062B80 , 32'hF3816D10 , 32'hFC561FC0 , 32'h00196E64 , 32'hFC0792E4 , 32'hF63EADB0 , 32'hE985E8A0 , 32'h00E83C67 , 32'h0B159A10 , 32'hF76133C0 , 32'h0012AAF7 , 32'hFF5763C6 , 32'hF0DBAD10 , 32'hFEB473B8 , 32'h05E78CF0 , 32'h11FC5D00 , 32'h019C5840 , 32'hF90E1B60 , 32'h06857440 , 32'h069A6638 , 32'h05B6AF48 , 32'h0731BA20 , 32'h07156890 , 32'h093C4E90 , 32'h05588C38 , 32'h095A8590 , 32'h02C43F84 , 32'hFC818C00 , 32'hF9725B48 , 32'h0112FCE0 , 32'hFA0D6498 , 32'hFC126E20 , 32'h05F49B70 , 32'h0283F5E4 , 32'h00980EA4 , 32'hFF2C0DC8 , 32'hFFFF9222 , 32'h0000B110 , 32'hFFFE83EA , 32'h00003BE9 , 32'hFFFAEBE0 , 32'h00030EF4 , 32'h0000FED0 , 32'hFFFCC8F7 , 32'hFFFD5BE9 , 32'h0002A0B4} , 
{32'h02ACF1B8 , 32'hFF4E4503 , 32'hFCCF9980 , 32'h018ADDB4 , 32'hFF7D822F , 32'hFD2BBB3C , 32'hFAB8E9A0 , 32'hFB33BFB0 , 32'hFD242BF0 , 32'h004D163E , 32'h03448B70 , 32'hFB453908 , 32'hFEC0921C , 32'hFCAEFB6C , 32'h021FE2C8 , 32'h00B70314 , 32'hFD5F4B10 , 32'h0825F140 , 32'hFF6F8B04 , 32'hFC9FEDEC , 32'h016B7FF4 , 32'h06EC38B0 , 32'h074C99E0 , 32'h010C989C , 32'hFF2A5138 , 32'hFD263250 , 32'hFFCDDAF7 , 32'h009DBCF1 , 32'hFA148520 , 32'hFAAB8738 , 32'h07372438 , 32'hFFF23176 , 32'h01E1E550 , 32'hFBF6DBD8 , 32'hF97A42E0 , 32'h01F971C0 , 32'hF89DAFE0 , 32'h054E48F0 , 32'hFDDEE9B4 , 32'hFB48AD38 , 32'h04DDF988 , 32'h072342C0 , 32'h0A56E570 , 32'hFE3A7578 , 32'h0008C20E , 32'h0271F578 , 32'hFAF45598 , 32'h0349DA24 , 32'h08B645E0 , 32'h0130FAF8 , 32'h0603C020 , 32'hFE569D44 , 32'hFFBE9B20 , 32'hFA3319A8 , 32'hF4552010 , 32'hFB51A568 , 32'h0131C6B4 , 32'hF9BDB410 , 32'hFCF42B08 , 32'hFBFBB358 , 32'h03C59BC0 , 32'hF9F36CE0 , 32'h02A27828 , 32'h045FE330 , 32'h0297FA50 , 32'h036DB520 , 32'hFC24F600 , 32'hFBCF9578 , 32'hFF1E10DA , 32'h00A61C35 , 32'hFA9A3E30 , 32'h015EDBB0 , 32'h0388BB4C , 32'hFC20F5FC , 32'hFB3DF038 , 32'h00F06981 , 32'h008266D0 , 32'h00CFD14E , 32'h038FD564 , 32'h000BD72B , 32'h02F240B0 , 32'hFF8C4E63 , 32'h00B23381 , 32'h0135D6FC , 32'hFCC2B244 , 32'hFF628B42 , 32'h01C7C928 , 32'hFD82A4B4 , 32'h0136BD68 , 32'hFFEB367D , 32'hFFF8DD3B , 32'h00000D46 , 32'hFFFA6F1F , 32'hFFF9E3B2 , 32'h0001B0FC , 32'h0004661A , 32'hFFFBDE12 , 32'hFFFD355C , 32'h000249D0 , 32'h0002D0A0} , 
{32'hFFFE8AE5 , 32'hFFFC064F , 32'hFFFAE2BF , 32'h0003E23D , 32'h000466F6 , 32'hFFFAD950 , 32'hFFFDC377 , 32'hFFFA89C6 , 32'h0000B917 , 32'h0002E073 , 32'hFFFF8586 , 32'hFFFE127E , 32'hFFFC631E , 32'hFFFDE6A8 , 32'hFFFDD1C4 , 32'hFFFEC480 , 32'h0008E315 , 32'h0007FE08 , 32'h000281E0 , 32'hFFFB19D3 , 32'hFFEEEAF9 , 32'h0000FA9E , 32'hFFFD627E , 32'h0000A018 , 32'hFFFFE25B , 32'hFFFC1276 , 32'h000092AF , 32'hFFFBCDC9 , 32'hFFFD28E0 , 32'h00033F9A , 32'h0001523A , 32'hFFFD7E00 , 32'h0009DBC9 , 32'h00045EA2 , 32'hFFFE0A7B , 32'h00035053 , 32'h00003879 , 32'hFFFEB36C , 32'hFFFBAEAB , 32'h00034B94 , 32'h0004F843 , 32'h0005A126 , 32'h0007A57A , 32'hFFFBA238 , 32'h000588CA , 32'hFFF8AB02 , 32'hFFFE0C32 , 32'hFFFB0655 , 32'h0000E04D , 32'h00049F79 , 32'h0001CF07 , 32'h0002D670 , 32'h0002DA90 , 32'h0003F8EA , 32'hFFFB9D90 , 32'h00040602 , 32'h00014740 , 32'hFFFF574A , 32'hFFFCC0A1 , 32'hFFFEFF46 , 32'h000894BD , 32'h0004579C , 32'h0006D2E3 , 32'hFFFF8001 , 32'h0003A63A , 32'h00008247 , 32'hFFFF5188 , 32'hFFF81260 , 32'h0005C4D9 , 32'hFFF60196 , 32'hFFFB0072 , 32'h0002F039 , 32'hFFFC91BF , 32'hFFFEEE32 , 32'hFFF5A994 , 32'hFFFA4E89 , 32'hFFFF1D80 , 32'h0005E5A6 , 32'hFFFF6EEC , 32'hFFFE4E43 , 32'h0003CFCC , 32'h0002CB3A , 32'hFFF76369 , 32'h000097EC , 32'hFFF8F52F , 32'h000694A8 , 32'h00003AFA , 32'h0003D873 , 32'h000206B1 , 32'hFFF9850A , 32'hFFF6D4B6 , 32'hFFF806A8 , 32'hFFFC4C25 , 32'hFFFF2428 , 32'hFFFDC9FA , 32'h0000B236 , 32'hFFFC98E0 , 32'hFFFB5571 , 32'hFFF8E772 , 32'h00064142} , 
{32'hE8418D00 , 32'hF73FB760 , 32'hE91C2BE0 , 32'h1ED2F080 , 32'hF7948710 , 32'h1BAD7C00 , 32'hF1677DD0 , 32'h0CAC40B0 , 32'h091DF140 , 32'hFD053008 , 32'hE5B44420 , 32'hF0800190 , 32'h00B165CC , 32'hF80A17A8 , 32'h09D86F20 , 32'hF2ACCA50 , 32'h134E58C0 , 32'hF775C810 , 32'hFE869000 , 32'h050E1568 , 32'h07703F58 , 32'h02E1D2A0 , 32'h09AA3EB0 , 32'hF7C153F0 , 32'h0FEE3310 , 32'h1291C9A0 , 32'hEE6B3720 , 32'h189A2560 , 32'hF21AE160 , 32'hEC429EE0 , 32'h10651680 , 32'h0F3B5DA0 , 32'h056BDCE0 , 32'h0F0C3D30 , 32'h03F90004 , 32'h0812B7B0 , 32'hFFA70626 , 32'hF6C692D0 , 32'hF94509E0 , 32'h16414640 , 32'hF5335260 , 32'h00C7FE79 , 32'hF9541AE8 , 32'h04841FB8 , 32'hED9CC040 , 32'h08A17020 , 32'h07252B20 , 32'hFBDD07E8 , 32'hF21CAC20 , 32'h0CEB5790 , 32'h153533C0 , 32'hFD151D14 , 32'hFAE380F8 , 32'hFCACA464 , 32'hFF2FBEA2 , 32'hEF245780 , 32'hF0FA7C30 , 32'hF19CDF90 , 32'hF1B961A0 , 32'h0B7B31D0 , 32'h03EEF580 , 32'hF96F6528 , 32'h0083B870 , 32'hF5F585B0 , 32'hFCC08B38 , 32'h0650A7E0 , 32'hFCDA3DC8 , 32'h0322A78C , 32'hF28CC550 , 32'h013E29C4 , 32'hFE6293C4 , 32'h050EC3B8 , 32'hFACCF7E8 , 32'hF53E2320 , 32'h06C629D8 , 32'hFE79C370 , 32'h04E838B8 , 32'h02AC268C , 32'hEF985BA0 , 32'h00AF980F , 32'hFCB741F8 , 32'h041B2548 , 32'h062B3548 , 32'h0158F3C0 , 32'hFEC46ED0 , 32'hF9ECC350 , 32'h06E45990 , 32'h01EEB430 , 32'hFD6E01C8 , 32'hFFAC4C95 , 32'hFFFDA2FE , 32'h0003E0F4 , 32'hFFFDEC5D , 32'h0003EF15 , 32'hFFFF2390 , 32'hFFFF5A0A , 32'h00028870 , 32'h00000270 , 32'h000255AD , 32'hFFFD6C3D} , 
{32'h14BA2040 , 32'h00AA5CBE , 32'h3CED8E80 , 32'hF58219A0 , 32'h236B7D80 , 32'h29454F00 , 32'hCC8ED2C0 , 32'hDE0E0080 , 32'hE6D6BAE0 , 32'hF3E59B90 , 32'hEC69C560 , 32'hED1D4F20 , 32'hF29221D0 , 32'hD981B680 , 32'hF70BE4C0 , 32'h029AFDD0 , 32'h07298A88 , 32'h1CFDD040 , 32'h0A5946A0 , 32'hEFE0C9E0 , 32'hF0372420 , 32'hEFB0CB00 , 32'h055102B8 , 32'h0A9AF400 , 32'hF2EF0550 , 32'h03576BF4 , 32'hEA805F00 , 32'h1F49EB80 , 32'h3312C280 , 32'hFEF9EFE8 , 32'hEFA36CA0 , 32'h025270F4 , 32'hFE48AC34 , 32'hF5DE8370 , 32'hF9F61190 , 32'hD70B7040 , 32'h2CC99C00 , 32'hD9C838C0 , 32'h05F9EEC0 , 32'h12DA3AC0 , 32'h101A47C0 , 32'h1BCC9500 , 32'h0560EEC0 , 32'hFD874958 , 32'h09F1DD30 , 32'h127F2C40 , 32'hFB6E9480 , 32'h020A6FA4 , 32'h0C8567F0 , 32'h0AE8CDF0 , 32'h0287CCF8 , 32'h24A5A3C0 , 32'h0EDD28E0 , 32'hEB219340 , 32'h0B4928F0 , 32'h0E44C770 , 32'h00ABF668 , 32'h080B6780 , 32'h0BF68C00 , 32'hECA324A0 , 32'hF7928630 , 32'h03DFBAC8 , 32'h053E0E38 , 32'h0293920C , 32'hFB4BE530 , 32'hFDBF87C4 , 32'hFD52462C , 32'hF50D2280 , 32'h03F2A0D0 , 32'hEAF17360 , 32'h024820D8 , 32'h05A52788 , 32'hFE3E00E0 , 32'hF9C692E0 , 32'hF6347130 , 32'h01FC0FD4 , 32'hF3B685A0 , 32'hF7D5E550 , 32'hF8532EB8 , 32'h08D39970 , 32'h0304DF54 , 32'h0138FDCC , 32'hFA7BE620 , 32'hF6AEF800 , 32'h093F7C50 , 32'hFFC32FDF , 32'hFEB90334 , 32'hFDF01554 , 32'hFF93A94E , 32'hFF23EC46 , 32'h0001C880 , 32'h00016E0A , 32'h0003786C , 32'hFFFD6251 , 32'h00024EBC , 32'h0003AF73 , 32'h00011AFA , 32'hFFFD3B91 , 32'hFFFE5C51 , 32'hFFFD298C} , 
{32'hF7623290 , 32'hF18739A0 , 32'hD01F68C0 , 32'h32341640 , 32'hE3B7C120 , 32'h25C66E40 , 32'hD3E1CCC0 , 32'h0D5BC8F0 , 32'hD2CCEBC0 , 32'h07415398 , 32'h0148D95C , 32'hD6C37440 , 32'h3EB76D80 , 32'h0CB0BDF0 , 32'h0B2C2050 , 32'h0AB55E90 , 32'hEE1BE5E0 , 32'hE95913E0 , 32'hF83BB958 , 32'hFF15837B , 32'hF5307770 , 32'h0417EDA0 , 32'h038085D4 , 32'hEE8714C0 , 32'h04D2B328 , 32'h21599640 , 32'h051F3EC0 , 32'h18780C60 , 32'hE5923DC0 , 32'hFA3035D0 , 32'hFCAE45BC , 32'hE891C1A0 , 32'h0A2523F0 , 32'hFFB690D4 , 32'hEC927BE0 , 32'h0118D898 , 32'h0A966F90 , 32'h015172E8 , 32'hFEF6B0FC , 32'hF8767400 , 32'hEA3EDC20 , 32'hF0ECD5E0 , 32'hFFA346EB , 32'h0431E660 , 32'hFFC42C96 , 32'hF55B7BB0 , 32'hFA54B5B8 , 32'hE0A76120 , 32'hD6EDA240 , 32'h0830FCC0 , 32'hF2D62EF0 , 32'h1672E5E0 , 32'h0025D674 , 32'hF78B1FB0 , 32'h030712E8 , 32'h003EA3C4 , 32'hFEC57004 , 32'hFDB3684C , 32'h018934E0 , 32'h04F03318 , 32'h01FDFA74 , 32'hFD4FCB0C , 32'h09F96220 , 32'h113A5B80 , 32'hF7B41F80 , 32'h0684B9B8 , 32'h07329E48 , 32'hFFCA2130 , 32'hFB17CE88 , 32'h06B1AEC0 , 32'hF591D2E0 , 32'h108E5880 , 32'hFC34D724 , 32'h08610C40 , 32'hFE35D130 , 32'hFB03D470 , 32'h0706C078 , 32'hFA9492B0 , 32'h07308188 , 32'hFC32170C , 32'h0152CDE4 , 32'hFEE89CE0 , 32'hF7A81B70 , 32'hFF164AC0 , 32'h035226B8 , 32'h067A9458 , 32'hF91187D0 , 32'hFDCDA788 , 32'hFF09B3CF , 32'hFEDE2AFC , 32'hFFFEE8E8 , 32'hFFFE0C9C , 32'hFFFC1963 , 32'h000252B7 , 32'hFFFBF986 , 32'hFFFF231A , 32'hFFFEDAC7 , 32'hFFF93F1B , 32'hFFFFF831 , 32'h0001DC30} , 
{32'hFFF8C1D2 , 32'hFFFD05E9 , 32'hFFF816CD , 32'h000461ED , 32'hFFFD66B4 , 32'hFFF8AA07 , 32'h0001B1D0 , 32'hFFFF7C57 , 32'hFFF5E0B9 , 32'h0005B89E , 32'h0005C38D , 32'h00024B0D , 32'h00034FB0 , 32'hFFFFA02E , 32'h00047661 , 32'hFFFC2E12 , 32'hFFF5BBCE , 32'hFFFF0141 , 32'hFFF508A1 , 32'hFFF8FAE2 , 32'h00022361 , 32'hFFFE7389 , 32'hFFFEF24B , 32'h0000D3C3 , 32'h0000E1F5 , 32'hFFFD9325 , 32'h00041871 , 32'h0001973D , 32'hFFFF99F9 , 32'hFFFE9406 , 32'hFFF4CFD0 , 32'hFFFF0EAE , 32'hFFFC508D , 32'hFFF5468A , 32'h0006DBFA , 32'h0005E685 , 32'hFFFBE2DF , 32'h0000CB02 , 32'h0009F07B , 32'h0007161E , 32'h000A8D87 , 32'h0002FCCD , 32'h0002D2C8 , 32'hFFFF7A89 , 32'hFFFB0080 , 32'hFFFE43C8 , 32'h0000AF4A , 32'hFFFCA4C1 , 32'h00056C66 , 32'h00021E81 , 32'h00032716 , 32'h0001B5EB , 32'hFFFE11D2 , 32'hFFFFFA8E , 32'hFFFD4CA6 , 32'hFFF88D9D , 32'h00043AF1 , 32'hFFFC030F , 32'hFFF7AC55 , 32'h00039630 , 32'h0005335B , 32'hFFF6C62D , 32'h00013DBD , 32'h00027143 , 32'h0000B4D3 , 32'hFFF9E22E , 32'h00088624 , 32'h00045AC9 , 32'h00031954 , 32'hFFFD105A , 32'h000081E3 , 32'h000967FB , 32'hFFFDA279 , 32'h00076727 , 32'h00055C06 , 32'hFFFAAC93 , 32'hFFFF1BA9 , 32'hFFFAA730 , 32'h0002430B , 32'h0003853A , 32'h0005CC12 , 32'h0005EB43 , 32'h00068536 , 32'hFFFAE769 , 32'hFFFAD210 , 32'hFFFA41D0 , 32'hFFFA1D3B , 32'hFFF822CB , 32'hFFFC7CBF , 32'h00009C1C , 32'hFFFB0B90 , 32'h00009C0D , 32'hFFFDE4B8 , 32'h0003F03B , 32'hFFFED286 , 32'hFFF7E770 , 32'hFFFF6D22 , 32'hFFFE9CCD , 32'h00032156 , 32'hFFF49BA4} , 
{32'h0CD48540 , 32'h0A58B940 , 32'h0B42EDB0 , 32'hF589EB70 , 32'hDE192D40 , 32'hFCA7FF78 , 32'hE51749E0 , 32'hFA574CC0 , 32'hF8BCA7E8 , 32'h03867C3C , 32'hFD2AC168 , 32'h0DD2DF70 , 32'hF11F4230 , 32'h0C7F96C0 , 32'h10AFF5C0 , 32'h12F6A600 , 32'hF7D81080 , 32'h0F37FD70 , 32'hF3F0F7A0 , 32'h078733D0 , 32'hF8FAF3F0 , 32'hEFCDF780 , 32'hF02AFA10 , 32'h1311E080 , 32'h069BEC90 , 32'hEF42D6E0 , 32'hE7BF95E0 , 32'h005F2D88 , 32'hF391CB40 , 32'hF9DBE280 , 32'h0B753000 , 32'hFDD95064 , 32'hEF18D4A0 , 32'h03D2D3F0 , 32'hFDAEB498 , 32'hFE097E0C , 32'hF3DCC0D0 , 32'h06C1FF68 , 32'h0E7C3C70 , 32'h039B2B6C , 32'hFA3D5660 , 32'h01DFB0E8 , 32'hF603F690 , 32'h00B5429C , 32'h05F09E30 , 32'hFD3063F8 , 32'h1E466B40 , 32'hEC959B40 , 32'hFA1B4B38 , 32'h141D3860 , 32'hFE75FBB4 , 32'hFFC54B86 , 32'hF9531230 , 32'h02254304 , 32'h10137420 , 32'hEF177080 , 32'hF70FD480 , 32'h0AB3D5F0 , 32'h026B4798 , 32'hECB38E40 , 32'h1646D820 , 32'hFFE4A679 , 32'hFCE99B74 , 32'h02DFF30C , 32'h0DA4A310 , 32'h0A5838B0 , 32'hF35F8810 , 32'hF3C5DC40 , 32'hFB43DBA8 , 32'hF8F6D240 , 32'hFF49C054 , 32'h00573331 , 32'hF1A19DC0 , 32'h0C5CD8B0 , 32'h02A12FF8 , 32'h0428E940 , 32'h02E27DC8 , 32'h0C0F31C0 , 32'hF41933A0 , 32'h02BC3A78 , 32'h0D82F670 , 32'h000F002B , 32'h03414310 , 32'hFE436B18 , 32'h0149474C , 32'hFD5E72A8 , 32'hF89379F8 , 32'hFEC894E8 , 32'h027B662C , 32'hFF9B72E7 , 32'hFFFEB2CA , 32'h0000652C , 32'hFFFD1833 , 32'h000059DC , 32'h000198EF , 32'hFFFE5C28 , 32'h00004364 , 32'h0000BD3B , 32'hFFFE957B , 32'hFFFE7CFA} , 
{32'hFFFDD91F , 32'hFFFE8650 , 32'h00035C01 , 32'hFFFFA21D , 32'h0006E950 , 32'hFFFD734C , 32'hFFFF6EF9 , 32'hFFFE6B41 , 32'hFFFFFF14 , 32'hFFFF2C8E , 32'h000373B0 , 32'hFFF5F551 , 32'hFFFBC23F , 32'hFFFF59C1 , 32'hFFFA2E40 , 32'hFFF79EED , 32'h0002AF37 , 32'h0000AFD5 , 32'hFFF569E9 , 32'hFFFE9C08 , 32'h00018253 , 32'h0002CA82 , 32'hFFFB7EDC , 32'h0006C5ED , 32'h0009CC00 , 32'h0007B63C , 32'hFFFCD894 , 32'h00029F2E , 32'h00072BDB , 32'h000454F3 , 32'hFFFC27FC , 32'h00076B2A , 32'h0004E3FF , 32'hFFFAC809 , 32'h000C3789 , 32'hFFFDD1C9 , 32'h0001B97F , 32'h0004784C , 32'h000405DA , 32'h00037E10 , 32'h00023FE5 , 32'h0007B52B , 32'h00099A18 , 32'hFFFFBD47 , 32'hFFFDE3FB , 32'hFFF768BE , 32'h00045CC0 , 32'h0000B38A , 32'hFFFE9FBC , 32'hFFFBE775 , 32'h00015214 , 32'h000208FC , 32'hFFF9EA07 , 32'h0001F6A5 , 32'h00037B37 , 32'hFFFFD698 , 32'hFFFDA08E , 32'h00027725 , 32'h0005F782 , 32'h0008580B , 32'h0002876B , 32'hFFFD6BA1 , 32'hFFFBF43F , 32'h0002FE6D , 32'hFFF9BE8A , 32'h0004E739 , 32'hFFFD70A0 , 32'h0002AD02 , 32'h0001BBDE , 32'hFFFBCAF0 , 32'hFFFFC41E , 32'hFFFBD39D , 32'h00066DD4 , 32'hFFFE3409 , 32'hFFFE7366 , 32'h00015B3B , 32'h0005B29E , 32'hFFFA9BA9 , 32'hFFFA210C , 32'h00073186 , 32'h000504F8 , 32'hFFFC8F53 , 32'hFFFB50FA , 32'hFFFF6980 , 32'h00078459 , 32'h0000F1BB , 32'hFFFBE4AB , 32'hFFFF0322 , 32'hFFFB2C5A , 32'h00039134 , 32'h00030827 , 32'hFFF92A57 , 32'hFFFEB691 , 32'hFFFE6C8E , 32'hFFF50796 , 32'hFFFFDFB7 , 32'hFFFD7CBA , 32'h0000FDFE , 32'hFFFE3BAB , 32'h0006E17C} , 
{32'h0000C465 , 32'hFFFC26EB , 32'h0000CA44 , 32'h0009627E , 32'hFFFA981A , 32'h0003E32C , 32'hFFFC345A , 32'hFFFBF44C , 32'hFFFC50CF , 32'h00001851 , 32'h0001EB71 , 32'hFFF50C27 , 32'hFFFD7A70 , 32'h0001182D , 32'h00081094 , 32'h000129C9 , 32'hFFFE51D9 , 32'hFFFD5E62 , 32'hFFFA242C , 32'hFFFF470B , 32'h000440B0 , 32'hFFFF0590 , 32'h0001802C , 32'h00004DA8 , 32'h00017468 , 32'h0001B15F , 32'h0007AFD1 , 32'h0003C311 , 32'hFFFA822C , 32'h0008C2F7 , 32'h000309D2 , 32'hFFFCB7F6 , 32'hFFFBBFEF , 32'h0000AB76 , 32'h00018081 , 32'h000BE790 , 32'hFFFCC3D8 , 32'hFFFD419E , 32'hFFFC5966 , 32'hFFFEC42C , 32'hFFFAAA4E , 32'hFFFA8208 , 32'h0007A55C , 32'h0004804D , 32'hFFF9F518 , 32'hFFFD2E6E , 32'h0000163A , 32'hFFFABD96 , 32'hFFFE344D , 32'hFFFC7B50 , 32'hFFF49952 , 32'hFFFD3FBE , 32'h000ED129 , 32'h0001FF9A , 32'hFFF52A14 , 32'h000BC2FF , 32'hFFFCE333 , 32'h0006FB78 , 32'h00026847 , 32'hFFFF9F93 , 32'h00061418 , 32'h000146CB , 32'hFFFEBB62 , 32'h000666F8 , 32'hFFFBE1C6 , 32'hFFFF3D92 , 32'hFFFF713B , 32'h00052833 , 32'h000181A5 , 32'hFFFCDA60 , 32'hFFFF864B , 32'h0001A5B6 , 32'h0001A40C , 32'hFFFAFBBF , 32'hFFFF6F7B , 32'hFFF6E910 , 32'h000354B2 , 32'h0000DEBE , 32'hFFFD23E7 , 32'hFFF2A03D , 32'h0003D3B6 , 32'h00068C35 , 32'h0005110B , 32'h0000C2BD , 32'h00000FB0 , 32'h00006C33 , 32'hFFFFF565 , 32'hFFF9B6D3 , 32'hFFFF9F02 , 32'h00059FC4 , 32'hFFFFD492 , 32'hFFFCA018 , 32'hFFFFDFBE , 32'h000588BA , 32'h0000D4AA , 32'hFFF90DA4 , 32'hFFFF5072 , 32'hFFFE12BC , 32'h0003A6E5 , 32'hFFFE69E0} , 
{32'h0BB27910 , 32'hEB495CC0 , 32'hFA0CEF98 , 32'h28398540 , 32'hEBA5FCA0 , 32'hFA8FDBE0 , 32'hFEDA5FA0 , 32'h14D23A20 , 32'hE38EF200 , 32'h11A9E300 , 32'h030CF910 , 32'h048B8798 , 32'h0E1834C0 , 32'h166031E0 , 32'hF5CBCB80 , 32'hFADF4F30 , 32'h03EA3060 , 32'h05DF4040 , 32'h127B84E0 , 32'h07588E48 , 32'hFB868FF0 , 32'h012B4CC4 , 32'hDDCB71C0 , 32'hF08FF1A0 , 32'hF3BC55F0 , 32'hEC6D2960 , 32'h0B3A3AF0 , 32'hF185CD10 , 32'hE1DBB6E0 , 32'h05CB9210 , 32'hEEE3AC40 , 32'h052F14D0 , 32'hFAE2D928 , 32'h04B00110 , 32'hF2298720 , 32'hFE16C4D0 , 32'hFA7E2AC8 , 32'hEEB93900 , 32'hFFF66BAC , 32'hFF0173E7 , 32'h03EFE388 , 32'h07EC1620 , 32'h0A068A90 , 32'hF4A9F580 , 32'hFD9184C4 , 32'h02EFBE8C , 32'hFB374C60 , 32'h01E93B2C , 32'h03623B64 , 32'hE860BF00 , 32'hF73FE270 , 32'hF6B26550 , 32'hFBEBDC60 , 32'h063E0830 , 32'hF9901588 , 32'hE808A940 , 32'hF25693A0 , 32'h06F4ABC0 , 32'hF795F5F0 , 32'hF90AA7E8 , 32'hEB888220 , 32'hEE884F40 , 32'hFB8D5A50 , 32'hEEF10500 , 32'hF5CBD8C0 , 32'hFC050820 , 32'h0943DB30 , 32'hF8F95298 , 32'h095D0070 , 32'hF9977C30 , 32'h0493E118 , 32'hFBC3AD88 , 32'hFB122D60 , 32'h018CBAC0 , 32'h00EF89C5 , 32'h058D8320 , 32'h008F2000 , 32'h04140798 , 32'hFC44D234 , 32'hF9D663E0 , 32'hFFFAAE06 , 32'h04570178 , 32'hFCC2F1C4 , 32'hF2EC6640 , 32'h05D4DDE0 , 32'hFEAA8F94 , 32'h03280FCC , 32'h02464D14 , 32'h0649FD60 , 32'hFFC4D339 , 32'h000A3EAE , 32'h0004D978 , 32'h00015D44 , 32'hFFFF7B6C , 32'hFFFC175C , 32'h0007FDEE , 32'h0000471E , 32'hFFFE3CCC , 32'hFFFC97CE , 32'hFFFE92C9} , 
{32'h032F199C , 32'hFB0C2098 , 32'hF7964850 , 32'hECEAC5A0 , 32'hFEC077D4 , 32'h01C8B8C0 , 32'h027165B4 , 32'hFDA397D8 , 32'hF5FB7140 , 32'h00D45AAC , 32'hF63032D0 , 32'h095C3B10 , 32'h095CA540 , 32'hFA9FA868 , 32'hFE3FA140 , 32'hFD9A4F88 , 32'hFC7472A0 , 32'h056E1468 , 32'hFA6BB8A0 , 32'h09A28510 , 32'h01F75810 , 32'h01EA7998 , 32'h032A1724 , 32'h00B5D067 , 32'hFE21AC04 , 32'hFA42E348 , 32'hF2034690 , 32'h04CCAC98 , 32'hF4F71780 , 32'h093F51C0 , 32'h042CDE00 , 32'hFB452E48 , 32'hFC9FE2BC , 32'hFC48B8F0 , 32'hFB217018 , 32'h06DAE370 , 32'h07B4EC00 , 32'h00CAFD37 , 32'h06F8AE50 , 32'hF8211268 , 32'hFFCA765F , 32'hFBF74498 , 32'h0DE12170 , 32'h021AC878 , 32'h012A457C , 32'hFE976EF8 , 32'hF55C9900 , 32'h062BD9C8 , 32'h0C80A580 , 32'h009587F5 , 32'h1168A200 , 32'h02C6B754 , 32'h03053E08 , 32'h0899C980 , 32'hF9470958 , 32'hFB422888 , 32'hFB5847D8 , 32'h029380F0 , 32'h06E817D8 , 32'hFD25FB24 , 32'hFD613248 , 32'hFD6F7CFC , 32'hF6F6B7F0 , 32'h0983A290 , 32'hFA7E4D08 , 32'h0A19E6F0 , 32'hFD76E338 , 32'h035C6344 , 32'h04558F78 , 32'hF875F400 , 32'h08612AB0 , 32'hF65B8B40 , 32'h062D5420 , 32'hF871E6B0 , 32'h0465C8C8 , 32'hFF8ADE06 , 32'h021CF2FC , 32'hFEC04F98 , 32'h0230BA5C , 32'h050D0638 , 32'hFA080338 , 32'hFB27EBA8 , 32'hF9B340E0 , 32'h005D0CBF , 32'h04CD2540 , 32'h00EEB4D7 , 32'h02737FD0 , 32'hF7FBF940 , 32'hFA646E70 , 32'h00018E68 , 32'h00045B3C , 32'h0001CC9D , 32'hFFF990F4 , 32'hFFFFFEDA , 32'hFFFEA4CC , 32'hFFFBF350 , 32'h000632F3 , 32'h00013EE9 , 32'h0002D675 , 32'h0005CC7A} , 
{32'hFCFBDC20 , 32'hFF49AABE , 32'hF24EF590 , 32'h1412E740 , 32'h02113BBC , 32'h38288180 , 32'hF4D38B90 , 32'hFCD2EF54 , 32'hF10A9310 , 32'h01DFCC98 , 32'h037E0DC0 , 32'h1A4E5340 , 32'h0A396770 , 32'hF793ED00 , 32'h0DCA6620 , 32'hFE3665D4 , 32'hE866A2C0 , 32'h07F3CBB0 , 32'hE0D86680 , 32'hEC5D1800 , 32'hF3CFBBB0 , 32'h201E2A40 , 32'hDF456D00 , 32'h01940FEC , 32'hEFADD040 , 32'hFA887378 , 32'h032878A4 , 32'hE2BDBA00 , 32'hF0590500 , 32'hE312AD00 , 32'hE47D0CA0 , 32'h00D27A3D , 32'hEDF460C0 , 32'hFC8342BC , 32'hF51248B0 , 32'hF3096C30 , 32'h1299A920 , 32'hFD03B6A4 , 32'hED020480 , 32'h01C70380 , 32'hE82F2F40 , 32'h12D930A0 , 32'hFDEF37D4 , 32'hEBD08BE0 , 32'hFEC88BAC , 32'hE6F0E7C0 , 32'hEFCA6C20 , 32'hF603B7D0 , 32'h0A91EA40 , 32'hF26F29B0 , 32'hF41A0C20 , 32'hFDD9D5C4 , 32'hE39AEEE0 , 32'hF2E8A470 , 32'h09B1B2F0 , 32'h0257CDCC , 32'hFE319470 , 32'h11C87440 , 32'h07CA6018 , 32'h118B5000 , 32'h054EF790 , 32'hF48DBB40 , 32'hF9F31508 , 32'hFBC99148 , 32'hF6288D50 , 32'h12C87F60 , 32'hF5E57F60 , 32'h0006489C , 32'h02DAE2F0 , 32'h02E8406C , 32'h02CD1048 , 32'hFCD0F898 , 32'hFE8BAD74 , 32'h074DD1C0 , 32'h00932D6B , 32'hFE6D4F84 , 32'h01FFB280 , 32'hFE9E9220 , 32'h08BAC060 , 32'hF5E36720 , 32'hFDF3FE38 , 32'h0525D098 , 32'h020C34C8 , 32'h05AD2A68 , 32'h0116EA44 , 32'h019245F8 , 32'hFDA1D458 , 32'hF9B55A80 , 32'hFE033FC0 , 32'hFFB5D1E3 , 32'hFFFE6559 , 32'h0000A763 , 32'h00020E56 , 32'hFFFC3ABF , 32'hFFFF66A1 , 32'h00000490 , 32'h0003AC99 , 32'h0002EFDA , 32'h000104FF , 32'hFFFD5D36} , 
{32'h3E74B8C0 , 32'hE53E1020 , 32'hD2CE0800 , 32'hD032D740 , 32'h4D36E600 , 32'hCB288900 , 32'h483C8080 , 32'hDA039780 , 32'hFB777418 , 32'h1078ACE0 , 32'h3EFCFFC0 , 32'h241888C0 , 32'h34E33500 , 32'h3ACF5640 , 32'h260A90C0 , 32'h089D0A30 , 32'hDA20C340 , 32'h15B34880 , 32'h19D6AB60 , 32'h0060567A , 32'h1C034020 , 32'hFE1C7818 , 32'hEFBD30E0 , 32'hDBE5BC00 , 32'hF0233C60 , 32'hF5DA2DF0 , 32'h10B8A120 , 32'hDF75B6C0 , 32'h030C9CFC , 32'h067B5A38 , 32'hE5C1F9A0 , 32'hEA0C47A0 , 32'h0244D4E0 , 32'hEA090BC0 , 32'hFF0874C8 , 32'hFFF312EA , 32'h116D59A0 , 32'h0296FB08 , 32'hF884A938 , 32'h07A2D648 , 32'h0501D8D0 , 32'hF85E2E78 , 32'h069D9AC0 , 32'h10F3B0E0 , 32'h04DF61F8 , 32'h14C14080 , 32'hEF2623C0 , 32'h103D8E00 , 32'hEC6AD420 , 32'h145FD8A0 , 32'hE4DBA620 , 32'h0424A138 , 32'h062B1518 , 32'h04688AC0 , 32'hFF8FF1B6 , 32'hEFCE6380 , 32'h024AF980 , 32'h04768C30 , 32'h0A4351D0 , 32'h01AFAEB0 , 32'hFD207090 , 32'hFADFEC98 , 32'h00F46D85 , 32'hFFE9B432 , 32'h04E1C7C8 , 32'h00F7F1A7 , 32'hF9A78D68 , 32'h07E3E850 , 32'h0B288A00 , 32'h00BEDFB7 , 32'hED082300 , 32'hFA834140 , 32'hFA465360 , 32'hF4652510 , 32'hFAA788E0 , 32'hFFA2F53B , 32'hF4AC4680 , 32'h02B7F034 , 32'hFA333AF0 , 32'hF6F68F90 , 32'h008F7C38 , 32'h05067368 , 32'h076DC148 , 32'h00902F7B , 32'h0187FA0C , 32'hFFF7D65A , 32'hFFDD3977 , 32'hFB9D0070 , 32'hFCB61478 , 32'hFF7F8424 , 32'hFFFFF41E , 32'hFFFF0BB4 , 32'hFFFD5302 , 32'h0005E26D , 32'h00013120 , 32'hFFFCF41A , 32'hFFFF8894 , 32'h00023FFA , 32'hFFFEE9BE , 32'hFFFCE67D} , 
{32'hFFFCE431 , 32'h00023CAA , 32'hFFF79794 , 32'h000073A7 , 32'hFFF93638 , 32'hFFFA2A94 , 32'h0000D50B , 32'hFFF5F55D , 32'hFFFE6824 , 32'h00035DA8 , 32'hFFFFE41F , 32'hFFFCA01C , 32'h000079DC , 32'h00022597 , 32'h0008CF5C , 32'h0003AE7D , 32'h0000A0B5 , 32'hFFFABDFB , 32'hFFFFC5EB , 32'hFFFFB47D , 32'h0003B98C , 32'h00062BE0 , 32'h000156AC , 32'h0005AF5C , 32'hFFFFA603 , 32'h0002B1BF , 32'hFFFD52FB , 32'hFFFD7D45 , 32'h0005254F , 32'hFFFCAA84 , 32'hFFFF2073 , 32'h00032493 , 32'h000470F9 , 32'hFFFCD702 , 32'h0000D463 , 32'h00044A51 , 32'h0000A404 , 32'hFFF9E279 , 32'hFFF919AD , 32'hFFF91452 , 32'h00094997 , 32'hFFFEE187 , 32'hFFFC948F , 32'hFFFE9CFE , 32'hFFFCEB9C , 32'h0009B7D8 , 32'hFFFD23AC , 32'hFFF721A0 , 32'hFFF87702 , 32'h00023B7C , 32'hFFFB5FE2 , 32'h00046313 , 32'h00010A22 , 32'h0002B64A , 32'hFFFDB9D3 , 32'hFFFD6483 , 32'h0008C78F , 32'h0002F815 , 32'hFFF74E4E , 32'h0001D6FB , 32'h0002CF86 , 32'hFFFDFEFE , 32'h000897A6 , 32'hFFFB3E29 , 32'hFFF92D0F , 32'hFFF82994 , 32'hFFF9FB75 , 32'hFFFF0FCF , 32'hFFFE2274 , 32'h0003DF01 , 32'h0003DD14 , 32'h0006020A , 32'h0000159F , 32'hFFFE37A8 , 32'hFFF76F52 , 32'h00068495 , 32'h000088C7 , 32'hFFFCE71B , 32'h0001AE60 , 32'hFFFD09B6 , 32'h00004AD3 , 32'h00051DCE , 32'h0002F31F , 32'h000382E0 , 32'h000E45EB , 32'hFFFEBB31 , 32'h000079DA , 32'hFFFBBC4F , 32'h0005D678 , 32'hFFFC01D1 , 32'hFFF859F0 , 32'h00051EB8 , 32'hFFFE7EF0 , 32'h0002B211 , 32'hFFF966CF , 32'hFFFBC527 , 32'h000396E6 , 32'hFFF82D28 , 32'h00022A1D , 32'h00074E3F} , 
{32'h8382D580 , 32'h34FD5140 , 32'hB5196380 , 32'h5B3DC100 , 32'hCD97AA80 , 32'h61EA8A00 , 32'hEE582FA0 , 32'h6EEFEB00 , 32'hF231A5E0 , 32'h1733D760 , 32'h5A08B900 , 32'h56868180 , 32'hE5602960 , 32'hE46F6BE0 , 32'h097C7030 , 32'hEE970120 , 32'hD2007C00 , 32'h150CB660 , 32'h0F3BA600 , 32'h2DD9D340 , 32'h25A85900 , 32'hE85DBA60 , 32'h0C140630 , 32'h15A41BC0 , 32'hF4652EA0 , 32'hFBFF8670 , 32'hF5DF1560 , 32'h0A26AAB0 , 32'hE1C88860 , 32'hE7EDE160 , 32'hFC244B8C , 32'hE68CFD00 , 32'hF92B5B60 , 32'h0304F68C , 32'hD48CFF80 , 32'h153761A0 , 32'hFA0D38E0 , 32'hF2914D90 , 32'h037115D4 , 32'h01D9AD14 , 32'h069F80C8 , 32'h06D92C58 , 32'hFBE7C0A0 , 32'hFC172C38 , 32'h09473450 , 32'h02A42090 , 32'hFDF37AE8 , 32'hFE3B4634 , 32'hF06C2D90 , 32'hECF91440 , 32'h0FA9AE90 , 32'hFAE20558 , 32'h1DFCB660 , 32'hFF330B68 , 32'hEF157DE0 , 32'hF9D66158 , 32'hF8A526A8 , 32'hFC6A67A8 , 32'hFDDBEE4C , 32'hFC70BDF8 , 32'hF6668A10 , 32'h0DC32AF0 , 32'h09EE4C30 , 32'h0284DB40 , 32'hF4E21960 , 32'h06B4A280 , 32'h04080160 , 32'hFC56BE24 , 32'h0A52A280 , 32'h00565A7A , 32'h04CBBF70 , 32'hF8F0A0E0 , 32'h0851AAF0 , 32'h07833BB0 , 32'hFB303C90 , 32'hFDE9FC00 , 32'hF64E30A0 , 32'h02BF9FE8 , 32'hFEC4E428 , 32'h087568F0 , 32'hFB5EFF28 , 32'h070ED3D8 , 32'h0062228F , 32'h03FB12F4 , 32'hF9F20248 , 32'hF97A8690 , 32'hFEE6ADC0 , 32'h00C98645 , 32'h01B2CD30 , 32'hFFD37EAB , 32'hFFFF9E7C , 32'hFFFABB0E , 32'hFFFEA8F1 , 32'hFFFD154C , 32'h0000110E , 32'hFFFECCEA , 32'hFFFBA9E9 , 32'hFFFF0C4A , 32'hFFFA221E , 32'hFFFE0E38} , 
{32'hFFFB5568 , 32'hFFF8639C , 32'hFFFFF245 , 32'hFFFC53B4 , 32'hFFF70987 , 32'h00032C64 , 32'hFFF4F863 , 32'hFFFFF17C , 32'h00049C38 , 32'hFFFEA6E4 , 32'h00060F6B , 32'hFFFBAA2E , 32'h0000DED5 , 32'hFFFB0124 , 32'h00004F99 , 32'h00015CBD , 32'h0008D340 , 32'h0004B7D5 , 32'h0005EBCE , 32'h000335A4 , 32'h0004F230 , 32'hFFFD2445 , 32'hFFFDBB95 , 32'h00059FD6 , 32'h000C5027 , 32'h0002B884 , 32'h00042208 , 32'h00054DE6 , 32'hFFFE2C22 , 32'h00028D55 , 32'h000257ED , 32'hFFFADCCD , 32'h00053550 , 32'hFFF98762 , 32'h00086FF7 , 32'h0005BBB5 , 32'hFFFC1020 , 32'h00020B86 , 32'hFFFDB6AF , 32'hFFFE920A , 32'hFFFFE5B5 , 32'hFFFF6B96 , 32'hFFFCB5F4 , 32'h0003EABD , 32'hFFF99B75 , 32'h0007D733 , 32'hFFFFCE15 , 32'hFFFBD9EB , 32'h0001C7CB , 32'hFFF7E886 , 32'hFFFFA031 , 32'h0001A1D2 , 32'h0009E828 , 32'h0007B833 , 32'h0002CA93 , 32'hFFFDBA05 , 32'hFFFED0A7 , 32'h0001A1A0 , 32'h00006323 , 32'hFFFE5D90 , 32'h0005D7B4 , 32'hFFFDCAEE , 32'hFFFEE30A , 32'hFFFDAF69 , 32'h00024EAB , 32'hFFFE05D8 , 32'h0000F542 , 32'h00061EB5 , 32'h00022D3E , 32'h00013CB8 , 32'h0004C0EB , 32'h000BE03E , 32'hFFFEB723 , 32'h0001A6AE , 32'hFFFBEA29 , 32'hFFF26754 , 32'hFFF9B341 , 32'hFFF50452 , 32'h0000EDD4 , 32'hFFFD6E1E , 32'hFFF6594B , 32'hFFFF4F8E , 32'hFFFB28F3 , 32'h00027A83 , 32'hFFFF8C65 , 32'hFFFF6763 , 32'hFFF8DF61 , 32'hFFF7A7CC , 32'hFFFFC4ED , 32'hFFFD5707 , 32'hFFF83558 , 32'hFFEF76B5 , 32'hFFF9F4B9 , 32'h0004EF67 , 32'hFFFAFCF6 , 32'h00023840 , 32'h0008A548 , 32'h0000ADF0 , 32'h00009427 , 32'hFFFF5F63} , 
{32'hE0649660 , 32'h5C55D380 , 32'h4E24F800 , 32'h7FFFFFFF , 32'hF6515E70 , 32'hEC67C100 , 32'h0706BC30 , 32'hACF9D680 , 32'hCED3CD80 , 32'h143BEB40 , 32'h0C2DDBF0 , 32'hF66DA110 , 32'hF071A9A0 , 32'hFB6FE668 , 32'h117CD920 , 32'h3821CF00 , 32'hD4F14840 , 32'h0118524C , 32'hEF5FF960 , 32'hF95029D0 , 32'hE8DC8140 , 32'hDA0D2780 , 32'h0AB04B60 , 32'h177C2840 , 32'h3D743400 , 32'hE7B2FC20 , 32'h0C7B28E0 , 32'hFC7E7958 , 32'h1A3F3600 , 32'hFBF325C0 , 32'h0A12E860 , 32'hDD104480 , 32'hEF99AC20 , 32'hE7253020 , 32'hFC4DE2E0 , 32'h12C1C6C0 , 32'h03F0958C , 32'hF494E140 , 32'hF0A48C70 , 32'hEFDCF080 , 32'h02C89518 , 32'hF2C803A0 , 32'hFB905760 , 32'hFD19D4E0 , 32'hF521A9C0 , 32'h0BDE6E90 , 32'hFC48C424 , 32'h1B72E900 , 32'hFCC1DBE4 , 32'hF959E1F8 , 32'hFE749AE0 , 32'hFA1ADC20 , 32'hF30429E0 , 32'h027BDE2C , 32'h065CB6B8 , 32'hFE109440 , 32'hF34533A0 , 32'h09A653E0 , 32'h04449530 , 32'h008A56BB , 32'hFB80B360 , 32'h0904A850 , 32'hFD61DA50 , 32'h01376BE0 , 32'h04E68800 , 32'hFE064A54 , 32'h09BCA920 , 32'hFAD1D960 , 32'h050D06E8 , 32'hF5AC0200 , 32'hFFD84707 , 32'h09F99290 , 32'hF9267AD0 , 32'h075157B8 , 32'h07FE36C8 , 32'h06AE2A60 , 32'h07F3BE80 , 32'hEE0833E0 , 32'h0235117C , 32'h063B70F0 , 32'hFB594F00 , 32'h060C1A30 , 32'h067208D8 , 32'h06A18AB8 , 32'hFAC75190 , 32'hFD33241C , 32'h0A78A370 , 32'h0254E5F8 , 32'hFED03748 , 32'h007942F0 , 32'hFFFC1CDC , 32'h0003584D , 32'h00008B13 , 32'hFFFDD985 , 32'h0000A49F , 32'h000131C0 , 32'h00012FCD , 32'hFFFBD729 , 32'h00014FBF , 32'h00029AC2} , 
{32'h052DF268 , 32'hF19809E0 , 32'h006491E7 , 32'h096B8ED0 , 32'hE99CC2C0 , 32'hFD5B9060 , 32'hDEDDF680 , 32'hF1E1F880 , 32'h1A3A3920 , 32'hE5F086E0 , 32'h0C14D430 , 32'hFF1E3240 , 32'hF2910250 , 32'hF2B2A1D0 , 32'hFAA28CD8 , 32'hF56E53B0 , 32'hFE2DA6BC , 32'h01445B84 , 32'hEE573640 , 32'h06616700 , 32'h01DF19EC , 32'hF88CFD90 , 32'hF6326E20 , 32'h08A87250 , 32'h020C8530 , 32'hF7A169A0 , 32'h0218EC3C , 32'h029A4BBC , 32'hFF3BA1D0 , 32'hFB925FA8 , 32'hFEBBF07C , 32'hF37D6210 , 32'hF0440340 , 32'h03339FD8 , 32'h035B0958 , 32'hFC842258 , 32'hF4E032F0 , 32'h021E9074 , 32'h0EE6DA00 , 32'hFD10E558 , 32'h0D52AC80 , 32'hF1BEFB60 , 32'hFD5744D0 , 32'hF574C670 , 32'h07349AF8 , 32'h044C66D8 , 32'h16841C20 , 32'hF760AF90 , 32'h15530F60 , 32'h0B2EFB00 , 32'hEE6A9AE0 , 32'hFA95FB78 , 32'h037F7638 , 32'h002891A2 , 32'hFE52FFE8 , 32'hF1D8BD90 , 32'h042CBFA8 , 32'h07BB0118 , 32'hF4439030 , 32'h06F7E0D0 , 32'h051F0058 , 32'h0B5CC620 , 32'hF67692A0 , 32'hF1D59320 , 32'h04A5DF18 , 32'h00E5B400 , 32'h01EF74D4 , 32'h07C15D90 , 32'h0946DB30 , 32'h0189E9F4 , 32'hFEB10F6C , 32'h05822528 , 32'hF118CC20 , 32'h06270DA0 , 32'hFF95764C , 32'h0F003B80 , 32'h098D24F0 , 32'hF7FA1680 , 32'h0384B3C0 , 32'h0211FD24 , 32'h02A7C8A8 , 32'h068386A8 , 32'h01AA1D18 , 32'hFD0A7050 , 32'h0042DB35 , 32'hFE4D77E4 , 32'hFCF0C144 , 32'hFEE8E36C , 32'hFE0941A4 , 32'hFF8A867A , 32'hFFFFF850 , 32'h0004EDAD , 32'h00003E63 , 32'h0003E8C4 , 32'h0001B3E4 , 32'h0001DD53 , 32'h0002573B , 32'h000013D4 , 32'h0002AAE4 , 32'hFFFE8551} , 
{32'hFFFFA5C2 , 32'h00039E23 , 32'hFFFAEF55 , 32'h00027D12 , 32'h0002F15D , 32'hFFFE1CC0 , 32'hFFFFEB5D , 32'hFFFCDF7E , 32'hFFF65D0A , 32'hFFFDEC08 , 32'hFFFED33D , 32'hFFFFD913 , 32'hFFFBBB77 , 32'h0000390E , 32'hFFF5D6CB , 32'h0000F4DF , 32'h000CAE0C , 32'h0000C847 , 32'hFFF77488 , 32'h00063160 , 32'hFFF98EC9 , 32'h0005EA23 , 32'hFFFFA1CE , 32'hFFFF518D , 32'h000206E3 , 32'h0004E585 , 32'hFFFA865D , 32'h000250EE , 32'h00054630 , 32'hFFFF0D9E , 32'hFFF64274 , 32'h00037B54 , 32'h00028E65 , 32'hFFFE6991 , 32'h000008C2 , 32'hFFFFD6E4 , 32'hFFFFDE4F , 32'h000A1BED , 32'hFFFECC4D , 32'h00008E56 , 32'hFFFB7F75 , 32'h0004E842 , 32'h00011004 , 32'hFFFFB857 , 32'h0008A12F , 32'h000688AF , 32'h0008F464 , 32'h00041C3C , 32'hFFFD27E3 , 32'hFFF816CA , 32'hFFFD2BE1 , 32'h000C5239 , 32'hFFF8663F , 32'h0002F2BA , 32'hFFF7739D , 32'h0002B315 , 32'h000025C5 , 32'hFFF8ACE2 , 32'h000037DF , 32'h0004453E , 32'h000727DD , 32'hFFFE948A , 32'hFFFE2ADB , 32'h0001C440 , 32'h0002C4A6 , 32'h0002762A , 32'hFFFC36F6 , 32'hFFFE7690 , 32'h00041075 , 32'hFFFA8583 , 32'h000793E6 , 32'hFFFDF125 , 32'h0004C85C , 32'hFFF3DBFB , 32'h000142D4 , 32'hFFFDBFA0 , 32'hFFFEC622 , 32'h0002ADB7 , 32'hFFFD1B61 , 32'h00017BB5 , 32'hFFFF9813 , 32'h0003FA56 , 32'h000620D9 , 32'hFFFE1BAE , 32'h0000AC53 , 32'hFFFA54C2 , 32'hFFFDD71B , 32'hFFFB3066 , 32'hFFFC284B , 32'h00009BE6 , 32'h00034FA2 , 32'h0007E141 , 32'h000131F5 , 32'h00023E7A , 32'h00020BAF , 32'h0001652E , 32'h0009B7F7 , 32'h00002104 , 32'hFFFBFE50 , 32'hFFFDB3AB} , 
{32'h7FFFFFFF , 32'hEB80B720 , 32'hC4A08580 , 32'hDE3CECC0 , 32'h358FFBC0 , 32'hB07FF680 , 32'h04483D48 , 32'h262B3780 , 32'h3BCB6A00 , 32'h3804C100 , 32'h08AB4B30 , 32'hF3C07490 , 32'hF4239B60 , 32'hEF462AA0 , 32'h0FC578A0 , 32'hEF1B7420 , 32'hEE3B59A0 , 32'h0963BAF0 , 32'hC40ECAC0 , 32'hF1364040 , 32'hF58E95F0 , 32'h00CD80A1 , 32'hF5233260 , 32'hE4B316C0 , 32'h162D4400 , 32'hFEAD5DE4 , 32'h4A987980 , 32'h11A811C0 , 32'hF6254FC0 , 32'hD5CF7E40 , 32'h0BFDA4E0 , 32'h004F1714 , 32'hFA90C580 , 32'h08CD7530 , 32'h01EBB840 , 32'hED164200 , 32'hFF40568E , 32'hECF0A660 , 32'hEC861760 , 32'hEB256420 , 32'h00F57E60 , 32'hFDF301E8 , 32'h0208DB8C , 32'hF9831D58 , 32'h24B559C0 , 32'h07FB57B0 , 32'h05C8A648 , 32'h02645758 , 32'h0351E73C , 32'h09276640 , 32'h00E8B465 , 32'hFFC1860A , 32'hFC0E01E4 , 32'h00DC2C96 , 32'hFAD2CB30 , 32'h0AD00480 , 32'h0188F05C , 32'h0A2213A0 , 32'hF694B760 , 32'h0838B900 , 32'h02754EDC , 32'h0202E63C , 32'hFFA42A65 , 32'hFF6F91DC , 32'h08300C40 , 32'hFC15EB1C , 32'h11537B80 , 32'h00B1D491 , 32'h0AFD9EA0 , 32'hF86C86F8 , 32'h08C8B8D0 , 32'hF35EA960 , 32'h00425CB5 , 32'h04B607B0 , 32'h0440B0B0 , 32'h037C4D4C , 32'hFD5EDA44 , 32'h02B74E4C , 32'h0DA511A0 , 32'h09A2FE20 , 32'h054C1D38 , 32'hF8F5CBA8 , 32'h026D8768 , 32'h03C865E4 , 32'h03C134D4 , 32'h01A407C0 , 32'hFEB86BB0 , 32'hFFB10938 , 32'hFD2151BC , 32'hFF16EA4D , 32'h0000C4B3 , 32'h0003AA2E , 32'hFFFF9E93 , 32'h0002FD98 , 32'hFFFF3A48 , 32'h00008FBC , 32'h0002782D , 32'hFFFF49E0 , 32'h0003974F , 32'hFFFE5066} , 
{32'hB3315200 , 32'hC1523080 , 32'h2F979980 , 32'hB5B9A700 , 32'hAC2C2F80 , 32'hD8E291C0 , 32'hCC870440 , 32'hEACCDA60 , 32'h46B92D00 , 32'h53286600 , 32'h2C8C0B40 , 32'hF7A7B330 , 32'hFF4A018B , 32'h2F4B8D80 , 32'h1B63B540 , 32'h250C8380 , 32'h053EC9C0 , 32'hEB64F440 , 32'h366E1540 , 32'h0C82AE00 , 32'hFCD46818 , 32'h0423DB50 , 32'h142ACCE0 , 32'h14B78C60 , 32'hFCFC0224 , 32'hD8553480 , 32'h00E70177 , 32'hECF2CDA0 , 32'h001E9E06 , 32'hEBC5BF20 , 32'hF2BDFD90 , 32'h12439DA0 , 32'h063CE2A8 , 32'hF9C073F0 , 32'h0B5ABF10 , 32'h14AE7140 , 32'hFBF7D780 , 32'hEE46FF80 , 32'h04CFB078 , 32'h0BF27760 , 32'hE2F308E0 , 32'hFC873CBC , 32'h0B471040 , 32'hFB9FBAE0 , 32'h07CAC868 , 32'hECAA40C0 , 32'h00AF2F8A , 32'h0C1BB680 , 32'h0CC20260 , 32'hFF6AE8F9 , 32'h0ACACAD0 , 32'h06647C00 , 32'hFDD807A8 , 32'hF99D2C50 , 32'h062865C8 , 32'hF769B240 , 32'hFA844278 , 32'hFD372B28 , 32'h042075E8 , 32'hF4058540 , 32'hFC94E2C8 , 32'hF67C2F40 , 32'hF5C4C370 , 32'hFEBB1300 , 32'hFB83E740 , 32'hFC7D5EDC , 32'hF01F0AB0 , 32'h09B2BB10 , 32'h08BB30E0 , 32'h05C16898 , 32'h099602F0 , 32'h059CDA18 , 32'hFF7649E2 , 32'h03FDF16C , 32'h03EAC2A0 , 32'h05BAD1E0 , 32'hF724D6A0 , 32'hFEE49018 , 32'hF62EC670 , 32'h0390292C , 32'hFBFAC448 , 32'hFAE8B190 , 32'hF9791500 , 32'h00BDEA35 , 32'h02CCFDAC , 32'hFD5CDCFC , 32'h01446FF8 , 32'hFEFF0C60 , 32'h02473230 , 32'h02A58A28 , 32'hFFFFDEBE , 32'h0001EA2C , 32'h0000663C , 32'hFFF7F4A4 , 32'hFFFCCF5D , 32'hFFFA3B6C , 32'hFFFBF346 , 32'hFFFE4714 , 32'hFFFE386F , 32'hFFFF6F72} , 
{32'hDA9478C0 , 32'hF20B3F40 , 32'hB21D1C00 , 32'hEDA17BC0 , 32'h31431FC0 , 32'h01E9DCE4 , 32'hE793C760 , 32'h0DCF09F0 , 32'h235862C0 , 32'hF8769898 , 32'hF284E640 , 32'hF9EA9AE8 , 32'h07FDF438 , 32'hDB52D380 , 32'h08852340 , 32'h02243C08 , 32'hF9416990 , 32'hEF08F180 , 32'hDFC78F80 , 32'h094622A0 , 32'h00B224FB , 32'h154ECF80 , 32'h0789F5E0 , 32'hF1DFCDF0 , 32'h0E184F20 , 32'hF1243A20 , 32'h1D118DE0 , 32'hE80D2C00 , 32'h0CD1FB00 , 32'hF2241960 , 32'hF9A25A00 , 32'hD54FBE40 , 32'hFD3995E4 , 32'h0189EA98 , 32'hFF5EFB8F , 32'hFC43F4A0 , 32'h1EC37D20 , 32'hFC456ACC , 32'h03992738 , 32'hFADC8840 , 32'h1A8D9B40 , 32'h008BC613 , 32'h05F893B8 , 32'h14972120 , 32'hF84A0738 , 32'h064C65D8 , 32'hFFC0EC0C , 32'hFF8AE877 , 32'h0BE519D0 , 32'hFB47E448 , 32'hF3AE4E70 , 32'hFCC3AAD8 , 32'hF2C83890 , 32'hF4937050 , 32'hF524A810 , 32'h060CA0B0 , 32'h0ADB2180 , 32'hF3970150 , 32'hF2C51640 , 32'h091581E0 , 32'hF9507570 , 32'hF29E5840 , 32'hF6027880 , 32'hF2926000 , 32'h06393AF0 , 32'h02014744 , 32'h06F29098 , 32'hF8443628 , 32'hFB9B6848 , 32'hFE612668 , 32'h028BC58C , 32'hFFD1BEA0 , 32'h00DB3701 , 32'hF9F0F190 , 32'h12CAE000 , 32'hF9835E88 , 32'hFE1EF128 , 32'h0671FA30 , 32'h0167B12C , 32'hFD781D5C , 32'hF79855A0 , 32'h0B795A90 , 32'h00F25AA5 , 32'hFF6F8A9B , 32'h01811498 , 32'h0FC5FC60 , 32'h034FE890 , 32'hFFF3D3E5 , 32'h01AB34A8 , 32'hFFB4CAA6 , 32'h00027551 , 32'h0002DE4E , 32'hFFF9DDEF , 32'hFFFDB00A , 32'h0001D3E0 , 32'hFFFA4706 , 32'hFFFD4F6F , 32'h00035252 , 32'hFFF75D15 , 32'hFFFD4C45} , 
{32'h000344D3 , 32'h0000F6D8 , 32'hFFFCE355 , 32'hFFFD29FC , 32'hFFFFB543 , 32'hFFFA4AB8 , 32'h0003B59B , 32'h000531F5 , 32'hFFFEE4B6 , 32'hFFFB32BA , 32'hFFFF3A3A , 32'h00071D23 , 32'h00014C4B , 32'h000057E0 , 32'hFFFE1936 , 32'hFFF9D3B6 , 32'h00008601 , 32'hFFF99E7E , 32'h00028196 , 32'hFFFE428E , 32'h0004F5E9 , 32'h00035C32 , 32'hFFFEB324 , 32'h00009633 , 32'hFFFE7CF7 , 32'hFFFFDC3A , 32'h00077EFA , 32'hFFF91244 , 32'h00031D8C , 32'h000187B4 , 32'h0000B9E4 , 32'h0000DBCF , 32'h00024DB6 , 32'hFFFE9A2C , 32'hFFF9C915 , 32'h0001BE3F , 32'hFFF45813 , 32'h000215C7 , 32'hFFFF8D3B , 32'h0005FBB7 , 32'hFFFD22C6 , 32'hFFF7AD3B , 32'h00059522 , 32'h0001EE63 , 32'h0001A545 , 32'hFFFD4F4F , 32'hFFF8FB28 , 32'h0002DC62 , 32'hFFFA9521 , 32'h0001761F , 32'h00016339 , 32'hFFFBDEC2 , 32'hFFFEA8CB , 32'h000213B2 , 32'h0003860F , 32'hFFFF5F87 , 32'hFFFEB28D , 32'hFFFC1B19 , 32'hFFFF4E52 , 32'hFFF2EE7D , 32'h0002BCB8 , 32'hFFFE6308 , 32'hFFFFB7C5 , 32'hFFF329FC , 32'hFFFDB355 , 32'h0004EB4C , 32'hFFFC6579 , 32'h000503C6 , 32'h00003680 , 32'hFFFC2EFB , 32'hFFFF985A , 32'h0004697E , 32'hFFFCAE96 , 32'hFFFDF9F9 , 32'h000515CF , 32'h0008EBE5 , 32'hFFFB3729 , 32'h0001FF5B , 32'h00001DD3 , 32'h00027766 , 32'h0007E038 , 32'h0001BCF6 , 32'h0002491C , 32'hFFF9C5FA , 32'hFFFF9233 , 32'h00023D65 , 32'h0007EEBE , 32'hFFFD3C65 , 32'h0002A552 , 32'hFFFCF30C , 32'h000A54C8 , 32'h00006BE9 , 32'hFFFA5995 , 32'hFFFE482B , 32'hFFF60B10 , 32'h000228BF , 32'hFFFBD112 , 32'hFFFEFAD8 , 32'hFFF96C8A , 32'hFFFB6818} , 
{32'h00002F0B , 32'hFFFFD1FE , 32'h00002693 , 32'h000156F7 , 32'hFFFCEFCD , 32'hFFFAAA39 , 32'hFFFDF97E , 32'h0007FAB9 , 32'hFFEF6559 , 32'hFFF7DAC0 , 32'hFFFA6F1F , 32'h000407B9 , 32'hFFFC5270 , 32'h0001F1C5 , 32'hFFFEA77D , 32'hFFFFE0F2 , 32'hFFFE22C4 , 32'h00054C30 , 32'hFFF714A1 , 32'h000546FE , 32'hFFFF2647 , 32'hFFFC707F , 32'hFFFAFF9A , 32'hFFFC3A63 , 32'hFFFFFF78 , 32'h00029778 , 32'h00062A85 , 32'h00019C0B , 32'hFFF20944 , 32'hFFFD0659 , 32'h0001E838 , 32'hFFF6ED0F , 32'hFFFB3716 , 32'hFFFA2FBA , 32'hFFFE5FD8 , 32'h000251EA , 32'hFFFBC377 , 32'hFFFCB8E5 , 32'hFFFDEF6E , 32'hFFF8ED30 , 32'hFFFAF3E9 , 32'h00071F78 , 32'h0005D50F , 32'h00003897 , 32'h00025FFD , 32'h0003C323 , 32'hFFF9999F , 32'h000278DE , 32'hFFFED689 , 32'hFFFED6ED , 32'h00008DB8 , 32'h0008835E , 32'h0000EA5A , 32'hFFF976DC , 32'hFFFC923E , 32'hFFFE353F , 32'hFFF838C2 , 32'h0002DF9F , 32'h000341B0 , 32'h00002FE2 , 32'hFFFB8D4B , 32'hFFF943F8 , 32'hFFFDFA95 , 32'h000028AA , 32'h00032B1F , 32'h000AD14E , 32'h00033372 , 32'h000435A2 , 32'hFFF96762 , 32'h00020B11 , 32'h00089B4F , 32'hFFF68BE0 , 32'hFFFE7FD9 , 32'hFFFD9BF6 , 32'h00075C6A , 32'hFFF848FC , 32'h00040840 , 32'hFFFE512A , 32'hFFFB50E3 , 32'h00057F35 , 32'h00005AC3 , 32'hFFFA83FE , 32'h0005D44A , 32'h000CC297 , 32'h00036FFC , 32'h00080C1C , 32'hFFF5BF34 , 32'h00020FE6 , 32'hFFFAAE66 , 32'h000152F4 , 32'hFFFF8C0A , 32'h00021DBA , 32'hFFFD7CD6 , 32'hFFFEE82F , 32'hFFFE720A , 32'hFFFFED9B , 32'h00005851 , 32'h00059879 , 32'h00011072 , 32'h0001D3EA} , 
{32'h00084D79 , 32'hFFFD809D , 32'h0001324E , 32'hFFFD9BD2 , 32'h0002569D , 32'h0002B082 , 32'hFFFBFB0A , 32'hFFFC82A4 , 32'h00016344 , 32'hFFFB181F , 32'h00018ED0 , 32'hFFF6318D , 32'hFFFD8B5B , 32'h00049746 , 32'hFFFB8594 , 32'hFFFCAB91 , 32'hFFFF43B4 , 32'h0004BC9F , 32'hFFFE77D0 , 32'hFFFED379 , 32'hFFFFCF90 , 32'h00027A56 , 32'hFFFF5D03 , 32'hFFF9E70A , 32'h000255DD , 32'hFFFFA777 , 32'hFFFCDAA6 , 32'h0000AD03 , 32'h00059F43 , 32'h0007DC4E , 32'h00038FBC , 32'hFFFCF902 , 32'hFFFC8D8B , 32'h00026469 , 32'hFFFE23F7 , 32'h0000CB6F , 32'h000020AD , 32'h000206C7 , 32'h0001CFE5 , 32'h0007C3E4 , 32'h00029369 , 32'hFFFC7D16 , 32'h000272D8 , 32'hFFFD05AF , 32'h0000DF08 , 32'hFFFF9B3C , 32'hFFF80ACC , 32'h0003B5C3 , 32'hFFFDCC37 , 32'h00041192 , 32'h0003B03D , 32'hFFFDE599 , 32'h0002611B , 32'hFFFA81FF , 32'hFFFDEE71 , 32'h0000F6C0 , 32'h000301B6 , 32'h0000DA2A , 32'h00091084 , 32'hFFFA8CFD , 32'hFFF959F0 , 32'h000019E4 , 32'h0000FE49 , 32'h0002022E , 32'h000483B3 , 32'hFFFB5435 , 32'hFFF9E038 , 32'h0005DB7F , 32'h00073ACD , 32'hFFFF4B98 , 32'h00033674 , 32'h00011D4C , 32'h0000E0BB , 32'hFFFCC507 , 32'h00048629 , 32'h00014281 , 32'h000367D5 , 32'hFFF3F46A , 32'h00018837 , 32'h000517EE , 32'h00000429 , 32'h00019ACE , 32'hFFFE2482 , 32'hFFFAFEF2 , 32'h00012A81 , 32'h000047C4 , 32'hFFF64A4E , 32'h0004AB16 , 32'hFFFFDF2F , 32'hFFFFEF22 , 32'hFFFDE9E8 , 32'h0001F56A , 32'h00029D7E , 32'h000671E1 , 32'h00041AA8 , 32'h00056E3A , 32'h00050331 , 32'h000357FD , 32'hFFFB08CC , 32'hFFF90FB6} , 
{32'h36600240 , 32'hBF4C4A00 , 32'h09E735F0 , 32'hA4F1FA00 , 32'hA02E0B80 , 32'hFAD957F0 , 32'h17A8B0C0 , 32'h11F689E0 , 32'hCDDC7480 , 32'h07705B58 , 32'h1270FB80 , 32'hC5D5E600 , 32'hD3A81000 , 32'hDC22D8C0 , 32'hFBBFDCF0 , 32'h2FE33980 , 32'hFC562A30 , 32'hC3745200 , 32'hE862B200 , 32'hF3A09660 , 32'hD3724D80 , 32'hFF168427 , 32'hDCB6AE00 , 32'h103B9C80 , 32'hF04A0430 , 32'hE4F3B680 , 32'hFE7F4F8C , 32'h10C4F320 , 32'hFB249E20 , 32'h047BD9D0 , 32'h0007060C , 32'h02046FA4 , 32'hFEB1F9E0 , 32'hE3789400 , 32'hCD9898C0 , 32'h19A72480 , 32'h0C48AD70 , 32'hFD1C4714 , 32'h090D1220 , 32'h1D5E0460 , 32'h1EC1A020 , 32'hED13FE80 , 32'hFD94CDA8 , 32'hFBCA9CB0 , 32'hF27AAB70 , 32'hFE8134FC , 32'h14127800 , 32'h0DC24010 , 32'hF2658890 , 32'hE4B6BC40 , 32'hFF4A6F73 , 32'h06BAAD98 , 32'hEA789880 , 32'hEB315EE0 , 32'hFB758970 , 32'h0C6B59D0 , 32'h003C2E90 , 32'hF7949BD0 , 32'hFA368E20 , 32'h0590C620 , 32'hFAFDD870 , 32'h05F0B330 , 32'h05D08D38 , 32'hFEA324D4 , 32'h0764CDC8 , 32'hFA46CAE8 , 32'h01F9EEC0 , 32'h01C7463C , 32'h00174776 , 32'h014654E8 , 32'hF9A071D8 , 32'hF65655D0 , 32'h0564FDC0 , 32'h0B122C00 , 32'hF8E474B8 , 32'h00F4DF86 , 32'hFC904AD8 , 32'hFC5410A0 , 32'hF8C5CCC0 , 32'hFA30AC08 , 32'hF9FCEE00 , 32'h00B2E85E , 32'hF9548550 , 32'h009D799F , 32'h079E39D8 , 32'h03CB6B9C , 32'h01D73008 , 32'hFE9CB010 , 32'hFB9382D0 , 32'hFF3A17B0 , 32'hFFFEABE1 , 32'h00019B8B , 32'hFFFB5CB5 , 32'h0003A95E , 32'h000166D6 , 32'h0000EF47 , 32'h000061D3 , 32'h00011778 , 32'hFFFDB106 , 32'hFFFDC661} , 
{32'h00B54C98 , 32'h18811760 , 32'hFE4F4BD8 , 32'h019EE840 , 32'h130B8C60 , 32'h11E32120 , 32'h1BA3FAE0 , 32'hF7FAFCA0 , 32'h39CAC740 , 32'hFE4C3C50 , 32'hF7859000 , 32'hF7260D60 , 32'h135E21C0 , 32'h1E836200 , 32'h00B16B5E , 32'h1487F6E0 , 32'hD63C2800 , 32'h0C64DF60 , 32'h1322E5A0 , 32'hF3C68360 , 32'hFC5B38A0 , 32'hF65738F0 , 32'h046EA440 , 32'hEADB39E0 , 32'h0165C82C , 32'hF44F6860 , 32'hDF189940 , 32'h06A84080 , 32'hF6095600 , 32'hF7085A80 , 32'h16A78260 , 32'h04AF1278 , 32'h25868E40 , 32'hFAAC2A60 , 32'hFB98CA08 , 32'hE7E9BF20 , 32'hF0A8B8D0 , 32'h0453C838 , 32'h14200B00 , 32'h01C13B08 , 32'h05C4DDC8 , 32'hFA65F028 , 32'hFC1F6994 , 32'h081851F0 , 32'hE2398E60 , 32'hF6CEBA70 , 32'h01FF93F0 , 32'h060CDCC8 , 32'hF2BE3DC0 , 32'h1757DF40 , 32'h0D0DBE30 , 32'hF2714E30 , 32'hF7688C10 , 32'h069F2100 , 32'hF5C17A50 , 32'h1036BA20 , 32'h0915F560 , 32'hFF796C8B , 32'hFED2F108 , 32'h03A02360 , 32'h04993DE8 , 32'h039706B4 , 32'hF7B304B0 , 32'hF3494670 , 32'hF6875F20 , 32'hF9849EC0 , 32'hFC230B18 , 32'h0265DD60 , 32'h05CCACB0 , 32'hF50441E0 , 32'hFB9E7530 , 32'hEF2D9120 , 32'h0A520400 , 32'h05E7FBD8 , 32'h08A8C9A0 , 32'h0ACEABA0 , 32'hFE003454 , 32'h03046E78 , 32'h02C3ACC0 , 32'hF514B9A0 , 32'hFEE9F22C , 32'h0168F53C , 32'hFD1265B4 , 32'h03F0CA9C , 32'hFD366358 , 32'hF8269D70 , 32'h0354D2C4 , 32'h03B7E8AC , 32'h042BF8A8 , 32'hFE7EFABC , 32'hFFFD840C , 32'hFFF9F389 , 32'h0002559A , 32'h0000CEB6 , 32'h00025A20 , 32'hFFFF5732 , 32'h0004D6E6 , 32'h00038766 , 32'hFFFE632C , 32'hFFFF717E} , 
{32'hFFFA5410 , 32'h000501E1 , 32'hFFF9F559 , 32'hFFFF2B57 , 32'h0005DF4E , 32'h0001F7BE , 32'h0005ED03 , 32'hFFFC586E , 32'h0000262A , 32'h000023E2 , 32'hFFFDCBEF , 32'h00039CAF , 32'h00004F73 , 32'h0002AFF7 , 32'h00020C6F , 32'hFFFD6CDE , 32'h0007C109 , 32'hFFFBF481 , 32'hFFFF2997 , 32'hFFFF802D , 32'h00004645 , 32'h0000BDDB , 32'h0003DDF7 , 32'hFFFFE856 , 32'h00049D7F , 32'h0005C62D , 32'h000151F4 , 32'hFFFF0D76 , 32'hFFFF1A9F , 32'h00029E63 , 32'h00088A6F , 32'h0003B78F , 32'h00006D87 , 32'h0002390D , 32'hFFFCAE2C , 32'h00061982 , 32'hFFFF5590 , 32'hFFF7BD2D , 32'h0000CEBF , 32'h00063FAF , 32'h00041278 , 32'hFFFABBA3 , 32'hFFFFF517 , 32'h0003AA60 , 32'h0001F5FA , 32'hFFFE4C5F , 32'hFFFF5BD4 , 32'hFFFCFF6E , 32'hFFFA8E1D , 32'hFFF743DB , 32'hFFFDB267 , 32'hFFFCB720 , 32'hFFFD8453 , 32'hFFFEC359 , 32'h00003E00 , 32'h00046696 , 32'h00036DAC , 32'hFFFEF5A2 , 32'hFFFA8CCE , 32'h0002AE93 , 32'hFFFC0C4D , 32'h00064155 , 32'hFFF9F786 , 32'hFFFDFCF8 , 32'h00039574 , 32'hFFFEF5F4 , 32'hFFFEC6C8 , 32'hFFFF7824 , 32'h000058FB , 32'hFFFD5E4D , 32'hFFFE5D0A , 32'h00026F55 , 32'h00070312 , 32'h0001A451 , 32'h0003C5D6 , 32'h0008CF16 , 32'hFFFDEEE8 , 32'hFFF93B2B , 32'h000710D4 , 32'h00019449 , 32'hFFFCAAE3 , 32'h00033137 , 32'hFFFE4D64 , 32'h0004361A , 32'h0001765B , 32'hFFFE6FAC , 32'hFFFD260F , 32'hFFFB70AF , 32'hFFF5E4CE , 32'h00059C74 , 32'h000099FA , 32'hFFFE8106 , 32'h0001C32D , 32'hFFFD8882 , 32'hFFEF96CE , 32'h00007CC6 , 32'hFFFF3C56 , 32'hFFFF7BC1 , 32'h00044B78 , 32'hFFF89B6D} , 
{32'h6FE4A700 , 32'h7FFFFFFF , 32'h78C9A280 , 32'h351666C0 , 32'h43B5C980 , 32'hC8571F80 , 32'hF8095D90 , 32'h43207080 , 32'hF3AADF40 , 32'h0B07FD10 , 32'hD3275140 , 32'hE0CB7700 , 32'hCF5EDE40 , 32'h01DDBA90 , 32'hBEB26F00 , 32'h36F61180 , 32'h1EC171E0 , 32'h045FC9B8 , 32'h062ED670 , 32'h0199B720 , 32'h03855434 , 32'h1D40BB60 , 32'h1CB7DEA0 , 32'hD86CEE00 , 32'hF3632520 , 32'h29039080 , 32'h2986A400 , 32'hF3D3A330 , 32'hFE724AB0 , 32'h0C5EA1D0 , 32'h15F10B40 , 32'h0FD3C260 , 32'hDD5E3340 , 32'hFF3B94E9 , 32'hE36A4760 , 32'hE4678220 , 32'h1A347D00 , 32'h0BFDECB0 , 32'hF33D7CA0 , 32'hF810C6D8 , 32'hEF217660 , 32'hE513B400 , 32'hFE6CFCCC , 32'h022830A0 , 32'hF2377030 , 32'hEF8130E0 , 32'h0D55D220 , 32'h055779E0 , 32'hFFD4DBFE , 32'h006F5A17 , 32'hFD968F50 , 32'hF0FD1AA0 , 32'h0F62FDD0 , 32'hFB771380 , 32'h04729DA0 , 32'hFCE4CEB0 , 32'h01C80F04 , 32'hF88D4F98 , 32'hF8D80BF8 , 32'hFE490DB4 , 32'hF69C3BC0 , 32'hF35E1A60 , 32'hF7038150 , 32'h001C5A45 , 32'hF31C9900 , 32'h04CBF940 , 32'hFB2EE2B8 , 32'h0AC86130 , 32'h0420A550 , 32'h022A32B0 , 32'hFB26EFB0 , 32'hFEDE98BC , 32'hFD8E3530 , 32'h02F7ABD4 , 32'h04896578 , 32'hF8422280 , 32'hFE5E2CB4 , 32'h00035936 , 32'hF892CC88 , 32'h00B2DC38 , 32'hFF5FFDB6 , 32'hFF3EEE56 , 32'h04983588 , 32'h003B3A30 , 32'hF5777450 , 32'hF8722888 , 32'hFD715158 , 32'h04C11DD0 , 32'h0172E384 , 32'hFF48E7DF , 32'hFFFE2BD1 , 32'h00008B8D , 32'h0002088A , 32'hFFFCDD81 , 32'h000279EA , 32'h000042D1 , 32'hFFFDD243 , 32'hFFFD0C57 , 32'hFFFDF033 , 32'hFFFF0B53} , 
{32'hFAEE44D8 , 32'h061CE338 , 32'h0157EB00 , 32'h02B09240 , 32'hF0043CB0 , 32'h051B8898 , 32'h00CF1D87 , 32'hE76E2AC0 , 32'h01DA0F64 , 32'hF73EC650 , 32'hF426CAA0 , 32'hF561AFA0 , 32'hF4DE8630 , 32'hFF066A32 , 32'hFBF05A40 , 32'h005FDA4D , 32'h0EECE860 , 32'hF85C1668 , 32'h02CCC8B4 , 32'h037B052C , 32'h020012F8 , 32'hF733A180 , 32'h0C51A590 , 32'hF9131C58 , 32'hFECAF468 , 32'hFDE4DEE0 , 32'h0F6E0710 , 32'hF4C1D000 , 32'hFC6896E4 , 32'hF31668F0 , 32'hF88F9208 , 32'h05358D48 , 32'hFFAAA305 , 32'hFF40C443 , 32'h11B93F60 , 32'h048244C0 , 32'hF6192460 , 32'h135569A0 , 32'h053EE428 , 32'hF2C94920 , 32'h05143110 , 32'hFBDC3078 , 32'hF472F100 , 32'hFE1797FC , 32'hF75F7230 , 32'h05CF8FA8 , 32'h04C1AF48 , 32'h0C344ED0 , 32'hFA9925E8 , 32'hF9B2BE90 , 32'h0E43BDA0 , 32'hF6C2B3E0 , 32'hFFBFB751 , 32'h076D1F48 , 32'h089E88C0 , 32'h07B67B00 , 32'hFF15816F , 32'h067FE258 , 32'h04021910 , 32'hFE7CDF7C , 32'h03FC1A18 , 32'hFBC7F208 , 32'h05F1F708 , 32'h136FCDA0 , 32'hFAA861E0 , 32'h08F32DA0 , 32'h095F01B0 , 32'hF40284B0 , 32'h05C9B440 , 32'hF6DF21F0 , 32'hF9A56DD0 , 32'hF6699A40 , 32'h01269998 , 32'h08D7B8D0 , 32'hFEBD8214 , 32'hF11EBA50 , 32'h0005DF04 , 32'hFD915E44 , 32'h097BFB20 , 32'h07360380 , 32'hF92012D8 , 32'hFC29D850 , 32'hFD3CBE6C , 32'hFDD86CE4 , 32'h04BA4FB8 , 32'h0700C658 , 32'hFEA0B0A0 , 32'h02BD9D10 , 32'hFE2390D8 , 32'hFF370DAC , 32'hFFFEF7E1 , 32'hFFFACB39 , 32'h0005337C , 32'hFFF867AC , 32'h0000DC90 , 32'h00084501 , 32'hFFFEF064 , 32'h00027B13 , 32'h0001A9B1 , 32'h00016751} , 
{32'hFFFCCE9A , 32'hFFFBC649 , 32'hFFFDDE85 , 32'hFFFED6AD , 32'hFFF9AA53 , 32'h00023C4D , 32'h000A1ABC , 32'hFFFD60DA , 32'hFFF86114 , 32'hFFFB64C8 , 32'h00042A06 , 32'hFFF972B2 , 32'h00046502 , 32'h0000FB5B , 32'h00036F5B , 32'h0006200D , 32'h00002448 , 32'h00054428 , 32'hFFFA6395 , 32'h0005ACE1 , 32'h0000A7D7 , 32'hFFFB9A02 , 32'hFFFD2749 , 32'h0001F72D , 32'hFFFBD1E4 , 32'h00021F18 , 32'h0004571D , 32'hFFFB86AC , 32'hFFFE36FC , 32'h00016712 , 32'h00003B32 , 32'hFFFDF994 , 32'hFFFEAE2A , 32'hFFFD9EDF , 32'h00020EB6 , 32'hFFF5BF7C , 32'hFFF8ED36 , 32'h000326B1 , 32'hFFFF55E3 , 32'h0003D735 , 32'h00045981 , 32'hFFFFDD8F , 32'hFFFA37B2 , 32'hFFFFC800 , 32'h00027AAD , 32'h0004F332 , 32'h0001BFD6 , 32'h00005E7A , 32'h0004CDA3 , 32'hFFF610F8 , 32'hFFFD51BF , 32'h00018C65 , 32'hFFF9E918 , 32'hFFFD52BA , 32'h00019C4E , 32'hFFFE9DA4 , 32'h00040C5E , 32'h00087087 , 32'h0000BD36 , 32'h0002D05B , 32'hFFFEA7EB , 32'hFFF9A681 , 32'h00052CDC , 32'h0004E15F , 32'hFFFD3DC1 , 32'h00024E00 , 32'h0002ED07 , 32'hFFF9466D , 32'h0001D783 , 32'hFFFB537F , 32'h00009146 , 32'h0002CB77 , 32'hFFFAFE0C , 32'h00001C64 , 32'h000326CD , 32'h00059F20 , 32'hFFFC32CF , 32'hFFFFB204 , 32'hFFFCF0CD , 32'hFFFF0B0A , 32'h0003F193 , 32'h00035219 , 32'hFFFD3EDE , 32'h000290A7 , 32'h00040A81 , 32'hFFFF2027 , 32'h0007DBE2 , 32'hFFFE6D8B , 32'hFFFC3A1E , 32'h00064605 , 32'hFFFBE8F1 , 32'h00029491 , 32'h0005BB2B , 32'h00016688 , 32'hFFFEB5DD , 32'h0001F92A , 32'h0002D8A5 , 32'hFFFA17B3 , 32'h00006E32 , 32'hFFFE01A0} , 
{32'hDAA46240 , 32'h7FFFFFFF , 32'h56AB4100 , 32'h184BD220 , 32'h371BEC40 , 32'h06AADB70 , 32'hCF520E40 , 32'hB7952A80 , 32'h13504A60 , 32'h1FE267C0 , 32'hEE8C8960 , 32'hE2CF2CC0 , 32'h17B4A120 , 32'hD2D4A0C0 , 32'h1ADACCA0 , 32'h1E9D7440 , 32'hEF727500 , 32'hEFCF5280 , 32'h292C4E00 , 32'h09D8ADF0 , 32'hFE3BE5C4 , 32'hD0D0D780 , 32'hFC90223C , 32'h04FC6310 , 32'hE525A920 , 32'h02409074 , 32'h0F9BBDE0 , 32'h23EED140 , 32'h0C8BE7F0 , 32'hDA327500 , 32'hE99519C0 , 32'h114A82E0 , 32'hE788F8E0 , 32'hFA0150E0 , 32'hFA5422A0 , 32'hFA0EB770 , 32'h05B343B0 , 32'hF1DE6AA0 , 32'h116B37A0 , 32'hFD9175EC , 32'hE80EEA80 , 32'h3049A440 , 32'h05457038 , 32'hFA0759E8 , 32'h182BAB80 , 32'h15112DA0 , 32'h11663C80 , 32'hFB063AC8 , 32'hEA2474C0 , 32'hFB4EF338 , 32'h09996910 , 32'hFA66E2F8 , 32'h153D7840 , 32'h00DBDBFC , 32'hFFC7EC0F , 32'h072E9CF0 , 32'h0906CF60 , 32'hF6B263C0 , 32'hF5A2C580 , 32'h0B9C4790 , 32'hFD4FD028 , 32'hF82F2438 , 32'hE601CAE0 , 32'h0D9586D0 , 32'h05F527F0 , 32'hFD5992E8 , 32'h07C55058 , 32'h05BFAD20 , 32'hFC8B6438 , 32'h0C725E40 , 32'hFCDCDD80 , 32'hFAEC1AE8 , 32'h0239424C , 32'h07295748 , 32'hFF0026F4 , 32'h01672CC4 , 32'h04B3CE18 , 32'hFF93D16F , 32'hFBAD60A8 , 32'hF2F6F920 , 32'h00472F87 , 32'hFB7DA1E0 , 32'h04DCCA50 , 32'h02A9B268 , 32'h019CB060 , 32'hFDA6DEC8 , 32'h00F9AF29 , 32'hFEB90348 , 32'hFEAB3844 , 32'hFF583521 , 32'h00002D99 , 32'hFFFD6FE2 , 32'h0001B1F7 , 32'h00022394 , 32'hFFFF4B82 , 32'hFFFED3FC , 32'hFFFFF26F , 32'h00014B69 , 32'h0001B52D , 32'hFFFF6750} , 
{32'hE5F55360 , 32'hFF8A52EF , 32'hB15A8180 , 32'hF9144128 , 32'hFDC17F68 , 32'hEA4D4060 , 32'hFD5516AC , 32'hF1464A80 , 32'hDDFF0BC0 , 32'hEDCB5500 , 32'h1AD275C0 , 32'hF9ED97B8 , 32'h116075E0 , 32'hEA6FDF60 , 32'hF3A30F90 , 32'hF59C2810 , 32'hF4C0BA10 , 32'h04C39F20 , 32'h0FBA81A0 , 32'h060BA790 , 32'h1E58F580 , 32'hF41AFE20 , 32'hE90E13E0 , 32'hF806B670 , 32'hEDC4A3A0 , 32'h0759D458 , 32'hFF57432F , 32'hFC29C9FC , 32'h1256ED00 , 32'h15BC8900 , 32'h099896F0 , 32'h029BFC28 , 32'h0A78B010 , 32'hFD98B45C , 32'hEE4359A0 , 32'hFB673F90 , 32'h01FC77BC , 32'hFEA231B0 , 32'hFC3200FC , 32'h0E1B3F70 , 32'hF4374290 , 32'hE7573CC0 , 32'hE4568FC0 , 32'hE6B0EC20 , 32'h0009E7E3 , 32'hEDFE2300 , 32'hE5F47C20 , 32'h070E99F0 , 32'hFF89DF86 , 32'hFD2C1CE4 , 32'hF57640B0 , 32'h05B40A98 , 32'hFAF91A80 , 32'h0CA95E50 , 32'hF7355A20 , 32'hF1022640 , 32'h0BFA8080 , 32'h015CC7F8 , 32'hF7AEF290 , 32'hF6715320 , 32'hFEADD75C , 32'hF099BB30 , 32'h026DCBA0 , 32'hF9B886B8 , 32'hFCE51B94 , 32'hF36C8F40 , 32'hF7E3D4C0 , 32'hFA8F23C8 , 32'hFCEB8570 , 32'hF5123240 , 32'hFA1EC850 , 32'hFA5425B8 , 32'h04E76370 , 32'h04F7EC78 , 32'h00A5C40C , 32'h0001CC68 , 32'h0ADF0C90 , 32'h01098308 , 32'hF7030ED0 , 32'h04A40108 , 32'hF9FBD618 , 32'hF3420BA0 , 32'h05DF4358 , 32'h00CB610C , 32'hFCEA5F58 , 32'h0163D368 , 32'h022D48F0 , 32'h0348B838 , 32'hFE4427AC , 32'h00962306 , 32'hFFFF9DCF , 32'h00039FE4 , 32'hFFF9A5D0 , 32'hFFFB5F56 , 32'h00036ACA , 32'hFFFED2DC , 32'hFFFCAF29 , 32'hFFFEFE23 , 32'h0002C634 , 32'hFFFA7C3A} , 
{32'h0003DE28 , 32'hFFFD8F6A , 32'hFFF7881E , 32'h0007A6C6 , 32'hFFFF36BF , 32'hFFF5FFAA , 32'h0005728A , 32'hFFF8ECD4 , 32'hFFF6C88C , 32'hFFFD78B9 , 32'hFFFA83BC , 32'hFFFF4184 , 32'hFFFCE3EE , 32'h000723DB , 32'hFFFE36C5 , 32'h00041A9C , 32'hFFFDC5BE , 32'hFFFF545D , 32'hFFFFCF1D , 32'h0001B0A9 , 32'h0009219E , 32'hFFFAEC97 , 32'hFFFF7C00 , 32'hFFFF2298 , 32'h00039AE0 , 32'hFFFF25F5 , 32'h0003E2B2 , 32'hFFF9010E , 32'h0008AFEE , 32'h00082B6C , 32'hFFFE799F , 32'h00019A23 , 32'hFFFEE0D3 , 32'hFFFE6B58 , 32'hFFFDB0D8 , 32'hFFFE0326 , 32'hFFFF9572 , 32'hFFFCF76F , 32'h00044601 , 32'hFFFE0BEA , 32'h000743EB , 32'hFFFC5F88 , 32'hFFFDDDC2 , 32'hFFF7C462 , 32'h000205A8 , 32'h00002F90 , 32'h0004200A , 32'h0002602D , 32'hFFF6665F , 32'hFFFC72C8 , 32'hFFFC310F , 32'hFFFD35F5 , 32'h000345D3 , 32'hFFF94BA9 , 32'hFFFE31BF , 32'h0002BCAD , 32'hFFFBA9E5 , 32'hFFFC20B3 , 32'h00014EDE , 32'h000872BA , 32'hFFFCF98C , 32'h00044E2C , 32'h00009B6A , 32'hFFFE243F , 32'hFFFFC850 , 32'h0001B584 , 32'h0000DA9E , 32'hFFFA0451 , 32'hFFFCD6C9 , 32'h0000C391 , 32'hFFF75AB0 , 32'h0005C535 , 32'hFFFD4FFA , 32'hFFFAE15E , 32'h0001A3D4 , 32'h0001E63F , 32'hFFFB5CBE , 32'h00069DD4 , 32'h0001DB3F , 32'h0003D3C7 , 32'hFFF6A7E0 , 32'hFFFDE4A2 , 32'hFFFD3D0F , 32'h0006B968 , 32'hFFFBBDD0 , 32'h0003A6F6 , 32'hFFFC9C54 , 32'hFFFAFB51 , 32'h0001D08D , 32'hFFFA4600 , 32'h00021AF0 , 32'h00029447 , 32'h0007C979 , 32'hFFFF2E70 , 32'h0007652A , 32'hFFFD4E37 , 32'hFFFDB92C , 32'h0002E54E , 32'hFFFCA370 , 32'h0001F0EB} , 
{32'hDD5BE780 , 32'h134D18C0 , 32'h2B3CA200 , 32'hC86DCC00 , 32'hF1759F80 , 32'hFF55E76A , 32'h0737A318 , 32'hE934F1E0 , 32'h39C3EF80 , 32'hEF58E6C0 , 32'hFDD4C68C , 32'h11F2B140 , 32'hF65273D0 , 32'hFD7EA894 , 32'h06FFB830 , 32'hFBC69DB0 , 32'hECE18A60 , 32'hFD9BB578 , 32'hFB557AF0 , 32'h03C83A64 , 32'hF4FEBE80 , 32'h168E9A60 , 32'hF67F0BF0 , 32'h0C9009D0 , 32'h071AB068 , 32'h1B461120 , 32'h02530FD8 , 32'h00C35612 , 32'h0472EEC0 , 32'hEC8A7F20 , 32'h0AD26110 , 32'h077CAF50 , 32'h03D13DB4 , 32'hE6F61BE0 , 32'hF213D5A0 , 32'h0D620850 , 32'hFA91E720 , 32'hF2B54320 , 32'hFF7B1E86 , 32'hF95AC278 , 32'h06622A70 , 32'hF2E112B0 , 32'hF11BB160 , 32'hEA8AA7E0 , 32'hF8CC6758 , 32'hF66D8980 , 32'hFCBF97A8 , 32'hFF031AAA , 32'h02DAB4C4 , 32'h013D8D28 , 32'h00387CAE , 32'h02A81664 , 32'hFFD5A6E5 , 32'hF1A22300 , 32'hFBD966D8 , 32'h0180BA90 , 32'hF4384980 , 32'hFBBAED18 , 32'h081CCD90 , 32'h014FCEF0 , 32'h059A3B68 , 32'hF555F200 , 32'h062DEA88 , 32'h05F533B8 , 32'h0E97C110 , 32'h0E335BE0 , 32'hF9EE3680 , 32'h06E43E28 , 32'h023F0264 , 32'hFA71A648 , 32'hFBAD1520 , 32'hF913AC38 , 32'h07095768 , 32'h125589C0 , 32'h057406D0 , 32'h0106B37C , 32'hEF723C80 , 32'h089B1AD0 , 32'hFD9BD46C , 32'h00379102 , 32'h017015CC , 32'h08194770 , 32'h080AFBA0 , 32'hFBB55C58 , 32'hF53305B0 , 32'h036587B8 , 32'hFB849630 , 32'hFCD0131C , 32'hFFE1D790 , 32'hFFCA8FC9 , 32'h0003EA50 , 32'h00049B28 , 32'h0005D3C5 , 32'hFFFDCF03 , 32'hFFFA832D , 32'hFFFAF57C , 32'h00016108 , 32'h0000A966 , 32'h0001CA26 , 32'h0004C7E7} , 
{32'hCBB31940 , 32'h35B7B200 , 32'hED99F180 , 32'h184440E0 , 32'h34FEC180 , 32'hD6A3F180 , 32'hDC4E6980 , 32'h0895F530 , 32'hE85D9740 , 32'hC2B021C0 , 32'h0988AD30 , 32'h12896D00 , 32'h1AA6BA60 , 32'h2FA80A40 , 32'h12626E00 , 32'h17DA5B40 , 32'h1B7779C0 , 32'hF58CD4B0 , 32'h0B2FEBF0 , 32'hEC78FAA0 , 32'hF0C24D60 , 32'h00B44011 , 32'h1E05E360 , 32'hF24A2270 , 32'hECFE9FC0 , 32'hE6B161C0 , 32'h1D153F00 , 32'h35341640 , 32'hF2753B10 , 32'h1FCE1060 , 32'h01856A24 , 32'h05B86380 , 32'hFED77564 , 32'h2385D000 , 32'hF4B323A0 , 32'h106F0620 , 32'h15ECBA60 , 32'h10A498E0 , 32'hEBF05D40 , 32'h0D9B3DB0 , 32'h07067EE8 , 32'h0714CA98 , 32'h0B9BA2C0 , 32'hF50F8A80 , 32'h0BE85AE0 , 32'h0FDF8450 , 32'h026537F4 , 32'hF4512550 , 32'h0749B500 , 32'h07148AA8 , 32'h179C3740 , 32'h021B5AE8 , 32'hF27CC220 , 32'h0BB49E50 , 32'h0C6FF7E0 , 32'h09885030 , 32'hF4336E50 , 32'h053BCB90 , 32'h100EF460 , 32'hF63CDBB0 , 32'hF73ECF90 , 32'hFAB80320 , 32'h16035500 , 32'h05D82650 , 32'hF9E77578 , 32'h02F2AF90 , 32'hFDFFD824 , 32'h0F72A210 , 32'h00C50A3D , 32'hF9826DB0 , 32'h03EF7738 , 32'hFDE90420 , 32'h07B2CCF0 , 32'h0808AF10 , 32'h0C9B2920 , 32'hF967A7C8 , 32'hF53B7F60 , 32'h07BEF810 , 32'h0AD2BCF0 , 32'hF839AEE8 , 32'h02590880 , 32'h05DB8180 , 32'hFA1602B0 , 32'hFC6D9A0C , 32'hFE0E2E74 , 32'h00F916F3 , 32'h01DCD498 , 32'hFD73486C , 32'hFF694D8E , 32'hFFDF18CB , 32'hFFF6369D , 32'h00021671 , 32'h00020BB1 , 32'hFFFB427F , 32'hFFFFE9B9 , 32'h00007A4D , 32'h00007797 , 32'hFFFF3AFC , 32'h0002F298 , 32'hFFFDD9F0} , 
{32'h11AF9D60 , 32'hFCD1EBC8 , 32'h1B1E6EE0 , 32'hE40543A0 , 32'h000C1948 , 32'hD3D562C0 , 32'hE8423A80 , 32'h0EDB4520 , 32'hF9E8B8C8 , 32'hEC033BC0 , 32'hFD2E76B4 , 32'hD7170680 , 32'h0292C7FC , 32'hFF2DA50A , 32'hF2FFC410 , 32'h085F4600 , 32'h160C0DA0 , 32'h069C8A88 , 32'hFC3A7B9C , 32'h0EB46C50 , 32'h062E0058 , 32'hD860D300 , 32'h152F8B60 , 32'hFD444A2C , 32'h07436170 , 32'hFE4CA4C8 , 32'h09C3DD20 , 32'h017746D4 , 32'h0F4E27A0 , 32'hF13E88E0 , 32'h0ABEFEF0 , 32'hED986FA0 , 32'h20EBA880 , 32'hFF0BA44F , 32'h001944D5 , 32'h0B1438B0 , 32'h107B51C0 , 32'h000BF347 , 32'hFFCC89DF , 32'hFC7B9210 , 32'h140BE7C0 , 32'hF62C7FA0 , 32'hF4E28EB0 , 32'h02E91184 , 32'h07B3B688 , 32'h041666C8 , 32'h0DB3B3C0 , 32'hFD8C0FC8 , 32'hDED38840 , 32'h0C8C2A60 , 32'hEDE545A0 , 32'hF677B980 , 32'hED75E980 , 32'h01989030 , 32'hF3B5FBC0 , 32'hECC09BE0 , 32'hFA4BD6F8 , 32'h002A2418 , 32'h11299EA0 , 32'hF6A44430 , 32'hFD03C59C , 32'hF302FC50 , 32'hF7F7C8C0 , 32'h00ED2232 , 32'hFF2B5DA3 , 32'hFB58C7A8 , 32'hFFD18A76 , 32'hF8B2A160 , 32'h08162AF0 , 32'h0A361CB0 , 32'h120494C0 , 32'hFBB8C498 , 32'h11C475A0 , 32'h052317D0 , 32'hF47ADCF0 , 32'h04A4AF38 , 32'hF8987010 , 32'hFB3B6A88 , 32'h05FE28D0 , 32'h00C4074B , 32'h004C8317 , 32'hF95DF710 , 32'h061C9600 , 32'h05F7FC00 , 32'hFC9D72BC , 32'h06D0C250 , 32'h02613E14 , 32'h006B9E03 , 32'h029319FC , 32'hFF5C8225 , 32'hFFFBE80F , 32'hFFFDD660 , 32'h0000A559 , 32'h0001DB2D , 32'h00068B23 , 32'hFFFB84DB , 32'h0002CF96 , 32'hFFFF9156 , 32'hFFFE0002 , 32'hFFFEA5B4} , 
{32'hFFFD571A , 32'hFFFE82E3 , 32'h00023C82 , 32'h0005B8C9 , 32'h000115CF , 32'h00019FA6 , 32'hFFFF0A97 , 32'hFFFE29B2 , 32'h0005C008 , 32'h0007F1A9 , 32'h0001BFA0 , 32'h000366D6 , 32'h00069B8C , 32'h00012B87 , 32'h00096755 , 32'hFFFB25D4 , 32'h0007472E , 32'hFFFF6EED , 32'hFFFC574A , 32'h00049177 , 32'hFFFA211A , 32'h0003CCEA , 32'hFFFDAD38 , 32'h00034BF4 , 32'hFFFD2A83 , 32'hFFFEEDFE , 32'h0005AB65 , 32'h000D6D4A , 32'hFFFA2337 , 32'hFFFB7F20 , 32'hFFFCB8AF , 32'hFFFC3B62 , 32'hFFFC8EA6 , 32'h000168AC , 32'hFFFE8CB1 , 32'h0003F3BC , 32'hFFFF8A11 , 32'h0009C053 , 32'h00001DF4 , 32'h0003813B , 32'h0002B816 , 32'hFFFE33CB , 32'h00065DA1 , 32'h000540C1 , 32'h0002FC2B , 32'hFFFDE42B , 32'h0002E2C9 , 32'hFFFC4300 , 32'hFFF8E9EB , 32'h00082E5E , 32'h0003C377 , 32'hFFFA58BB , 32'hFFF78765 , 32'h00030823 , 32'h000008DC , 32'hFFF8C76A , 32'hFFFC4EDF , 32'h0002C7CB , 32'h00002037 , 32'hFFFB2B86 , 32'hFFFEA63D , 32'hFFFA9F97 , 32'h000106B9 , 32'hFFFB9C86 , 32'hFFFC2F29 , 32'h00041E00 , 32'h000053ED , 32'hFFFD1F06 , 32'h0003CAAB , 32'hFFFD335D , 32'hFFF80A1F , 32'hFFFD2E1F , 32'h000429DE , 32'h00011FBF , 32'h0000AFEC , 32'h0001F281 , 32'h00032288 , 32'hFFF5D1F6 , 32'hFFF8D156 , 32'hFFFCDCC8 , 32'h00027FA3 , 32'hFFFCF05C , 32'hFFFF00D8 , 32'h0007598E , 32'h00028C4B , 32'h00014B3E , 32'hFFF9E650 , 32'hFFFF5A87 , 32'hFFFD7CAA , 32'hFFFE3188 , 32'hFFFFB782 , 32'h00040E79 , 32'h00006A6A , 32'hFFFA39BD , 32'h00006244 , 32'hFFF9A818 , 32'h00029271 , 32'h0008A2C4 , 32'hFFFEBCA4 , 32'h00016103} , 
{32'h00085ED0 , 32'hFFFEB7C1 , 32'h00025F4F , 32'hFFFF3F28 , 32'hFFFFC707 , 32'h00063313 , 32'hFFFA6952 , 32'hFFFCE746 , 32'h0000D9F7 , 32'h000768CB , 32'hFFFF30EF , 32'hFFFF1B7B , 32'h0000B448 , 32'h000124F1 , 32'hFFF9DC7B , 32'hFFFF3080 , 32'hFFFBE75F , 32'h0004C9F3 , 32'h0001D4C6 , 32'hFFF7550F , 32'h00040FA3 , 32'h00049231 , 32'hFFFDBC76 , 32'h0006ECFB , 32'h0008F88F , 32'h0003715B , 32'hFFFC6915 , 32'hFFFCD84D , 32'h0007873A , 32'h00078481 , 32'hFFFB6E39 , 32'hFFFF9B74 , 32'hFFFE20AC , 32'h0008445F , 32'h00078426 , 32'hFFFE234D , 32'h00000B43 , 32'hFFFE0B2B , 32'h00028340 , 32'hFFFD4409 , 32'hFFFFC093 , 32'h0001E236 , 32'hFFFCA58F , 32'h00006E95 , 32'hFFFD0E63 , 32'h0000BA67 , 32'hFFFD29C3 , 32'hFFFD101E , 32'h0001FE26 , 32'hFFFD04AD , 32'hFFFAD38E , 32'h00033553 , 32'h0001CA57 , 32'hFFFBD911 , 32'h00008919 , 32'hFFFE3303 , 32'h00002E3D , 32'hFFF6C8D6 , 32'h00025CBB , 32'hFFFFD657 , 32'h00045638 , 32'h00009291 , 32'hFFFE22CE , 32'h0007DB63 , 32'h000474BD , 32'h00021DE1 , 32'hFFFF8DCB , 32'h0007C843 , 32'hFFFA1D09 , 32'hFFF8B537 , 32'hFFF73413 , 32'hFFFEB581 , 32'h00063F6B , 32'h00023645 , 32'h00031590 , 32'h0009E26C , 32'h00065EBA , 32'hFFF814EA , 32'h000518AC , 32'hFFFAA7B0 , 32'hFFFBBA58 , 32'h000AD271 , 32'h0002F0C9 , 32'hFFFE2559 , 32'hFFFEC1FC , 32'hFFFD488C , 32'hFFFED391 , 32'h0005CD1B , 32'hFFFAED01 , 32'hFFFF2E8B , 32'h0006BFAC , 32'hFFFF0AA9 , 32'hFFFB27D0 , 32'hFFF878AC , 32'hFFFBFC72 , 32'hFFF78DF9 , 32'h00034278 , 32'h000177B6 , 32'h000967B7 , 32'hFFFF9BF3} , 
{32'hEF7B2420 , 32'hD890D340 , 32'hD66B78C0 , 32'h70F1DD00 , 32'h99522500 , 32'h15A90320 , 32'hA560F100 , 32'hDB52ED80 , 32'hC23B0EC0 , 32'h2812DB40 , 32'hE24E2920 , 32'hCFECA1C0 , 32'h276A3E80 , 32'h0AF02270 , 32'hFA6EE730 , 32'hDC65B5C0 , 32'h070D41B8 , 32'h1C783520 , 32'h14A77640 , 32'hF50F6160 , 32'hE13F26A0 , 32'h235116C0 , 32'h0EA78830 , 32'h17D2AC40 , 32'h05CAB908 , 32'h29F5CFC0 , 32'hEF054980 , 32'h16FE1220 , 32'h089262C0 , 32'hF656BF90 , 32'hEFAFCA60 , 32'h11D9A920 , 32'h23403CC0 , 32'hEDE9BCA0 , 32'h03A824BC , 32'hF5125F20 , 32'h1E362700 , 32'h119415C0 , 32'hD8BE5BC0 , 32'h020BD6CC , 32'h0952CC40 , 32'h04D81980 , 32'h12ACE0E0 , 32'h0ED24490 , 32'hFFAB721F , 32'h117B8AA0 , 32'h110476C0 , 32'h11C0E120 , 32'h0074F31F , 32'h03447968 , 32'hF5DB5BF0 , 32'hE07C0700 , 32'hE6B34C20 , 32'h08772E70 , 32'hFA9573B0 , 32'hE4BCDCC0 , 32'h07711B48 , 32'h099A53A0 , 32'hFDA139CC , 32'hF3F1CF30 , 32'h09616D20 , 32'h008540C2 , 32'h0ED25EB0 , 32'h0923CC90 , 32'h04DE8970 , 32'h09353A00 , 32'hF7353560 , 32'h00EA0C1C , 32'h0AC27650 , 32'h021F51E8 , 32'hFFD3B63C , 32'h03573028 , 32'h08AA8B00 , 32'hFFE88959 , 32'hFC4963E4 , 32'h03B347B0 , 32'hFC2F02FC , 32'h054E80D0 , 32'h016A9AC0 , 32'hFFB24205 , 32'hFAFB3400 , 32'h07F601E8 , 32'h035D9EBC , 32'h003895DD , 32'h02B26EBC , 32'hFEB7DBAC , 32'h0157B350 , 32'h0066C211 , 32'hFFDD0BF4 , 32'h009A65F0 , 32'h0001D2C7 , 32'hFFFBEAC1 , 32'h0002E036 , 32'h0004665A , 32'hFFFFCF73 , 32'hFFFC9341 , 32'hFFFFAFF1 , 32'h00024A88 , 32'hFFFF715B , 32'h00005E4E} , 
{32'hFFF7EA20 , 32'hFFFCD805 , 32'h0005A6D8 , 32'hFFFC2A62 , 32'hFFFDA918 , 32'h0005CA54 , 32'hFFFA2B4A , 32'h00002518 , 32'hFFFD70B9 , 32'h0007555F , 32'h0001E2A6 , 32'h0004212B , 32'h000356EC , 32'h0003C7EA , 32'hFFFECFA3 , 32'h00041A9C , 32'h00045047 , 32'h00083226 , 32'hFFFC75DC , 32'h0004AB03 , 32'h00011F2D , 32'hFFFD5278 , 32'hFFFE3C62 , 32'h0005698F , 32'h00014DCB , 32'hFFFAF43B , 32'h0000228C , 32'h000122EC , 32'hFFFD1355 , 32'h0005C5CB , 32'hFFFF03FA , 32'h000209A0 , 32'hFFFE937F , 32'hFFF70D1F , 32'h000102B7 , 32'hFFFA66A4 , 32'h0007B66D , 32'hFFF9EB08 , 32'hFFF9ED3D , 32'h00032951 , 32'hFFF5921A , 32'h000641E9 , 32'h0009E31C , 32'h00061ADB , 32'h00023A46 , 32'hFFF9C62E , 32'h0009189C , 32'hFFFF0870 , 32'h00031C36 , 32'h00021DE1 , 32'h000464BC , 32'h00038803 , 32'h000337CF , 32'hFFF867D3 , 32'hFFFE5DDE , 32'hFFFF77DE , 32'hFFFF02B4 , 32'h0002ED25 , 32'h00035A39 , 32'hFFFB353D , 32'h0001F645 , 32'hFFFE6F9D , 32'hFFFC4DDE , 32'h0002A811 , 32'h00035F98 , 32'hFFFDE607 , 32'h00031AE5 , 32'hFFFB2135 , 32'hFFFF6AEA , 32'hFFFFACA1 , 32'hFFFFF5C4 , 32'hFFFFF523 , 32'h0000851C , 32'h0002CED7 , 32'h0001A46D , 32'h00034758 , 32'hFFFA1237 , 32'h000134E4 , 32'h0007C55B , 32'hFFFD1CF8 , 32'hFFFD937D , 32'hFFFE7852 , 32'h000B4294 , 32'hFFFCADB7 , 32'h000411C3 , 32'hFFF7459B , 32'hFFFC3C98 , 32'h0003208B , 32'hFFFBD1B2 , 32'h00041B8E , 32'h000608C2 , 32'h000ECF1D , 32'hFFFDFACD , 32'hFFF7ED63 , 32'h0000C043 , 32'h00050BDA , 32'h0006B53B , 32'hFFFA1468 , 32'hFFFDBB9C , 32'hFFFF1689} , 
{32'hD8614080 , 32'h09189E40 , 32'h1042D440 , 32'hE380F5E0 , 32'h211039C0 , 32'h33E0D000 , 32'hF96E4960 , 32'hE0BEFF20 , 32'h217F3EC0 , 32'hF599FE40 , 32'h175ED280 , 32'h0E34C890 , 32'hEC87B020 , 32'h112845E0 , 32'hE55ECFE0 , 32'hFAD79FA8 , 32'h01007894 , 32'hEC99E180 , 32'hEFAD1C20 , 32'hEFD076A0 , 32'h014ECF6C , 32'hF66CFB70 , 32'h2535CCC0 , 32'h0CBFBF00 , 32'hF3604160 , 32'hFC263E34 , 32'hE3250E20 , 32'hEF04FB40 , 32'hF55D10D0 , 32'hED5EB4A0 , 32'h171CA840 , 32'h0C413870 , 32'h0F704AA0 , 32'hF30A9670 , 32'hEDE1F900 , 32'hFD5BD4D4 , 32'h12486780 , 32'hF2AF19C0 , 32'hF3649400 , 32'hF7981DA0 , 32'h1068FB40 , 32'hFA7298E8 , 32'h07034A50 , 32'h012CBEA0 , 32'h0BC8E630 , 32'hFA3F4D98 , 32'h0D8484B0 , 32'hDA2D1640 , 32'hF60D9190 , 32'hF91DE4A0 , 32'hFE9C53F4 , 32'h0FD4E6D0 , 32'hF7DD56D0 , 32'hFB8237C8 , 32'h0D7ECAF0 , 32'hF9AD7AE8 , 32'h08DB9640 , 32'hF3000CE0 , 32'hFC51F13C , 32'h027E6218 , 32'h04B48A60 , 32'hEF460D40 , 32'hF1E46CB0 , 32'hFE79CCC0 , 32'h00177221 , 32'h06FB32C8 , 32'h027C8958 , 32'hFB0D57B0 , 32'h046B08A0 , 32'hF74F1840 , 32'h03539164 , 32'hFDA0535C , 32'hFF8F54C8 , 32'hFAA389C0 , 32'h040E8698 , 32'hEAB03D00 , 32'hFD201C5C , 32'hF66660E0 , 32'hFD0D8FAC , 32'hFCA7C100 , 32'hFFFBF01B , 32'h014C7EB8 , 32'h04F13210 , 32'h05D300E0 , 32'hFD8AC784 , 32'hFFFE5FC8 , 32'hF95C1550 , 32'h00A7402C , 32'h01402574 , 32'hFFA002EC , 32'h0002A4D7 , 32'hFFFFAED0 , 32'hFFFC6502 , 32'h000018AB , 32'hFFFEA7F8 , 32'h0007D425 , 32'hFFFFFE5B , 32'hFFFE9676 , 32'hFFFDAF43 , 32'h000545BB} , 
{32'h0000B526 , 32'hFFFFED84 , 32'hFFFC9BAC , 32'h00058DC4 , 32'hFFFDB4F2 , 32'hFFFDA72C , 32'h0003242D , 32'h0005B828 , 32'h00044DAF , 32'h0002A9F9 , 32'h000024B3 , 32'hFFFC3FCA , 32'hFFFEAB94 , 32'hFFFB3670 , 32'h00022F51 , 32'h000068AD , 32'h0000CA5A , 32'h0004D614 , 32'hFFF95A35 , 32'h00008AE4 , 32'h0004A13A , 32'h00005915 , 32'h0007914E , 32'h0001023B , 32'h0000F86B , 32'h0005903F , 32'h00025F71 , 32'h0003A541 , 32'hFFF6DB08 , 32'hFFFFE6F3 , 32'h0002F04C , 32'hFFFE3674 , 32'hFFFB9CD6 , 32'hFFFA0E72 , 32'hFFF51D7F , 32'h0009AAD4 , 32'h0004A1BF , 32'h0009B6B3 , 32'h0005EA62 , 32'hFFFE201C , 32'hFFFC652F , 32'h00071963 , 32'hFFFECB28 , 32'hFFFAE08B , 32'h0004016B , 32'hFFFA8DCF , 32'h0000C6B3 , 32'h0007630E , 32'h000608CB , 32'h00031A2A , 32'h0004C139 , 32'hFFFA4776 , 32'h0003B842 , 32'hFFFF0417 , 32'hFFF987C2 , 32'h0005CE1D , 32'h0006EBC0 , 32'h00017968 , 32'hFFF7E323 , 32'h0001B320 , 32'hFFF9689A , 32'hFFFDD2FE , 32'hFFFCA220 , 32'h0006A476 , 32'hFFFEBC8A , 32'hFFFAA6A6 , 32'h0004B1AA , 32'hFFFFFA7F , 32'h0000E72C , 32'h00039622 , 32'h00053775 , 32'hFFFA5625 , 32'hFFFD183F , 32'h0001CB01 , 32'h00022F43 , 32'hFFFD8316 , 32'h00068AFB , 32'hFFFA3523 , 32'h00046091 , 32'h00006AED , 32'hFFFEA4C0 , 32'hFFFA1C2B , 32'hFFFEDA5D , 32'hFFFAD01F , 32'hFFFEEE3F , 32'hFFFE78CC , 32'hFFFAC5FC , 32'h0007F054 , 32'hFFFBCDE8 , 32'h00013911 , 32'hFFFB8893 , 32'hFFFC7101 , 32'hFFF95892 , 32'h0000B2BB , 32'hFFFF5853 , 32'hFFFFD402 , 32'h00041020 , 32'hFFFDE38B , 32'hFFFE7C0A , 32'hFFFD3A95} , 
{32'hE41EB760 , 32'hF3EB9B50 , 32'hD1CC3040 , 32'h25019900 , 32'h35F95980 , 32'h117FBDC0 , 32'hF203B5F0 , 32'h07D2C798 , 32'hD96B2D80 , 32'hFFAD372C , 32'hF36D62C0 , 32'h198888C0 , 32'hF60DF400 , 32'h10713640 , 32'hEA050180 , 32'hF71B8A90 , 32'hE0B68020 , 32'hF90DB898 , 32'h1DFBCD00 , 32'h0B5536A0 , 32'hE5F23160 , 32'hF49A9810 , 32'h066D8570 , 32'h1435E980 , 32'h199799C0 , 32'hF245AA90 , 32'hF676C540 , 32'hFD9CC360 , 32'h038B2608 , 32'hF5224E80 , 32'h33941040 , 32'h02441D30 , 32'hF4AB3210 , 32'hFFE32D93 , 32'hF4E3CC70 , 32'hF4995FD0 , 32'h17DB2FC0 , 32'h0CECF070 , 32'h0EE32720 , 32'h04F124B0 , 32'h08C9C340 , 32'h0FD10120 , 32'h01C45604 , 32'h0F6C5D00 , 32'hFBDBDFF8 , 32'h08B7CFC0 , 32'h0D9B69A0 , 32'h0223D81C , 32'h009436B8 , 32'hED619180 , 32'hFF12B78E , 32'h045F1AD0 , 32'h094B0DA0 , 32'hFFAC20BD , 32'h12065720 , 32'h0C2D87B0 , 32'h0C0B6510 , 32'hFDE39818 , 32'hF3E07350 , 32'h054628B0 , 32'h0B2AA9D0 , 32'hFB24D168 , 32'hFC47FB8C , 32'hFA461028 , 32'hF7767520 , 32'hFAC096F0 , 32'hF9B97AE0 , 32'h100D35C0 , 32'h0262745C , 32'h02D57330 , 32'hE839DF00 , 32'hFB259398 , 32'hFF723599 , 32'h002DFA8B , 32'hF7218520 , 32'h0D33A720 , 32'hF662ABA0 , 32'h02C3D1B8 , 32'h0C7A0310 , 32'h0A15F7C0 , 32'hF2A30780 , 32'h00866290 , 32'h06C73B78 , 32'h03553E44 , 32'h04A78658 , 32'h02C467A4 , 32'hF5259230 , 32'hFDEC0408 , 32'h071B9580 , 32'h00AC2A94 , 32'h00022F0A , 32'h0006F81D , 32'h0003F3DA , 32'hFFFA3237 , 32'hFFFE0C5D , 32'hFFFD932D , 32'h00071861 , 32'hFFFE9E11 , 32'h00030BAD , 32'hFFFCDC2C} , 
{32'h032ED5E8 , 32'h03188490 , 32'h02DE0768 , 32'h02DB5FB4 , 32'h05D3DBF8 , 32'h07A4F390 , 32'h02CFEB10 , 32'h00C73920 , 32'hFEBC106C , 32'hFFCBF48F , 32'hFF34B9D2 , 32'h0211C950 , 32'hFF9F5402 , 32'h014E3FAC , 32'h0385E41C , 32'h034D80D0 , 32'h039D1684 , 32'hFE727A40 , 32'hF849F508 , 32'h051F90E8 , 32'hFE5AFCE8 , 32'hFBA1B6B8 , 32'hFCCEF7D0 , 32'hFD902A28 , 32'h03C2AFEC , 32'hFFB21426 , 32'h023BA4FC , 32'h028E2F3C , 32'h011EE65C , 32'hFBF23270 , 32'hFB6BC7F0 , 32'hFE7E3FEC , 32'h04263260 , 32'hFDD187C0 , 32'hFC10ED24 , 32'hFEA7BA80 , 32'hFFA803F9 , 32'h012F5144 , 32'h00E6D48C , 32'h0110A158 , 32'h0269220C , 32'h00E7484F , 32'h03CDBF8C , 32'hFC4BCFD0 , 32'hFD5389DC , 32'h04051D00 , 32'hFF3F8822 , 32'h033CE220 , 32'h00D5937E , 32'hFD92EA5C , 32'hFEDE38F0 , 32'hFFFB795A , 32'h00E8042F , 32'hFF62E024 , 32'hFEB0C338 , 32'hFE9B9FEC , 32'hFDA106F8 , 32'h01381874 , 32'hFF73B08F , 32'hFF52EAD3 , 32'h00EE33E6 , 32'h05516E38 , 32'hFF94F114 , 32'h006235FA , 32'h026EABF0 , 32'h05146538 , 32'hFAF70930 , 32'h03290EA0 , 32'h01B3AFC4 , 32'h025009F8 , 32'h00C0CC17 , 32'hFEAE4628 , 32'hFDEA750C , 32'hFF4372A7 , 32'hFBFA7700 , 32'hFE35206C , 32'hFD34787C , 32'hFD4AE8DC , 32'hFF59AAD4 , 32'hFF6CE1E4 , 32'h037CEA3C , 32'hFD53B744 , 32'h012514E4 , 32'hFD5A5324 , 32'hFFC6B6FB , 32'h01BCE0E8 , 32'hFCB35CA4 , 32'hFEDFA9CC , 32'hFE945E00 , 32'hFFC63D7A , 32'hFFFFFBC6 , 32'h0002A9EA , 32'hFFF81504 , 32'h00021367 , 32'h00053311 , 32'hFFF9FBBB , 32'hFFFB934D , 32'hFFFF8FC2 , 32'hFFFEC2C9 , 32'h000139CE} , 
{32'hFFFF07A7 , 32'hFFFF18F9 , 32'h000019BC , 32'h0006A15C , 32'h0005AEDF , 32'hFFFD66D0 , 32'h0002952F , 32'hFFFBDC5D , 32'h00039C44 , 32'hFFFAD311 , 32'h0003848A , 32'h00036101 , 32'h00036D96 , 32'hFFFBB6ED , 32'h000589FE , 32'h00003B17 , 32'h0001E6CF , 32'h000023E4 , 32'h00051585 , 32'hFFFCE233 , 32'hFFFE842A , 32'h0000BE0B , 32'h0002BC2B , 32'hFFFE6D24 , 32'h0001A6AC , 32'hFFFD7B7C , 32'hFFFE2BA1 , 32'h00004645 , 32'h0001E648 , 32'hFFFF2A4C , 32'hFFF9810A , 32'h0001A288 , 32'h00048503 , 32'h00025EEC , 32'hFFF76387 , 32'h0007098B , 32'h00004752 , 32'hFFFE7EE9 , 32'hFFF28B2C , 32'h000705A7 , 32'h00088D06 , 32'h00035E3B , 32'h0001FAB3 , 32'hFFFB3B7A , 32'hFFFBC32D , 32'hFFFD5351 , 32'h000002BF , 32'h000529BF , 32'h00037735 , 32'h00054922 , 32'hFFFF43DB , 32'h0004438C , 32'hFFFA4FBF , 32'h000168FE , 32'h0006B6E2 , 32'hFFF8A09F , 32'h000479F8 , 32'h00004016 , 32'h00007154 , 32'h0001F889 , 32'hFFFF2EFD , 32'hFFFF93A4 , 32'h000729A0 , 32'hFFFFFBD5 , 32'hFFF81510 , 32'h0006FFB5 , 32'h00012C52 , 32'hFFFCA515 , 32'h000756FA , 32'hFFFA711F , 32'hFFFB8E1F , 32'h00013F3C , 32'h000A07E0 , 32'hFFFA706A , 32'h000698E7 , 32'hFFFC1003 , 32'hFFF94D72 , 32'hFFFE47BB , 32'h00013708 , 32'hFFF9B0BB , 32'h000954A3 , 32'hFFFEF6B7 , 32'h0002BD40 , 32'h000C4454 , 32'hFFFDDF57 , 32'hFFFB8CEC , 32'h0001456F , 32'h0000751E , 32'h000142D9 , 32'hFFFFD389 , 32'hFFF95E32 , 32'h0001C5D6 , 32'h000191A7 , 32'hFFFC6F85 , 32'hFFFE6CAC , 32'hFFFA6E89 , 32'hFFFFA559 , 32'h00003E77 , 32'h0003ED5C , 32'hFFFA352E} , 
{32'h00076394 , 32'hFFFF0EE1 , 32'hFFF8AB6C , 32'hFFFD65D0 , 32'hFFF62D29 , 32'h0008F740 , 32'hFFFD14E9 , 32'h0000C6DB , 32'hFFFA548F , 32'hFFFC80F4 , 32'hFFFDAF13 , 32'h0001640C , 32'hFFFFEAF9 , 32'hFFFD8FE1 , 32'h0002116B , 32'hFFFDF576 , 32'h0005B7C9 , 32'h000578F5 , 32'hFFF965F9 , 32'hFFFCAB99 , 32'h00069324 , 32'h000AAAB2 , 32'hFFFF4007 , 32'hFFFC0942 , 32'hFFFD12D7 , 32'hFFF57D84 , 32'hFFFD2E98 , 32'hFFFAFE02 , 32'hFFFC0C21 , 32'h00000744 , 32'h000154C3 , 32'hFFFEE717 , 32'h00046581 , 32'hFFFE7834 , 32'hFFFA30AC , 32'hFFFBEFF2 , 32'hFFFEB3A7 , 32'h00075D57 , 32'h0002124C , 32'h0005C324 , 32'hFFFE246A , 32'h0002FC0E , 32'hFFFCC0AF , 32'hFFF82640 , 32'h000192B5 , 32'hFFFCF12F , 32'hFFFE0765 , 32'hFFFB5BD1 , 32'hFFFF0617 , 32'h000A2CDE , 32'h00014F8B , 32'h0005CB85 , 32'h0001C232 , 32'h0001CA0F , 32'hFFF9D62E , 32'h0003CB82 , 32'hFFFE2CE4 , 32'h00015769 , 32'hFFFF38BB , 32'hFFFE4F8E , 32'h0000D376 , 32'h0004A0E1 , 32'hFFFD0F52 , 32'h00060F13 , 32'h00008564 , 32'h0003E815 , 32'h00027F09 , 32'h0000D9EC , 32'hFFFD0CC8 , 32'hFFFF1DEA , 32'h00052773 , 32'h0004B94E , 32'hFFFEB219 , 32'hFFF5E2C6 , 32'h00048170 , 32'h00072C20 , 32'h00040A24 , 32'hFFFD0DF2 , 32'h00082654 , 32'hFFF7F1BB , 32'hFFFFFB05 , 32'hFFFC01D7 , 32'hFFFF835E , 32'hFFF1B63A , 32'hFFFEDDCB , 32'h00018160 , 32'hFFFBAC8A , 32'h00048610 , 32'hFFF3B6C3 , 32'hFFFAEBD3 , 32'h00069BAC , 32'hFFFFB23A , 32'hFFFE87ED , 32'hFFFDA06E , 32'h00042A18 , 32'hFFFD3A52 , 32'hFFF8CE36 , 32'hFFFC712F , 32'hFFFB5A5A , 32'hFFFC6787} , 
{32'hFFFA69ED , 32'h00085056 , 32'hFFFA3AF1 , 32'h000045ED , 32'h0002C6F2 , 32'h00022F14 , 32'h00066EE9 , 32'hFFF6C96A , 32'hFFFF9FD5 , 32'h0001475D , 32'hFFF97AD4 , 32'hFFFC86A5 , 32'hFFFE8AF7 , 32'h0001E846 , 32'h000274DC , 32'hFFFAB16F , 32'hFFFE603F , 32'hFFFDB249 , 32'h0002C0C5 , 32'h00047D53 , 32'h00025FDC , 32'hFFF7EB9C , 32'h00034FAE , 32'hFFFBE969 , 32'h0002E885 , 32'h0001A873 , 32'hFFFFB4F5 , 32'h0004F019 , 32'hFFFBF9E7 , 32'hFFFD9057 , 32'hFFFE1032 , 32'h0001EF52 , 32'hFFFC4301 , 32'h0003B260 , 32'hFFFFC0AF , 32'h00027D34 , 32'hFFFF93A7 , 32'h0006800C , 32'h0002EB00 , 32'hFFFE6FB7 , 32'h0000D555 , 32'h00020BF5 , 32'hFFFFE1D2 , 32'h00039EAB , 32'h00031557 , 32'hFFFA33A2 , 32'hFFFD4655 , 32'h000027A5 , 32'hFFFE52ED , 32'hFFFD2755 , 32'h00058960 , 32'hFFFFABB2 , 32'hFFFD55EE , 32'hFFFCCDF4 , 32'hFFFC77EC , 32'h00095766 , 32'h00005349 , 32'h0002F1A3 , 32'hFFFDBD91 , 32'hFFFCFBC5 , 32'hFFFB11B6 , 32'hFFFDA0F2 , 32'h00034694 , 32'h0000DC60 , 32'hFFFEF972 , 32'hFFFFE6FD , 32'hFFFC86A0 , 32'hFFFF5800 , 32'h00026A71 , 32'h00045301 , 32'hFFF8F221 , 32'h00005736 , 32'hFFFD9DEC , 32'hFFF9F259 , 32'h00029743 , 32'h00023B55 , 32'hFFFB560B , 32'hFFFF11BA , 32'h000787E5 , 32'h00087ABB , 32'hFFF73225 , 32'hFFFC63FA , 32'hFFFDE893 , 32'h0004EB71 , 32'hFFFF3656 , 32'h00039201 , 32'hFFFB816A , 32'hFFF02A65 , 32'h0001D4D2 , 32'hFFF9A33B , 32'hFFFE29F3 , 32'hFFFAA7F5 , 32'h0002083D , 32'hFFFE68AD , 32'hFFFACD42 , 32'h000895A3 , 32'h0005B721 , 32'hFFF9DAD8 , 32'hFFF8233C , 32'hFFFF9824} , 
{32'h0004D8D1 , 32'h000A6C31 , 32'h000AE784 , 32'h000227D9 , 32'h0002E5DE , 32'h00025C2B , 32'h0004C978 , 32'hFFFCF2ED , 32'hFFF9F2DB , 32'hFFF7D031 , 32'hFFFCAC2A , 32'hFFFF975D , 32'h00091CDA , 32'h0003550E , 32'h00034771 , 32'hFFFFD02D , 32'hFFF88D29 , 32'hFFFD4123 , 32'hFFFD2114 , 32'h00063D0E , 32'h0003EAAA , 32'h00051DBA , 32'h0001EF4D , 32'h0002505D , 32'h00006181 , 32'hFFFFA611 , 32'hFFF727D6 , 32'h00024717 , 32'hFFFEA867 , 32'hFFFF6476 , 32'h00074EBF , 32'h0003DC15 , 32'hFFFDF88C , 32'h000152CF , 32'hFFFD9052 , 32'hFFFE936D , 32'hFFFD9CFF , 32'h0005D041 , 32'hFFFC6D0C , 32'hFFF8CF1C , 32'h00034E9B , 32'h00026206 , 32'h0002F5E1 , 32'h000448AC , 32'h0000EBFA , 32'hFFF5E94B , 32'h0004466E , 32'h0007C8B9 , 32'h0001747B , 32'hFFF8974F , 32'h0004161F , 32'h00037007 , 32'h0001525C , 32'hFFFED457 , 32'hFFF9FD35 , 32'hFFFEB95F , 32'h0002F7CB , 32'h000A650F , 32'h00011E51 , 32'h0004DA40 , 32'hFFFC16A5 , 32'h0004BD32 , 32'h0004C11B , 32'h00085416 , 32'h00054C05 , 32'h000105E3 , 32'h0000D365 , 32'h00056767 , 32'hFFFE9CCF , 32'hFFF5F265 , 32'hFFFD2E83 , 32'hFFFD2ECA , 32'h00077FEB , 32'h00030C14 , 32'hFFFFA60F , 32'h0005321D , 32'hFFFB494F , 32'hFFF9E452 , 32'hFFFD1406 , 32'hFFFE7E3B , 32'h000074CB , 32'hFFFE887F , 32'hFFFECFD3 , 32'hFFFE8AB6 , 32'hFFFDCFF6 , 32'h0001C9D7 , 32'h0002B761 , 32'h0003518E , 32'hFFFD2A77 , 32'hFFFF4B16 , 32'h00032EF8 , 32'hFFF7D809 , 32'h00026D0B , 32'hFFFD7176 , 32'h00037C93 , 32'h00023E70 , 32'h0005E67A , 32'h000438C5 , 32'h000164FE , 32'hFFFCD36B} , 
{32'hF7EAD570 , 32'h188BF1E0 , 32'h22954400 , 32'hD799B4C0 , 32'h1996E280 , 32'h1E0AE700 , 32'h183F70A0 , 32'hE1349760 , 32'h25002AC0 , 32'hF1A2BE20 , 32'h3F0CAB00 , 32'hDE2206C0 , 32'hED74FF40 , 32'h1C5BE7A0 , 32'hFCACC848 , 32'h181A1540 , 32'hD1854980 , 32'hFF3B2390 , 32'hEF633260 , 32'h03DC98BC , 32'hF833FA90 , 32'hF22CDA70 , 32'h074C8530 , 32'h0E262830 , 32'hF96E6040 , 32'h29F14880 , 32'hFC38CBA4 , 32'hEA3483C0 , 32'hE95E4840 , 32'h14A49920 , 32'h1917CD80 , 32'h0954A0A0 , 32'h0D9C6A10 , 32'h11BD1460 , 32'hF13621B0 , 32'h0E79DBD0 , 32'h0D7BA630 , 32'h00DCE25C , 32'h0ACCC4E0 , 32'hFD0AB480 , 32'h02BEE0B8 , 32'hFF6E8858 , 32'hFFE81744 , 32'hE86E5920 , 32'hF7067530 , 32'hEB4DD520 , 32'h06347360 , 32'h0A72BDB0 , 32'h0FB12E60 , 32'hF7B7FF50 , 32'hED1ED700 , 32'h0E0C98B0 , 32'h13AA5240 , 32'h0F8E3BA0 , 32'h096A9BC0 , 32'hFC9745A4 , 32'hFD6C5C28 , 32'h0068CB4E , 32'h145F4A00 , 32'h0F9D7650 , 32'hF3D1EFA0 , 32'hE57A12E0 , 32'hF3CC1B80 , 32'h0ED2EC30 , 32'h01BDF084 , 32'h051764F0 , 32'h01197BC8 , 32'hFE48C948 , 32'hFBF9FD98 , 32'hFE174600 , 32'hF1E02A20 , 32'hFE1A4690 , 32'h03EB34F0 , 32'hFEE946B4 , 32'h0056BD47 , 32'h0B948430 , 32'h018AEF44 , 32'h0070EE61 , 32'hFEF95538 , 32'h0156EE98 , 32'h00F96210 , 32'h0C766ED0 , 32'hFD806604 , 32'hFBCB1940 , 32'h01EA3CA0 , 32'hFF128D45 , 32'h05C51488 , 32'h00B57883 , 32'hFD4A62E4 , 32'hFFC0849B , 32'h00036910 , 32'hFFFB7D85 , 32'hFFFE7FDD , 32'hFFFF21C1 , 32'hFFFCD6B0 , 32'h0000BFCE , 32'h000102AC , 32'hFFFEEA61 , 32'h000370C6 , 32'h0000CC0C} , 
{32'h19A18080 , 32'h055DE4C0 , 32'h0D275480 , 32'hCDD78480 , 32'h0C38FE20 , 32'hEB2B91E0 , 32'hFB79BFA0 , 32'hFE5C3294 , 32'h0E7DE8E0 , 32'hF3E12520 , 32'hFDB8FE0C , 32'hF8D2FFB8 , 32'h0D95A770 , 32'hF5D18EF0 , 32'hFF2E2837 , 32'h0ACF25C0 , 32'h0D2AA7B0 , 32'h253872C0 , 32'hE428BBA0 , 32'h0F894C70 , 32'hE60D3AA0 , 32'hECCCB560 , 32'h199CD0A0 , 32'h13783160 , 32'h03775718 , 32'hFDC2EF38 , 32'h01BD61A8 , 32'h01770FF0 , 32'h042610B8 , 32'h28DB40C0 , 32'hFB8C4EA0 , 32'h0612C028 , 32'h14E93400 , 32'hEBE22EE0 , 32'hEFC831E0 , 32'h15BE92A0 , 32'hFFCA38FA , 32'hEB38F8C0 , 32'h02F1F140 , 32'h0A757330 , 32'hF39265A0 , 32'hEDF7EFC0 , 32'h02E4ACBC , 32'h048A3F20 , 32'h0F28EEB0 , 32'h09752370 , 32'h038A0184 , 32'hF27B7A90 , 32'hFC1290EC , 32'h0085B4B4 , 32'hFACD4EF0 , 32'hFDD4826C , 32'h0087B250 , 32'hF6777220 , 32'hD67CD2C0 , 32'hFB98E108 , 32'h022670EC , 32'hEDC8EE00 , 32'h10FBA660 , 32'h0691A8C8 , 32'h0014DFB3 , 32'hFF8B20E9 , 32'hFAF614D0 , 32'hFB57E780 , 32'h005BEED3 , 32'h01D92A20 , 32'h0E122400 , 32'h05A9E160 , 32'h001ACE10 , 32'h069A0D58 , 32'hFEB1D1B8 , 32'h0D7D1A40 , 32'h06FA92E0 , 32'h008D9F03 , 32'h072E8A00 , 32'hFF8B4F25 , 32'hF7B01E90 , 32'h031E7668 , 32'hFB28CE50 , 32'h01B3A520 , 32'hFC7147F8 , 32'hFFADF58D , 32'h024526C0 , 32'h05D98CB0 , 32'hFDD05300 , 32'hFD268E84 , 32'h02A8CAEC , 32'hF6F5D0E0 , 32'h06DA4A60 , 32'h011B5D30 , 32'h00049245 , 32'h00035894 , 32'h000461B5 , 32'hFFFEA973 , 32'hFFFF4C96 , 32'h00029C25 , 32'h0000FE80 , 32'hFFFB725B , 32'h0000781C , 32'hFFFFFAE4} , 
{32'h0002E602 , 32'hFFF977E0 , 32'hFFF960B5 , 32'h000404F1 , 32'hFFFDDA9E , 32'hFFFC6352 , 32'h00056FD4 , 32'h0001E1A6 , 32'h0004BD74 , 32'h0000E401 , 32'hFFFF94FD , 32'hFFFE9B07 , 32'hFFFDEE79 , 32'h0007EBAC , 32'hFFFF1D1F , 32'h0003D739 , 32'hFFFA9578 , 32'h0000124B , 32'hFFFDB2CE , 32'hFFFF3FD3 , 32'h00015BA6 , 32'h0003737C , 32'hFFF993F8 , 32'h00013AE4 , 32'hFFF9FAFC , 32'h000B4E50 , 32'hFFF73EFA , 32'hFFFC0BDA , 32'h000F6BAA , 32'h00048BBD , 32'hFFF529FF , 32'hFFFAE32F , 32'h000421A3 , 32'h0005AA43 , 32'hFFFF1804 , 32'h000700CD , 32'h0001BAC8 , 32'hFFFC0220 , 32'hFFFDEFED , 32'hFFF800DE , 32'h0003FAD4 , 32'h0002E95B , 32'hFFF9DDD6 , 32'hFFF8F73E , 32'h00009717 , 32'hFFFFBB9B , 32'hFFFC435C , 32'hFFFF9C20 , 32'hFFF8A3C4 , 32'h0001C737 , 32'h00001D3A , 32'hFFFC6090 , 32'h000BA356 , 32'h0002313A , 32'hFFFC6486 , 32'hFFFBE296 , 32'hFFFD7346 , 32'hFFFAF4EB , 32'h00034F6D , 32'h000031D3 , 32'h000736A1 , 32'h00054308 , 32'h00042AD1 , 32'h0008B1B3 , 32'hFFFBCC5D , 32'h0000A29A , 32'h0001A90A , 32'h0002F429 , 32'h00057C45 , 32'h00008DC8 , 32'h000B386D , 32'hFFFE6B10 , 32'h000528F6 , 32'h000065AA , 32'h0001E50F , 32'h0000B002 , 32'hFFFB93FD , 32'hFFFCF6A8 , 32'h0001BFDF , 32'hFFF9F88A , 32'h00055E89 , 32'hFFFB9C19 , 32'h0004769F , 32'h00022782 , 32'h00021109 , 32'h000A1D69 , 32'h000733BE , 32'h00032930 , 32'h0004F471 , 32'hFFFC8CB0 , 32'h0000E643 , 32'hFFFB7EB4 , 32'hFFFEACDC , 32'hFFFDA5EC , 32'h00015371 , 32'h0004A281 , 32'hFFF6E793 , 32'h00065E78 , 32'h00055EB0 , 32'h0002B2B8} , 
{32'h13D8D560 , 32'hEE18AF20 , 32'h02457A64 , 32'hD6225640 , 32'h4DBE3680 , 32'h4841A700 , 32'h17E7EEA0 , 32'hF880C4C8 , 32'hF7FE9DC0 , 32'hF6E35290 , 32'h44B1FA00 , 32'hDB6F2B40 , 32'h0F7178E0 , 32'h2B41B0C0 , 32'hFAE12158 , 32'h078B3CF8 , 32'h0FBAE340 , 32'h146E3940 , 32'hF8BCE888 , 32'hE994C2A0 , 32'h06AA8950 , 32'hD6663340 , 32'hFA7652B8 , 32'hF3FE6090 , 32'hE895F2A0 , 32'hF0C0B670 , 32'hFB5A8440 , 32'hF30C8340 , 32'hF91B0228 , 32'h08D73770 , 32'hF89EB980 , 32'h059C1F18 , 32'hED2D6FA0 , 32'hEF3D19C0 , 32'h0F61C8B0 , 32'hF26118B0 , 32'hEC43F580 , 32'hE8801980 , 32'h0A2463E0 , 32'hE6F873A0 , 32'hF2A36890 , 32'h1AD148E0 , 32'h1AD8F740 , 32'hFEA5C1A0 , 32'hF38DC040 , 32'hF1B27250 , 32'h082DDC60 , 32'hEAD16140 , 32'hF794D660 , 32'hFAF82390 , 32'hFC9AEB88 , 32'hE2D01FA0 , 32'hEA3FC100 , 32'hF7857340 , 32'h083F7580 , 32'hF9F3D410 , 32'h0DB079B0 , 32'h0EB2B960 , 32'h00C85C2F , 32'hF9E9AFA0 , 32'h027FA798 , 32'h07FC2668 , 32'h100619E0 , 32'h07D88B00 , 32'hEE9E2680 , 32'hF4427A70 , 32'hF4105670 , 32'hF9D74D68 , 32'h013917B4 , 32'h06776530 , 32'hFAA21F60 , 32'hFAD5A300 , 32'h0150F7A8 , 32'h00A737C8 , 32'h08227320 , 32'hFEC17B98 , 32'hF5EFCF20 , 32'h0303B984 , 32'hFCD31780 , 32'h0DD8CA90 , 32'hF3F38130 , 32'h0AB684F0 , 32'h031371F4 , 32'hFCE50124 , 32'h06285FB0 , 32'h00B08291 , 32'h0297EEC4 , 32'h01888748 , 32'hFAF83AF8 , 32'hFF24CCCD , 32'hFFFFB896 , 32'h00018CA1 , 32'hFFFEA2A3 , 32'h0003E01F , 32'h00032A96 , 32'h00005E14 , 32'h000080ED , 32'hFFFDFA0A , 32'hFFFFEF88 , 32'h000208A1} , 
{32'hB36A8900 , 32'hA9839880 , 32'hB325A300 , 32'hEB8C3220 , 32'h398E78C0 , 32'hEADDC200 , 32'hED4F2900 , 32'h08847760 , 32'hF3BB4D00 , 32'hDD723DC0 , 32'h07F65C78 , 32'hDA583D40 , 32'hD89749C0 , 32'h20734AC0 , 32'h92A5B800 , 32'h05DDFCB0 , 32'hF64320C0 , 32'hFAE4ADD8 , 32'hD7C1F400 , 32'hFAF81408 , 32'hF9F8D478 , 32'hE8256B60 , 32'hEA436E60 , 32'hEE561240 , 32'h12FC92A0 , 32'hE536D900 , 32'h11F2F5C0 , 32'hF4A833E0 , 32'h2C4652C0 , 32'hF07ACFD0 , 32'hE466C9A0 , 32'h10EF3C00 , 32'hFEF84BBC , 32'h0D64CA60 , 32'hE664FE00 , 32'h26714800 , 32'h06EAE998 , 32'hF35AED50 , 32'h04D346B8 , 32'hF0665370 , 32'h00360EC4 , 32'hFAAC9838 , 32'h02E63F58 , 32'h011693D4 , 32'hEB498760 , 32'hFFF8472D , 32'h07975318 , 32'h1056F720 , 32'hFC3D0B48 , 32'h1742FCC0 , 32'h0D0B1DC0 , 32'hF8CF8078 , 32'h1A04A100 , 32'hE4F04EE0 , 32'hF56F7370 , 32'hFF0BFC3C , 32'h086227B0 , 32'h0A4870F0 , 32'h02337014 , 32'hE5D21860 , 32'hFD79D264 , 32'h0670A238 , 32'h0C8DB060 , 32'hFDE4AA30 , 32'h01848368 , 32'h072C77D0 , 32'hF71E5C60 , 32'h083F0640 , 32'hFA257CA0 , 32'hFE92C384 , 32'hFBB7C518 , 32'hFAB1FB20 , 32'hF82E06F0 , 32'h007992EE , 32'hFC730C1C , 32'hF98DEE58 , 32'h03549820 , 32'hFD521518 , 32'h095B97B0 , 32'hF3DB0540 , 32'h05A0B0B0 , 32'h05A31F10 , 32'hFB647B88 , 32'hFDA53708 , 32'h053F0E40 , 32'h0212E7B4 , 32'h010EE398 , 32'h0247C434 , 32'hFF3D34DE , 32'h023AC72C , 32'h0004A891 , 32'hFFFAB6AC , 32'hFFFE28D0 , 32'hFFFE5C01 , 32'hFFFC4CD3 , 32'hFFF97491 , 32'hFFFE53FB , 32'hFFFE31B0 , 32'h0001934D , 32'h00020D98} , 
{32'h1B243DC0 , 32'h08B84620 , 32'h353C5180 , 32'hEB9D4540 , 32'h0F597400 , 32'hE1A1D960 , 32'hED103040 , 32'hFA022780 , 32'hE8496300 , 32'hE94D0B60 , 32'h2550BC80 , 32'h034FB150 , 32'h0ED64010 , 32'h161DB7A0 , 32'hF630EB30 , 32'hF3884990 , 32'hFA7F08B0 , 32'h07ACC328 , 32'hF32DDCE0 , 32'hFB2D06C8 , 32'hF8F802B8 , 32'hF9F4DE80 , 32'hDF810B00 , 32'h0B0BE1B0 , 32'h01B59604 , 32'hF14C1D90 , 32'h19AFB620 , 32'hE4738E20 , 32'h00038A04 , 32'hFD2D3EE0 , 32'hF4FD4A90 , 32'h03DA4DE0 , 32'h265F0380 , 32'h0141F1B4 , 32'h0C872FE0 , 32'h082B9400 , 32'h029A2A5C , 32'hF89A0DB8 , 32'h0112B1AC , 32'hEEE05580 , 32'hF0F36600 , 32'hF7031A20 , 32'hF3D30ED0 , 32'h0E5D8850 , 32'h156D8FA0 , 32'h0055127F , 32'h0B82DF70 , 32'hF928DB58 , 32'h041D6DE0 , 32'hF7BB3000 , 32'h04541540 , 32'hF341B080 , 32'h096DD230 , 32'hF8163A20 , 32'hF90F6750 , 32'h0E5DB880 , 32'hFA8339E8 , 32'h08AD68D0 , 32'hFD8B1424 , 32'h064133C0 , 32'h07035FE0 , 32'hEE540A20 , 32'hFA0C91C0 , 32'h02C83AFC , 32'h014BE7F4 , 32'h06E89230 , 32'hFE095F44 , 32'hFABEC520 , 32'h023C28BC , 32'h03A074B8 , 32'hF7422CC0 , 32'h07EF0580 , 32'h0663FA30 , 32'hFFB0EF4A , 32'h00D2F4F8 , 32'hFB0C6BC8 , 32'hFFE3895B , 32'hFE2D1E3C , 32'hFB420278 , 32'h0AAF7000 , 32'hFF18BCAB , 32'h0610CFF0 , 32'h02A258E4 , 32'hFB12F618 , 32'hF7770690 , 32'h0278D2F8 , 32'h00C48F52 , 32'hFDE544A8 , 32'hFD67E4D8 , 32'h02376954 , 32'hFFFF691E , 32'hFFFC6886 , 32'h0000D935 , 32'h00052981 , 32'hFFFEFA21 , 32'h000308FA , 32'hFFFD7FB3 , 32'h0004EA49 , 32'hFFFFDFCD , 32'hFFFDCD3C} , 
{32'h000A12A1 , 32'h000436AE , 32'hFFFFCD0A , 32'hFFFDDF9A , 32'hFFFB3B72 , 32'hFFFCA02C , 32'hFFFBDBE7 , 32'h00015B7F , 32'h000019B2 , 32'hFFFBFBAF , 32'hFFFC0881 , 32'h000384E5 , 32'h00017434 , 32'h0001F47B , 32'hFFFC6BDC , 32'h0002EA93 , 32'h0003E266 , 32'h00013AC4 , 32'h0005D003 , 32'h00084416 , 32'hFFFE7459 , 32'h0004805A , 32'h00069409 , 32'h0000C47B , 32'hFFFC4198 , 32'hFFF6BF20 , 32'hFFFE6F12 , 32'h00003792 , 32'hFFF580EB , 32'hFFFB0339 , 32'h0001D61E , 32'h00028BFD , 32'hFFFD5A9B , 32'hFFFEB06A , 32'h000105BF , 32'hFFFE5861 , 32'h0006D412 , 32'hFFF8C5F3 , 32'hFFFC4AE1 , 32'hFFFB518D , 32'h000466EB , 32'hFFFF8097 , 32'h0000F324 , 32'h00069D67 , 32'h00042BD0 , 32'h00055104 , 32'hFFFF227E , 32'h0000546B , 32'h0004BC97 , 32'hFFFBF6C4 , 32'h000312B6 , 32'h00004F5F , 32'h0005D77D , 32'hFFFC083D , 32'hFFF91E86 , 32'h0004CB59 , 32'h000083E5 , 32'h0009DFD2 , 32'h00045963 , 32'h00038AB6 , 32'hFFFA7EE4 , 32'hFFF79C65 , 32'hFFFE15C8 , 32'hFFFED617 , 32'h000836B1 , 32'h00029DB4 , 32'h0000C478 , 32'hFFFBBAC9 , 32'h00036C5D , 32'h00018D87 , 32'hFFFDE176 , 32'h00046A36 , 32'hFFF88FDF , 32'hFFFDC5D6 , 32'h00004BDA , 32'hFFFA9F19 , 32'h00022108 , 32'hFFFEDF03 , 32'h000079F9 , 32'h0002FE10 , 32'hFFFD2E6E , 32'hFFF8E627 , 32'hFFFD1AF6 , 32'h00027AF7 , 32'hFFF8EAAE , 32'h00011923 , 32'h00034B40 , 32'h00036977 , 32'h000DE63C , 32'h00055CB6 , 32'hFFFCE62E , 32'h00004041 , 32'hFFFD0D32 , 32'h00031EA9 , 32'hFFFF0D6A , 32'h00071B3C , 32'h000049EF , 32'hFFFB239E , 32'hFFF9AAF7 , 32'hFFF513E6} , 
{32'hFFFF523D , 32'hFFFE69B9 , 32'h0001A639 , 32'hFFFDE76B , 32'hFFFE1379 , 32'hFFFD08D1 , 32'hFFFE4CC3 , 32'hFFFF8051 , 32'h0002E98D , 32'h00019BA7 , 32'hFFFE0181 , 32'hFFFB95FA , 32'hFFFFB614 , 32'h0000C67B , 32'hFFFFA67D , 32'hFFFFD23A , 32'h0000E72E , 32'h000044A4 , 32'hFFFF0C2C , 32'hFFFC5BDE , 32'h00009DAC , 32'h0003A47D , 32'hFFFF4720 , 32'hFFFD25E1 , 32'hFFFE8FE7 , 32'h00000F24 , 32'hFFFB17D9 , 32'hFFFDBAC7 , 32'h00019311 , 32'hFFFDA301 , 32'hFFFD39A3 , 32'h00046311 , 32'h000416C3 , 32'hFFFE0CE2 , 32'hFFFAE63F , 32'h000064E9 , 32'hFFFB642E , 32'h000058F3 , 32'hFFFEE7E4 , 32'hFFFFFD94 , 32'h0000C479 , 32'h00011109 , 32'hFFFAE3F9 , 32'h00004456 , 32'h00022784 , 32'hFFFF7B0B , 32'h000103D0 , 32'h0001A443 , 32'h0001EC86 , 32'hFFFF947A , 32'h00038B84 , 32'hFFFF6D0D , 32'hFFFD635B , 32'h00004B79 , 32'hFFFBBCF4 , 32'h0004A5FC , 32'hFFFC004A , 32'h00008E81 , 32'h0000F4DD , 32'hFFFDD6A9 , 32'h0002873A , 32'h00004E2D , 32'hFFFD407E , 32'h00022D83 , 32'h00016778 , 32'hFFFEB574 , 32'hFFFEE5BE , 32'h00014BD4 , 32'h00012F0E , 32'h00028E52 , 32'hFFFB9746 , 32'hFFFD71D7 , 32'hFFFE85EF , 32'h00020B63 , 32'hFFFFF04C , 32'hFFFA807E , 32'h000010E1 , 32'h0000D693 , 32'h000152FF , 32'h0000E166 , 32'h0001D5C8 , 32'h00018D0E , 32'hFFFADE4F , 32'h0001BA66 , 32'hFFFFA708 , 32'h00020B34 , 32'hFFFC8C1E , 32'h0000B09C , 32'hFFFDECDF , 32'h000286A6 , 32'h00012F77 , 32'hFFFA13F8 , 32'h000CAF9A , 32'h0003CEA4 , 32'hFFFB8CF7 , 32'hFFFC1EF4 , 32'hFFFEF54E , 32'hFFFAB3A6 , 32'hFFFFED5D , 32'hFFFBCD61} , 
{32'hFFF9BC19 , 32'hFFF9564A , 32'h0000F908 , 32'h000112EB , 32'hFFFEA601 , 32'hFFFF000E , 32'hFFFEC247 , 32'hFFFE5A8A , 32'hFFFE9B4A , 32'hFFFDE957 , 32'hFFF8B77C , 32'hFFF8327E , 32'h0000585E , 32'hFFF587C1 , 32'hFFFB5364 , 32'hFFFD2C32 , 32'h00038354 , 32'h0002517E , 32'hFFFDB044 , 32'hFFF81E72 , 32'h00043808 , 32'hFFFB638D , 32'hFFFE787F , 32'hFFFD1877 , 32'hFFFFEE40 , 32'hFFF874AA , 32'h0003844C , 32'h000335E9 , 32'h00033105 , 32'hFFFF0185 , 32'hFFFB2616 , 32'h0005F486 , 32'h00034244 , 32'hFFFE1A94 , 32'h00049E69 , 32'hFFFE0D15 , 32'hFFFF9246 , 32'h00095F34 , 32'hFFFCA61C , 32'hFFFD8884 , 32'hFFFDB635 , 32'h000790BE , 32'h00033943 , 32'hFFFCFADD , 32'h000A08C6 , 32'h0000CB33 , 32'hFFFF67C4 , 32'h0003F326 , 32'h0004C607 , 32'hFFFCFFBD , 32'h000198FC , 32'h00024E19 , 32'hFFF8B561 , 32'h000403AB , 32'h0004F425 , 32'h0009BF59 , 32'hFFFC4716 , 32'hFFF72764 , 32'hFFFA34AA , 32'hFFF79EB8 , 32'hFFFB37D4 , 32'h0005669F , 32'h000388C6 , 32'h0005FBE9 , 32'hFFFAE9F8 , 32'hFFF81B5D , 32'hFFFE2FF7 , 32'hFFFDD31E , 32'h0002F7B9 , 32'h0006CD68 , 32'hFFFDAECF , 32'h000034D0 , 32'h00089B3A , 32'h0000689F , 32'hFFF80CF2 , 32'h00022D29 , 32'hFFFD68F9 , 32'hFFEE3646 , 32'hFFFE777E , 32'h0006E633 , 32'h00014C41 , 32'hFFFE6DB3 , 32'h0005F73D , 32'hFFFD19B1 , 32'h0004FA96 , 32'h0005B94D , 32'h000948CB , 32'hFFFB2155 , 32'hFFF86388 , 32'h0002EB8C , 32'hFFFE0DD5 , 32'h00019B63 , 32'hFFFA082E , 32'hFFFF0677 , 32'hFFFB827B , 32'hFFFD6F87 , 32'hFFFDA84C , 32'hFFFD7399 , 32'h00018150 , 32'h000083CB} , 
{32'hDF9CC000 , 32'h07127320 , 32'hFAF5F040 , 32'hECBAD280 , 32'hCCF20CC0 , 32'hFB4ED868 , 32'h2CE4A200 , 32'hEACE1500 , 32'h1DCB5AC0 , 32'h082BC390 , 32'hECD6BA40 , 32'h220C38C0 , 32'hE0205000 , 32'h17EACC40 , 32'h0FBF2FB0 , 32'hE6BBBA00 , 32'h0B395FA0 , 32'hEBF77700 , 32'hE827A440 , 32'hFBA35CA8 , 32'h101812A0 , 32'hE123A1E0 , 32'h108D6460 , 32'hD5D2FA00 , 32'hF1677850 , 32'h0BC521C0 , 32'h00099B47 , 32'h054B3318 , 32'h03952134 , 32'h0E795AE0 , 32'hE9C5DC40 , 32'h1D105B60 , 32'hE3E0B060 , 32'hC3159C40 , 32'h008712F7 , 32'hF4691BB0 , 32'hF7BFC0D0 , 32'h16955980 , 32'h060314B0 , 32'hF9721D88 , 32'h0F9838C0 , 32'hE5DBF6C0 , 32'h05351708 , 32'h00DF86B6 , 32'h085C7680 , 32'hF955B5D0 , 32'h032689E0 , 32'hFDB30EAC , 32'h0BC7ED50 , 32'hFF7B6AAC , 32'h1BD67AC0 , 32'hFA3077D0 , 32'hF9AA4F10 , 32'hEDC98620 , 32'hF1B9D040 , 32'hFDEC8C84 , 32'hFB37D2B0 , 32'hF4F57980 , 32'h09959A60 , 32'h11075760 , 32'hFFFE3E7D , 32'hF7BC1730 , 32'h04CA4750 , 32'h0F818A40 , 32'h01894228 , 32'h05117548 , 32'hF7F30290 , 32'hF7C81E40 , 32'hF206E770 , 32'hF94A1FF0 , 32'hF6B22F00 , 32'h0525E100 , 32'h029F3C84 , 32'hF5BB5C10 , 32'hFE909B2C , 32'h07C78BB0 , 32'h0014EE23 , 32'hFCE849B0 , 32'h041EE420 , 32'h00D0E7AD , 32'hFFA29A5D , 32'h06396880 , 32'h02F4A3E0 , 32'hFF54804E , 32'h050E5690 , 32'hFE22F7E8 , 32'h00503CB8 , 32'hFFEE372A , 32'h04CEF428 , 32'h00A41F13 , 32'hFFFC9DA8 , 32'hFFFE7BCF , 32'h00010F33 , 32'hFFFF2831 , 32'h0003A9B4 , 32'hFFFE9F1D , 32'h0006547E , 32'h00039DE4 , 32'hFFFC9347 , 32'hFFFC8003} , 
{32'hF87D4870 , 32'h38BA5680 , 32'hD7A8D880 , 32'hF6312CE0 , 32'hCBAACF80 , 32'h2CB92200 , 32'h0DEAD8A0 , 32'h99EEA900 , 32'h4D209000 , 32'h09E16A20 , 32'hE0CA12A0 , 32'hFB3B2568 , 32'h31261540 , 32'hF3A80F00 , 32'h1096CE20 , 32'hFFF1E17B , 32'h0C148ED0 , 32'h3BC48340 , 32'hDA199840 , 32'hEF768960 , 32'h18DACB00 , 32'hE5F1BB40 , 32'hD9B5B740 , 32'h15F514A0 , 32'hCFAA8740 , 32'hE5FE1680 , 32'h04C4D5C0 , 32'h08E627F0 , 32'hD63F3340 , 32'h02448B74 , 32'h037820CC , 32'h3D075A80 , 32'hEF150080 , 32'h15800B40 , 32'h001548AF , 32'hF6DD4CD0 , 32'h2806F200 , 32'h040E78E8 , 32'h056E1048 , 32'hD5F92940 , 32'hF92B0F40 , 32'hF6DE73D0 , 32'h07A96978 , 32'hFE54F050 , 32'hF87E5288 , 32'hF17915D0 , 32'hEDE42F00 , 32'h1E660180 , 32'hEC5BB320 , 32'h0266CD54 , 32'hEE48CC20 , 32'h02077110 , 32'h047982D8 , 32'hF78A7960 , 32'h028C4858 , 32'h0EF497F0 , 32'hE5670320 , 32'hE5650D00 , 32'hF4470A20 , 32'hE8F09E40 , 32'h04850E68 , 32'h0F1C3130 , 32'hF7A254E0 , 32'hFE4D90E4 , 32'hFF2A46D1 , 32'h05D8CBB8 , 32'h0911AFE0 , 32'hF87D23F8 , 32'hFC405150 , 32'h03E6F768 , 32'h04369F18 , 32'h000DC0FC , 32'h0129526C , 32'h02E92810 , 32'hFF317F27 , 32'hF7D20FD0 , 32'hFAC42540 , 32'hF98BB918 , 32'hFC7CFD98 , 32'hFF565C02 , 32'h02A2B29C , 32'h07107868 , 32'hFBE6EA20 , 32'h02D86820 , 32'hFC8CBD28 , 32'h03FF8C34 , 32'hFFCD62B4 , 32'h05466FC0 , 32'hFEF60894 , 32'h0117ED70 , 32'hFFFF3E86 , 32'h0003BCFE , 32'h0001BC93 , 32'hFFFFC08D , 32'hFFFFEFCB , 32'hFFFD4714 , 32'h0000E04B , 32'h0000896E , 32'h0000F12D , 32'hFFFE1E98} , 
{32'hFFFF239C , 32'h0002B402 , 32'hFFFCC99E , 32'hFFF9E9C3 , 32'h0005EFDA , 32'h00010C81 , 32'h000680B0 , 32'hFFF98DFB , 32'hFFFC7D98 , 32'h00034156 , 32'h0005CE6E , 32'h0001C20C , 32'hFFF8DDBE , 32'h00015712 , 32'hFFFBE13A , 32'h00005FA6 , 32'h00022175 , 32'h000301CB , 32'hFFFEEFCE , 32'hFFFBE4F9 , 32'h00043822 , 32'h00022705 , 32'hFFFDC1C6 , 32'h0006A62C , 32'hFFFA2467 , 32'h00007B5D , 32'h0002E2E6 , 32'hFFFFF859 , 32'hFFFAF59E , 32'h0005683F , 32'hFFFE06CA , 32'hFFFA3E52 , 32'h00028712 , 32'h0003D373 , 32'h0002F2F2 , 32'hFFF8F09E , 32'h00049EAE , 32'h0002F1D0 , 32'hFFFD022F , 32'h00027AF6 , 32'h0004391E , 32'h00012636 , 32'hFFFF0948 , 32'hFFFE3755 , 32'h000301E6 , 32'h00031770 , 32'hFFFDC4EC , 32'h0008FC46 , 32'h000331C9 , 32'hFFFF50C5 , 32'h000086B3 , 32'hFFFE992D , 32'h0005D104 , 32'h00044F4C , 32'h0005BAE7 , 32'h0002A88F , 32'h0000B80C , 32'hFFF97994 , 32'h0000CA8D , 32'hFFFAF547 , 32'h000385F5 , 32'hFFFE4295 , 32'hFFFFE209 , 32'hFFFCC3B8 , 32'hFFF62AA7 , 32'hFFF68597 , 32'hFFFBADF2 , 32'h0001A6C5 , 32'hFFF8E016 , 32'hFFFDF09A , 32'h0000D56C , 32'hFFFE7974 , 32'h000763F0 , 32'hFFF566BB , 32'hFFFAE29C , 32'h0004C7DB , 32'h0002DB0B , 32'hFFF6CF81 , 32'hFFFC3AAB , 32'h0005CA3D , 32'h0007B3CA , 32'hFFFBDBE3 , 32'hFFFD21F3 , 32'hFFF8EF3D , 32'h0003F166 , 32'h00024BB6 , 32'hFFF72B26 , 32'hFFFECEED , 32'hFFFDB172 , 32'hFFFD5857 , 32'h0001D234 , 32'hFFFE337E , 32'hFFFDAE37 , 32'hFFF6051B , 32'h0008D29C , 32'hFFFE9CF5 , 32'h0003F348 , 32'h0000D969 , 32'hFFFEA028 , 32'hFFFD577A} , 
{32'h90261D00 , 32'h11758E80 , 32'h4F8A2B00 , 32'h541EC880 , 32'h6AE63C80 , 32'hBA6E1600 , 32'h0A355320 , 32'hFB7C5700 , 32'h0BDB5860 , 32'h069206A0 , 32'h5BEB6900 , 32'h403CE080 , 32'hF4ADC530 , 32'h1B7839A0 , 32'h040D0960 , 32'h0EECFA40 , 32'h2C47AF00 , 32'hE738D760 , 32'h0EF1D080 , 32'h39B88580 , 32'hCB55E480 , 32'hF5429A00 , 32'hF5EA66B0 , 32'hF58DCAD0 , 32'hE36429A0 , 32'h1230D9E0 , 32'hF1D0BD10 , 32'h01AEEEE0 , 32'hFF6B30E9 , 32'h081F4F20 , 32'hD8EFF000 , 32'h2504BD80 , 32'h07A96BE8 , 32'hF505CB40 , 32'hF6BB2570 , 32'h14B68200 , 32'h096AB1C0 , 32'h15389E40 , 32'hE8974880 , 32'h0E0C0BD0 , 32'h05F41D00 , 32'hF8218DC8 , 32'hF1235150 , 32'hF364FD30 , 32'hF05EA6C0 , 32'h0D3E47B0 , 32'hED3A15C0 , 32'hF87B0B88 , 32'h037E0488 , 32'h064A8110 , 32'h0D234CE0 , 32'h06D91330 , 32'hF65B9F60 , 32'h06354A88 , 32'h03113E98 , 32'hFB0441C8 , 32'h01CB148C , 32'hEDEA5B00 , 32'hFDA6652C , 32'hF1CD2910 , 32'h05523E70 , 32'h0617A408 , 32'hE35B1860 , 32'hFD1CAD74 , 32'h0C2D6FC0 , 32'hF74D8220 , 32'hF8D761F0 , 32'h069B9660 , 32'hFA877ED0 , 32'hF84D2478 , 32'h0227C0AC , 32'hFCE1CC9C , 32'hF86CEE40 , 32'hFF8C1722 , 32'hFC488D00 , 32'h032DEBF4 , 32'h069960F0 , 32'h0137B830 , 32'h04BB7D00 , 32'h058CD7A8 , 32'h04A7C9B8 , 32'h04401AE0 , 32'h05304680 , 32'hFB979168 , 32'h01031970 , 32'h05FF8BB0 , 32'hFD01A07C , 32'h01D06F18 , 32'hFB6A63B8 , 32'h01334050 , 32'hFFFC9680 , 32'hFFFF9747 , 32'h0000D69E , 32'h0001F382 , 32'h000077DE , 32'h000440DA , 32'h0000AFAE , 32'hFFFF5BB6 , 32'hFFFEB200 , 32'hFFFE969B} , 
{32'h0006D5E2 , 32'h000462B9 , 32'hFFFC7E00 , 32'hFFFDBED4 , 32'h00008308 , 32'h0003FE94 , 32'hFFFD5A02 , 32'hFFFC681D , 32'h00003304 , 32'hFFFC51E6 , 32'h0006DB35 , 32'hFFFC77FE , 32'h0000030F , 32'hFFFE0234 , 32'hFFFDF2D6 , 32'h0004F8E5 , 32'h00000835 , 32'h0004B904 , 32'h0003B7E5 , 32'hFFF75C0A , 32'h00004560 , 32'h00028F5A , 32'h0000FC62 , 32'hFFFAFCC8 , 32'hFFFC49FF , 32'hFFFA8453 , 32'h0005C076 , 32'h0005A73A , 32'h0002CD69 , 32'h0003F31F , 32'h0002AA4F , 32'hFFFEB471 , 32'hFFF8AD54 , 32'hFFFDC127 , 32'h00000FE6 , 32'h0002E991 , 32'hFFF93160 , 32'h00031541 , 32'h0002CA31 , 32'hFFF968FB , 32'h00076C09 , 32'h000155A4 , 32'hFFF71E5D , 32'h00013C18 , 32'hFFFCFAB7 , 32'h00003B1A , 32'hFFFC0698 , 32'h00001B72 , 32'hFFFCFC36 , 32'h00041F05 , 32'h00056790 , 32'hFFFF0E13 , 32'hFFF694FB , 32'h0006B3E7 , 32'h0005F0C0 , 32'h0000AE38 , 32'h00008461 , 32'hFFFB21BF , 32'hFFF7683F , 32'h0002FA19 , 32'hFFFE8E74 , 32'hFFFAB56C , 32'h000A497C , 32'hFFFE54C0 , 32'hFFFA9BF9 , 32'h0007AF5B , 32'h0002B788 , 32'h00046ECE , 32'hFFFD0F99 , 32'h000AA9FA , 32'hFFFD3375 , 32'h0000636B , 32'hFFFD6DBC , 32'h0003728D , 32'hFFFFA448 , 32'hFFFE3BC0 , 32'h00007D8A , 32'hFFFF0C47 , 32'hFFF5EE13 , 32'h0000A528 , 32'hFFFCB8B3 , 32'h00061EC6 , 32'hFFF8B322 , 32'h000088A7 , 32'hFFFE2B92 , 32'hFFFE46DD , 32'hFFF66C4F , 32'h00013639 , 32'hFFF8BEF8 , 32'h00043D13 , 32'h000A7DBC , 32'h0002216B , 32'h00054B0F , 32'h000AAFFE , 32'hFFFD4803 , 32'h0002B820 , 32'hFFFEB53A , 32'h000371D5 , 32'h0006C8C3 , 32'h000237D6} , 
{32'hFFFBEFAF , 32'h0000A031 , 32'hFFF745D5 , 32'hFFFF794C , 32'h0000A945 , 32'hFFF98C2B , 32'hFFFCD4AF , 32'hFFFA43CA , 32'hFFFB1F4F , 32'h00017EDD , 32'hFFF8ADFE , 32'hFFFBC68D , 32'hFFFE21FB , 32'h00011AAB , 32'hFFFEDB28 , 32'hFFFF7163 , 32'h00031A4F , 32'hFFF8A128 , 32'hFFFCF7B9 , 32'hFFF92BEF , 32'h000832CB , 32'h0005A3D8 , 32'h00020246 , 32'hFFFA26A4 , 32'hFFFFFD5E , 32'hFFFFAC6A , 32'h00019949 , 32'h0001C52D , 32'h0003412D , 32'hFFFF3432 , 32'hFFFB9481 , 32'h0004749C , 32'hFFFDD77C , 32'hFFF9D2E1 , 32'h0004E35D , 32'hFFFE6E2E , 32'h0001B3DB , 32'h00023293 , 32'hFFFCE43A , 32'hFFFD810E , 32'h0001ECC2 , 32'hFFFD7FBB , 32'h00004EAB , 32'h00016D47 , 32'h000AB459 , 32'hFFFB1A03 , 32'hFFFB787E , 32'h00017DA7 , 32'hFFFD05F9 , 32'hFFFEBB5B , 32'hFFFD54BF , 32'hFFFEAA8C , 32'h0005867C , 32'h00002DD4 , 32'hFFFDCC21 , 32'hFFFBB7D9 , 32'h0000B604 , 32'h00028EC0 , 32'hFFFE5103 , 32'h0000FAD0 , 32'hFFFD77A7 , 32'h0002E33C , 32'hFFFD564E , 32'h0005283F , 32'hFFFBC01A , 32'h00032B55 , 32'hFFFDF61D , 32'hFFFFCE93 , 32'hFFFEC7D9 , 32'hFFFEA767 , 32'hFFFB94FF , 32'h0001B305 , 32'hFFFE98FF , 32'h0007462D , 32'h000970EF , 32'hFFF9E73B , 32'hFFFDA7E3 , 32'h0003C7E9 , 32'hFFFCE7F2 , 32'h0001E39F , 32'h000523C8 , 32'hFFFDDE63 , 32'hFFF92AAE , 32'h0006068F , 32'hFFFA9B41 , 32'h00012937 , 32'h00010097 , 32'h00020377 , 32'h00010C7F , 32'h0000D1D7 , 32'h000CCB52 , 32'h00023267 , 32'h00045CC1 , 32'h0008D1F5 , 32'h00042A40 , 32'h000482F9 , 32'h000185B1 , 32'h0004EC43 , 32'h00015021 , 32'h0001C59B} , 
{32'hDD8047C0 , 32'h498B8980 , 32'hE2DA87A0 , 32'h0DDB95D0 , 32'h0D41A800 , 32'h3DCFDF40 , 32'h305B0980 , 32'h25B266C0 , 32'h1A348F40 , 32'h0A0BB080 , 32'hE88FA5A0 , 32'hE814DDA0 , 32'hD92286C0 , 32'h1C685120 , 32'hE955E500 , 32'h574C4A00 , 32'hE83D4DE0 , 32'h12A21980 , 32'hFF51E4E8 , 32'hD668EAC0 , 32'h19553B00 , 32'hDF397440 , 32'hEB938AC0 , 32'h027E821C , 32'hEC270CC0 , 32'hE33B2C80 , 32'hEC0B64A0 , 32'h2295B0C0 , 32'hF07C13B0 , 32'hFE471E34 , 32'h18068AC0 , 32'h144EE2C0 , 32'h24C70B40 , 32'hEE3B9EE0 , 32'h2CEDD5C0 , 32'hEC904A80 , 32'hF4514340 , 32'hFB0BDD98 , 32'hFFBF530C , 32'hFFB8875F , 32'h0552FB60 , 32'h077FE7D8 , 32'hEA0097A0 , 32'hF03E46D0 , 32'hF28C16D0 , 32'h12376400 , 32'hEB19DD80 , 32'hF8FF9F58 , 32'h0DA4E450 , 32'hFF317FDB , 32'h1E7872C0 , 32'hFEACB4C4 , 32'h04AB6080 , 32'hEAB66D40 , 32'hF43A8D30 , 32'hFBE3F3B8 , 32'h077B8578 , 32'h02FE7F18 , 32'h04B433F0 , 32'hFF8B8511 , 32'h077E1F98 , 32'h0AF3E810 , 32'hFFB00F8D , 32'hFC8393EC , 32'h05FAA7E0 , 32'h05E71968 , 32'hF94559C8 , 32'h03CEB9DC , 32'h0DDEC020 , 32'h02792138 , 32'hFE2F972C , 32'h05E78760 , 32'h0B1036C0 , 32'h08132950 , 32'hFDEF0D44 , 32'h00B6B426 , 32'h09E95960 , 32'hFE4FD6DC , 32'h01F9C958 , 32'hF8904BC8 , 32'hF8E6E2D0 , 32'hF5F1E4E0 , 32'h05C53768 , 32'hFD162504 , 32'hFB0F1BF8 , 32'h042E51A8 , 32'h0172EDA8 , 32'h0087ED86 , 32'h011CE574 , 32'hFFC30D74 , 32'h00019D10 , 32'hFFFF510A , 32'hFFFDD8AB , 32'h00029984 , 32'hFFFD0574 , 32'hFFFE7085 , 32'hFFFE2B09 , 32'hFFFED536 , 32'hFFFE24BB , 32'h00002BD8} , 
{32'h1D51BD80 , 32'hE95EBD40 , 32'h098287C0 , 32'hEA65AB80 , 32'h11502340 , 32'hFA607FA8 , 32'hEE3DC300 , 32'h159FA980 , 32'hF9FBCE68 , 32'hFC7DA950 , 32'hF8A9CD78 , 32'hE279B100 , 32'hE63EA5C0 , 32'hFED078B4 , 32'hEF3B6460 , 32'h0062B67F , 32'h0162695C , 32'h0CAD7FE0 , 32'hF7E68B60 , 32'h0625EB40 , 32'h06575420 , 32'hFDE011A0 , 32'hFFDB83A0 , 32'hFD5C52A0 , 32'hFE73B0F0 , 32'hEEEE77E0 , 32'h028C37E0 , 32'h1B9525C0 , 32'hF8584C80 , 32'hF333EA00 , 32'h015F812C , 32'h05C7D018 , 32'hF882B448 , 32'hFE4E36B4 , 32'hF32C3880 , 32'hF8535BD0 , 32'h1535DAA0 , 32'hFF0CED16 , 32'h08EE0740 , 32'hFA87B700 , 32'h0570CF18 , 32'h00E28AF4 , 32'hF515D7F0 , 32'hFE543640 , 32'h06B78768 , 32'hFB7245F0 , 32'hF003D680 , 32'hF03919D0 , 32'h0341CCE4 , 32'h0E573F60 , 32'hFAB19C60 , 32'hF1AE0650 , 32'hF31A0340 , 32'h01B6ED14 , 32'hF7EC4D70 , 32'hFB9506B8 , 32'hF6BDFA10 , 32'hFD0B5210 , 32'h16EC1980 , 32'h0D864D90 , 32'h05218240 , 32'hF462EB20 , 32'h004D618A , 32'h02A89C5C , 32'hFFB39C9D , 32'h106380C0 , 32'hFCF2ED30 , 32'hFC5C9330 , 32'h08574E70 , 32'hFE6B4B50 , 32'h0B0427D0 , 32'hEAB7A6C0 , 32'h0308E16C , 32'hF73510B0 , 32'h0DF4DE80 , 32'h08C51170 , 32'h07022E28 , 32'hFE5E40FC , 32'hF99B2068 , 32'h0290A4DC , 32'h028420C4 , 32'hFE622D20 , 32'h043F7BF0 , 32'h05843678 , 32'h07BC3190 , 32'hFC209678 , 32'hFF745CD6 , 32'h03F399F4 , 32'hFDD8AADC , 32'h004C676A , 32'h0004FCBE , 32'h00045A3C , 32'hFFFBA273 , 32'hFFFFA56F , 32'hFFFD7EAF , 32'h00027EDC , 32'h00006F66 , 32'hFFFC93BF , 32'hFFFFD95C , 32'h00009048} , 
{32'hFCC80E5C , 32'h0057A3B2 , 32'hF0FF6370 , 32'hFE405D64 , 32'hF5DE7A50 , 32'hFDA65F8C , 32'h13F6C580 , 32'h0038B55E , 32'h03495DB0 , 32'hFBDA6048 , 32'h06449820 , 32'h066A6D60 , 32'hFB5715B8 , 32'h0E53CBA0 , 32'hF09FB0A0 , 32'h0A301870 , 32'h015CFD2C , 32'h1303D740 , 32'h03EB15AC , 32'hFD3047E8 , 32'hFBE67E40 , 32'hECD5A580 , 32'hFAA529F8 , 32'h07074E40 , 32'h0CB17510 , 32'hFF031777 , 32'h0A0F20C0 , 32'h09BF4B60 , 32'hF7499880 , 32'hFA609590 , 32'h00982546 , 32'h06A12D40 , 32'hF8AD04C0 , 32'hF71C2530 , 32'hF7A599D0 , 32'hEF925A60 , 32'h072A9B68 , 32'h0CA380D0 , 32'hF6DE0B50 , 32'hEF100D20 , 32'hF6995BA0 , 32'hF51F09D0 , 32'h00DDB151 , 32'h0A9A6440 , 32'h0D17D7E0 , 32'hF65CA010 , 32'hEF946660 , 32'h006666CF , 32'h0AA66E90 , 32'h07E75F40 , 32'h056542C0 , 32'h0486CC88 , 32'hF71ACBA0 , 32'hFF467632 , 32'h0BADFAE0 , 32'hF5DF43C0 , 32'hFE8A0B84 , 32'hF872D118 , 32'hF75EA510 , 32'h04E53C48 , 32'hF6613900 , 32'h06FD9430 , 32'h0CF1D690 , 32'h043C3FD8 , 32'h00531CD7 , 32'h0AE09800 , 32'h042EDC08 , 32'h0D9A8780 , 32'hF7911900 , 32'h0AD41FC0 , 32'hFB80CA98 , 32'hF6A3C5B0 , 32'hF21EEDF0 , 32'h01D06ED4 , 32'hFAD11E48 , 32'h088DCFB0 , 32'hF844B608 , 32'hF7E5A890 , 32'hF7BEDEB0 , 32'h01F08840 , 32'hF18854E0 , 32'hFFA8DC18 , 32'hFCE1C680 , 32'hFFB68FBC , 32'hF654AE00 , 32'hFDBB8628 , 32'h0056131A , 32'hFC23C904 , 32'h00632668 , 32'h01E5B248 , 32'h0000A7C8 , 32'h000060B0 , 32'hFFFAB1F2 , 32'h000690F3 , 32'h000095F5 , 32'h0001761C , 32'hFFFF9F3B , 32'hFFFDEA2C , 32'h00014C76 , 32'hFFFE6CD2} , 
{32'hFFF330BE , 32'h00012F37 , 32'hFFFD5C6B , 32'hFFFE1A4E , 32'hFFF2E67E , 32'h00068189 , 32'h0008BA83 , 32'h00006F2C , 32'h00077440 , 32'hFFF50906 , 32'hFFFE9A79 , 32'h00034BE5 , 32'hFFFC33AA , 32'h0004BE1D , 32'hFFFFAAE4 , 32'hFFFF0A66 , 32'hFFFEA6D6 , 32'hFFF7C9FC , 32'hFFFB28CB , 32'hFFFDBE44 , 32'hFFFEBD0C , 32'hFFFE6FD8 , 32'h0000A10D , 32'h00054FE1 , 32'hFFFD8740 , 32'h000237F3 , 32'h00086FD4 , 32'hFFFE930B , 32'h00005C56 , 32'hFFFD2E4D , 32'hFFFDC66C , 32'hFFFE7BBE , 32'hFFF8896C , 32'hFFFD01BE , 32'h000170C3 , 32'h00010569 , 32'h0000B1D5 , 32'hFFF60695 , 32'h00051605 , 32'hFFFAB058 , 32'hFFFAB772 , 32'h0003B05B , 32'h00006AF6 , 32'h00033670 , 32'hFFF5C4F7 , 32'hFFFA07C7 , 32'hFFFEFB07 , 32'hFFFADEAE , 32'hFFF9A1C3 , 32'h0001E677 , 32'h0003F1F6 , 32'hFFF9E773 , 32'hFFFD424F , 32'h0004DC00 , 32'hFFFCB783 , 32'hFFFAC233 , 32'hFFFFCA6A , 32'hFFFBF166 , 32'h0000A504 , 32'hFFFF3AE8 , 32'hFFFD7A6F , 32'hFFF9FB52 , 32'hFFFB32F5 , 32'hFFF2CC1A , 32'hFFFD8E09 , 32'h000AA53E , 32'hFFFFFFE8 , 32'hFFF5E6C0 , 32'hFFFC4790 , 32'hFFFD66A0 , 32'hFFFCBDDD , 32'hFFFF7379 , 32'h0005F4E4 , 32'h00068146 , 32'hFFFEA2A9 , 32'h00035492 , 32'h000D029C , 32'h00013B02 , 32'h00046155 , 32'h000931BE , 32'h000B09DF , 32'hFFFE4B39 , 32'h000301B2 , 32'h000010AD , 32'h00037DEE , 32'h000CDD29 , 32'h00035C03 , 32'hFFF79C9D , 32'h00068E32 , 32'h0005E7B7 , 32'h0002EAAD , 32'h0002A1BE , 32'h00002B29 , 32'hFFF5CB54 , 32'h000E5106 , 32'hFFFE486E , 32'h0002261C , 32'h00003CDF , 32'h00008995 , 32'h0001A115} , 
{32'h11561540 , 32'h0ECC33E0 , 32'h226F69C0 , 32'hF03B66D0 , 32'h55B4F200 , 32'h213494C0 , 32'hD40A51C0 , 32'h1FBF25A0 , 32'hE2B9E9A0 , 32'hF62BB760 , 32'hF40664D0 , 32'hF208B920 , 32'hF7288110 , 32'h0E072C60 , 32'h2AD1A700 , 32'hF6E70C40 , 32'hFAF4CB68 , 32'h04186CD8 , 32'hFBC2F1B8 , 32'h12B507E0 , 32'h19B963E0 , 32'hDE7FB140 , 32'hF8345758 , 32'hDEEBF740 , 32'h033F6078 , 32'h1C821860 , 32'hE97002A0 , 32'h24C87DC0 , 32'hF9DDD040 , 32'hF58CA420 , 32'hF5CAE6B0 , 32'h01A59444 , 32'h095545D0 , 32'hF3EAE460 , 32'hECDB0CC0 , 32'hF00902B0 , 32'hF0A17C30 , 32'hF04E0800 , 32'h00A9719F , 32'hF2F16AD0 , 32'h14CD1380 , 32'hDF58EA40 , 32'hFBC192C0 , 32'hF77E1120 , 32'h13DD7940 , 32'h0CC76490 , 32'hF4C9BD70 , 32'h06E4A120 , 32'h1CE4D420 , 32'h0672AC48 , 32'hF11A52A0 , 32'h11B46F40 , 32'hE75C3700 , 32'hFF91EE15 , 32'hFF34A352 , 32'hF6477320 , 32'hFF5E8E60 , 32'hFE0503B8 , 32'h036015D0 , 32'hF2380310 , 32'h13E9AAC0 , 32'h01F83480 , 32'hF6207B90 , 32'hF5A27A10 , 32'hF9709F20 , 32'h03247AC4 , 32'h18AE6A20 , 32'h07148EA0 , 32'h0551C308 , 32'h01A9791C , 32'hFAFB3658 , 32'hFF640EA8 , 32'hF1E99340 , 32'h03190BF8 , 32'hF46AEC00 , 32'h03003A04 , 32'hF9940F10 , 32'h05D54488 , 32'hFACD4A20 , 32'hF49A1CE0 , 32'hF74DC8F0 , 32'h0A762BE0 , 32'hFB666D28 , 32'hFA4BB9E8 , 32'hFC6E5764 , 32'hFF5AC7F9 , 32'h02E63E20 , 32'h0282BCFC , 32'h013E0ACC , 32'hFE51CE3C , 32'h00042D5C , 32'hFFF827FD , 32'hFFFEC343 , 32'hFFF94617 , 32'h0002FDED , 32'hFFFE179B , 32'hFFFF6E76 , 32'hFFFFCC5D , 32'h00014BFD , 32'h0000DBCF} , 
{32'hFFFDE397 , 32'h00003337 , 32'hFFF8CF91 , 32'h00078AE1 , 32'h0000736B , 32'hFFFE37A8 , 32'h00024721 , 32'hFFFF2D27 , 32'hFFFF85AB , 32'h00083952 , 32'hFFFDC79B , 32'h000087BF , 32'h000BE7C2 , 32'hFFFA656E , 32'h000101E1 , 32'hFFFB4E04 , 32'h0001FC2B , 32'h00008005 , 32'h00016F99 , 32'hFFFC7F1E , 32'hFFFF567A , 32'hFFF918B2 , 32'hFFFDD623 , 32'h0002BDDC , 32'h0002C8AE , 32'h000B4499 , 32'h000243E7 , 32'h00072254 , 32'hFFF6AB69 , 32'hFFFC42A7 , 32'hFFF96B4E , 32'hFFFF7DD9 , 32'h0001272D , 32'h000906FB , 32'hFFFFC28D , 32'h000C5289 , 32'h000187C2 , 32'h0001A41D , 32'h0004A04B , 32'h00030119 , 32'hFFFEDFD9 , 32'h00017205 , 32'hFFFADEA7 , 32'hFFFBC9FA , 32'h0004AF1B , 32'h0003301E , 32'hFFFEAA10 , 32'h00020140 , 32'h00064C11 , 32'hFFF9083C , 32'hFFFCD0F5 , 32'h000296B0 , 32'h00089236 , 32'hFFFC7366 , 32'hFFFB7051 , 32'hFFFFE8DB , 32'hFFFF51A0 , 32'h0005FE75 , 32'h0004B115 , 32'hFFFDB140 , 32'h0000E827 , 32'hFFFC1F5C , 32'h00007B10 , 32'hFFFE52FD , 32'hFFFAFDD6 , 32'hFFFF38BA , 32'h00021B41 , 32'h0001BE65 , 32'h00011606 , 32'hFFF96FEB , 32'h0000B390 , 32'hFFF9C4E6 , 32'hFFFC49A1 , 32'h000405C9 , 32'hFFFF4AEF , 32'hFFFFB4AE , 32'hFFFDDF2E , 32'h0003986B , 32'hFFFE4675 , 32'hFFFAFF4A , 32'h0008D044 , 32'hFFFD4CA9 , 32'hFFFB666A , 32'hFFFB2DC0 , 32'h000112F3 , 32'h000156B3 , 32'h0002A94B , 32'hFFF9AF09 , 32'h0002AFD9 , 32'h000007CD , 32'h00044037 , 32'h0000F301 , 32'hFFFE5DB9 , 32'h0001D052 , 32'hFFF820CD , 32'h0003EFD3 , 32'h0000FF7D , 32'h0001962E , 32'h0003621A , 32'hFFFFFC71} , 
{32'h0007B2B3 , 32'hFFFC9259 , 32'h00007920 , 32'h0000FCE8 , 32'hFFFBF731 , 32'h0002DCD5 , 32'h000289AB , 32'h0007DDF8 , 32'hFFF9893C , 32'hFFFE2B37 , 32'hFFFE3B7B , 32'hFFFD0807 , 32'h000109D5 , 32'hFFFB4AB8 , 32'hFFF9919C , 32'hFFFDA31B , 32'h00024B1D , 32'h00063D4C , 32'hFFFD9155 , 32'h0002D675 , 32'hFFF8581B , 32'h0002DA3F , 32'hFFFD3D54 , 32'hFFF84D9C , 32'h000046DE , 32'h00019392 , 32'h00082A9A , 32'h00029B02 , 32'hFFFE1C32 , 32'hFFFBA736 , 32'hFFFBE66D , 32'hFFF93CB7 , 32'h000471A2 , 32'hFFFFFDD2 , 32'h0001A63A , 32'h00057BEB , 32'h0004BFD8 , 32'h00081E7B , 32'h000521B9 , 32'h00022960 , 32'h0002BD8C , 32'h00024EF4 , 32'hFFFB136B , 32'hFFFDE2AB , 32'h0001BB3C , 32'h0001331B , 32'hFFFE9901 , 32'h00074569 , 32'h00018718 , 32'hFFFAFCD3 , 32'h000442D3 , 32'hFFFE2431 , 32'hFFFFE382 , 32'h00002883 , 32'h000136E0 , 32'hFFF91B71 , 32'hFFFE643A , 32'h00065EB6 , 32'hFFFFD7F5 , 32'h00011DAE , 32'h00035E84 , 32'h0000E0CD , 32'h0000A0CE , 32'hFFFEFEAE , 32'hFFF8B2A8 , 32'hFFF9884A , 32'hFFF8121A , 32'h000AAB53 , 32'hFFFD08D5 , 32'h00040A55 , 32'h0000A515 , 32'h000437C5 , 32'hFFFFE7D7 , 32'hFFFD9824 , 32'hFFFEA2FE , 32'hFFFCCA25 , 32'hFFFF9708 , 32'h00003075 , 32'h00085F53 , 32'h0006AD28 , 32'hFFFC7B71 , 32'h0004086E , 32'hFFFED51B , 32'h0000B59E , 32'h0005CBB8 , 32'h0001422A , 32'h00049B7A , 32'h00002D48 , 32'hFFF859BB , 32'h0005C3C0 , 32'hFFFB9BEF , 32'h0001258E , 32'hFFFD2E87 , 32'h0003BA3D , 32'h000B2CAC , 32'hFFFF036F , 32'hFFFC79AC , 32'h0002A364 , 32'h00045A8D , 32'hFFFD77F6} , 
{32'hF9CFE5D8 , 32'h081FB830 , 32'h07B2A8E0 , 32'h18D88320 , 32'h1032C4C0 , 32'h00DB120F , 32'h1F0096C0 , 32'hDF6A6E00 , 32'h1C9B2DE0 , 32'h1DB7BA60 , 32'h10ED4000 , 32'h09080340 , 32'h213E5B40 , 32'h010FC2C0 , 32'h003AA163 , 32'hEFFA0B40 , 32'h033642CC , 32'h115B3240 , 32'hFA1ABA78 , 32'h032AAC78 , 32'h18B7E440 , 32'hF5832190 , 32'h14370DA0 , 32'h11ED61E0 , 32'hEFD99E60 , 32'hF2E7BEF0 , 32'hEBDE6DE0 , 32'hF14CF5C0 , 32'hF8C68930 , 32'hFB4B70D8 , 32'hF915F2F0 , 32'h0B770EF0 , 32'h0DBB7EA0 , 32'h1168D9C0 , 32'hFCA32B44 , 32'hFA2A5318 , 32'h0B1E9770 , 32'hEFB38E80 , 32'h0C513310 , 32'h13D4CCC0 , 32'h039F5B20 , 32'hF72BCA30 , 32'h0468EAD8 , 32'h062AEF98 , 32'hFE04C808 , 32'h1D826A00 , 32'h08EE58D0 , 32'h02C63C98 , 32'h04CF23A8 , 32'h04D68188 , 32'h089CD1C0 , 32'hFF250845 , 32'hF4F15730 , 32'h0A3DC010 , 32'h01AB4C30 , 32'h0ADF5BF0 , 32'h20CE9080 , 32'h0E439590 , 32'hDB7B8340 , 32'h0692AC08 , 32'h01C40AA0 , 32'hF1865310 , 32'hFB5505B8 , 32'h08BBD180 , 32'h027D4764 , 32'h002DFEA5 , 32'h036CB318 , 32'h09EBA670 , 32'h08C76A40 , 32'hF5F24EF0 , 32'hF981A110 , 32'hFD04DFC4 , 32'h05E462D8 , 32'h075C54F0 , 32'h02712FDC , 32'h0C3A43F0 , 32'h0146E6AC , 32'hFE6BA0CC , 32'hFF1A41B4 , 32'hFE79D2D8 , 32'h0DC8DE90 , 32'h015CD5EC , 32'hFAC07DD0 , 32'hFF010051 , 32'hFF72F84A , 32'h03E670CC , 32'h0249A484 , 32'hFE759054 , 32'h0417C388 , 32'hFF3FC5AF , 32'hFFF9C0BB , 32'hFFFF692B , 32'hFFFB5684 , 32'h00037B80 , 32'hFFFFAF74 , 32'hFFFF096A , 32'hFFFB8010 , 32'hFFFCA46D , 32'h0003994B , 32'h00032181} , 
{32'h0002AFE2 , 32'h000063AC , 32'hFFFC12FF , 32'hFFFE5442 , 32'h00055C8F , 32'h0000F8A8 , 32'h0001AEB8 , 32'h000762AF , 32'h0005E9E7 , 32'hFFFEB393 , 32'hFFFEA7BF , 32'h0007D2F5 , 32'h0002D40B , 32'hFFFBC9D2 , 32'hFFFFCD70 , 32'hFFFC3EE5 , 32'h00030B94 , 32'h0002FD47 , 32'h0000B8D4 , 32'h0002A462 , 32'hFFFD9120 , 32'h00027738 , 32'h0000DD5C , 32'hFFFBE475 , 32'hFFFCF70F , 32'h0006A262 , 32'h0004C866 , 32'hFFFCF4CF , 32'h0000BAC7 , 32'hFFFC2707 , 32'hFFFBC3A9 , 32'h000308BB , 32'h00006646 , 32'h00022123 , 32'h00022056 , 32'hFFF72C00 , 32'h00068F12 , 32'h00021E7A , 32'hFFFE9598 , 32'hFFFE8064 , 32'hFFFB2B9E , 32'hFFF8BDEE , 32'h0003679A , 32'hFFFF5FE7 , 32'hFFFF402E , 32'h0004AD9D , 32'hFFFB6220 , 32'hFFFE1DB7 , 32'h0000D81A , 32'hFFFE4D0A , 32'hFFFACF21 , 32'h0004B5C1 , 32'h0001328F , 32'hFFFEE6C7 , 32'hFFFECB8D , 32'hFFF6553E , 32'hFFFC611D , 32'h000821C2 , 32'h0009767E , 32'hFFFCA950 , 32'hFFFB340C , 32'h0004E534 , 32'h0002E9C3 , 32'h00037E5F , 32'h0002A519 , 32'h0007C2C7 , 32'h00006608 , 32'hFFFDCAFC , 32'h0000CE74 , 32'h000536B8 , 32'hFFFD78F1 , 32'h00055B9A , 32'h000412A3 , 32'hFFFF04F8 , 32'h0009DB7C , 32'h00043F42 , 32'hFFF93AAB , 32'h0004180F , 32'h0005F384 , 32'h0000BDAA , 32'h0003369E , 32'h00016C6D , 32'hFFF94C5C , 32'hFFFD1FFA , 32'hFFFC4FD8 , 32'hFFFE0020 , 32'hFFFEAED6 , 32'hFFFD97BF , 32'h00073AA6 , 32'h00078E77 , 32'h00083CFE , 32'hFFF894E2 , 32'h0006D2D2 , 32'hFFFC9C3B , 32'hFFFF7734 , 32'h00000D5D , 32'h00011178 , 32'hFFFF4356 , 32'h0003FCFE , 32'h00057966} , 
{32'h00050642 , 32'h000334FF , 32'hFFFC15F0 , 32'hFFFC9EFE , 32'h000584B8 , 32'h0000A540 , 32'h0002B733 , 32'hFFFB9CFA , 32'h000236E0 , 32'h0001C568 , 32'h00059288 , 32'h0001891C , 32'h000049BB , 32'h0001B046 , 32'hFFFAF755 , 32'hFFFBB968 , 32'hFFFFF2C5 , 32'h0002D47F , 32'h00044690 , 32'hFFFB6ADA , 32'hFFFE7685 , 32'h0000881A , 32'hFFFCC406 , 32'h000037ED , 32'hFFFDBF92 , 32'hFFFB74D7 , 32'hFFF65378 , 32'h0003C025 , 32'h0001200A , 32'hFFFA3EAC , 32'hFFF92EDF , 32'h00052019 , 32'h0003024B , 32'h00060662 , 32'h00058EB7 , 32'h000028F8 , 32'h0006009D , 32'hFFFF1D4D , 32'h0001D9B5 , 32'h000564C4 , 32'h00008809 , 32'h00039FD0 , 32'hFFFFF86C , 32'h000589BA , 32'h000646AA , 32'hFFFB70B7 , 32'h00029038 , 32'h0004E123 , 32'h0004BD75 , 32'hFFFE5700 , 32'hFFFAD008 , 32'h0002E32A , 32'hFFFB3894 , 32'h0001D43E , 32'hFFFC89DE , 32'hFFFDBBF6 , 32'hFFF70EAC , 32'hFFFF2BEB , 32'h00010D82 , 32'h00056935 , 32'h000229B2 , 32'hFFFED65E , 32'hFFFA559B , 32'hFFFB97D3 , 32'hFFF734B6 , 32'hFFFD3E51 , 32'h00070D58 , 32'hFFFF663D , 32'h0001075B , 32'h00003B4D , 32'hFFFDDB7A , 32'hFFFE7EC1 , 32'hFFFCDC86 , 32'h0003394F , 32'hFFFD3793 , 32'h0007218A , 32'h0003D4D4 , 32'hFFFA05CA , 32'h00005357 , 32'h00001DFA , 32'hFFFA2344 , 32'hFFFF553A , 32'h000543C3 , 32'h000ABFF9 , 32'hFFFF6AF6 , 32'hFFFA95C4 , 32'hFFFE92FE , 32'h00047B3D , 32'h00058C65 , 32'hFFF8E618 , 32'hFFFFC9DC , 32'h000698A7 , 32'hFFFD669A , 32'hFFFFE8CC , 32'hFFFC2D39 , 32'hFFFB9445 , 32'hFFF8B04E , 32'hFFFBA86B , 32'hFFFEAB8B , 32'hFFFD90C3} , 
{32'hCCE14700 , 32'h4989F680 , 32'h118B2CE0 , 32'h143A78E0 , 32'h2905E640 , 32'h0594ACB8 , 32'h3F95D4C0 , 32'h70C79500 , 32'hE57ECB60 , 32'h03B899F4 , 32'h063498C0 , 32'hF564FA20 , 32'h18D91560 , 32'hF65E7AE0 , 32'h1898F360 , 32'h0F1349B0 , 32'h01BB63F8 , 32'h129A52A0 , 32'h21212300 , 32'h01714840 , 32'hFAA30FC0 , 32'h0F31C1E0 , 32'hFB5DF680 , 32'h16A3CA40 , 32'h1DD218E0 , 32'hEA9F5AC0 , 32'h1CE215E0 , 32'h09C56A90 , 32'hEB3B3A20 , 32'hFF63171E , 32'h0935BFD0 , 32'h0AEE8490 , 32'hF69D5D00 , 32'hE7556240 , 32'hF6FE8000 , 32'hF99869A0 , 32'h052219B0 , 32'h059A8880 , 32'hF5033DE0 , 32'h0DEEC580 , 32'h1D30E820 , 32'h1A2287C0 , 32'hFA030D90 , 32'h16BF7A60 , 32'h00F8CD56 , 32'hE993D360 , 32'hF73A0030 , 32'hEC449C40 , 32'hF8690190 , 32'h0DEA8210 , 32'hFBF49C38 , 32'h027D76C4 , 32'h10472160 , 32'hEA635340 , 32'h040169D0 , 32'hF9D7ACB8 , 32'h00ED6578 , 32'hF9DDFA40 , 32'h03B015CC , 32'h083B67C0 , 32'hFBB4FD70 , 32'h0A4608B0 , 32'hF5FD5B00 , 32'h106EE9E0 , 32'hFD2FADD4 , 32'hEAA170A0 , 32'hFEC2AA1C , 32'h03C07F5C , 32'hF8FF77D0 , 32'h058F84B8 , 32'h0AB345B0 , 32'hF99EBFD0 , 32'h00046DC4 , 32'hFD45CFA0 , 32'hFCA21080 , 32'hFE526944 , 32'hFFCEEB75 , 32'hF445E0E0 , 32'hFF9BC768 , 32'hFBFFD670 , 32'h038AF6C8 , 32'h05A72F58 , 32'h0349CD34 , 32'h006B7583 , 32'h035655E4 , 32'hFB5F55F0 , 32'h0201E2E0 , 32'hFEC7322C , 32'hFD8D397C , 32'hFECADF34 , 32'h000150F5 , 32'hFFFFD8D8 , 32'h0001F33F , 32'h0000F49C , 32'hFFFD2B4D , 32'hFFFF800B , 32'hFFFD0B04 , 32'h00017EE3 , 32'h00038D71 , 32'hFFFF698A} , 
{32'h0753C820 , 32'h16551EC0 , 32'h013D80F0 , 32'hD9147740 , 32'h053B8DE8 , 32'hDA030200 , 32'h53DCEF80 , 32'hBC497F00 , 32'h27413840 , 32'h24E75DC0 , 32'hEC2F1BC0 , 32'hFCA2A00C , 32'h069234A8 , 32'hF9186F08 , 32'hDB3636C0 , 32'hF586F720 , 32'h15D28340 , 32'h23EE16C0 , 32'hDE794080 , 32'h0D5D3630 , 32'hFECE99C4 , 32'hFA297430 , 32'hEED05D60 , 32'h1DD6C1A0 , 32'h05C208C0 , 32'h1A0CB320 , 32'h10085C60 , 32'hE6AC3B60 , 32'hE6E55740 , 32'h145BA260 , 32'h0E6A25E0 , 32'h0E599E20 , 32'h074B73A8 , 32'h27BBBE80 , 32'hE9F07240 , 32'h03DF55C0 , 32'hF0949460 , 32'hF775A560 , 32'hF86966B8 , 32'h00DE1AE3 , 32'h1B9583C0 , 32'h10EBED80 , 32'h18AFEF00 , 32'h0D098860 , 32'hEDFA9300 , 32'h0BD075E0 , 32'h07274890 , 32'hEAF65B80 , 32'hF6B3C4A0 , 32'hE9D99FE0 , 32'h17B59920 , 32'hF9D75EF8 , 32'hF6BF3C40 , 32'hE95A9B00 , 32'h1C41C100 , 32'hF3440B00 , 32'h09405EC0 , 32'h0D1A06A0 , 32'h1471C6A0 , 32'h05799360 , 32'h01E5B730 , 32'hFB8D0978 , 32'hFB527098 , 32'hFEB89D80 , 32'h00E70B21 , 32'h0881BAA0 , 32'h0854DC30 , 32'h044922D8 , 32'hF921B5A8 , 32'h03E9CF3C , 32'h0F4BEBF0 , 32'hFCD7C344 , 32'hEDA98D20 , 32'h05F8B8E8 , 32'hFD563F70 , 32'h0589D328 , 32'h00A1375E , 32'h01E335A4 , 32'hFE568430 , 32'hFF86512F , 32'hF973BDF0 , 32'hF806CF70 , 32'h019D79C8 , 32'hFF09E789 , 32'hFF0A820E , 32'h011A65F4 , 32'h06CC8F78 , 32'hFB29B3E8 , 32'h04790C38 , 32'hFE979D84 , 32'hFFF8B299 , 32'hFFF9802A , 32'h00022B11 , 32'hFFFC4117 , 32'h00020CB8 , 32'h0000B878 , 32'hFFFBC20D , 32'hFFFDD454 , 32'hFFFDF724 , 32'hFFFB0AF9} , 
{32'hFFFFC896 , 32'h0005EC1E , 32'hFFFE96D5 , 32'h00021E14 , 32'h0005A102 , 32'hFFFAB165 , 32'hFFF9CCC6 , 32'hFFFEBD1F , 32'hFFFDE739 , 32'hFFFD1E06 , 32'hFFFC8D8C , 32'hFFFC5245 , 32'h00013A9D , 32'hFFFC6C7E , 32'hFFFFE0EE , 32'h00005589 , 32'hFFFEE09B , 32'h00056D93 , 32'hFFFDE7F5 , 32'hFFFBA077 , 32'h000522BC , 32'hFFFFA28E , 32'h00016220 , 32'hFFF6EC58 , 32'h000058FB , 32'h000593F5 , 32'hFFFFE5D5 , 32'hFFFF4543 , 32'h000062CA , 32'h0002AB5A , 32'h000005B9 , 32'hFFF8B014 , 32'h00063F1F , 32'hFFFFF8EB , 32'h0001E02B , 32'hFFFC9742 , 32'hFFFDAD99 , 32'hFFFE04AD , 32'h0003C426 , 32'h0001F563 , 32'hFFFE0A9A , 32'h0003A3BF , 32'h000C0D9F , 32'h0003F4D8 , 32'h00078921 , 32'hFFFF43AF , 32'hFFFFCE84 , 32'h0000EED0 , 32'hFFFE6C36 , 32'hFFFF1B56 , 32'hFFFD4CDC , 32'hFFF060D1 , 32'h00011522 , 32'hFFFF29B4 , 32'hFFFC6583 , 32'h00029C88 , 32'hFFFD0091 , 32'hFFFC7EDE , 32'hFFF38883 , 32'hFFFFEF23 , 32'hFFF94BE4 , 32'h00047056 , 32'h000433C3 , 32'h000788AA , 32'h00020F7B , 32'h0009A88B , 32'hFFF76024 , 32'h00017F26 , 32'hFFFE07CD , 32'hFFF60049 , 32'hFFFFBE23 , 32'h0004C4DD , 32'h00015B25 , 32'h00015E10 , 32'hFFFCA162 , 32'h00053C82 , 32'hFFFE5665 , 32'hFFF734E5 , 32'h0008CAC7 , 32'hFFF94F49 , 32'hFFFDE111 , 32'hFFFED6E3 , 32'hFFFE2DCB , 32'hFFFE4389 , 32'hFFFB24CB , 32'h0001E5F2 , 32'hFFFC3677 , 32'h0001CF76 , 32'h00079886 , 32'hFFF5FD21 , 32'hFFFF7E1C , 32'hFFFFA8EF , 32'hFFFCEB23 , 32'hFFF9F848 , 32'h000231CD , 32'h00018A94 , 32'h0003784F , 32'hFFFB5698 , 32'hFFF5C28E , 32'h00000C83} , 
{32'hFFFD3725 , 32'hFFFDF024 , 32'h00090FE5 , 32'h0004C9C4 , 32'hFFFE12B2 , 32'hFFFD795F , 32'hFFFEBFAA , 32'h000A94AE , 32'h00095954 , 32'h0002B408 , 32'hFFFAB73C , 32'hFFFE2544 , 32'hFFFD8493 , 32'h0007D0C1 , 32'hFFF9DD17 , 32'h00039537 , 32'hFFF6BB70 , 32'h0000FE70 , 32'h00001AC1 , 32'h00040241 , 32'hFFF5582A , 32'hFFFD06D7 , 32'hFFFA37B9 , 32'hFFFC663F , 32'h0000451C , 32'h00047B75 , 32'hFFFA8C82 , 32'hFFFC5A37 , 32'h000382D9 , 32'hFFFF5C1D , 32'h000168BE , 32'h00072EAB , 32'hFFFD00AE , 32'h0001D417 , 32'h00047A02 , 32'hFFFAF318 , 32'h0002A05D , 32'h0004E85C , 32'hFFF5BFAB , 32'h0002C98D , 32'hFFF84E89 , 32'h000111B7 , 32'hFFF31D70 , 32'hFFF44F57 , 32'h000132D6 , 32'h0009FDAC , 32'hFFFE2E5A , 32'hFFFCBD38 , 32'hFFFD406D , 32'h0000950C , 32'h0005A592 , 32'h0000DAD0 , 32'hFFF5C187 , 32'hFFFA9C30 , 32'h00069916 , 32'hFFF71CA0 , 32'h00018445 , 32'h000C3611 , 32'h0004F826 , 32'hFFFF21F3 , 32'hFFFE0B50 , 32'h000540A2 , 32'h00049137 , 32'hFFFE4EAC , 32'hFFF8AF73 , 32'hFFFE32D3 , 32'hFFF656D7 , 32'hFFFBD58C , 32'hFFFE6DB8 , 32'hFFFA6B98 , 32'hFFFE7C65 , 32'h00028B99 , 32'hFFFE7645 , 32'hFFFEE6C8 , 32'hFFFC401E , 32'hFFF97842 , 32'hFFFB921C , 32'h000928FE , 32'hFFFCAD7B , 32'h00017A4C , 32'h00038CB5 , 32'h000AA842 , 32'h00071396 , 32'hFFFD0193 , 32'h00020754 , 32'h000726C4 , 32'h00033D04 , 32'h0005519D , 32'h000005EE , 32'hFFF97864 , 32'hFFFB8DF6 , 32'h00008C70 , 32'h000E005A , 32'h0006DAEB , 32'hFFFFA91A , 32'hFFFC3D93 , 32'h000366DB , 32'hFFFE7BA2 , 32'h0002145F , 32'hFFFF6B05} , 
{32'hFFFB976C , 32'h0006CF8E , 32'hFFFF025C , 32'hFFFE22A6 , 32'hFFFD1010 , 32'hFFFD8BF9 , 32'h00043E53 , 32'h0000B70D , 32'hFFFD9E17 , 32'hFFFBBA9D , 32'h00050740 , 32'hFFFF6E74 , 32'h00035373 , 32'h0006A4B4 , 32'hFFFFB69C , 32'h00028009 , 32'h00013EDB , 32'hFFFC1FE5 , 32'hFFFE2408 , 32'hFFFDFEAF , 32'h00062993 , 32'h000109F1 , 32'h0002A9F3 , 32'h0001444F , 32'hFFFC3EC6 , 32'hFFFB8DD8 , 32'hFFFAD4F9 , 32'hFFFE34AD , 32'h0003B6D4 , 32'hFFFE8AA2 , 32'h0004C013 , 32'hFFF9ED95 , 32'hFFF95526 , 32'h00001928 , 32'h00037461 , 32'h00049676 , 32'hFFFFAD15 , 32'h000302F4 , 32'hFFFEB796 , 32'h00025D5E , 32'hFFFCBE2A , 32'hFFFEA3EE , 32'h0003B1A8 , 32'h0001FFF7 , 32'hFFFDB8FA , 32'hFFF99F77 , 32'h000240B9 , 32'hFFF9E367 , 32'h00097ABC , 32'hFFFE9C0E , 32'hFFFCB59B , 32'hFFFC748F , 32'hFFFC24E7 , 32'h00024360 , 32'h00014CAB , 32'hFFFE4131 , 32'hFFFACA63 , 32'hFFFA706C , 32'h00084DA1 , 32'hFFFF95E2 , 32'h0000DCF1 , 32'hFFFB547B , 32'hFFFD6151 , 32'h0001005B , 32'h00054A47 , 32'h0003C096 , 32'hFFFDC6B1 , 32'hFFFC026A , 32'h00022D63 , 32'h00008A05 , 32'h00076EFF , 32'hFFFE1383 , 32'h00044F87 , 32'h0006AA7C , 32'h0004987F , 32'hFFF8AA41 , 32'h0002A56C , 32'h0004DF1B , 32'hFFF8D4CB , 32'h0008EAD9 , 32'h0003F377 , 32'hFFFBB28F , 32'h00022494 , 32'h00141057 , 32'hFFFA0570 , 32'h000051F4 , 32'hFFFDC5B3 , 32'hFFFFE74C , 32'h0000657D , 32'h000294F2 , 32'h00017185 , 32'hFFFF3C94 , 32'hFFF7511C , 32'hFFFE5EF5 , 32'h000389CA , 32'h000427ED , 32'hFFFA65E6 , 32'h00090E05 , 32'h00047875 , 32'h0003332A} , 
{32'h00080C0C , 32'h0002FBEA , 32'h0004740A , 32'hFFF9F28E , 32'hFFFDF084 , 32'h000497BE , 32'hFFF96479 , 32'hFFFB13FB , 32'hFFFB8345 , 32'hFFFC0A6B , 32'h00055358 , 32'hFFFD1790 , 32'hFFF81814 , 32'h0002450D , 32'hFFFD824A , 32'h00007C82 , 32'h00045FC0 , 32'hFFFD16F2 , 32'h00015BF8 , 32'h00057C85 , 32'hFFFE5FD8 , 32'h0004B49F , 32'h000036D6 , 32'h000009A8 , 32'h0002FFE1 , 32'hFFFB24F0 , 32'h0001170B , 32'hFFFF260C , 32'h000352CD , 32'hFFFF3B79 , 32'hFFFA67BF , 32'h00018217 , 32'hFFFE0027 , 32'h00005734 , 32'h0004A84D , 32'h000251C4 , 32'h0003D77C , 32'h000387C8 , 32'hFFF5F839 , 32'h000AA675 , 32'h00020AD2 , 32'h000342D1 , 32'hFFFD1942 , 32'h00030E9E , 32'h0003D145 , 32'hFFFFB1A4 , 32'h00004DA6 , 32'hFFF8BD05 , 32'h00035085 , 32'hFFFC7FBD , 32'h0006FD51 , 32'h00062410 , 32'hFFFD563A , 32'hFFFDDA73 , 32'h0000306B , 32'h0006BA46 , 32'h00016B8F , 32'hFFF9A3A3 , 32'hFFFA690A , 32'h00013EE0 , 32'h00061AE3 , 32'h00002491 , 32'h0005E7C6 , 32'h0000722D , 32'h0003EDE8 , 32'h00037017 , 32'hFFFB804C , 32'h000153EB , 32'hFFFE7C50 , 32'h00006651 , 32'hFFFA2C84 , 32'h0002FE3D , 32'h0003B682 , 32'h00028FFA , 32'h0005E002 , 32'h00049255 , 32'h000609EE , 32'hFFFE91D5 , 32'h00063E88 , 32'h00023A6D , 32'h00023313 , 32'hFFF7777B , 32'h000174BC , 32'h0001EBFB , 32'h00071702 , 32'h0005F087 , 32'hFFFE93D7 , 32'h000351EF , 32'hFFFB689C , 32'hFFFED31B , 32'h00013360 , 32'hFFFC2EC6 , 32'h000822B2 , 32'hFFFFDFFE , 32'h00099FA4 , 32'h00021455 , 32'h00015412 , 32'hFFFC0B12 , 32'hFFFCA2BA , 32'hFFFFB158} , 
{32'hFFFB5940 , 32'hFFF71314 , 32'h0006A07D , 32'hFFFB7FBD , 32'hFFFD8D34 , 32'h00059C9F , 32'hFFFBF325 , 32'h0002FB0B , 32'hFFFEDE6A , 32'h00077059 , 32'hFFFFEFE5 , 32'hFFFE2827 , 32'h0005B8B2 , 32'h00016B7F , 32'hFFFFE1C5 , 32'hFFF8CA45 , 32'hFFFF9CCB , 32'h0004AA1A , 32'hFFFF8162 , 32'hFFFE0A80 , 32'h00051769 , 32'h00020DF1 , 32'hFFFE9931 , 32'h00002993 , 32'hFFFB35E5 , 32'hFFFC85DC , 32'hFFF7C1F7 , 32'h0006EF99 , 32'h00009C05 , 32'h00027412 , 32'hFFFAAB7F , 32'h00046144 , 32'h00021F7E , 32'hFFFCEDA4 , 32'hFFFF11CE , 32'h00005680 , 32'hFFFE7274 , 32'hFFFD6D8F , 32'h0008E40E , 32'h000162D5 , 32'h00011E0B , 32'h0004D69D , 32'h00048646 , 32'hFFFD7A8E , 32'hFFFED378 , 32'h00035127 , 32'h00036009 , 32'hFFFF9254 , 32'hFFFF16AF , 32'hFFF7D5FD , 32'hFFFFDE4E , 32'h00009880 , 32'hFFFEC5D4 , 32'hFFF035C9 , 32'hFFFD31F0 , 32'hFFF84C8D , 32'hFFF46F4C , 32'h0000F1BB , 32'hFFFB672F , 32'hFFFF68AF , 32'hFFF9EBA5 , 32'hFFFD1616 , 32'hFFFAC20C , 32'hFFFEEBE1 , 32'h000364B7 , 32'h0000D498 , 32'hFFFD62AD , 32'h00038361 , 32'h0000ADE5 , 32'h0008F52A , 32'hFFFF0981 , 32'h000373FB , 32'h00022326 , 32'hFFF74766 , 32'hFFF95395 , 32'h0005495E , 32'h0003374F , 32'hFFF8783E , 32'hFFFF0D33 , 32'h0000978B , 32'hFFF51B1A , 32'h0004856F , 32'hFFFD356B , 32'h00040600 , 32'hFFFE9EA0 , 32'h0001D176 , 32'h0003697B , 32'h0003AA2B , 32'hFFFEA537 , 32'hFFFF76CE , 32'h00031729 , 32'hFFF7EEAD , 32'hFFFE328C , 32'h00019D0C , 32'h0005C8A1 , 32'hFFFDCB1C , 32'h0001FAAE , 32'hFFFD4B83 , 32'h00050E47 , 32'hFFF9C408} , 
{32'hDA686A40 , 32'h0028ED90 , 32'h13A50A80 , 32'hF8456420 , 32'hF02B3EA0 , 32'h24506EC0 , 32'hE6BF5960 , 32'h169B9A00 , 32'hDAFACA40 , 32'h0449AEA0 , 32'hEBA5C260 , 32'h2B640400 , 32'hE16884C0 , 32'hDD1D8800 , 32'hFC1C4D38 , 32'hFEE8E4C4 , 32'hE54D9500 , 32'hFCF800B0 , 32'h1C6E7B40 , 32'hF58BC9A0 , 32'hFFD3CAD4 , 32'h0A0FB900 , 32'hF8B8CC08 , 32'h0B861260 , 32'h0E3A0560 , 32'h02C59A68 , 32'h15A8C1C0 , 32'h0CFE29F0 , 32'h00CB6855 , 32'hF15D1380 , 32'hE1F31CE0 , 32'h0C995180 , 32'hFB9E3C60 , 32'h0E6B4580 , 32'h09EE3340 , 32'h07E429A0 , 32'hE985B020 , 32'h06F7DD48 , 32'h0C4DADE0 , 32'hFC66F438 , 32'hF2CC2A20 , 32'hFFBE2209 , 32'h0C59CF40 , 32'hFB31F438 , 32'h0CFF0430 , 32'hF80FF5E8 , 32'hF1398930 , 32'hFAE5F800 , 32'h083A2A80 , 32'h02339B3C , 32'hF7214620 , 32'hFC92E034 , 32'hFD285514 , 32'hED6E04E0 , 32'hFF028B56 , 32'h03F24DA4 , 32'h008694AF , 32'h0426EA20 , 32'h11AD6860 , 32'hF77927E0 , 32'h0AA89810 , 32'hF5DD8F00 , 32'hF4DBDF90 , 32'h04B09DE8 , 32'h1031D3E0 , 32'h02E19784 , 32'h107187E0 , 32'h111972A0 , 32'h00AB2EBD , 32'h0ACCFD90 , 32'hF68E2B80 , 32'hFA187240 , 32'h02A2370C , 32'h090F1690 , 32'hFCB1DB14 , 32'hFB0D5878 , 32'hFB71C3A8 , 32'hFCB30A88 , 32'hFE5D7AB4 , 32'h0526E958 , 32'hFF23AC79 , 32'hFD9C3834 , 32'hF6096D20 , 32'hFD41E9EC , 32'hFE236300 , 32'hFFCF3988 , 32'hFDFA3DA4 , 32'h023540C8 , 32'h00457433 , 32'hFFF04C08 , 32'hFFFDC05E , 32'h000294DF , 32'hFFF88EE6 , 32'h00063A85 , 32'h0005214F , 32'h00059F72 , 32'h00014D8F , 32'h00034D42 , 32'hFFFDD35D , 32'hFFFE079B} , 
{32'hDC91B500 , 32'h1834E260 , 32'h0158E638 , 32'hE4825A40 , 32'hCF960C80 , 32'hEA36A9A0 , 32'h1858B380 , 32'hE7B84F60 , 32'h00850A9F , 32'h17CF2A40 , 32'hFBACD1B0 , 32'h21A9B840 , 32'hC75F4A00 , 32'h08C76EC0 , 32'h1BED9160 , 32'hDF4D0280 , 32'hE2F66180 , 32'h2192B340 , 32'hE5FF67C0 , 32'h120BB700 , 32'h0B895EF0 , 32'h058371B0 , 32'hEA8BC2A0 , 32'hF2518EF0 , 32'hDC6C1700 , 32'hE8A22340 , 32'h22D263C0 , 32'h0846B800 , 32'h0859EC60 , 32'h1D9155E0 , 32'h0F647750 , 32'hD00F8D00 , 32'h139A9960 , 32'h0F960F30 , 32'hF75EDDE0 , 32'hEA43AAC0 , 32'h1530B620 , 32'h1D9AEBE0 , 32'h0658B5F8 , 32'hFBE9F718 , 32'h06C88ED8 , 32'h0564ADE8 , 32'h13C3A380 , 32'h0628B140 , 32'h0727C230 , 32'hF11D7400 , 32'h16B54020 , 32'hF563C2C0 , 32'hF7073240 , 32'hF3444000 , 32'h123CE9C0 , 32'h0F82C7E0 , 32'hDA59A500 , 32'hFBED4440 , 32'hF73B11D0 , 32'hFE4B9C34 , 32'hF69BAD10 , 32'hF8694818 , 32'hFCB0A6EC , 32'hFBD18050 , 32'h01179D7C , 32'hFBCE41D8 , 32'h0520C890 , 32'h0F7B7750 , 32'h108EEC20 , 32'hF7195FC0 , 32'hF250EDA0 , 32'h0F0863A0 , 32'hFD9ECF90 , 32'h066EC798 , 32'hFAE242F8 , 32'h03AE3A44 , 32'hFCDA2E84 , 32'hFDDA5220 , 32'hFDF92E90 , 32'hFBE93F68 , 32'h0033117B , 32'h04F12E90 , 32'h006204C7 , 32'hFCD195BC , 32'h06F7BC10 , 32'hF8A11590 , 32'h08732540 , 32'hF44FADA0 , 32'h0351DA1C , 32'hFAE123D0 , 32'h004FDF42 , 32'h060588F8 , 32'h02E384DC , 32'h0131C6A8 , 32'h00084DC4 , 32'h00017D60 , 32'hFFFD34E3 , 32'h000211F8 , 32'h0001131B , 32'hFFFD05C3 , 32'hFFFF2421 , 32'hFFFC59A1 , 32'h0001CB24 , 32'h000341C0} , 
{32'hFFFC70B0 , 32'h0000F45F , 32'hFFFEAF2E , 32'hFFFE824A , 32'h000000EF , 32'h0000EF5E , 32'h00071477 , 32'h000078B9 , 32'h0003CA35 , 32'hFFF517BC , 32'h000089E6 , 32'hFFFDE3BF , 32'h0002ECFA , 32'h0000B43E , 32'hFFFE99B8 , 32'hFFF7D881 , 32'h000999EA , 32'h000F66EF , 32'hFFFFE381 , 32'h00067522 , 32'h0000CCD0 , 32'hFFF88704 , 32'h0003B861 , 32'h0001F411 , 32'h00017CBD , 32'hFFFF5A51 , 32'h0000F889 , 32'h00013B40 , 32'h0005DC96 , 32'hFFFED829 , 32'hFFF84A23 , 32'hFFFE1374 , 32'h0009D836 , 32'h000599A1 , 32'h00012C11 , 32'hFFF75F37 , 32'h00017A1E , 32'hFFF5E56C , 32'hFFFE7C06 , 32'h00085C2C , 32'h00070023 , 32'h000181AE , 32'hFFFFA034 , 32'h0004620A , 32'h000306C3 , 32'h0002064E , 32'hFFFA96DF , 32'hFFFFB1F4 , 32'hFFFB507D , 32'h00026395 , 32'hFFFEE311 , 32'hFFFC851F , 32'h000448BB , 32'h0004794D , 32'hFFF0A388 , 32'hFFFE21D5 , 32'h0008693B , 32'h00065F2B , 32'hFFFEA8D7 , 32'h000389B3 , 32'h000AA5E7 , 32'hFFFC5524 , 32'h0003B6F2 , 32'hFFFC2151 , 32'h0002D791 , 32'hFFFE2BF7 , 32'h00016244 , 32'h0000B2BE , 32'hFFFDB215 , 32'hFFFF4F45 , 32'hFFF8FB2A , 32'hFFFC3F41 , 32'h00027C5F , 32'h000095EE , 32'h00014781 , 32'h000282EF , 32'hFFFE4277 , 32'hFFF826A1 , 32'h0007B92C , 32'h00076113 , 32'h00002DCC , 32'hFFFCEE41 , 32'hFFF40086 , 32'h00028B4A , 32'hFFFD315E , 32'hFFFFF2BE , 32'h000052D0 , 32'h0000A155 , 32'hFFFCC535 , 32'hFFFBC44A , 32'hFFFF639C , 32'h00000C73 , 32'h0007321F , 32'h00002CD3 , 32'hFFFF32B6 , 32'h0003E143 , 32'h000638DF , 32'h00096351 , 32'hFFFF33DB , 32'hFFF723F9} , 
{32'h0002D39E , 32'hFFFDDBCD , 32'h0001304C , 32'h00017C81 , 32'h000259D8 , 32'hFFFD2139 , 32'h0008F37C , 32'hFFFF807F , 32'h00098384 , 32'h000031F2 , 32'h0002A8F9 , 32'h00070D0C , 32'hFFFF6C46 , 32'h0001788B , 32'hFFFDC495 , 32'hFFFC354C , 32'hFFF81364 , 32'hFFFB98BC , 32'hFFFFD4E5 , 32'h0000404E , 32'h0005AF11 , 32'hFFFC2BC8 , 32'hFFFFD462 , 32'hFFFF819F , 32'h00064493 , 32'hFFFD4067 , 32'hFFFE2F78 , 32'h0001CD70 , 32'hFFFAF6ED , 32'hFFFFDE39 , 32'h0005FC33 , 32'hFFFDC26B , 32'hFFFCE822 , 32'hFFFD3D90 , 32'hFFFC6D5F , 32'h00071BB6 , 32'h000079C7 , 32'hFFFD3B1D , 32'h00074C94 , 32'hFFFC6CF4 , 32'h00034F1B , 32'h0000541B , 32'h00012368 , 32'h00003BD8 , 32'h00038201 , 32'hFFFEA259 , 32'h00027749 , 32'h0009A0F0 , 32'h0002F35F , 32'h0002AABF , 32'h00047718 , 32'hFFFB197B , 32'h0001B636 , 32'h00074E9A , 32'h0004C5C6 , 32'h0004547E , 32'h00009E0C , 32'h00021CE7 , 32'h0001DA99 , 32'h0002B529 , 32'h00017AFD , 32'hFFF88BC3 , 32'hFFFCCAB2 , 32'h00009832 , 32'hFFFF0333 , 32'h000105CF , 32'hFFFC7892 , 32'hFFFE0160 , 32'h0004148B , 32'hFFFF8036 , 32'hFFFEAD4E , 32'h0009FAD1 , 32'hFFFE12E6 , 32'hFFFDE5D4 , 32'hFFF8AAFA , 32'hFFFEC3B7 , 32'hFFFD5D4F , 32'h0002562E , 32'h00040C1A , 32'h0003277C , 32'hFFFFF0A9 , 32'hFFFE5057 , 32'h00032A78 , 32'h00065DE9 , 32'hFFF8A7CA , 32'hFFFBA7D8 , 32'hFFFC32AA , 32'hFFFF1090 , 32'hFFFDFE16 , 32'h0004EA5B , 32'h0004304B , 32'hFFFA2337 , 32'h000459AB , 32'h000144EC , 32'hFFFDC38D , 32'hFFFF03AD , 32'h000017D2 , 32'hFFFB9036 , 32'h00009033 , 32'hFFFED36A} , 
{32'h7FFFFFFF , 32'h25C6D1C0 , 32'h76415A80 , 32'h3273C600 , 32'h9609C000 , 32'hFA15AD18 , 32'h17573680 , 32'h3A755E80 , 32'h14DFB5A0 , 32'hFE7982B0 , 32'h01EEFEB0 , 32'h0AFDE0A0 , 32'h25AEB5C0 , 32'h26AE6440 , 32'hFD4C6880 , 32'h078E5818 , 32'hD4931540 , 32'h0EEE2F80 , 32'hE53BE660 , 32'hE76F04E0 , 32'h03425E10 , 32'h0F864EE0 , 32'h07999CA8 , 32'hE3C6D0E0 , 32'h07D61C60 , 32'h0E4A8CC0 , 32'hF6179780 , 32'h0FE5AF00 , 32'h1DA0BCC0 , 32'hEAA1DF00 , 32'hE60A7640 , 32'h1E913C20 , 32'h1A7FC640 , 32'h01DC4B84 , 32'hE2BFB480 , 32'h0E51A1B0 , 32'h05F279E8 , 32'h1AC8A6E0 , 32'h0DDA1110 , 32'hE02D2400 , 32'h1235BE40 , 32'h1226E580 , 32'h01864ED4 , 32'h1D63F280 , 32'h033D9B18 , 32'hF9619AB0 , 32'hFBB2BEF0 , 32'h05A587A8 , 32'h0E840A00 , 32'h03991600 , 32'h03B11E70 , 32'h0D3790F0 , 32'h085D2A00 , 32'hFBE9E390 , 32'h10FFA000 , 32'h06AEAB10 , 32'h0C56E680 , 32'h03DA25D0 , 32'h04E658A0 , 32'h095D6FB0 , 32'hFA7FF918 , 32'h0D35DB20 , 32'hF69C21E0 , 32'hF2F9DAB0 , 32'h0914F2E0 , 32'h0561D320 , 32'hFF12F983 , 32'hFBE547B0 , 32'h04784068 , 32'h08ED65F0 , 32'h023260F4 , 32'hFCDDCF58 , 32'hF231EC00 , 32'h03967004 , 32'h04F74E28 , 32'hFB74E6F0 , 32'h00FF17E0 , 32'h0590BEA0 , 32'h01465FD8 , 32'h099F5500 , 32'h022261A4 , 32'hFA897E18 , 32'h03C28EDC , 32'hFFB60BDF , 32'h02516480 , 32'hFF105757 , 32'h01D6B81C , 32'hFB487868 , 32'h01D4EE60 , 32'h0134D7BC , 32'hFFFBE491 , 32'h00012DB5 , 32'hFFFBCCCB , 32'hFFFD228D , 32'hFFFDBF64 , 32'hFFFAD977 , 32'hFFFEF5BF , 32'hFFFED209 , 32'hFFFFBFEE , 32'h0001FCEA} , 
{32'h261A8680 , 32'h1ABB8020 , 32'h3FC566C0 , 32'h18A8A800 , 32'hD8FFDE00 , 32'h1390D940 , 32'hE90698C0 , 32'h0E2F3660 , 32'h18A3C9E0 , 32'hFC91BA28 , 32'h0B49F2E0 , 32'h18657320 , 32'hF5514C20 , 32'h11D79E40 , 32'h2D484980 , 32'h04C9EC40 , 32'h09B5BA40 , 32'hF8E16718 , 32'h0A5DE320 , 32'h188031C0 , 32'hE9635C20 , 32'hF76A69C0 , 32'h02DCC49C , 32'h18546940 , 32'h07AE7968 , 32'hE81BFB20 , 32'h016A56B4 , 32'hFB5D5A00 , 32'hF49FBC00 , 32'h15DF04A0 , 32'h22073A00 , 32'h06F662A8 , 32'hE2E51BC0 , 32'hF8F43290 , 32'hF99C3A90 , 32'hF24E4110 , 32'h0507B0A8 , 32'h0C463520 , 32'h081EE7B0 , 32'h04BB3128 , 32'hF837AA60 , 32'hF2E5B370 , 32'hF2C5A770 , 32'h03FB86A8 , 32'h08F19A00 , 32'hF7848840 , 32'h03ADC1A8 , 32'hF3D33AB0 , 32'h00CE8915 , 32'h22FE6E80 , 32'h13AF9740 , 32'hF82C9700 , 32'hFCDA8F80 , 32'hFBD4F9C8 , 32'hF7A4EFD0 , 32'hFC5AACB0 , 32'h086516D0 , 32'h01836960 , 32'hED112B80 , 32'hF45F6D80 , 32'h13174320 , 32'hEE6EFC00 , 32'h02D8D528 , 32'hEEE38400 , 32'hF976BB98 , 32'hFCC21408 , 32'hF95BD730 , 32'hF9D03F00 , 32'hF7BAA1A0 , 32'h0825A3C0 , 32'h01CBEE70 , 32'hFAF5A348 , 32'hF5430840 , 32'hFCB12D18 , 32'h044239F0 , 32'hF8045908 , 32'hF2F45EF0 , 32'hFC7AACA4 , 32'h116A6260 , 32'hFFD16C4E , 32'hFA30E230 , 32'hFF2C5667 , 32'hFAA7BBB8 , 32'h02DCA6AC , 32'h0791A5B8 , 32'h06C07850 , 32'h07B27BC0 , 32'hFC2F8608 , 32'hFD08291C , 32'hFE460A4C , 32'h0001CE3B , 32'h00015A54 , 32'h00025AA0 , 32'hFFFF5B97 , 32'hFFFE7832 , 32'h0000D46C , 32'hFFFA75A2 , 32'hFFFEF426 , 32'hFFFEAFD3 , 32'h00005615} , 
{32'h00030599 , 32'h00007EFB , 32'h00013249 , 32'h00029B75 , 32'hFFFE5BB3 , 32'h0002E2FE , 32'h0008056C , 32'hFFFF5BC5 , 32'hFFFCCDB0 , 32'hFFFDA17D , 32'h0003C41C , 32'hFFFFD356 , 32'hFFF58B6D , 32'h000A1722 , 32'hFFFC748E , 32'hFFF9A147 , 32'h000052ED , 32'hFFF812E7 , 32'h0004451E , 32'hFFF8F030 , 32'h000201F2 , 32'h0002669D , 32'hFFFB05C5 , 32'h000036B7 , 32'h00038FAB , 32'h000585FB , 32'h0000BDC7 , 32'h0004054E , 32'hFFFD213E , 32'hFFFD5BFA , 32'h0005D416 , 32'h0007AB73 , 32'h00030A2A , 32'h00009930 , 32'h0004B089 , 32'h0000086E , 32'hFFFF081C , 32'hFFFA8E45 , 32'h00054BBB , 32'hFFFFD3FE , 32'h0001E6A3 , 32'hFFFFB9B1 , 32'hFFFBBD5D , 32'hFFF933F9 , 32'hFFFA259E , 32'h0002F430 , 32'h0004C702 , 32'hFFF96717 , 32'hFFFC57A5 , 32'hFFFCFF15 , 32'hFFFE4590 , 32'hFFFCA966 , 32'h00000ABB , 32'hFFFB4B5C , 32'hFFFF976B , 32'h00024B27 , 32'hFFFC18EC , 32'hFFF3E400 , 32'h0003EB09 , 32'hFFF960C0 , 32'hFFF9E387 , 32'h00065F14 , 32'h000733D5 , 32'hFFFCB7BA , 32'hFFFAECC1 , 32'h00064331 , 32'hFFFE4F8E , 32'hFFFC4880 , 32'hFFF8CFBE , 32'h00004917 , 32'hFFFFD15F , 32'hFFFE7F5B , 32'hFFFF9055 , 32'h0004AE3D , 32'h00012E12 , 32'h00032B5A , 32'h00064BED , 32'hFFFD3BE5 , 32'hFFFF55C2 , 32'hFFF6D0D3 , 32'h0003625A , 32'hFFFEAC94 , 32'h0004CE2B , 32'h0004F4D1 , 32'h0007F8FF , 32'h0002C817 , 32'h00007151 , 32'h00018646 , 32'h000249FA , 32'h0003666A , 32'h00014A87 , 32'h0000CC5E , 32'h0001B523 , 32'hFFFE18FE , 32'hFFFE191F , 32'h0005DEAD , 32'h000254E5 , 32'hFFFE950A , 32'h0000A94F , 32'h00003574} , 
{32'hFFFFC714 , 32'hFFFF3C5C , 32'hFFFA9CB0 , 32'hFFFF8CB1 , 32'h00002E40 , 32'hFFF9BB97 , 32'h000602B6 , 32'h0002F968 , 32'hFFFBB308 , 32'h00022B52 , 32'h00037C85 , 32'h00066B75 , 32'hFFFC6328 , 32'hFFFCD80D , 32'h0006EF3A , 32'hFFFCDB90 , 32'hFFFCA7EA , 32'hFFF8F18F , 32'h0004F3BA , 32'hFFFC8073 , 32'hFFFF8F58 , 32'hFFFAD0BB , 32'hFFFBFBB3 , 32'h00011A3C , 32'h0001143B , 32'hFFFB1DFC , 32'hFFFFC820 , 32'hFFFBA7DD , 32'hFFFB96F4 , 32'hFFF9D482 , 32'h0006EFC6 , 32'h00003FAB , 32'hFFFBFFB5 , 32'hFFFF7E9C , 32'hFFFFB20A , 32'hFFFA39A5 , 32'hFFFE4087 , 32'h0006E4EB , 32'hFFFF4EB1 , 32'hFFF86112 , 32'hFFFF81E3 , 32'h00051142 , 32'h0006A129 , 32'h00005BFE , 32'hFFFFE560 , 32'hFFFA8E24 , 32'hFFF60F38 , 32'h0003A6FF , 32'h000279AD , 32'h000974C1 , 32'h0002FE05 , 32'h00079F1F , 32'hFFFD7BA6 , 32'h000680EC , 32'hFFFC7AE0 , 32'h0007F0B1 , 32'h0000F3FC , 32'h0002B507 , 32'hFFF7EC22 , 32'hFFF5BA2A , 32'h00042BB8 , 32'hFFFB0862 , 32'hFFFB716A , 32'hFFFD03E4 , 32'hFFFCAFB5 , 32'hFFFABFF0 , 32'h0002DC93 , 32'h0003A4FB , 32'hFFFA736B , 32'h00086A85 , 32'h00050853 , 32'hFFFC1636 , 32'h00056553 , 32'h0002374E , 32'h0003C78C , 32'hFFF8C759 , 32'hFFFFFAF8 , 32'hFFFE2610 , 32'h0000C476 , 32'h0003DE61 , 32'hFFF3F719 , 32'hFFFC3F24 , 32'h0004DB6C , 32'h00003F4E , 32'hFFFF9B57 , 32'h00004FE9 , 32'hFFFBAACA , 32'h00041523 , 32'h0001747B , 32'hFFFDAAAE , 32'hFFFDD5C4 , 32'hFFFD52CB , 32'hFFFCD399 , 32'hFFF88FBF , 32'hFFFDD8D1 , 32'h00001B32 , 32'h00058CB4 , 32'h0001D22A , 32'hFFFC1B5D , 32'hFFF9909A} , 
{32'hD20E62C0 , 32'h1E70AA40 , 32'h030A938C , 32'h47949F80 , 32'hEA0C6F00 , 32'h0BD70B70 , 32'hF6F849A0 , 32'hF44BAC60 , 32'h10D1B120 , 32'hF4BB6A90 , 32'hF2827A00 , 32'h1771B240 , 32'h1D7EB7E0 , 32'hEABC06A0 , 32'h266E6100 , 32'hF17D5450 , 32'hF7C42950 , 32'h1E81EB80 , 32'hF1675D70 , 32'h05D4F8F0 , 32'hE4A44740 , 32'hF0C9F440 , 32'h0D7A21B0 , 32'h14B65F80 , 32'hF5A49D30 , 32'h20D54500 , 32'hF780C6E0 , 32'hDE0CCAC0 , 32'h01502240 , 32'h10035F40 , 32'hFCA49810 , 32'hEB48DA00 , 32'h18380E80 , 32'h01B7B2F8 , 32'h092D2BA0 , 32'hFF0768F0 , 32'h1F3AF600 , 32'h0906B4D0 , 32'hF9E92280 , 32'hE7992060 , 32'hEB5D1AE0 , 32'hFFB87714 , 32'hFF6CE906 , 32'h194F2FE0 , 32'hF80CA780 , 32'hFF47D3D2 , 32'h005A6F30 , 32'h021CCB34 , 32'hFC18963C , 32'h005FCF69 , 32'h0CC110B0 , 32'hF0E5E7A0 , 32'h0B2B05C0 , 32'hEF4383E0 , 32'hFA982BF0 , 32'h0970DBA0 , 32'h13FE39A0 , 32'h041D06D8 , 32'hF5545B40 , 32'hF5B68430 , 32'h0147C6EC , 32'hF5D63F70 , 32'hF4FF3A70 , 32'h0A8E90C0 , 32'h0C2018D0 , 32'h0A515290 , 32'hFF52A3D0 , 32'h094D3100 , 32'hF9E91AF8 , 32'hF786E9F0 , 32'h06E38338 , 32'hEFC9DFA0 , 32'h06416DE8 , 32'h052349B8 , 32'hF591C860 , 32'h01E471B4 , 32'h005E9064 , 32'hFEC9ABD8 , 32'hFC697FB4 , 32'hFCE58F0C , 32'hFCC886E8 , 32'hFF746926 , 32'hFC3F1764 , 32'hFD4DE368 , 32'h020BBC58 , 32'hFC0B5530 , 32'h017C9B2C , 32'hFF2C90F5 , 32'h0066DBAA , 32'h007624E9 , 32'h00066ADF , 32'h00024631 , 32'hFFFB0C25 , 32'hFFFCE054 , 32'h000465B6 , 32'h00073740 , 32'hFFFCAA4C , 32'hFFFF012F , 32'hFFFC9B10 , 32'hFFFECB66} , 
{32'h00011E36 , 32'hFFFB9A38 , 32'h0006B8D3 , 32'h00064B34 , 32'hFFFA7273 , 32'h0000D833 , 32'hFFFDF2F4 , 32'h00025DC9 , 32'hFFFB84BB , 32'hFFFB4614 , 32'h00031A86 , 32'h0006DC8F , 32'h00052734 , 32'hFFFB81C8 , 32'h0000AA06 , 32'hFFFDE5AB , 32'h0004E191 , 32'hFFFD56E5 , 32'h0004D1C8 , 32'h00010FEB , 32'hFFFBC2FA , 32'hFFFA21B8 , 32'h00031B46 , 32'hFFFE49E5 , 32'h000B0D68 , 32'h0007B3DE , 32'hFFFD58DE , 32'hFFFC0066 , 32'hFFFDFBD4 , 32'h00038243 , 32'hFFFCB3CE , 32'hFFFA759B , 32'hFFF442FD , 32'h00020A4C , 32'h0006B4EF , 32'h00018867 , 32'h0001592B , 32'h00014426 , 32'hFFFE61D9 , 32'hFFFE88E5 , 32'hFFFA3009 , 32'hFFF81AD2 , 32'h00081E3E , 32'h0002E2DF , 32'h000246D9 , 32'h0006549B , 32'hFFFB9C37 , 32'hFFFEBEDA , 32'h00040668 , 32'h0000D130 , 32'h00035D4A , 32'h0006DC87 , 32'h000028D4 , 32'hFFFD14E8 , 32'hFFFDF8FA , 32'h00009445 , 32'hFFFF83AC , 32'hFFFED167 , 32'hFFFB8BA6 , 32'hFFFDEB8C , 32'hFFFFC83F , 32'hFFF9128D , 32'h00028564 , 32'h0000A9F2 , 32'hFFFB0A04 , 32'hFFFEBB3C , 32'h000035EF , 32'h00000F63 , 32'h0001AE70 , 32'hFFFF428F , 32'hFFFB2E83 , 32'hFFFFDA32 , 32'h0003E198 , 32'hFFFB0384 , 32'hFFFB4107 , 32'h00053533 , 32'h000531DA , 32'h0004D89D , 32'h0000D4EE , 32'hFFFB2799 , 32'hFFF8E7CA , 32'hFFFDEFEB , 32'h00002D4A , 32'h0006FD93 , 32'h0005AE44 , 32'h000138AD , 32'hFFFFC844 , 32'hFFFF34D2 , 32'h000BD885 , 32'h000015AF , 32'hFFFBF82F , 32'h0006CDEF , 32'h00001C43 , 32'h00022D89 , 32'hFFFD7914 , 32'hFFFEC162 , 32'h0000E693 , 32'h0004778C , 32'hFFF94CD4 , 32'h00026916} , 
{32'hFFFE03D0 , 32'hFFFC9412 , 32'hFFFD9EEF , 32'h00030D89 , 32'hFFFED1CE , 32'h0003570D , 32'hFFF80B34 , 32'h0002C32C , 32'h00018948 , 32'h00002A76 , 32'h0004E7A1 , 32'h0001E326 , 32'hFFFCF9AF , 32'h000422BC , 32'hFFFC9245 , 32'hFFF476C9 , 32'h00050690 , 32'hFFFDC2DA , 32'hFFFC3F59 , 32'h0001D209 , 32'h00043C64 , 32'h0003F1B0 , 32'hFFFB9B7F , 32'h0000F3D5 , 32'h000217FD , 32'h0001BBB6 , 32'hFFFFCCDD , 32'hFFFDAE99 , 32'hFFFA26D4 , 32'hFFFE60AE , 32'h0005A251 , 32'hFFFB11ED , 32'h0001C3D3 , 32'hFFFD587E , 32'hFFFEEE4F , 32'hFFFCF553 , 32'hFFFD7ADE , 32'h000A6F61 , 32'hFFFCB9DA , 32'h0002D2CE , 32'hFFFA8918 , 32'hFFF6ECAA , 32'hFFF7B82C , 32'h00025589 , 32'h0008032D , 32'h00010827 , 32'h00064DCA , 32'hFFFD698B , 32'h000335AB , 32'hFFF8123E , 32'hFFFEB13A , 32'hFFFA69D6 , 32'h0003C2F5 , 32'h00046047 , 32'h000D99C3 , 32'hFFF0EF5B , 32'hFFF38187 , 32'hFFFC9DB4 , 32'hFFF647EC , 32'h0007163C , 32'hFFF6035F , 32'h0008B428 , 32'h00031350 , 32'h0002187C , 32'hFFFE3C16 , 32'h000073B1 , 32'h000237F8 , 32'hFFFB11CB , 32'h0004C582 , 32'h0000519B , 32'h00049D66 , 32'hFFF86B9B , 32'h00098B33 , 32'hFFF7D8B2 , 32'hFFFB176B , 32'hFFFB183C , 32'hFFFD4113 , 32'h00039E4D , 32'hFFFF8CCE , 32'h0002C328 , 32'h0008F0E3 , 32'h00034AB7 , 32'hFFFAEFD0 , 32'hFFFEB30B , 32'h00039D78 , 32'hFFFA88C4 , 32'hFFFE16E9 , 32'h0001B1EA , 32'h000110B1 , 32'hFFF834BC , 32'hFFF26D31 , 32'hFFFEF91C , 32'hFFFCFA69 , 32'h00090F4E , 32'hFFFEE5DF , 32'hFFFC38A7 , 32'hFFFB2A88 , 32'hFFFA66EC , 32'h00005E0E , 32'hFFFD1139} , 
{32'h049A3CF0 , 32'hE7982C80 , 32'h0A5EB4F0 , 32'h0166EF34 , 32'hF45FB8F0 , 32'h0E27ED50 , 32'h1CE10920 , 32'hED689020 , 32'hEF5FE300 , 32'hECAE5440 , 32'h11C16520 , 32'hFDE45FBC , 32'h009F5592 , 32'h0F393F00 , 32'hF67C7F10 , 32'hF9D26C88 , 32'h06446408 , 32'h2AF4C740 , 32'h165C4680 , 32'hF58BB6C0 , 32'h049EE2D8 , 32'hF013C470 , 32'h046E1E70 , 32'hFE83CFA0 , 32'h10AF31E0 , 32'h1B4B2200 , 32'hFC2BFC74 , 32'hF889DCF0 , 32'h026AA7E8 , 32'hFF77C033 , 32'hF7E282F0 , 32'h09B017A0 , 32'hF2322A10 , 32'h07ED1CC0 , 32'h062443A8 , 32'h018F8F60 , 32'h1535F9A0 , 32'hFEB22F8C , 32'h063036C0 , 32'h1674E180 , 32'h05CAD4A0 , 32'h0C188F30 , 32'hF8BCD6B8 , 32'hF449EDC0 , 32'hFCE0A9B8 , 32'h040E21D8 , 32'h0E14A5D0 , 32'hFE61BE64 , 32'h121321A0 , 32'h050329B0 , 32'h0B062710 , 32'h0696C980 , 32'hF13FC680 , 32'hF74B45A0 , 32'h02BAA2E0 , 32'hFBBE9600 , 32'hFF8DB7C5 , 32'hFA317900 , 32'h070B8F78 , 32'hF80453A8 , 32'hF8044F90 , 32'h09C4FC20 , 32'h00374735 , 32'h1267AA40 , 32'h07CF5FD0 , 32'h04F7D458 , 32'hFE1EAC84 , 32'h0B323A20 , 32'hF93A2B60 , 32'h06A0A090 , 32'hFFFD0144 , 32'hFD37F660 , 32'h08AF8D80 , 32'h03881C74 , 32'h048D89E8 , 32'h01569560 , 32'h041AF8C0 , 32'hF2E25110 , 32'h0044C7B6 , 32'h080211A0 , 32'h04945A78 , 32'h022FAD84 , 32'h09100250 , 32'hFF38A9DD , 32'hFEB150B0 , 32'h0602D578 , 32'hFEC49AF0 , 32'hFBC048F8 , 32'h042E4008 , 32'hFEE87874 , 32'h000965E2 , 32'hFFFEA704 , 32'hFFFA7954 , 32'h00040170 , 32'h00016160 , 32'h000200CD , 32'h0000EAB1 , 32'h00027D8D , 32'hFFFE4C6C , 32'h0001755E} , 
{32'hEBA64D00 , 32'hA4661D00 , 32'h154BFE80 , 32'h0C7114F0 , 32'h04641978 , 32'h1E507A40 , 32'h1F5D9DE0 , 32'h016D3A78 , 32'hE2B320A0 , 32'hEC9B7300 , 32'hEF88EB00 , 32'h2BE37380 , 32'h15F0CB00 , 32'h0A974330 , 32'h0A126F00 , 32'hFF50B397 , 32'hED7F0300 , 32'h10B3A0A0 , 32'hE4B4FF60 , 32'hEF8AE880 , 32'hF5C40C90 , 32'hE82B7A60 , 32'h15159680 , 32'hFDE77CAC , 32'hEEBD7140 , 32'hF6919790 , 32'h0A07EC10 , 32'h14878AA0 , 32'h0648CAA0 , 32'h0BBB58A0 , 32'h0E7C4000 , 32'hF4A1B200 , 32'h1A803560 , 32'h13CEEBC0 , 32'hE82CD5C0 , 32'h00957ED9 , 32'hFB498F08 , 32'h00E82D63 , 32'hFD470F74 , 32'hFD72CB14 , 32'h17B4BBC0 , 32'hF9624D30 , 32'hF3A82E50 , 32'hEA559A20 , 32'hEBF4FCC0 , 32'h0942B8C0 , 32'h0B1FE450 , 32'hF819D1F0 , 32'h0E548D70 , 32'hF60BAB10 , 32'hF8A419B0 , 32'hF8744670 , 32'h0166DF48 , 32'hF8248990 , 32'h0D807BE0 , 32'hFB953F90 , 32'h0D3BC450 , 32'hF08AF070 , 32'h0F4C2B20 , 32'hFCC58404 , 32'hFCEC5454 , 32'hFFAD9225 , 32'h01676278 , 32'h0C7870C0 , 32'hF614A940 , 32'hEFD76DC0 , 32'hF169EE00 , 32'hF3845160 , 32'hFD1BB430 , 32'h09D90910 , 32'h0841D2B0 , 32'hFE91AB94 , 32'hFEA473CC , 32'h0518C650 , 32'hF46AEB00 , 32'h0525A780 , 32'hFCEDB7D8 , 32'hFF8D4604 , 32'hF9B840E8 , 32'h04F40E58 , 32'h03BA1EA0 , 32'h018D6264 , 32'hFB6863A0 , 32'h05AF9B88 , 32'hFD1B8084 , 32'h026D9C60 , 32'h01C0E44C , 32'h083ABEF0 , 32'h045BBC78 , 32'h00B9752B , 32'hFFFDD9FB , 32'h000A44A5 , 32'hFFFF3437 , 32'hFFFEFCB5 , 32'hFFF892C0 , 32'h00016EB8 , 32'hFFFFC399 , 32'h00031967 , 32'h00021969 , 32'hFFFE3907} , 
{32'h0FFE9A20 , 32'hF4AFD630 , 32'h0F562750 , 32'hFBAEAE90 , 32'h00CD77D7 , 32'h09130BB0 , 32'hF7A70560 , 32'h028F5EFC , 32'h04440F48 , 32'h07F322B8 , 32'h08E704C0 , 32'hFCD5FAC4 , 32'hF90E15A8 , 32'hFF4B9F94 , 32'h09C0B8B0 , 32'hFEC025EC , 32'h0BB1D470 , 32'h0E9B9040 , 32'h0A936F90 , 32'hFE029A54 , 32'hF948D3C8 , 32'hFF0500BD , 32'h0C140C90 , 32'hF860B690 , 32'hF9F33A90 , 32'hF540DC60 , 32'hFF4874F3 , 32'h06C808A8 , 32'h048E2460 , 32'hFFC4CB8E , 32'hFA3D3D00 , 32'h01A9B464 , 32'hF3E8BD40 , 32'h0838EFE0 , 32'h033A10FC , 32'hFD3F2B28 , 32'h04609A50 , 32'hFF4211A1 , 32'hF8D30930 , 32'hFD775FB8 , 32'h00FB9544 , 32'hFE2353C4 , 32'hFA4E1D88 , 32'h032A28EC , 32'hF39CA420 , 32'h0AD01CC0 , 32'hFF0287F9 , 32'hFC432CE0 , 32'h0D6801A0 , 32'hFFCF187F , 32'hFFE711DC , 32'h0B0AAE40 , 32'hFE580414 , 32'h0861F1F0 , 32'h0178E084 , 32'h0B65B2C0 , 32'hF829CCC0 , 32'hF94489A0 , 32'h086428A0 , 32'h022E7A88 , 32'hFD96046C , 32'hFA31EC00 , 32'h047D8B10 , 32'hFAB855D0 , 32'h03ED3410 , 32'h096FD510 , 32'h03A2B780 , 32'h041E74C8 , 32'hFDE247D4 , 32'hFFA9AD34 , 32'h0355BCDC , 32'hFD226B84 , 32'h0579CE68 , 32'hFB2842E0 , 32'h0704C650 , 32'hFA8765C0 , 32'h002C507C , 32'hFC713100 , 32'hFA175768 , 32'h025DFDF8 , 32'h02392B54 , 32'h03A3CDD8 , 32'hFEE93978 , 32'hFC3A5CF4 , 32'h045D7A88 , 32'hFEFF2EEC , 32'hFCC4EAF0 , 32'h067FA448 , 32'h04AB5410 , 32'h00532B78 , 32'hFFF9132C , 32'hFFFE01AD , 32'hFFFF7791 , 32'h0003E820 , 32'h000670B4 , 32'hFFFE8C08 , 32'hFFFD5D4A , 32'hFFFC00ED , 32'h0003870F , 32'h00003E7D} , 
{32'h08BE6470 , 32'h0E6A1A60 , 32'hF1C30770 , 32'h06D0EAC8 , 32'h025992C8 , 32'h0D630860 , 32'hF7DE4D30 , 32'hFBC48448 , 32'h03E1CB80 , 32'h05079E88 , 32'hF7972F80 , 32'hFA961368 , 32'hF8E138D0 , 32'hEE1B4F20 , 32'hFF8D8337 , 32'h04E74738 , 32'h0CED2C40 , 32'h0268D994 , 32'h04F36258 , 32'h0DFEAEE0 , 32'h10D79720 , 32'hF6C7F500 , 32'hF8843218 , 32'hF498E740 , 32'h0D9761B0 , 32'h04BB5700 , 32'h0020FD59 , 32'hFC8A76EC , 32'hF6537A90 , 32'hF59051A0 , 32'hFE169CCC , 32'hFFB2AB66 , 32'hFB61D648 , 32'hF6749980 , 32'h00B95816 , 32'hFFD2527E , 32'hFDF7C52C , 32'hFD223AF0 , 32'hFDC7D7C8 , 32'h01C8BA34 , 32'hF7DFFF30 , 32'hFA5A6CF8 , 32'h046F0F58 , 32'hFF187A78 , 32'hFDA3F3DC , 32'h06E92950 , 32'h09E49E50 , 32'h020302E8 , 32'h0157D7C8 , 32'h00D8F2F6 , 32'h0B720EE0 , 32'hFD2558D0 , 32'hFE94E7E8 , 32'h01004EA8 , 32'h01014E44 , 32'h01DAAC54 , 32'hF56672E0 , 32'h078480C8 , 32'h0083AA54 , 32'h06809080 , 32'hFFB30A5A , 32'hFB2D3748 , 32'h07C15838 , 32'h067EBAD0 , 32'hF6387C20 , 32'hFA4C73F8 , 32'hFD283EB8 , 32'h0E23B520 , 32'hF7868520 , 32'h0AAC54B0 , 32'h056643E8 , 32'hFE158458 , 32'h012EB76C , 32'hFD85DDDC , 32'hF813E350 , 32'hFE888D00 , 32'hFAD98180 , 32'hFF6EF26D , 32'hFE6B3908 , 32'hF054AAA0 , 32'h03C099B0 , 32'h049170C0 , 32'h09BB6370 , 32'h02E68E0C , 32'hFE3EB80C , 32'h05CDF8A8 , 32'hFF3F1811 , 32'h032438C8 , 32'hFD43A1DC , 32'hFFC74CCD , 32'hFFFF7DDC , 32'h00073940 , 32'hFFFF2DE8 , 32'hFFFC7DFD , 32'hFFF970DA , 32'h00056BD4 , 32'hFFF9B801 , 32'hFFFCBA62 , 32'hFFFB6240 , 32'h0006819A} , 
{32'hFFFF0943 , 32'hFFFB6F0B , 32'hFFFD3B9B , 32'h0000C870 , 32'h00040C82 , 32'h00060B47 , 32'h00062848 , 32'hFFFD0318 , 32'hFFFE95EC , 32'hFFFB5729 , 32'hFFFF2081 , 32'hFFFF8F7E , 32'h0001D375 , 32'h00023A02 , 32'h0005FF8E , 32'h00016062 , 32'hFFFDEE00 , 32'h0002A135 , 32'hFFFF2A0E , 32'hFFFD7014 , 32'h000063EA , 32'hFFF88A07 , 32'h00070D9B , 32'hFFFA6269 , 32'hFFF8D5EE , 32'hFFFCE773 , 32'h0000BF3D , 32'h0004F91A , 32'h0001D38E , 32'h0003FC8E , 32'hFFF2886F , 32'h0005E173 , 32'h00065125 , 32'h00028231 , 32'hFFFF0988 , 32'h0005221E , 32'hFFFFBDDB , 32'hFFFF2126 , 32'hFFFEE997 , 32'hFFFF5464 , 32'h00027A10 , 32'h0000668D , 32'hFFFCB7C6 , 32'h00080F16 , 32'hFFFC3A9A , 32'h00018ECF , 32'hFFFE5E2C , 32'hFFF81C0D , 32'h000251F2 , 32'hFFFAE6DE , 32'hFFFC1153 , 32'h0004F4D5 , 32'h000122C6 , 32'hFFFFA3C0 , 32'h0004BCD2 , 32'hFFFE342B , 32'hFFFE38D7 , 32'hFFF87193 , 32'hFFFCC219 , 32'h0002EDA5 , 32'h0000E71D , 32'hFFFB3E19 , 32'h0005D108 , 32'hFFFE3101 , 32'hFFFC7CD1 , 32'hFFFE6260 , 32'hFFFC5E92 , 32'hFFFEC74D , 32'h0005803E , 32'h00007824 , 32'h000104D7 , 32'hFFF7626F , 32'hFFFE8A2E , 32'hFFFFF1E3 , 32'h0006DA3A , 32'hFFFB0E26 , 32'hFFFD36B0 , 32'hFFFD005E , 32'hFFFE3980 , 32'hFFFB05CE , 32'hFFF9BA56 , 32'hFFFE3EE1 , 32'hFFFF3666 , 32'h0002B709 , 32'h0004954A , 32'h0000755B , 32'hFFF8F5CF , 32'hFFF5D5F1 , 32'h00052896 , 32'h0006409D , 32'h00026544 , 32'hFFF93378 , 32'h00035463 , 32'h00014CCA , 32'hFFFAB80B , 32'hFFF9A431 , 32'hFFF78A0D , 32'hFFFCFF50 , 32'h0002D457 , 32'hFFFDD1D7} , 
{32'h0001A716 , 32'h0005BE62 , 32'hFFFB8C6B , 32'h0007E4FE , 32'h0003DE28 , 32'h0001B4D0 , 32'h000221B4 , 32'h000823EB , 32'hFFFAC442 , 32'h00008F8C , 32'hFFF9B66A , 32'hFFFCC37B , 32'hFFFB1024 , 32'h00039874 , 32'hFFF66F20 , 32'hFFFDD750 , 32'h0003B0B1 , 32'h00075E00 , 32'hFFF997FB , 32'h0001122C , 32'hFFFED87D , 32'h00044BD8 , 32'h0001A3E2 , 32'hFFFE32E0 , 32'h0000B6B1 , 32'h00026287 , 32'h00026F27 , 32'h00010A86 , 32'hFFF9BA62 , 32'hFFF18BF6 , 32'h0001487C , 32'hFFF4B66F , 32'h00028016 , 32'h00043663 , 32'h000029EB , 32'h0003C26B , 32'h00013438 , 32'hFFFF9F79 , 32'h0002D26A , 32'h0002EBC7 , 32'hFFFC9048 , 32'hFFFF996F , 32'hFFFE0BDD , 32'hFFFBC619 , 32'hFFFA509F , 32'hFFF4F369 , 32'hFFFA114B , 32'h00024B41 , 32'h0008AE3B , 32'h00075188 , 32'h0001FA9E , 32'hFFF9D2A4 , 32'hFFFEEE28 , 32'hFFFB9804 , 32'h000B2C57 , 32'hFFFAC334 , 32'hFFFCF074 , 32'hFFF21F2E , 32'h00043029 , 32'h00010345 , 32'h000474A4 , 32'h0003324F , 32'hFFFECB37 , 32'hFFFF8A51 , 32'h000812FB , 32'h000163E7 , 32'hFFFD2D8C , 32'hFFFEC79F , 32'h00053C4D , 32'hFFFF380D , 32'h000297ED , 32'h0003F1B6 , 32'hFFF96042 , 32'hFFF5522D , 32'hFFF7E1D6 , 32'hFFFA209F , 32'h000232BC , 32'h00028DC7 , 32'h0004446B , 32'hFFFFD8F2 , 32'hFFF881F3 , 32'h0004A1A9 , 32'hFFFC5863 , 32'h00075409 , 32'hFFFD751B , 32'h0001F489 , 32'hFFFE2A40 , 32'hFFFB07B2 , 32'h00041312 , 32'h0003B105 , 32'hFFFEEED0 , 32'h0004135B , 32'hFFFF1614 , 32'h0005D4E0 , 32'hFFFDA64C , 32'hFFF97A0B , 32'hFFFEC3D4 , 32'h0004991D , 32'h00080F28 , 32'hFFFE2408} , 
{32'hEE1BE800 , 32'hF2C4DEB0 , 32'hEE28CDE0 , 32'h105DDF20 , 32'h037317F8 , 32'hFAC6A858 , 32'hEE26B000 , 32'h0A65EFB0 , 32'hE43360E0 , 32'h08E3D4E0 , 32'hF7ED0FF0 , 32'hFB0F7970 , 32'h06FBF5B0 , 32'hF2F58400 , 32'h02383A0C , 32'h0BF7F900 , 32'h0FA43AD0 , 32'h09E3E960 , 32'hE74A8D80 , 32'h08E60260 , 32'h07F20318 , 32'hF8821228 , 32'h06ED5848 , 32'hF40E5F50 , 32'hFDF01220 , 32'h02DEABE8 , 32'hEE6B3F60 , 32'h0BD0B9F0 , 32'hFCBF063C , 32'hF41E7150 , 32'h05757DC8 , 32'hF7DBEC20 , 32'hF097BCE0 , 32'h06EA3038 , 32'h17B88E60 , 32'hFDB73284 , 32'hFACAD4D0 , 32'h0DAD8B20 , 32'hFF1AE424 , 32'h12896380 , 32'hFB67EC60 , 32'hF68DC680 , 32'h006E7051 , 32'hFEC72C4C , 32'h10A8AB20 , 32'h0506E108 , 32'hEFAD0C00 , 32'h09C02E40 , 32'h03943748 , 32'h107E6000 , 32'h03723B6C , 32'h1A12C060 , 32'hF953A3C0 , 32'hFBF20968 , 32'h0B378690 , 32'h17569FC0 , 32'h00E64B91 , 32'h0C9F2D20 , 32'hFFBF553C , 32'hFDDB3E98 , 32'h0204A620 , 32'h01F0F638 , 32'hFD290EC4 , 32'h0EA11330 , 32'hEF6300C0 , 32'h051166C8 , 32'hEC528520 , 32'hFFDF483A , 32'hF9AB6EA0 , 32'hF73328E0 , 32'h0CBAF140 , 32'h0353EB10 , 32'hFE344DCC , 32'hFD911084 , 32'h0087EC9A , 32'h055759F8 , 32'hFF36D1B4 , 32'h05875E30 , 32'hF6BA6860 , 32'h04794400 , 32'hFCF398B0 , 32'h08D3F3D0 , 32'h041EF7A0 , 32'h08127A50 , 32'hF7F2D0C0 , 32'h06820970 , 32'h051B4A40 , 32'hFD28F124 , 32'hFE211C68 , 32'h014595B4 , 32'h0005435C , 32'h0003D6BB , 32'hFFFD092D , 32'hFFFF58ED , 32'hFFFC4E9D , 32'hFFFF8311 , 32'h0000544E , 32'hFFFE7D21 , 32'hFFFB03F3 , 32'h000111EB} , 
{32'h0001C61A , 32'h00039570 , 32'hFFFE892F , 32'h0005E106 , 32'hFFFB9833 , 32'hFFF92644 , 32'hFFFE684C , 32'h00031E44 , 32'hFFFEDDC6 , 32'h0004BA98 , 32'hFFFE461A , 32'hFFFC5A30 , 32'h00026E5A , 32'h0004CCB4 , 32'hFFFB8271 , 32'hFFFE122E , 32'h0005B329 , 32'hFFFBA30A , 32'h0000C0BE , 32'h00019F97 , 32'hFFFE83CF , 32'h00033C21 , 32'h00013167 , 32'h0000C942 , 32'h00026170 , 32'h0004F7EF , 32'h00058E62 , 32'hFFFD5A8E , 32'h000043C4 , 32'hFFFEF823 , 32'h00013B1C , 32'h0006B480 , 32'h000302A7 , 32'hFFFB5BCE , 32'hFFFEB4AC , 32'h00002F2F , 32'hFFFF8B99 , 32'hFFF65E35 , 32'h000255F1 , 32'h0004FE6E , 32'h00003998 , 32'h0004CFD0 , 32'h0003E99F , 32'h000E4D00 , 32'hFFFC9980 , 32'hFFFC354D , 32'hFFFE9C5A , 32'h00052088 , 32'h0000E659 , 32'h0007BA6C , 32'h00009350 , 32'h000829EA , 32'hFFF6FC37 , 32'hFFF98D9C , 32'h0000178C , 32'hFFFBAE5F , 32'h0004D9BD , 32'hFFFCCF3F , 32'h0004D48D , 32'h0002F154 , 32'h00030F57 , 32'h000562FE , 32'h00031B5D , 32'hFFFD1E82 , 32'hFFFF1FF3 , 32'h00040373 , 32'h000100C2 , 32'hFFFCBA53 , 32'h0002D5FD , 32'hFFFB57D3 , 32'h00002F1F , 32'hFFFACF21 , 32'h0000631C , 32'hFFF86C6E , 32'h00045D14 , 32'hFFFDDF26 , 32'h0001EC71 , 32'h00023DF8 , 32'hFFFCA6DD , 32'hFFF8B493 , 32'hFFF7B49A , 32'hFFF9D6F9 , 32'hFFFEBC54 , 32'hFFFE6AB5 , 32'h00027274 , 32'h000182EF , 32'hFFF72308 , 32'hFFF6BC3D , 32'h0002C208 , 32'hFFFEB23E , 32'h0001CD97 , 32'h0003A79A , 32'h00011F6D , 32'hFFFD6495 , 32'h0006A8D1 , 32'h00024812 , 32'hFFF7E588 , 32'h000194CD , 32'h0002A2DE , 32'hFFFE52B6} , 
{32'hFFFAA0D8 , 32'hFFF9F6D4 , 32'hFFFCA6E9 , 32'h0003D884 , 32'h0003391C , 32'hFFF9365E , 32'hFFFFC3AE , 32'h00047670 , 32'h0001CAB1 , 32'h00000F5B , 32'h0003AB72 , 32'h0004C343 , 32'h000029DD , 32'hFFFDF2CF , 32'h000514AA , 32'h00010DEF , 32'hFFF86EE3 , 32'hFFFED0A9 , 32'hFFFE5E5A , 32'h00068453 , 32'h00022EAE , 32'hFFF54A5B , 32'h00025B32 , 32'hFFFF94C7 , 32'h0004050B , 32'h0000A013 , 32'hFFFFCA05 , 32'hFFFC5AC5 , 32'hFFF7EF63 , 32'h00048E8D , 32'hFFFA4E80 , 32'h000AC59A , 32'hFFFFF1A8 , 32'h00004118 , 32'hFFF8832B , 32'h0001F04E , 32'hFFFE776D , 32'h0003A18A , 32'h000335DA , 32'h000635A7 , 32'hFFFE63B6 , 32'h00048101 , 32'h0007003E , 32'h00048F0E , 32'hFFFD3256 , 32'hFFFF6BC5 , 32'hFFFE48B4 , 32'h0002610F , 32'h000316F4 , 32'h00028998 , 32'hFFFB9710 , 32'h000643E5 , 32'hFFF92000 , 32'hFFF985A7 , 32'h000135EB , 32'h0002681D , 32'hFFFB722F , 32'h00068B79 , 32'hFFFBD91E , 32'hFFF96E1E , 32'h00003D79 , 32'hFFF8287C , 32'h0001C1CA , 32'hFFFCD6FA , 32'h00046A64 , 32'h0001CB75 , 32'hFFFF979A , 32'h00064193 , 32'h0009757A , 32'h00043291 , 32'hFFFFD13C , 32'h00028E61 , 32'hFFFF2410 , 32'hFFFB19FA , 32'h00061159 , 32'h000981AC , 32'hFFFC5700 , 32'h00044433 , 32'h00044326 , 32'hFFFBF7EF , 32'h00015415 , 32'h0002D573 , 32'hFFFD79E7 , 32'hFFFD725B , 32'h00061EB1 , 32'h000280D0 , 32'hFFFD7564 , 32'hFFFE8824 , 32'h00017B31 , 32'h000099B0 , 32'hFFF82F1F , 32'h00075095 , 32'hFFFE4D5D , 32'h000A160F , 32'hFFFCBDED , 32'h0001E5B9 , 32'hFFFB98BE , 32'hFFFA0169 , 32'hFFFD818C , 32'h0002CCC8} , 
{32'h080810F0 , 32'hE7A70160 , 32'h0BA2DE80 , 32'hDB40E400 , 32'h182C32C0 , 32'hE7ABBBE0 , 32'hFD7224D8 , 32'hFF8A8476 , 32'h146106C0 , 32'hF977B510 , 32'h03B1146C , 32'hFE6C6648 , 32'hEA95DB40 , 32'h09156050 , 32'hFE99FE54 , 32'hF955CED8 , 32'hEAD0FCE0 , 32'hF83EE1E8 , 32'h0192D088 , 32'hF07D8470 , 32'hF782ECE0 , 32'h08155990 , 32'hF0824090 , 32'h0BB34C00 , 32'h14896280 , 32'hF89100B8 , 32'hF6D6C000 , 32'hF85E5F28 , 32'h0C882320 , 32'h0B56D1C0 , 32'hF11F66B0 , 32'h072B8C68 , 32'h01784A0C , 32'hF8286130 , 32'hECFCF580 , 32'hFE4F0E6C , 32'h0D21BF20 , 32'h0F847940 , 32'h039BEB18 , 32'hFA2E3F70 , 32'h0C142A60 , 32'h0F463DD0 , 32'hFBAA1F50 , 32'hF0F0D2C0 , 32'h0B789B80 , 32'hFC70E888 , 32'h00A045DF , 32'hF6F8EB10 , 32'hF761AA00 , 32'h05D15CB8 , 32'hF77CB300 , 32'hF8A5E710 , 32'hF6180CC0 , 32'h01CA37F0 , 32'h0B187CE0 , 32'hF7B72890 , 32'hF4F108F0 , 32'hFFE8837F , 32'hFA7D98B0 , 32'h05FE8E90 , 32'h0B2D28D0 , 32'h01D5B574 , 32'hFA4DB880 , 32'hF83707C8 , 32'hFECA85D8 , 32'h0BF2BE10 , 32'hFC4F211C , 32'hFC710E98 , 32'h07B622C8 , 32'hF434F380 , 32'h03D37800 , 32'hFEE779D8 , 32'h0DC64350 , 32'hF42BA760 , 32'hEA5D0500 , 32'hF22D1BE0 , 32'hFB2E6750 , 32'hF69E8B90 , 32'h02110A84 , 32'h04F2DBB8 , 32'hFA00C570 , 32'hFEA07FF0 , 32'hFC08E56C , 32'hFBDE79A0 , 32'hF9A6AE38 , 32'hFC3C446C , 32'h0101708C , 32'hFA4EACA8 , 32'h084341B0 , 32'h0062170E , 32'hFFF95801 , 32'hFFFD34DD , 32'h0004362D , 32'hFFFF1F4A , 32'hFFFF0D16 , 32'hFFFD7736 , 32'hFFFDC7E2 , 32'hFFFF25D0 , 32'h00004E73 , 32'h00021946} , 
{32'hFFF9993C , 32'h0005292A , 32'h0002959A , 32'h00075CE6 , 32'h00011102 , 32'hFFFE4A53 , 32'hFFFF7947 , 32'hFFFA7A6B , 32'h00019426 , 32'hFFF62E13 , 32'h0003F148 , 32'h00024DD6 , 32'h00066499 , 32'hFFF7E60F , 32'h0001AF30 , 32'h0001F1F1 , 32'h00014F70 , 32'h0006346F , 32'hFFFE2214 , 32'hFFFFEACE , 32'h00070AC2 , 32'h000A22F3 , 32'h00028765 , 32'hFFFF57DD , 32'h0008F40E , 32'h000320CF , 32'h00003782 , 32'hFFFD6149 , 32'h00007DFC , 32'hFFFE7054 , 32'h00092B72 , 32'hFFFF81AA , 32'hFFFF6B60 , 32'h00006DE3 , 32'hFFFF0A98 , 32'hFFFCC9E1 , 32'hFFFB98E6 , 32'hFFF85A73 , 32'h00079BA3 , 32'h00055F47 , 32'h00040A94 , 32'h00017C25 , 32'h0000C561 , 32'hFFFDE328 , 32'hFFFCAA15 , 32'hFFFCF70A , 32'h00030894 , 32'h0004070B , 32'hFFF94F75 , 32'hFFFCBD34 , 32'h0000116D , 32'hFFF9BE42 , 32'hFFFD9B3E , 32'h00005C05 , 32'h0003ED04 , 32'hFFFEDCC7 , 32'hFFFD57F3 , 32'hFFFAC43B , 32'hFFFC3A1B , 32'hFFFB2454 , 32'hFFFEDBE4 , 32'h0002D7E8 , 32'hFFFC84CC , 32'hFFFE2C91 , 32'hFFFEACB5 , 32'h00027455 , 32'h0002961D , 32'hFFF5110F , 32'hFFFDA28F , 32'h00023328 , 32'h0003D3D4 , 32'h00005096 , 32'h00039325 , 32'h0000BFF3 , 32'h0002DD6B , 32'hFFFB9E0D , 32'h0006ED86 , 32'hFFF7C71D , 32'h000DF1AF , 32'h00024798 , 32'h0002AE82 , 32'h0003CE6A , 32'h000539AF , 32'h0007AD0D , 32'h0000E894 , 32'h00017D63 , 32'h000036A0 , 32'hFFFD86AA , 32'h00027F89 , 32'hFFFA2472 , 32'h0008AF43 , 32'h00053B08 , 32'h0000FEF0 , 32'hFFFF69B4 , 32'h000394C4 , 32'h000208CA , 32'h0004E5A7 , 32'h00053254 , 32'hFFFF419B , 32'hFFF820E4} , 
{32'hFFF8CA72 , 32'h00055EFB , 32'h0000E6C7 , 32'h00062C99 , 32'hFFFF7722 , 32'h00017A24 , 32'hFFFDA511 , 32'hFFFF00F5 , 32'h00013AC5 , 32'hFFFD1B4B , 32'h00018217 , 32'hFFF8F13A , 32'hFFFDFBE1 , 32'h00085FB6 , 32'h0006BC30 , 32'h0000A93B , 32'h00047766 , 32'h0001AC59 , 32'hFFFE5895 , 32'h000604D2 , 32'h0002D2D4 , 32'h00031277 , 32'h00064E61 , 32'hFFF81BFF , 32'hFFF4C4F7 , 32'h0002AC9C , 32'h00014119 , 32'h0000905B , 32'hFFF47A9B , 32'h0003B28E , 32'h00027DEA , 32'hFFFF1827 , 32'hFFFFB6CE , 32'hFFFD1CCF , 32'hFFFDC081 , 32'h00000B35 , 32'h00012819 , 32'hFFFD5C09 , 32'hFFFE1999 , 32'h00008892 , 32'hFFF8B207 , 32'h00048B41 , 32'h0002A6AB , 32'hFFFBEE28 , 32'h000B4CC9 , 32'hFFFCEE25 , 32'hFFFDCF5A , 32'hFFFE7A6C , 32'hFFFDB99A , 32'h00001EEF , 32'hFFFEA398 , 32'h00068FF9 , 32'h00083A22 , 32'hFFF6AFD8 , 32'h00008D42 , 32'h00003DE7 , 32'h0000FE13 , 32'hFFFF0C23 , 32'hFFFBA386 , 32'h00035C29 , 32'hFFFC32AC , 32'hFFFAA314 , 32'h0001A10D , 32'h00040AB0 , 32'hFFF7D5AF , 32'h0002AD89 , 32'h00071069 , 32'hFFFB18BA , 32'hFFFE76A0 , 32'hFFFE4006 , 32'hFFFDA5C4 , 32'hFFF8A4ED , 32'hFFFEEF70 , 32'hFFFD52A9 , 32'h0006945B , 32'h0008E93E , 32'hFFFC11F2 , 32'hFFF8B0CE , 32'hFFF949E2 , 32'hFFFD8291 , 32'hFFF6BF03 , 32'hFFFE7AAE , 32'h00074B2D , 32'h0000E554 , 32'hFFFE87B2 , 32'h0008CCCC , 32'hFFFB3322 , 32'hFFFBE390 , 32'hFFFE504C , 32'hFFFFEC7D , 32'hFFFE282D , 32'hFFF6CF93 , 32'h00078CF4 , 32'hFFFF23DE , 32'hFFF5DAE3 , 32'hFFFF5487 , 32'hFFFFFB3A , 32'h0001F1AD , 32'h00006336 , 32'hFFFD4556} , 
{32'h1AFDEA80 , 32'hF9F75B50 , 32'hEBC80A80 , 32'hA3056080 , 32'h35255600 , 32'hFCA648F0 , 32'hF8E0CF78 , 32'h1A6E35A0 , 32'h025F6844 , 32'hF8713F40 , 32'hFE7B68A0 , 32'h183628C0 , 32'hF258B970 , 32'h0F833D70 , 32'hF1BF5A60 , 32'h319C03C0 , 32'hE78D5200 , 32'h02D89168 , 32'h23D15300 , 32'hF481C0B0 , 32'hF49F52D0 , 32'hED149800 , 32'hFEC128C8 , 32'hF921A528 , 32'hE60DED60 , 32'hEB1304C0 , 32'hF9582C58 , 32'hFE6877FC , 32'h0CB1CF70 , 32'hF81149F0 , 32'h1A61A880 , 32'hF6C19550 , 32'hF2B622F0 , 32'h036C726C , 32'h0314448C , 32'h12683C60 , 32'h13CC6720 , 32'h1DD6E1C0 , 32'h10F9E6C0 , 32'hDEFFD880 , 32'h0E2FE450 , 32'h1DE4DF40 , 32'h0108BBC8 , 32'hEE4FA580 , 32'hF189FAE0 , 32'h1A8DC3E0 , 32'hF87C5888 , 32'h06230C20 , 32'hEE5683E0 , 32'hFF417045 , 32'hF4DDCFA0 , 32'h0168B38C , 32'hF7D912D0 , 32'hF5AD0AA0 , 32'hFE89D268 , 32'hECE07380 , 32'h04932CF0 , 32'h0C39F690 , 32'hF1F7DF00 , 32'h0627DEB8 , 32'h0DA7D640 , 32'h00362BF3 , 32'h05230018 , 32'hFF329CBD , 32'hF51333C0 , 32'h03BCA9A4 , 32'h065509B8 , 32'h0C178AE0 , 32'h0BCBED70 , 32'h06D6A7E8 , 32'h1365EE60 , 32'h073D74F8 , 32'hFEAFEAC8 , 32'hFA52CCB8 , 32'h0838E8D0 , 32'h097C37D0 , 32'h024D5A70 , 32'h03D45150 , 32'hFB3B1730 , 32'h04006600 , 32'h00EB6087 , 32'hFDDF7568 , 32'hFD7AC8D8 , 32'hFD3B5A9C , 32'h039020BC , 32'hFC5D02F8 , 32'hFFC13C5C , 32'hFE72A064 , 32'hFA35F718 , 32'h01630850 , 32'h00035F91 , 32'hFFFD1F94 , 32'hFFFDDED0 , 32'hFFFF0BB0 , 32'h0003B4DA , 32'h0003CA07 , 32'h0001C0E4 , 32'h00026679 , 32'h0001DA3E , 32'h0002C9E8} , 
{32'h00015F25 , 32'hFFF9A6BF , 32'hFFFBD49B , 32'hFFFFF62C , 32'hFFF63773 , 32'h0001BE09 , 32'h00077BAD , 32'h0005CA59 , 32'hFFFF0C98 , 32'h00048E03 , 32'hFFFFFBAA , 32'hFFFB77FC , 32'h0007B1AF , 32'h000079DC , 32'hFFFD8DF6 , 32'h0002B742 , 32'hFFFFEE0F , 32'h00048901 , 32'hFFF3098F , 32'h00009470 , 32'h0001B912 , 32'h00016A1B , 32'hFFF3B4B8 , 32'hFFFFEBA8 , 32'h0004A5D7 , 32'hFFF69647 , 32'h00037C48 , 32'hFFF8D55D , 32'hFFFF07F9 , 32'h0004F10D , 32'hFFFDADB1 , 32'hFFFDB22D , 32'hFFFAE0AF , 32'hFFFC666F , 32'h000DE1D2 , 32'h0006C939 , 32'h000134D5 , 32'h000059FE , 32'hFFFDD713 , 32'hFFF91C8C , 32'hFFF76AD4 , 32'hFFFFA20B , 32'hFFFFAF6F , 32'hFFF594F1 , 32'hFFFE009D , 32'hFFFD9A8F , 32'hFFF4B0B4 , 32'h0004D727 , 32'hFFFFFF4F , 32'h0007A386 , 32'hFFFC63DF , 32'h000504DA , 32'h0003683D , 32'hFFF92133 , 32'h0008A632 , 32'h000218FF , 32'h0004393F , 32'h00012485 , 32'h0007DD6F , 32'hFFF8860D , 32'hFFFA5174 , 32'h0001F094 , 32'h0008053B , 32'hFFF8D628 , 32'hFFF9D0C0 , 32'hFFFB715E , 32'hFFF965AE , 32'hFFFB8BEE , 32'hFFF5015C , 32'h0003ECAD , 32'h00064DAD , 32'hFFFB9DFB , 32'h00049FA4 , 32'h00008029 , 32'hFFF99B8C , 32'hFFF93B3F , 32'hFFFD9F0A , 32'h000372BD , 32'h00010B42 , 32'hFFFFA53B , 32'h000AF738 , 32'h00000170 , 32'hFFFF30F3 , 32'hFFFA04AF , 32'hFFFE4ACD , 32'h00031D33 , 32'h000123EB , 32'h0008E95C , 32'h000788DF , 32'h00069D25 , 32'h0001E895 , 32'hFFFC8E2C , 32'h0000D2C8 , 32'hFFFECC1B , 32'h0006476A , 32'hFFFBB12F , 32'h000030BD , 32'hFFFE267A , 32'hFFFEC5FD , 32'h0006EE21} , 
{32'h3CA7C180 , 32'h135FEBC0 , 32'hFCF88580 , 32'hEDC2BFE0 , 32'h00040A2F , 32'hC6AE7940 , 32'hEE775340 , 32'h0E780CD0 , 32'h2BD5D7C0 , 32'hF0757BE0 , 32'hF495D650 , 32'h0ACE8A80 , 32'h037CC5A8 , 32'hD7565180 , 32'hE3EBF980 , 32'h08476860 , 32'hEA0A4800 , 32'h377F4540 , 32'h0795BE88 , 32'h2839E980 , 32'h1E4F8D40 , 32'hE5694700 , 32'h17543400 , 32'hFFA6A31B , 32'h123277C0 , 32'h0B283CF0 , 32'h05A64AC8 , 32'h11811640 , 32'hE65AAFC0 , 32'hF88E5328 , 32'hFF637D09 , 32'hF9C13A18 , 32'h1A32CDC0 , 32'h06F5D4A0 , 32'h009DDAD0 , 32'h0568D4F8 , 32'h08B4A530 , 32'hFD44E4EC , 32'h07C6ABD0 , 32'hFF15DC7E , 32'h13516300 , 32'h00CE33C7 , 32'hFD1BCEA4 , 32'h036ED4FC , 32'h02FC4854 , 32'h04A27680 , 32'h03D59228 , 32'h2D182500 , 32'h014FB074 , 32'hFD6BA98C , 32'h08802100 , 32'h0217D740 , 32'hF56C20F0 , 32'h12E81E40 , 32'h05D6EC80 , 32'hFC95568C , 32'h08797A30 , 32'h083290E0 , 32'h19225CE0 , 32'h005C279C , 32'hF72E5A90 , 32'h06022070 , 32'hE9473A40 , 32'h047CEC70 , 32'hF9353588 , 32'h0129097C , 32'hFA4893D8 , 32'hFF421196 , 32'h08B80510 , 32'h0C21CE00 , 32'hFCE39DF0 , 32'h10477E60 , 32'hFD486F28 , 32'hFAF05C60 , 32'h00BE4D74 , 32'hF7BD39D0 , 32'hFE5628A0 , 32'h08FC94E0 , 32'h055BFE38 , 32'hF7AFFE80 , 32'hFDBE0D8C , 32'hFD47C618 , 32'hFC015004 , 32'hFBA41728 , 32'hFEA31194 , 32'h045C6C80 , 32'hFA9A3D78 , 32'hFDED4FC0 , 32'hFD2E4A78 , 32'hFF130B41 , 32'h0001D511 , 32'h00058321 , 32'h00010C56 , 32'h0003DD68 , 32'hFFFBA1C8 , 32'h0003FA3E , 32'hFFFDC54D , 32'h000178D9 , 32'hFFFFD912 , 32'hFFFFAFDE} , 
{32'h05AE8910 , 32'h04A64510 , 32'hFEA8ABC0 , 32'h00EE3162 , 32'h09544640 , 32'h0B02AF20 , 32'h044141A0 , 32'hF3B9A040 , 32'h077D3228 , 32'h03B3B6AC , 32'h04A32AE8 , 32'hFBCD6028 , 32'h04A260D8 , 32'h06520418 , 32'h00E50591 , 32'h01B875D8 , 32'h00F7C565 , 32'h0093C61E , 32'hF0E349C0 , 32'h00278638 , 32'h06C418A8 , 32'hEF506E20 , 32'hFE5E417C , 32'hFD70462C , 32'hFE9248FC , 32'h00C9EEDA , 32'hFAB9A910 , 32'h00856B33 , 32'hF67FE420 , 32'h00CCC852 , 32'h03BB8BF4 , 32'h03058D18 , 32'h093C1890 , 32'h00C36702 , 32'hF3C07170 , 32'hF57F1C90 , 32'h012734B0 , 32'hF63F8010 , 32'hFD5734CC , 32'h00D771C9 , 32'h045A9FD0 , 32'hFFC0B7E5 , 32'h02A821E8 , 32'hFBBBB3C0 , 32'hFBEE47D8 , 32'h0BB92250 , 32'hFF9E56FD , 32'h06A20D40 , 32'hFEDA5BE4 , 32'hFE6A9F50 , 32'hFEF6F568 , 32'h02DE7168 , 32'hF6D7BE20 , 32'h005CEEA8 , 32'h05688070 , 32'h024BC9DC , 32'h0318E32C , 32'h08AB0970 , 32'hF8264B38 , 32'h03CC0444 , 32'h04D0E0A0 , 32'hFE75A354 , 32'h02C6719C , 32'hFB7A9718 , 32'hFE1E9428 , 32'h02526F8C , 32'hF7853D80 , 32'h01369E14 , 32'h036D13BC , 32'hFF2F16B1 , 32'h0127D03C , 32'hF743EC70 , 32'h017777C4 , 32'hFEB81640 , 32'hFF823517 , 32'hFBD60100 , 32'hFE07FDB8 , 32'h011CD44C , 32'h07376FA8 , 32'hFD0267F4 , 32'h04AB3F70 , 32'h048FA130 , 32'hFF026DAB , 32'hFD2BFF30 , 32'h0029BCC2 , 32'h007E90C5 , 32'hFB909C28 , 32'h033F7010 , 32'h0065B12F , 32'hFF3A16FA , 32'hFFFCA311 , 32'h00020AA8 , 32'hFFFEA322 , 32'hFFFE67FB , 32'hFFFAED1A , 32'hFFFDCBA0 , 32'h0005431C , 32'hFFFD5F7C , 32'h000045A8 , 32'hFFFD137E} , 
{32'hFFF8C60A , 32'hFFFAF382 , 32'hFFFBDC21 , 32'h00070A09 , 32'hFFFC7D57 , 32'h00032A9D , 32'h000079ED , 32'hFFFD7FF7 , 32'h000AF98C , 32'h00016FE5 , 32'hFFFC0465 , 32'h000028BA , 32'h0002B8E6 , 32'hFFFCFF1B , 32'hFFF9B20D , 32'h000030C1 , 32'h000592C6 , 32'h000323BA , 32'h0005E86B , 32'h0000F7D8 , 32'hFFFE3625 , 32'h00012C87 , 32'h00021B04 , 32'h00031322 , 32'hFFF91C1D , 32'hFFFC6AE8 , 32'hFFFE1297 , 32'h0000DA0F , 32'h0000F442 , 32'hFFFD55DA , 32'hFFFE3E04 , 32'h0009935D , 32'h00062E4B , 32'h0000ACDE , 32'h00087CBF , 32'h00004A9C , 32'hFFFD3A33 , 32'h00031E42 , 32'hFFFB1B1D , 32'hFFF9692D , 32'h0002614D , 32'h000523B9 , 32'hFFFD7C49 , 32'hFFFE7987 , 32'h000021DC , 32'h00038443 , 32'h0006515F , 32'h00024213 , 32'hFFFFD2CC , 32'hFFF9EA39 , 32'h00023291 , 32'h0005EF0A , 32'h0005BFFA , 32'h0002FCBA , 32'h0001F112 , 32'hFFFD6944 , 32'h000451CB , 32'hFFFF39F8 , 32'h0002A129 , 32'h00010E3B , 32'hFFFCD846 , 32'hFFFCC83B , 32'h00025F8A , 32'h00036DE3 , 32'h0003C93D , 32'h0002C824 , 32'hFFFD029C , 32'h0000C16A , 32'h000344BB , 32'h000415E3 , 32'hFFFCD290 , 32'h000216A9 , 32'hFFF6C25C , 32'h0000AB60 , 32'h0001C105 , 32'hFFF5D483 , 32'hFFFAAD2C , 32'h00041CD2 , 32'hFFFDEA4B , 32'h0000A22D , 32'h0004B9B8 , 32'hFFFD471E , 32'hFFFD471C , 32'hFFFD6240 , 32'hFFFC3645 , 32'h0003F75F , 32'h00040A75 , 32'hFFFC2DAA , 32'hFFFCB0DD , 32'h0003C5C9 , 32'h00073C9C , 32'hFFFCC642 , 32'h0000CE8F , 32'h0000627F , 32'hFFFD97C3 , 32'h0006A8AC , 32'hFFF8593A , 32'hFFF8A6D6 , 32'h0003570D , 32'hFFFE9B78} , 
{32'h00031A99 , 32'hFFFC1B48 , 32'hFFFB1330 , 32'h00005F26 , 32'h000551F7 , 32'hFFFD376A , 32'hFFFD24EA , 32'hFFFCF943 , 32'hFFFCA5E1 , 32'hFFF77CA9 , 32'h00001BD5 , 32'h000438DC , 32'hFFFC8495 , 32'h0000EFA4 , 32'h0004CE50 , 32'hFFFF1ADF , 32'h0004C723 , 32'hFFFC36A7 , 32'hFFF926EC , 32'hFFFFBEA1 , 32'h00058210 , 32'hFFFFAE13 , 32'h000491FC , 32'h00029894 , 32'h00064A4B , 32'h0003362B , 32'h0005A7EA , 32'h0002A2E5 , 32'h000147BF , 32'hFFFBD139 , 32'h00004DCE , 32'hFFFE426F , 32'hFFF7EE67 , 32'h0006FB49 , 32'hFFFA4A67 , 32'h000353A0 , 32'hFFFA0CF6 , 32'hFFFF8B2F , 32'hFFFCECEA , 32'h00003AC9 , 32'hFFF87539 , 32'hFFFCB66A , 32'h0003E46A , 32'hFFFE969F , 32'h00015925 , 32'hFFFCE570 , 32'hFFFE2680 , 32'hFFFAD6B7 , 32'h000100A0 , 32'h0004D57E , 32'h00000107 , 32'hFFFEFFA5 , 32'hFFFE9019 , 32'h00013A0D , 32'h00017DBF , 32'h00073D84 , 32'h000476B0 , 32'hFFF847A1 , 32'h0000E8B1 , 32'h0002DFDA , 32'hFFFF1EE5 , 32'h000928F0 , 32'hFFFC1E41 , 32'hFFFCCE2F , 32'h00014497 , 32'h000987DA , 32'hFFFC7D3B , 32'hFFFF3849 , 32'h00020452 , 32'hFFFC9E08 , 32'hFFF69A4F , 32'h0000D4F2 , 32'hFFFE9C29 , 32'hFFFD29AB , 32'hFFF23697 , 32'hFFFC79B4 , 32'h00023FC0 , 32'h00000263 , 32'hFFF993E5 , 32'h0000D919 , 32'h0003125F , 32'hFFFC54B5 , 32'h00070985 , 32'h0002AA1F , 32'h00004410 , 32'hFFF8838A , 32'hFFFF6EA4 , 32'hFFFF0372 , 32'h0005AAF7 , 32'h000135E0 , 32'h0006BCD7 , 32'h000228DA , 32'h00037152 , 32'h000413D5 , 32'h000189B9 , 32'h0001586C , 32'h00072BA3 , 32'hFFFCE983 , 32'h0004DAB2 , 32'hFFFE3B36} , 
{32'hFFFBF37D , 32'hFFF8E9D4 , 32'hFFFE0B39 , 32'h0003A208 , 32'h0009693B , 32'hFFFF3E3D , 32'hFFFF48DD , 32'hFFFB55B3 , 32'hFFFDC230 , 32'hFFFF182E , 32'h000908B2 , 32'hFFFDC49E , 32'hFFFB5ECE , 32'hFFFC7EF5 , 32'h0002B11E , 32'h0000BDEF , 32'h0004F798 , 32'h0002EC1A , 32'hFFFD2FA4 , 32'h00053C98 , 32'h000243AC , 32'hFFFE4C90 , 32'hFFFF4AAE , 32'hFFFBFABE , 32'h00063177 , 32'h000140E0 , 32'hFFFBC9B9 , 32'hFFFFF07E , 32'hFFF5F4BE , 32'h0004C54B , 32'hFFFC398E , 32'h000118B5 , 32'hFFFF70C6 , 32'hFFFFBE7C , 32'h0001B4A7 , 32'h0001C26A , 32'hFFFE1586 , 32'hFFFED11E , 32'hFFF6292E , 32'hFFFF2196 , 32'h00041CA5 , 32'h00012827 , 32'hFFFF139A , 32'hFFFEBF1A , 32'h0000B2A2 , 32'h000412A6 , 32'h0001C830 , 32'hFFFC8DA6 , 32'h000267A1 , 32'hFFFDDEE5 , 32'hFFFF6477 , 32'h000243A1 , 32'h0005444C , 32'h0001A05C , 32'hFFFDA49F , 32'hFFFF24D1 , 32'h0003FD0D , 32'hFFFE4CBE , 32'hFFFCD383 , 32'hFFFD416C , 32'hFFFDE809 , 32'hFFFD7495 , 32'hFFF9AD60 , 32'h000505CD , 32'h000E218A , 32'h000735E3 , 32'hFFFC811C , 32'h0003C08C , 32'h0007C131 , 32'h0006863F , 32'h0004BF9A , 32'h0005E1AE , 32'hFFF698AF , 32'h0007441C , 32'h000198A1 , 32'h0000987C , 32'h0001D6EC , 32'hFFFF82B0 , 32'h00006689 , 32'h00017C41 , 32'h00010F89 , 32'h00013C7B , 32'hFFFF9994 , 32'hFFFC37FE , 32'hFFFF952C , 32'hFFFF4606 , 32'hFFFD7FA9 , 32'hFFFF5F7A , 32'h0001DABA , 32'hFFF5DF73 , 32'h000C80D1 , 32'h0000CEF1 , 32'h0007C3C9 , 32'hFFFBE863 , 32'h0001F37D , 32'h0008500C , 32'hFFFFC72A , 32'hFFFB2D32 , 32'hFFFBE7A7 , 32'h0002BE78} , 
{32'h56674000 , 32'h16F288A0 , 32'h2BCD8300 , 32'hBE0C0A00 , 32'h325398C0 , 32'hE6671820 , 32'hE0DAF5E0 , 32'hD2935E00 , 32'h06C02D08 , 32'hF401FE30 , 32'h14D08C00 , 32'h3AF36F00 , 32'hF80F1B48 , 32'h037704AC , 32'h0879D620 , 32'h12390940 , 32'hDE30C140 , 32'h1288C300 , 32'h09827540 , 32'hFA5B9C70 , 32'hFE17F540 , 32'hFD19C4FC , 32'h2A52CF40 , 32'hFE178688 , 32'h13520BC0 , 32'h071BFFD8 , 32'hF9528180 , 32'hFEA2FFE4 , 32'h003FFA40 , 32'hDE5BD5C0 , 32'hFA575270 , 32'h01858EC8 , 32'hFD22E478 , 32'h0B048E60 , 32'h12A66700 , 32'h0658E5C8 , 32'h2D3CBF00 , 32'h0D470BE0 , 32'h0C776B50 , 32'h0AE989F0 , 32'hE9C286C0 , 32'hEC4D2D40 , 32'h023970FC , 32'hE8A91CA0 , 32'hEAFC4540 , 32'hF424FA30 , 32'h09F0CFF0 , 32'hF55ECCB0 , 32'hFDCD04B8 , 32'hFDA3FD50 , 32'hFD819EEC , 32'hF93F4018 , 32'hFF81D9CB , 32'hF9306050 , 32'h008E2DBA , 32'h099FDC50 , 32'hF2892F10 , 32'h05774938 , 32'h102CFB80 , 32'h0D5DE080 , 32'h103C5EE0 , 32'h06A6EAA8 , 32'h14750E00 , 32'h002C2041 , 32'hFBB70E28 , 32'hFC4725BC , 32'h1A65BE40 , 32'hFCD366D0 , 32'hF0E7EF60 , 32'hFFCBEF3E , 32'h02657324 , 32'hFD3CE5B4 , 32'h01F74078 , 32'hFBEE9BB8 , 32'hFFD3A2C0 , 32'h09045CD0 , 32'h058E3458 , 32'hFDD5D2A4 , 32'h018AFBDC , 32'hFDF720C0 , 32'hFC9D76A8 , 32'hFC3DF058 , 32'h04E3E8B0 , 32'h027873CC , 32'h0751A000 , 32'hFF1E6645 , 32'h013C033C , 32'h01349E74 , 32'h03B0B854 , 32'h018D74CC , 32'h000507C9 , 32'hFFFDA7E8 , 32'hFFFEB10B , 32'hFFFF4466 , 32'hFFFC539F , 32'hFFFDDF13 , 32'hFFF9777A , 32'h00021B63 , 32'hFFFCA84F , 32'hFFFF23A7} , 
{32'hD70AE940 , 32'h111140C0 , 32'hE32102A0 , 32'h0D5E7570 , 32'hDB5FDB80 , 32'h2B602640 , 32'hFF44A894 , 32'hFA1FF840 , 32'h1DA8D2A0 , 32'hE2C786E0 , 32'hD45D7080 , 32'h0E425B90 , 32'hD58B2500 , 32'hE58140E0 , 32'hF1EF4130 , 32'hD9ABFD40 , 32'hF7C21040 , 32'h056C6470 , 32'hE630BDC0 , 32'hFDD98C90 , 32'h00F7A94C , 32'hF28C1B90 , 32'h0AB5CCE0 , 32'hF309F5B0 , 32'hEBD21C80 , 32'hF5F1C160 , 32'hECC8C9E0 , 32'hF552CE90 , 32'h00A14ABE , 32'h1FCDABE0 , 32'hEB769BC0 , 32'hFF9045CE , 32'hF2BAF180 , 32'hF43D7FA0 , 32'h004B90BB , 32'h049903E0 , 32'h1D913E80 , 32'h04780D18 , 32'h150F6800 , 32'hFCF83A40 , 32'hFBBF16C8 , 32'hFEABB4A4 , 32'hEF5AF3C0 , 32'hED322340 , 32'h0B2B6150 , 32'hFCEE2E74 , 32'h0CE52D80 , 32'h103DB9E0 , 32'hE6A40140 , 32'h00A17D24 , 32'h06AE01D8 , 32'h0BA1FEF0 , 32'hF8AA5690 , 32'h06F3E428 , 32'hF4C43C20 , 32'hF0727ED0 , 32'h06649950 , 32'h037ED860 , 32'h06902740 , 32'h0556EAB0 , 32'h03394D48 , 32'h0206641C , 32'hFAB82478 , 32'h07002238 , 32'hF580D710 , 32'hFAC63AE0 , 32'hF866C200 , 32'h0BF0D350 , 32'h0D2353D0 , 32'hFCB84C30 , 32'h03374EF4 , 32'hFFC50F80 , 32'hFE957B44 , 32'hF36FD710 , 32'h0CE2D050 , 32'h06AC9308 , 32'hFAC4F9D0 , 32'hFE4B590C , 32'h052923F0 , 32'hFDCE9E3C , 32'hFCB61154 , 32'hF9A11D88 , 32'h00B0B779 , 32'h025B8BFC , 32'hFFA1616D , 32'h00F78C06 , 32'hFEAC937C , 32'h0203BC08 , 32'hFB29ADF0 , 32'hFFFCC8DE , 32'hFFF8B57A , 32'h00019198 , 32'h00028FF6 , 32'hFFFF1745 , 32'hFFFEC638 , 32'h00035F3A , 32'hFFFD3CF2 , 32'hFFFFC37F , 32'hFFFF960F , 32'hFFF95B5C} , 
{32'hE83807A0 , 32'h028B107C , 32'h11DCECA0 , 32'hE13C22E0 , 32'hE70FA640 , 32'hFD21A38C , 32'hFDE59860 , 32'hF57FF930 , 32'h15C45640 , 32'hE9874B00 , 32'hF4F0B220 , 32'h2113F600 , 32'hEE088D80 , 32'hE8B86C20 , 32'hE3B76D40 , 32'h2854C280 , 32'h125E1D60 , 32'h011B7FEC , 32'hDF569A00 , 32'hEEF17240 , 32'h11915160 , 32'h0EA85090 , 32'h0B8FFC40 , 32'hF10A38A0 , 32'h15EA3B00 , 32'h0209DAC4 , 32'hD2E4B9C0 , 32'h0998A700 , 32'hF5092CC0 , 32'hEA85EDC0 , 32'hF6CF3660 , 32'hF0725110 , 32'h0D9EF130 , 32'hFB4E7090 , 32'hEE8B1AE0 , 32'h0EA49F60 , 32'h0BB19770 , 32'h0A2766D0 , 32'hF9BE8428 , 32'h02D85914 , 32'h06B12CD8 , 32'h06EE4CA8 , 32'h09BA6A20 , 32'h02862C0C , 32'hF9CC9FF0 , 32'hEAD61860 , 32'h03DFBC84 , 32'h09C09F20 , 32'hFCF138B8 , 32'h17645C80 , 32'h14D181E0 , 32'h0E2CA4A0 , 32'h02FE027C , 32'h12EED200 , 32'h10626380 , 32'hF3B50510 , 32'h04502B10 , 32'h0DA97AD0 , 32'hF684B6B0 , 32'h02D0099C , 32'h0388CA50 , 32'hF8D5FBA0 , 32'h05EF2670 , 32'hFEFB73CC , 32'h04727DD8 , 32'hF2B5BC70 , 32'h0594B948 , 32'h0E8B5E20 , 32'hFC0F1B64 , 32'h06533628 , 32'h00E0F71E , 32'h06C77BC0 , 32'h07043890 , 32'h0BB675A0 , 32'h08EC22D0 , 32'hF9825560 , 32'hFBB45F50 , 32'hFEC0BF88 , 32'hF718EA70 , 32'h08012140 , 32'h004EA311 , 32'h069E8F78 , 32'hFCFE314C , 32'hFFA4CF7F , 32'h01F6CB38 , 32'hFD2F9524 , 32'h003268C0 , 32'hFC5357D8 , 32'hFB3C66B0 , 32'hFF4600C3 , 32'hFFFFE623 , 32'hFFFD5C81 , 32'hFFFDD190 , 32'h0003D4E0 , 32'h0003306B , 32'h0003F6E0 , 32'h0001DA63 , 32'h000421ED , 32'hFFFD7F94 , 32'hFFFC1DB4} , 
{32'h131E4DC0 , 32'h00A8A10D , 32'h2706BAC0 , 32'hBD069280 , 32'h1972CD40 , 32'hF6DD32E0 , 32'h376DF840 , 32'hF9460080 , 32'hDB3E4380 , 32'h02813550 , 32'h0E3B55A0 , 32'h12920280 , 32'hF6EC3180 , 32'h158A9B40 , 32'hF66F45A0 , 32'h0CA48510 , 32'h03BEB0E8 , 32'hF213EFE0 , 32'h12E7BE80 , 32'h06E127A8 , 32'h2C49EC00 , 32'h0ABC7AD0 , 32'hFE38DC28 , 32'hE8AAE1A0 , 32'h22557000 , 32'hF665BB30 , 32'hFAF43A60 , 32'hF604C940 , 32'hF499DDC0 , 32'h03A86B9C , 32'hF30CF740 , 32'h16600E60 , 32'h0793F070 , 32'hE75F1700 , 32'hFC2107A4 , 32'hE2A72220 , 32'hF53D5730 , 32'hF684BA00 , 32'h053A5268 , 32'hEC606F80 , 32'h03A3A3E4 , 32'h1D982A40 , 32'h0B24B7F0 , 32'hF5D3C660 , 32'hF93AFD80 , 32'h036E1C98 , 32'h0EC8CCE0 , 32'h06200978 , 32'h065256A8 , 32'hE30977E0 , 32'h0051AF19 , 32'hF8766638 , 32'hF3F55BF0 , 32'h0F152030 , 32'hFD9D8F74 , 32'h0CD25CF0 , 32'h04B7EC60 , 32'hF1A9ED00 , 32'hFCDE0398 , 32'hFE6A56D4 , 32'hFBD80320 , 32'h092F3900 , 32'hF625D600 , 32'h08511950 , 32'hFE3012FC , 32'hFFF8B209 , 32'h068BFAA8 , 32'h06A72A20 , 32'hF9EA6330 , 32'hEEA88D20 , 32'hFE0EF974 , 32'h0F780A80 , 32'hFCB1F0C0 , 32'h0A93DF00 , 32'hF64D4050 , 32'hF52ECCF0 , 32'hF4A23230 , 32'h0D6DCA20 , 32'h09C50DC0 , 32'h03255354 , 32'h09478470 , 32'h02455B28 , 32'h00EE8B32 , 32'h0E1739A0 , 32'h01D5BFFC , 32'h00718EE5 , 32'h09CA7610 , 32'h03948CE0 , 32'h005E55A2 , 32'hFF568EAA , 32'h0002D40D , 32'h0000FC10 , 32'hFFFD06BA , 32'h00039247 , 32'h0001ABFA , 32'h00006E4E , 32'hFFFDB007 , 32'hFFFDD2E7 , 32'hFFFE6269 , 32'hFFFEE391} , 
{32'hFFFC9ABE , 32'hFFFD145D , 32'hFFFE8082 , 32'h000680CE , 32'hFFF7D2B3 , 32'h000529CA , 32'h0005B0FF , 32'h0001D174 , 32'hFFFB7B59 , 32'hFFF0AE95 , 32'h00085F1C , 32'h00001448 , 32'h0001BCE0 , 32'h0005EECB , 32'hFFF8ED07 , 32'hFFF7E948 , 32'h0006EE25 , 32'h000079EA , 32'hFFFED17B , 32'h00047FEE , 32'hFFFCEFD0 , 32'h00027456 , 32'h0000B8A9 , 32'h0008B59B , 32'h000634C3 , 32'hFFFAD507 , 32'hFFFF2C75 , 32'h0005AAAD , 32'h00019368 , 32'h00006C71 , 32'h0005B19A , 32'hFFFB1569 , 32'h0005E910 , 32'hFFFE761E , 32'hFFFD34AA , 32'hFFFE3671 , 32'h0003226B , 32'hFFFB6D4E , 32'hFFF07DAB , 32'hFFF88E52 , 32'hFFFE99A2 , 32'hFFFB80EB , 32'hFFFF68F4 , 32'hFFF678F1 , 32'h0001D457 , 32'hFFF7253B , 32'hFFFB7E3D , 32'hFFFDD91D , 32'hFFFA57DA , 32'hFFFE895B , 32'h0005CF8F , 32'hFFFC0894 , 32'h0008DF28 , 32'hFFFF04DA , 32'hFFFCB19B , 32'hFFF9C03A , 32'h0005AF43 , 32'h000011ED , 32'hFFF6E092 , 32'hFFFB55FB , 32'hFFFD8C54 , 32'hFFFE4D30 , 32'h0002F1F4 , 32'h000426FD , 32'h00023626 , 32'h0001FC62 , 32'hFFFEAC16 , 32'h00036FE5 , 32'h0001FBEB , 32'hFFFE2AC5 , 32'h00026B54 , 32'hFFFB4D06 , 32'hFFFDAA28 , 32'hFFFA8FF3 , 32'hFFFF8624 , 32'h000525AE , 32'hFFF9B8DA , 32'hFFF71016 , 32'hFFFFAE0A , 32'h00051DD5 , 32'h000285DB , 32'h00099124 , 32'hFFFD08C6 , 32'h0007C4F3 , 32'hFFFC9364 , 32'h0006AB3D , 32'hFFF89DEC , 32'h00049679 , 32'h00016D1A , 32'hFFFEDAC0 , 32'hFFFF3050 , 32'hFFFF0CE5 , 32'h00023EA0 , 32'h0000CD6A , 32'hFFFA2A14 , 32'h00053511 , 32'h0001D537 , 32'h0002DEF5 , 32'hFFFE23DD , 32'hFFFC9DBC} , 
{32'hD3AE7FC0 , 32'h6D35AC00 , 32'h7071B780 , 32'h7FFFFFFF , 32'hEDDA7EA0 , 32'hA34F4C00 , 32'h7FFFFFFF , 32'h0A2AFAB0 , 32'hE60154E0 , 32'hFEFE3500 , 32'h1668E9A0 , 32'hDFB17B00 , 32'hBB1E6580 , 32'h2907CB00 , 32'h1AE20420 , 32'hE8375000 , 32'hEF4BA380 , 32'h0A1768D0 , 32'hE48A5180 , 32'hE6DCD920 , 32'h1985BB60 , 32'h01F77BAC , 32'h21F35640 , 32'hF153EA60 , 32'hCD084E00 , 32'h04AA3370 , 32'hEE2E3EA0 , 32'hD385DB80 , 32'hEB380EE0 , 32'h0CB87130 , 32'h1132C800 , 32'hF2C0E060 , 32'hF4C09C60 , 32'hEA3363E0 , 32'h0545B730 , 32'h09BB4110 , 32'hE84B1B40 , 32'hFBCE0428 , 32'h0A651730 , 32'h0B91E3E0 , 32'h168843A0 , 32'h2E744680 , 32'h04615020 , 32'hF502BF10 , 32'hFCD80978 , 32'h07F5CE88 , 32'hF5900A20 , 32'h01DE78B8 , 32'hFF3A5A85 , 32'hFEFB0608 , 32'hF4A88C80 , 32'hF50D0590 , 32'h07D36AE0 , 32'hF31EC610 , 32'h01EEBE20 , 32'h12C6F860 , 32'h005CA88A , 32'h030E8234 , 32'h00E42843 , 32'h01B20BB0 , 32'hFD711174 , 32'hF4315160 , 32'h06730100 , 32'h01D9FEBC , 32'hFC3327A0 , 32'h001E1BD3 , 32'h10DA4B80 , 32'h0A9A4000 , 32'hFCC45A58 , 32'hFB936350 , 32'h04C572D8 , 32'hF9990828 , 32'hFF6D3324 , 32'hFC1F9AD8 , 32'hFE71D4C4 , 32'hF53C4890 , 32'hFF740E6D , 32'h04661CA0 , 32'hF15BFDD0 , 32'hFBE74F98 , 32'hFC1827A0 , 32'hF753ECF0 , 32'h00D799E4 , 32'hFBBC1208 , 32'hFCCF00D8 , 32'h09CCEE90 , 32'h00DBF082 , 32'hFFBECCDA , 32'hFCF82344 , 32'h00D4A570 , 32'hFFFDAD71 , 32'h0003D86D , 32'h0001474E , 32'h000337AE , 32'hFFFF672C , 32'hFFFAB0AD , 32'h00017DCD , 32'h00004064 , 32'h0002075E , 32'hFFFDBD73} , 
{32'h0008FDAA , 32'h0006D5A5 , 32'hFFFC0B44 , 32'hFFFB5A1B , 32'h000199F1 , 32'h00026A78 , 32'hFFFB1183 , 32'h0005CCCB , 32'hFFF740D6 , 32'hFFFC5F48 , 32'hFFF71A2B , 32'h0008B81A , 32'hFFFA475F , 32'h0002F13B , 32'h00065EBA , 32'hFFF9EDEE , 32'hFFFEFEA0 , 32'h00009C81 , 32'h00085E7B , 32'h00024036 , 32'hFFFAAC37 , 32'h0004D1CF , 32'h00023019 , 32'h0003D307 , 32'hFFFAA8D1 , 32'h0002CB02 , 32'h0005A82F , 32'hFFFBE743 , 32'hFFF70385 , 32'h000769FA , 32'hFFFEE29E , 32'h0005E538 , 32'h00037807 , 32'h0001CF85 , 32'h00048B3B , 32'hFFFABEA8 , 32'hFFFDC9A2 , 32'hFFF689C5 , 32'hFFF3FC69 , 32'hFFFD26AC , 32'hFFFD8A71 , 32'h0000B5CE , 32'h00053462 , 32'hFFF5ED5F , 32'h0002E0B0 , 32'hFFFF7080 , 32'hFFFFC140 , 32'h00015231 , 32'hFFFDD588 , 32'hFFFDD9B8 , 32'hFFFCE9C0 , 32'hFFFE224F , 32'hFFFD5D62 , 32'h00030874 , 32'hFFFE76CE , 32'h00048CA1 , 32'h00051E82 , 32'hFFFF5479 , 32'h0002EF50 , 32'h00038121 , 32'hFFFFF102 , 32'h0005D6B5 , 32'hFFFD973F , 32'hFFFD2BAE , 32'hFFFBAF97 , 32'hFFFFF5E3 , 32'h00069162 , 32'h00045B1E , 32'hFFFFFE62 , 32'h0006AE27 , 32'h0002A01D , 32'hFFFDAFB0 , 32'hFFFA488A , 32'hFFFCA82F , 32'h0004BA57 , 32'h0000BC3A , 32'hFFFCE8A1 , 32'hFFFB9276 , 32'h00016AA6 , 32'h0007CBC4 , 32'h00034BAA , 32'hFFFD0013 , 32'h000006ED , 32'h0003C13D , 32'h00032697 , 32'h00044892 , 32'h0001227B , 32'hFFFD2C06 , 32'h00031D96 , 32'hFFF794D0 , 32'hFFFD3384 , 32'h000B738B , 32'h0000A70F , 32'hFFF7EB9A , 32'hFFFF7402 , 32'h0001A385 , 32'hFFFEE22E , 32'h0005A053 , 32'h00011FFB , 32'h0005A8BD} , 
{32'hFFFE92C1 , 32'h0001CC23 , 32'h000AFC9F , 32'hFFFAE689 , 32'h0000835D , 32'hFFFA007A , 32'hFFFBFF25 , 32'h00048C83 , 32'h0008B730 , 32'hFFF4DDEE , 32'h0000C6FB , 32'h00005B56 , 32'hFFFF8CE4 , 32'h00002BD1 , 32'hFFFFB384 , 32'hFFFFE553 , 32'hFFFF01C8 , 32'hFFFDBD7D , 32'h000366B4 , 32'h00029C01 , 32'hFFFCCFCE , 32'h0004FB29 , 32'h0000C255 , 32'hFFFF2C6C , 32'hFFFB5B4F , 32'hFFFB8A04 , 32'h00065764 , 32'h00038ABD , 32'hFFFD89AA , 32'hFFFAE502 , 32'hFFFA6285 , 32'hFFF57D13 , 32'hFFFFFBC8 , 32'hFFFB0905 , 32'h0006C85E , 32'hFFF7C3A6 , 32'hFFF75A94 , 32'h00055F84 , 32'h00005DA0 , 32'h00003019 , 32'hFFF3D84D , 32'hFFFDF0B8 , 32'hFFF7B8A1 , 32'h000465D7 , 32'hFFF91C84 , 32'hFFFC732E , 32'hFFFF1351 , 32'h0003BB6A , 32'h00024FA8 , 32'hFFFFC6CE , 32'h00057E31 , 32'hFFFD293E , 32'hFFFE723F , 32'h0001566B , 32'hFFF6D0F4 , 32'hFFFFD26A , 32'h0005DC08 , 32'hFFFEC952 , 32'hFFFE1308 , 32'hFFFE428B , 32'h00004781 , 32'h00086181 , 32'hFFFDE889 , 32'h00006501 , 32'h0004FD84 , 32'hFFF9944E , 32'hFFFBE999 , 32'hFFFD1880 , 32'hFFFD1D78 , 32'hFFFD00C0 , 32'hFFFFD4E3 , 32'h00069CB6 , 32'hFFFD676C , 32'h000316AD , 32'hFFFF84D0 , 32'hFFFC7415 , 32'h0005E847 , 32'hFFFB25B2 , 32'hFFFBB79E , 32'hFFFA9C30 , 32'h0004EBFE , 32'h0003BC23 , 32'h00004B1F , 32'hFFFB97DA , 32'hFFFCACC0 , 32'h00028D2F , 32'hFFF56AD3 , 32'hFFF97A6B , 32'hFFFED504 , 32'h00026E39 , 32'hFFFBA2C1 , 32'h0000956C , 32'h000471A1 , 32'hFFF5AF76 , 32'hFFFE420C , 32'hFFFF0BE7 , 32'h00078385 , 32'h000553B7 , 32'hFFFA7388 , 32'h00025A37} , 
{32'h56AD7600 , 32'hE8DA92C0 , 32'h00E8D800 , 32'hD5857D40 , 32'h64925100 , 32'h25AD7740 , 32'hDB8317C0 , 32'hFB033088 , 32'hE2A338E0 , 32'h272EC9C0 , 32'h19644A40 , 32'hF3187640 , 32'hFEB5E2CC , 32'hC053F900 , 32'h20C3D080 , 32'hFF364759 , 32'h1158DD60 , 32'h154E11C0 , 32'hFEEEC00C , 32'hD99E0E40 , 32'h13CCB960 , 32'h0E924A40 , 32'h1637AEA0 , 32'h0A22F4C0 , 32'hEF144D20 , 32'h22D74980 , 32'h091EDDF0 , 32'hFDB5DB10 , 32'hEE11F100 , 32'hFA08EE58 , 32'h071886D0 , 32'hE70D4F20 , 32'hF8EA5820 , 32'h0F9D6B30 , 32'hF3275800 , 32'hEB7514A0 , 32'hD477C540 , 32'hF6F152E0 , 32'hF71B3310 , 32'h12478700 , 32'h0B7A3470 , 32'hF847FDB0 , 32'hEF215160 , 32'h08E9C3C0 , 32'hFCD588F8 , 32'hED95AA20 , 32'h0632DB18 , 32'h0BD6A280 , 32'hFBF33428 , 32'h0C3A92A0 , 32'h15210CA0 , 32'hEF1B98E0 , 32'hFA09A2C0 , 32'hFF66027B , 32'h1E9EDF40 , 32'hF71CA970 , 32'h010EEBC4 , 32'hE65011A0 , 32'h0AB7B190 , 32'hFDB18F20 , 32'h03E1A238 , 32'h08982570 , 32'hF776D140 , 32'hF42BF810 , 32'hF9EBDBC8 , 32'h089F8E00 , 32'hFC631A28 , 32'h0A562090 , 32'h0F628780 , 32'hFCEC6B08 , 32'hF88E1D60 , 32'hFB69A5B0 , 32'h0516C930 , 32'h0936C050 , 32'hFD352580 , 32'hFE2E7C94 , 32'hFD7BA784 , 32'hFD457118 , 32'h0A2EC790 , 32'hFC71EE04 , 32'h02CB93A0 , 32'hFCAE30F0 , 32'h00986BDB , 32'h02A5A980 , 32'h0A0AF220 , 32'h05073638 , 32'h036F848C , 32'hFFC218B2 , 32'hFDCAE588 , 32'h076D4E00 , 32'h000248A9 , 32'hFFFEE6CB , 32'hFFFE3ACE , 32'hFFFFE1E2 , 32'h00026A89 , 32'h0000735E , 32'h00003F17 , 32'h000188A3 , 32'hFFFEF3FA , 32'hFFFECE6B} , 
{32'h0F66E1F0 , 32'hF936D590 , 32'hEF9CA360 , 32'hDD08F380 , 32'hF0F7BE50 , 32'hF4C96750 , 32'h0353510C , 32'hEE004DC0 , 32'hE99A8A80 , 32'h0B5F59F0 , 32'h142B2CE0 , 32'h0CD76B30 , 32'h0745D390 , 32'hE0E76020 , 32'hFEF323D4 , 32'h0F9892C0 , 32'h03708440 , 32'hFBD5B158 , 32'hE8AF5D20 , 32'h07D53890 , 32'hE468E200 , 32'h06B5E960 , 32'hF1798EB0 , 32'h0147EFFC , 32'h08331F90 , 32'h17C4D220 , 32'hFA6D6D58 , 32'h0426F068 , 32'hF3240600 , 32'h07372920 , 32'hFC3D6510 , 32'hFCEB706C , 32'hFD82A5AC , 32'hFCD47EB8 , 32'h0CCFEDB0 , 32'hFCB0CF18 , 32'h08376270 , 32'hF8F7FF88 , 32'hFEB837C4 , 32'h015A2E80 , 32'h0223AE44 , 32'h04581CF8 , 32'hF4F910F0 , 32'h0EC2A130 , 32'hFB3CF920 , 32'h00F5328D , 32'hFB84D058 , 32'hFD0962F0 , 32'hF65622D0 , 32'h04751FF0 , 32'h01C04D0C , 32'h0099D7FA , 32'h08A118F0 , 32'hFD7438E8 , 32'hF4B3CCB0 , 32'h08986FC0 , 32'h052A8CF0 , 32'h041D9F08 , 32'hFDDE5FE8 , 32'hF677E750 , 32'h05C35228 , 32'hF663FCD0 , 32'hFF31BAC7 , 32'hF6ACA530 , 32'h00D0340A , 32'h07D3D828 , 32'hF62485F0 , 32'h18847740 , 32'h0C70D000 , 32'hFF77515D , 32'h01F5A380 , 32'hFDE2835C , 32'h0BEC5E30 , 32'hF4CBA520 , 32'hF9884308 , 32'hF8A005E8 , 32'h05F92DB0 , 32'h025AF5B4 , 32'hF868E670 , 32'h0A20B250 , 32'hFC108250 , 32'hFE1E91E4 , 32'hF5EDCF80 , 32'hFFECEE27 , 32'hFBC07DA8 , 32'h018F37E0 , 32'h06EA1EC8 , 32'h000408BD , 32'h0075BFB4 , 32'hFFAAC2EE , 32'h0004ACD6 , 32'hFFFCEF5A , 32'h0000389A , 32'hFFFFE9EB , 32'hFFFAB518 , 32'h0000E81B , 32'h00048C2F , 32'hFFFD0517 , 32'h0001E371 , 32'h0001DFDC} , 
{32'h1094AA60 , 32'hF3A72ED0 , 32'hFBFF0EA8 , 32'hE2B794C0 , 32'h102D38A0 , 32'hE0184B80 , 32'hFA525718 , 32'hE5B7CF00 , 32'h0CFC69B0 , 32'h07B18E70 , 32'hFC76C210 , 32'h10F297E0 , 32'h156A2560 , 32'hE63F3E60 , 32'hF310EC60 , 32'hE74B3100 , 32'h0AF7CDC0 , 32'hF5994D50 , 32'hE7BCDA80 , 32'h067461C8 , 32'hF1D52290 , 32'hEEC5ACA0 , 32'h16887C20 , 32'hFFCDB038 , 32'h07106738 , 32'hFAE401C0 , 32'hFFD30DBA , 32'hFE34B5AC , 32'h0E511DC0 , 32'h13EB0F20 , 32'hEB1D1A00 , 32'h0246878C , 32'hEEFF1080 , 32'hE1412AA0 , 32'hF4CFA730 , 32'h148B9DE0 , 32'hDE3FAFC0 , 32'hFF71182C , 32'h0316DF24 , 32'hFD0E4FD8 , 32'h04C7ED90 , 32'hFC80C6B0 , 32'h022F63B8 , 32'h1013D6A0 , 32'hF17D1A10 , 32'h06979250 , 32'hFFF6551D , 32'hF5BA92D0 , 32'hF807E638 , 32'hFF831E5F , 32'hF9FFAC18 , 32'hF2E3AE40 , 32'h11A66E60 , 32'hF870ECC0 , 32'h03A1A118 , 32'hFFDD5BFC , 32'hF3EF07D0 , 32'h09264930 , 32'h09CE74C0 , 32'hF5AE9820 , 32'hFF44298E , 32'h01362D68 , 32'h03DD9D0C , 32'hF9292460 , 32'hFA5D9670 , 32'hFC581CAC , 32'hFDDAF8BC , 32'hF3E11FE0 , 32'h04185C50 , 32'hFBD9B300 , 32'h021CB208 , 32'hF7785B30 , 32'hFCFBED68 , 32'hFDCFF0AC , 32'h06EAAE00 , 32'h0ADF1D30 , 32'hFBD3A750 , 32'h02FE4308 , 32'hFED72F4C , 32'hFDD58730 , 32'h015D4BF4 , 32'hFA90BEA8 , 32'hFF2438F6 , 32'hFC2580BC , 32'hFE0384B8 , 32'h0415E088 , 32'hFE71DE34 , 32'h00AD516F , 32'h0168DFA4 , 32'hFFD8CA5B , 32'hFFFFA351 , 32'hFFFFA81B , 32'hFFFECFA9 , 32'h00074A43 , 32'hFFFCBF1E , 32'h000442D5 , 32'hFFFFD4A4 , 32'hFFFF0A49 , 32'hFFFF5C3A , 32'h00013416} , 
{32'hFFF86F7D , 32'hFFFF00EA , 32'hFFFE4AB0 , 32'hFFFF2C03 , 32'hFFFFA408 , 32'h00067A9C , 32'h0001C376 , 32'h00002997 , 32'h00014B5A , 32'hFFFE6E3F , 32'hFFFACC72 , 32'h0001E808 , 32'hFFFA478C , 32'hFFFCF40E , 32'hFFFDA96D , 32'hFFFB3DC1 , 32'hFFFB2ECB , 32'hFFFE5A3F , 32'h0001795D , 32'h0005EF97 , 32'hFFF92CC2 , 32'hFFFF138A , 32'hFFFA3301 , 32'hFFFC1E2C , 32'h000703C6 , 32'hFFFB2753 , 32'h0002ACE0 , 32'hFFFAE880 , 32'h0002315B , 32'hFFFEDC12 , 32'hFFF95FA7 , 32'hFFFC3BE4 , 32'h0004138B , 32'hFFFE11CD , 32'hFFFBFF27 , 32'hFFFFD442 , 32'h0006F5ED , 32'h0004B8FB , 32'h0003BCAB , 32'hFFFD9EE6 , 32'h0000CF42 , 32'h00004A4A , 32'h0004230A , 32'h0002F769 , 32'h0005221C , 32'h0001396B , 32'h00021859 , 32'hFFFE52FB , 32'h00018E38 , 32'hFFFD5F8D , 32'h000FC341 , 32'h00047336 , 32'hFFFD4E35 , 32'h00004DCD , 32'hFFF4EE50 , 32'hFFFF0527 , 32'hFFFCBBFA , 32'h0002ADB7 , 32'h00017957 , 32'hFFFE2243 , 32'hFFFA1C6F , 32'h0000D31D , 32'hFFFB83A3 , 32'hFFFC6ED3 , 32'hFFFCF168 , 32'h0001CF42 , 32'h000A5653 , 32'h00025AAC , 32'hFFFC83F9 , 32'hFFF87BA5 , 32'hFFFB011C , 32'hFFF72AE4 , 32'hFFF6CB91 , 32'h00060A58 , 32'hFFFC3877 , 32'h00012C31 , 32'hFFFDDF67 , 32'hFFFF70A5 , 32'h00015FF7 , 32'hFFFF8C26 , 32'h0004B2A1 , 32'h00027919 , 32'hFFFE2E04 , 32'h00019086 , 32'hFFF9DE54 , 32'h0000C057 , 32'h0003FBE4 , 32'hFFFE3B51 , 32'hFFFAF709 , 32'h000023B7 , 32'hFFFD4EF7 , 32'h000219EB , 32'hFFF6CAF1 , 32'h0004B9B9 , 32'hFFF740F6 , 32'h000191D8 , 32'h00009E96 , 32'h00030710 , 32'hFFFF83AD , 32'h0003FB34} , 
{32'h6886B400 , 32'h2FE32580 , 32'h7FFFFFFF , 32'h1A3487A0 , 32'hCBEE5B80 , 32'h018FE6F0 , 32'hFBB7EE60 , 32'h3A8FD680 , 32'hFB9A3488 , 32'h9187DA80 , 32'h263D1000 , 32'hCE1FE980 , 32'hFB511BE8 , 32'h16738940 , 32'h085C4110 , 32'hFD9CFFF0 , 32'h206CD5C0 , 32'hE1416540 , 32'hE3EEEAE0 , 32'h1222D3E0 , 32'h27BD3CC0 , 32'h21353C80 , 32'hE4C0A440 , 32'h1235CE40 , 32'hD66B06C0 , 32'hE81413E0 , 32'h04243980 , 32'h07341738 , 32'hE2367800 , 32'hEBF27CE0 , 32'h1EFCD000 , 32'hFBB6ECE0 , 32'hF82B7BC0 , 32'h0EBEA0F0 , 32'h24465B00 , 32'h03F19CE4 , 32'h033F1AFC , 32'hE2105FA0 , 32'hF0CFAF90 , 32'h0E6E82C0 , 32'h0A6FBEC0 , 32'hEF0EA500 , 32'h0BB92CB0 , 32'hFD7203D4 , 32'hFEA865B4 , 32'h014ACCF8 , 32'h114961C0 , 32'h164DB700 , 32'hF3DD6390 , 32'hFA9DBEF0 , 32'hF84D4740 , 32'hEDC54860 , 32'h08AC5470 , 32'h044D21D0 , 32'hF99B1538 , 32'h00CA86EB , 32'h0A3AF230 , 32'h03E23170 , 32'h02F5FCDC , 32'hF28560E0 , 32'h0AD67750 , 32'h052029C8 , 32'hF2FA0420 , 32'h0B8B0150 , 32'h05E11C88 , 32'hFD343C54 , 32'h05F59CF0 , 32'h01E8B1C0 , 32'hF6D2D2A0 , 32'h0658E740 , 32'h008AA911 , 32'hFC044E68 , 32'hFE093E4C , 32'hF6EEE720 , 32'hF8CF27A8 , 32'h0F7F6670 , 32'hFBEA0D78 , 32'hFA8C2190 , 32'h08822030 , 32'h06941FE8 , 32'h02A2581C , 32'h026FE7AC , 32'h01A69744 , 32'hFCC134FC , 32'hFFDC49E1 , 32'h01600358 , 32'hFD189644 , 32'hF9F10E68 , 32'h02CF4EDC , 32'h00605F42 , 32'h00018960 , 32'hFFFD993F , 32'hFFFC678E , 32'hFFFB93AE , 32'hFFFE2C58 , 32'h00006DEF , 32'h000022AE , 32'h000393AE , 32'hFFFFF7CB , 32'hFFFF4B8D} , 
{32'h1FE4A1E0 , 32'h0024AF7E , 32'hF31AAFC0 , 32'hE1074A80 , 32'h115DA940 , 32'hEDC18E60 , 32'h07A07328 , 32'hFBF9D7C0 , 32'h119AF800 , 32'h08BFAA60 , 32'h203FC140 , 32'h1190A100 , 32'h023011E8 , 32'hE464E1A0 , 32'hFB32FD60 , 32'h183624E0 , 32'h021F4F84 , 32'hFC7DE994 , 32'h03406D34 , 32'hFBF8F4E0 , 32'hF52E0370 , 32'hF94FBA08 , 32'h0CAA8710 , 32'h09A79410 , 32'hFF4DAFB5 , 32'h16D722A0 , 32'h086608F0 , 32'hF84F7248 , 32'hFEFC90D8 , 32'h141F1E60 , 32'hFB68C1C8 , 32'hF588DDF0 , 32'h111AC780 , 32'hF84A07D0 , 32'h07088E90 , 32'h02BEF2B0 , 32'h01DC0858 , 32'hFBBF34D8 , 32'hFFCB2AAC , 32'h03CFFB0C , 32'hFE676418 , 32'h048E5240 , 32'hFB34EE88 , 32'h0719EEB8 , 32'hFD2D14E8 , 32'h0EDFCEE0 , 32'h023D6874 , 32'hF19E32A0 , 32'hF5C3B300 , 32'h10E172C0 , 32'hFC339F10 , 32'hF692E900 , 32'h11779F60 , 32'hEFE14AA0 , 32'hFF3BB0A9 , 32'hF01E0800 , 32'hF844E878 , 32'hFD8F6858 , 32'h06CDA370 , 32'hFED737CC , 32'h03EF16B8 , 32'h0438A790 , 32'hFC2D7E30 , 32'h0422CD68 , 32'h03CBECDC , 32'h0420EF18 , 32'h07054D38 , 32'h00DCA426 , 32'hFFA1413F , 32'h04BC1C90 , 32'hFF8799A1 , 32'h01A4E080 , 32'h00F4FF8D , 32'hFFE1CA2B , 32'hFEE26874 , 32'h016A0B30 , 32'hF9BC8F38 , 32'h01F6B3DC , 32'h02B17F14 , 32'h07DB50E0 , 32'h02C1F2BC , 32'h08445250 , 32'h0546C0B0 , 32'h027AF6A0 , 32'h024E0794 , 32'h00AE5AF0 , 32'hFBAB1500 , 32'hFECC1428 , 32'hFC644CC4 , 32'hFF0C84D1 , 32'hFFF74E24 , 32'h00069941 , 32'hFFFBC3D9 , 32'h000476EC , 32'hFFFFD291 , 32'hFFFACCC8 , 32'h000991F9 , 32'hFFFC6BA9 , 32'h00046AA9 , 32'h00007F2F} , 
{32'h3741F380 , 32'h0BFF33D0 , 32'h367A1F00 , 32'h16B67F80 , 32'h4321A780 , 32'hFD613AA0 , 32'h28025500 , 32'hEFA24C40 , 32'h0C3DB180 , 32'h057D6868 , 32'hE660B9A0 , 32'h04D5FA50 , 32'hF7CD3F40 , 32'hEA92B0A0 , 32'h06651CC0 , 32'hF4C8D720 , 32'h3374C680 , 32'hDF72BE40 , 32'h058FF4B0 , 32'h0C70CF70 , 32'hC626CE00 , 32'hFED47D54 , 32'hE4468A60 , 32'h02A008B8 , 32'hE79865C0 , 32'hF5B77970 , 32'hDDF8A940 , 32'hDF4D5E80 , 32'hEA2ABE20 , 32'hF9FEF488 , 32'h2B3B67C0 , 32'h12E48460 , 32'hF63753C0 , 32'h0961C7E0 , 32'hFA9993B8 , 32'h15D654E0 , 32'h0BB42F70 , 32'h08B72F60 , 32'hD02D9A40 , 32'hF22171B0 , 32'hFCA06440 , 32'h12446AE0 , 32'hF6992790 , 32'hF6FC37C0 , 32'h297D62C0 , 32'h1110A280 , 32'hFE3BED78 , 32'h1119D400 , 32'h10DE21A0 , 32'h0A8D7060 , 32'hFF90AD53 , 32'hFE9B42C8 , 32'hF8780D58 , 32'hFCDD118C , 32'hEDC6ABA0 , 32'hF552E910 , 32'hFEEFFC58 , 32'h0FD09040 , 32'h0CE69A30 , 32'h1F9D05A0 , 32'h02BE8ED0 , 32'h0DC6BD40 , 32'h002351A7 , 32'h07C00388 , 32'h04BBB298 , 32'hFE6F28D4 , 32'hFF93D090 , 32'hFCDC88FC , 32'h03EDAE4C , 32'h02ECEAF8 , 32'h03EC3C78 , 32'hFDC13B90 , 32'h00A6146F , 32'h0304F64C , 32'hF6C5B390 , 32'hF9A5CE30 , 32'h06045F90 , 32'h06E78AC0 , 32'h052264B0 , 32'hFDE0FC4C , 32'hF8419870 , 32'h039E0E14 , 32'hF704DC90 , 32'hFEA22748 , 32'h0148835C , 32'hF6667D40 , 32'h00E568A0 , 32'h0639FF58 , 32'h014C8D04 , 32'h00B6527D , 32'h000159F4 , 32'h00020ACA , 32'hFFFB415E , 32'h00016CEB , 32'hFFFEB8E3 , 32'hFFFB0DFD , 32'h00010339 , 32'hFFFCE16D , 32'hFFFD24ED , 32'h000039F7} , 
{32'hF69C3FB0 , 32'h35525080 , 32'h7AA12B00 , 32'hB4AAAD80 , 32'h1155E200 , 32'hCFE2A740 , 32'hF2F00270 , 32'h0B747A00 , 32'hE4DEF5E0 , 32'hD7CA0540 , 32'h0A512E80 , 32'h24B40A00 , 32'h047FC528 , 32'hFAFADDD0 , 32'hE11651C0 , 32'h06B01898 , 32'hD12FEC80 , 32'h470C7E80 , 32'hF4177A50 , 32'h1A40D8A0 , 32'hD96E1F40 , 32'h05CEB608 , 32'hF9AB6298 , 32'h283F5900 , 32'h04819FA8 , 32'hF1BDC910 , 32'hE3B885C0 , 32'h0BDB8D80 , 32'h02159B98 , 32'h0FAE5320 , 32'hECBC5AE0 , 32'hFD909490 , 32'h13B4A8E0 , 32'hF67A8FA0 , 32'hE84D6220 , 32'hDED4B740 , 32'hE7D72260 , 32'hF050F1D0 , 32'hE78C3A40 , 32'h0856BA30 , 32'hED523A60 , 32'hE02AC180 , 32'h1D95F860 , 32'h0741F590 , 32'h193A1760 , 32'hFA5829F8 , 32'hFFCFA604 , 32'h0FFA6980 , 32'hF7071DF0 , 32'hEF3735E0 , 32'h0BE60E10 , 32'hF7DA7360 , 32'h0174DE48 , 32'h006C1E46 , 32'hF9DCC200 , 32'h121479A0 , 32'h0D65AD10 , 32'h035E1F58 , 32'hF1B38F30 , 32'h048812F8 , 32'hED85E7C0 , 32'h02F43734 , 32'h064F7B48 , 32'hF509B270 , 32'hECD56CC0 , 32'h010269B8 , 32'h076616E0 , 32'hFBB2E3E8 , 32'hFBFFDCC8 , 32'hFFCD4669 , 32'h0B3C3620 , 32'hF8BBE140 , 32'hFCB7FBB8 , 32'hFB592BD0 , 32'h06F15FB0 , 32'hFEB2079C , 32'h072350D8 , 32'hFE3E3D88 , 32'hFFBF62DE , 32'hFF997664 , 32'h015B5644 , 32'h012234AC , 32'h0703B360 , 32'hFCE6FE44 , 32'h05E5B280 , 32'hFD8A5054 , 32'hF8FE6220 , 32'h01EFC398 , 32'hFD611F54 , 32'h01109BA0 , 32'hFFFF574B , 32'hFFFEF6A4 , 32'hFFFEB8B1 , 32'h0001552F , 32'hFFFF6676 , 32'hFFFC84EE , 32'h00059FC7 , 32'hFFFDA8E2 , 32'hFFFF51DF , 32'h0001606E} , 
{32'hF7715710 , 32'hBA071F80 , 32'hEB997360 , 32'h177CB100 , 32'h1F75B640 , 32'h1C900320 , 32'hC267CE00 , 32'h554DAE80 , 32'h16E00940 , 32'h1F515F80 , 32'h18CF84A0 , 32'hF4051800 , 32'h10411440 , 32'h08676A60 , 32'hF6345130 , 32'hEB136EA0 , 32'h14B12040 , 32'h0A923750 , 32'hDA9EF400 , 32'hDD4973C0 , 32'hBD33A400 , 32'hEF5758A0 , 32'hEFB52B60 , 32'hC6A27E80 , 32'h238C8B40 , 32'h0E7900E0 , 32'h1187D360 , 32'hD8D20100 , 32'h0854C880 , 32'h0F1544A0 , 32'hFC87208C , 32'hEA62E520 , 32'h1A1AD120 , 32'hEF04E700 , 32'h17A554A0 , 32'hFDC53558 , 32'h006AE295 , 32'hDC873B40 , 32'h13B62BE0 , 32'h15EBE4A0 , 32'h184AB860 , 32'h11C1B220 , 32'h09F915C0 , 32'hEDF9D3A0 , 32'hFB9DE3C0 , 32'hEE007BA0 , 32'hE79611E0 , 32'h05D89238 , 32'h03716804 , 32'h07C9A898 , 32'h1A4C4200 , 32'h053169E0 , 32'hF0652100 , 32'h05560320 , 32'hFCADD3CC , 32'h056B5000 , 32'h05B5DFA8 , 32'hF6849590 , 32'hF7DD3500 , 32'hF201C910 , 32'h1B09D420 , 32'h05A74370 , 32'hF65C9C80 , 32'h0F53DE90 , 32'hF67CC870 , 32'h0746FCD8 , 32'h0C69FFD0 , 32'hF64E9000 , 32'hF85F32F0 , 32'h09978D90 , 32'h0517E630 , 32'h0189DED8 , 32'h0075C517 , 32'h02CD67E4 , 32'hFE96FBD0 , 32'h07505D40 , 32'h0443E7E0 , 32'h01F740B8 , 32'hFF6706D2 , 32'h0160CB90 , 32'h036F5938 , 32'h05267868 , 32'hFC8C7958 , 32'h04AF4FB0 , 32'hFB566C50 , 32'hF724F7D0 , 32'hFB9D0D10 , 32'h0017553D , 32'h03D86424 , 32'h0124DFCC , 32'hFFFEFE10 , 32'h0003899B , 32'hFFFFA76D , 32'h0001D4CB , 32'hFFFEC3E7 , 32'h00000488 , 32'hFFFD3B3D , 32'hFFFF7CFD , 32'h00001F12 , 32'hFFFE3C20} , 
{32'h7FFFFFFF , 32'hF4B95590 , 32'h5EDCC580 , 32'h993F7980 , 32'hB11C2F00 , 32'h1904E140 , 32'hD7D75F00 , 32'h1BF2E040 , 32'h35FA7F40 , 32'h212CD700 , 32'hFBFDF718 , 32'hE9AA79C0 , 32'h312F8980 , 32'h19C21B20 , 32'hE8CDA1C0 , 32'h20A8F000 , 32'hFA20C2F8 , 32'h22977440 , 32'h30FB70C0 , 32'h03796BFC , 32'h14E988C0 , 32'h4CD67600 , 32'h030D9F4C , 32'hD6B43180 , 32'h02F1F690 , 32'h03199564 , 32'hEC9946A0 , 32'hF5F4C610 , 32'hEC103D60 , 32'h14D6DF00 , 32'hF7939FC0 , 32'hE2418440 , 32'hD45ECD80 , 32'h0D319F20 , 32'hE6047640 , 32'hF6518030 , 32'hF040EAE0 , 32'h0E3914D0 , 32'hEE9FF140 , 32'hF37F3190 , 32'h05363440 , 32'hF76DAAB0 , 32'hF51C4310 , 32'hF705A810 , 32'hE5498240 , 32'h1C37BEC0 , 32'h0C170460 , 32'h0B7DF9A0 , 32'h0EA6D520 , 32'h0C907DB0 , 32'hF34DA150 , 32'hFEA313D4 , 32'h0B309ED0 , 32'h022E6778 , 32'hF2AB21E0 , 32'h046C0E60 , 32'h0B2C0040 , 32'hF30E86B0 , 32'hFF79729E , 32'h08D18ED0 , 32'h0B8AC080 , 32'h07275C20 , 32'h04DD9F20 , 32'hFEC37738 , 32'h02507B50 , 32'h0C5D7B50 , 32'hFB6060E8 , 32'hFEDDBA5C , 32'hFBDFA718 , 32'hF98D4298 , 32'h0A190200 , 32'h016B4858 , 32'h04CAF928 , 32'h03115648 , 32'hFD2CDA0C , 32'h049CCB40 , 32'h00F8E718 , 32'hF6F62550 , 32'h07189940 , 32'h0516C630 , 32'hFDD43488 , 32'hFE0C89E4 , 32'hFDC46760 , 32'hFEC248C8 , 32'h00BF69D9 , 32'h03BFD92C , 32'h025B2F68 , 32'hFE18EEC0 , 32'h01703E2C , 32'hFFCAE780 , 32'hFFFFF032 , 32'h00030B36 , 32'hFFFCE0F2 , 32'h0005F383 , 32'h00002428 , 32'h00036B76 , 32'h00012722 , 32'hFFFBC3CB , 32'hFFFF7FEF , 32'hFFFEEAD6} , 
{32'h01AD7814 , 32'h0EA00650 , 32'hFADF03C0 , 32'h066A9360 , 32'hFADF7260 , 32'h031925A8 , 32'hFA35F4A0 , 32'h084AB110 , 32'h05207658 , 32'h075236B8 , 32'h04B87D80 , 32'hFAD5CF50 , 32'hFB9E6490 , 32'hFACE3C08 , 32'hF8CFDFB0 , 32'h09F22220 , 32'hFA2448E8 , 32'h0221F288 , 32'h05EF3FF0 , 32'h0C04A190 , 32'h0FCF0D90 , 32'hFD68F004 , 32'hF40D27F0 , 32'h02113FEC , 32'h06338580 , 32'h01F50664 , 32'h065812B8 , 32'hFAF1F8E0 , 32'h03945C80 , 32'h03A50984 , 32'h0270A448 , 32'hFE651F20 , 32'h032B693C , 32'hF674F420 , 32'h0A9C5CF0 , 32'hFCAABF60 , 32'h09A208C0 , 32'h0038C218 , 32'hF8184418 , 32'hFAF9F968 , 32'h07894A58 , 32'hFE3D285C , 32'hFC3F6BDC , 32'h00F41A9A , 32'hFF49F734 , 32'hFB4AD838 , 32'h00917C8C , 32'hF8C5C6E8 , 32'h07DA7AC0 , 32'hFCF3B87C , 32'h0FD13B70 , 32'h0A1F27F0 , 32'hFD5F55F8 , 32'hFEA2EC38 , 32'hFDE45C40 , 32'h007811C6 , 32'h09E74F70 , 32'hFD503364 , 32'hFC8AAEA0 , 32'hFD13EE50 , 32'hFDB9BBC4 , 32'hF8F12488 , 32'h0332576C , 32'hFB1F18B0 , 32'h05D412A0 , 32'h061F0EC0 , 32'hFE153C84 , 32'h07364970 , 32'hFCBFCCEC , 32'h02FF4870 , 32'h0803C210 , 32'hFD8A54E8 , 32'hFD52B6E0 , 32'h00881E1E , 32'hFF17B442 , 32'hFDB0E56C , 32'h00FA6D14 , 32'h0009B1D3 , 32'h007D0F12 , 32'h031FF974 , 32'h025B424C , 32'hFEEEA174 , 32'h00C2514D , 32'h01E00E58 , 32'h024AC0C4 , 32'h02EABFE4 , 32'h04EEC188 , 32'h000B5C0F , 32'hFF19EC0C , 32'hFFE1B69A , 32'h00080074 , 32'hFFFFAAB9 , 32'h000D4D9D , 32'hFFFEEB79 , 32'h0001D522 , 32'hFFFFAC8C , 32'h0003BE61 , 32'hFFFE6E44 , 32'h0004E450 , 32'hFFFE0927} , 
{32'hB65BDB80 , 32'h310EE100 , 32'hEF17D6C0 , 32'h19F820C0 , 32'h0B4ECBF0 , 32'hE0FA4460 , 32'hEE186660 , 32'hEC686F40 , 32'hFD9A30DC , 32'hFC1E38A4 , 32'hE5271240 , 32'hFC4B825C , 32'hD9376CC0 , 32'hF3DD4920 , 32'hFB06E5C8 , 32'hFD01F3CC , 32'h0E07D980 , 32'h0E29C3A0 , 32'hE754A340 , 32'h24ECADC0 , 32'h0B2DC380 , 32'hF09D5090 , 32'hE88F7A60 , 32'h0F4C9A10 , 32'h00933050 , 32'h0ECFF000 , 32'hFC1B1F78 , 32'hF18DA570 , 32'hE7C60720 , 32'h0F5F8920 , 32'hF2E755B0 , 32'h0BEC1070 , 32'hE772F7C0 , 32'hE3F8D1A0 , 32'hF7560860 , 32'hFB351710 , 32'h079320A0 , 32'h14A59F00 , 32'h0CBD5820 , 32'h12915660 , 32'hE9E26E60 , 32'h19D35620 , 32'h0D1073D0 , 32'h0CB611F0 , 32'hF7998F70 , 32'h06238848 , 32'hF8EC5248 , 32'h1639C5A0 , 32'h00CD58E0 , 32'h0D4BDAF0 , 32'h02BC77A0 , 32'hF04FCCC0 , 32'h0B69C280 , 32'h0AF552F0 , 32'h068E02D8 , 32'hFBBC5AE8 , 32'h10697940 , 32'h0AFA0EE0 , 32'h15F801A0 , 32'hF34A8A60 , 32'h015844D4 , 32'h0244EE28 , 32'h0264A38C , 32'h06264498 , 32'hFC6BE9B4 , 32'hF9BA6740 , 32'h0396D56C , 32'hF45E2AB0 , 32'hFD104738 , 32'h042F1158 , 32'hF7409550 , 32'h0373AC8C , 32'h07C3E570 , 32'h044CA990 , 32'h07B14448 , 32'hF79C96E0 , 32'h05174038 , 32'hFE11B9EC , 32'h08A66F30 , 32'h0060AA1B , 32'h04FA02B8 , 32'h073FC2B0 , 32'hFFAA2B95 , 32'h0739CA90 , 32'h02D8B134 , 32'hF6BBEE70 , 32'h0311651C , 32'hFEADF1B0 , 32'h03B3A7D4 , 32'hFFA39E3C , 32'h00066A17 , 32'h0002D506 , 32'hFFFA5937 , 32'hFFFF9925 , 32'h0001CAC4 , 32'hFFFAF1D3 , 32'h0000A12C , 32'hFFFFE277 , 32'hFFFFD3CA , 32'hFFFEF86E} , 
{32'h0002C357 , 32'h000501F2 , 32'h00011CD1 , 32'h000369C1 , 32'hFFFEA9CB , 32'hFFFA9BD2 , 32'h000052D4 , 32'h0005F3D6 , 32'h0005E6AB , 32'h00001E7E , 32'hFFFF8115 , 32'h00014080 , 32'h0000F932 , 32'h0003E8DD , 32'h0002252A , 32'hFFF86C00 , 32'h0002318E , 32'hFFFB470B , 32'hFFFB8558 , 32'h00037797 , 32'hFFFE5F49 , 32'h00001122 , 32'hFFF540EF , 32'h0006A300 , 32'hFFFD7932 , 32'hFFFF9EA3 , 32'h00034348 , 32'hFFF9DE66 , 32'hFFF703F1 , 32'hFFFDB2EF , 32'hFFFA9043 , 32'hFFFE234C , 32'hFFFB7A0C , 32'h000373B2 , 32'hFFFFA6E7 , 32'h00059800 , 32'hFFFF952D , 32'hFFF98F99 , 32'hFFF719DF , 32'hFFFF82B2 , 32'h00098C72 , 32'h0000DCBE , 32'h0002E3D2 , 32'h0004B672 , 32'h000295F6 , 32'h0004371E , 32'hFFFF9CD0 , 32'hFFFFB7D8 , 32'h0006B7A6 , 32'h000693CB , 32'hFFFA3D52 , 32'hFFFDE169 , 32'h00007B6E , 32'hFFFFDBAE , 32'hFFF9EC06 , 32'h000214A0 , 32'h00004855 , 32'hFFF92807 , 32'hFFFA0E94 , 32'h00065E4D , 32'h000297E9 , 32'hFFFED1A4 , 32'hFFF7B264 , 32'h000288EA , 32'h0005C256 , 32'hFFFE9C36 , 32'h0008313B , 32'h000505D4 , 32'hFFF993D3 , 32'hFFFAF149 , 32'hFFFA6194 , 32'h00015620 , 32'hFFFD912F , 32'h00030316 , 32'h00068B23 , 32'hFFFA3DD0 , 32'hFFFC06A8 , 32'h0005F7FE , 32'hFFFF7162 , 32'hFFFCEFDF , 32'hFFFCF048 , 32'h0003455D , 32'h0000ECEB , 32'hFFFFA2B3 , 32'hFFFFD099 , 32'hFFF96C40 , 32'h000052FF , 32'hFFFDBA96 , 32'hFFFFAF24 , 32'hFFFCE463 , 32'h0000A6D9 , 32'hFFFF4E1F , 32'h0003F327 , 32'h000277C5 , 32'h00025F8C , 32'hFFFEF21D , 32'hFFF95A04 , 32'h0001009C , 32'hFFFF3BD9 , 32'h00009262} , 
{32'h00017675 , 32'hFFFD1D10 , 32'hFFFF9268 , 32'h00018067 , 32'hFFFE5F3B , 32'h00024E2C , 32'h00044356 , 32'hFFFDADA3 , 32'hFFFDC74B , 32'h00030286 , 32'h00026983 , 32'hFFFBF821 , 32'hFFF8DDF8 , 32'h0001D99A , 32'h00063FF6 , 32'hFFFD474E , 32'hFFFC5420 , 32'hFFFE058C , 32'h0002EE27 , 32'hFFFD3326 , 32'hFFFD182F , 32'h000A8331 , 32'h0000446B , 32'hFFFB5DF3 , 32'h00090DE4 , 32'hFFF88003 , 32'hFFFA54A0 , 32'h00081A29 , 32'hFFFAC3C8 , 32'h000098C8 , 32'hFFFEDC76 , 32'hFFFE54EF , 32'h00023482 , 32'h0003B770 , 32'hFFFF527A , 32'h000105C9 , 32'hFFFE1625 , 32'h00013839 , 32'h000A5F09 , 32'hFFF7CB03 , 32'h0005A2D6 , 32'h000128F7 , 32'hFFFB95C9 , 32'hFFFEDA1A , 32'hFFFBEE2F , 32'h00006A47 , 32'hFFF82BC9 , 32'h00098E7E , 32'hFFFA8E1C , 32'hFFFD52EB , 32'h00022184 , 32'hFFFBD4F5 , 32'hFFFB0228 , 32'h00026E32 , 32'hFFF7F360 , 32'hFFF76DB1 , 32'h00024DA6 , 32'h000162B4 , 32'h0001CFF7 , 32'hFFF8AB98 , 32'h0007107A , 32'hFFFFAD6B , 32'hFFFF53AE , 32'h000095FB , 32'hFFFB7D9E , 32'h0002DECC , 32'h00089C6A , 32'h00028024 , 32'h000798BD , 32'h0007BA19 , 32'h0003E45C , 32'h000514BC , 32'hFFFE5965 , 32'hFFFAAAE7 , 32'h00048807 , 32'h0005BE24 , 32'hFFFD6C02 , 32'hFFFC2617 , 32'hFFFE9051 , 32'h0003D20A , 32'h00014A84 , 32'hFFFF8A0D , 32'h0006A0E2 , 32'hFFFFC640 , 32'h00001975 , 32'h00071CA9 , 32'h0005A27F , 32'hFFFC9B92 , 32'hFFFA1D97 , 32'hFFFD94A4 , 32'hFFFF20A4 , 32'hFFFE35AC , 32'hFFFF1FAB , 32'h00007D85 , 32'h00047275 , 32'h00050E34 , 32'h0002560A , 32'h00017A34 , 32'hFFFFC8CC , 32'hFFFC6746} , 
{32'hFFFFBBA1 , 32'hFFF75946 , 32'hFFFF6063 , 32'h0003F65B , 32'h00028EE0 , 32'h00013C87 , 32'h00006036 , 32'hFFF91669 , 32'hFFF896CF , 32'h000ACDDE , 32'h000BC7E5 , 32'h00019E3A , 32'h000052C4 , 32'h00046BB9 , 32'h0001FD35 , 32'hFFFF748D , 32'h00018147 , 32'h0004D99D , 32'h000174B2 , 32'h0007DD89 , 32'hFFFBFB55 , 32'hFFFC88A9 , 32'hFFFD4AF7 , 32'h00007DA6 , 32'hFFFF032D , 32'hFFFA418A , 32'h0000231E , 32'h0003EF46 , 32'hFFFAB41F , 32'hFFFD8DC8 , 32'hFFFDE3DF , 32'h0008152E , 32'hFFF97B8E , 32'hFFFD1E13 , 32'hFFFFD28B , 32'hFFFF9507 , 32'h0001D93C , 32'hFFFBF6FC , 32'hFFFACD35 , 32'h0001C8B3 , 32'h00026E78 , 32'hFFFE3E90 , 32'hFFFF850A , 32'hFFFA639A , 32'h000B4C4B , 32'h00001588 , 32'hFFFD7EBD , 32'h000108DE , 32'h000015A5 , 32'hFFFD92AE , 32'hFFFD020A , 32'hFFFD0299 , 32'h00039C83 , 32'h000291BA , 32'hFFF99523 , 32'h0001C67E , 32'hFFFF5CFF , 32'h0003FF1F , 32'hFFF92CFB , 32'h0001568A , 32'hFFFE729B , 32'h00043589 , 32'h0000A6A3 , 32'hFFFC20D8 , 32'hFFF7B56A , 32'h0004A38A , 32'hFFF7E944 , 32'hFFFAB02F , 32'h0005AAC9 , 32'h0004B9D9 , 32'h0007BEEB , 32'h00006121 , 32'h00043BDF , 32'hFFFA8EDA , 32'hFFF5A513 , 32'hFFF88BD1 , 32'hFFF78F2C , 32'h00013B58 , 32'h000360F8 , 32'hFFF67764 , 32'hFFFC2B10 , 32'h00048CD1 , 32'h0000A921 , 32'h00080316 , 32'hFFFDFA2B , 32'hFFFA5FCF , 32'h00076DC6 , 32'h00073D41 , 32'hFFFE8ECC , 32'h0000AB95 , 32'h0006518F , 32'h000218AB , 32'h000B58C9 , 32'h00024375 , 32'h000175BA , 32'h0003ABE5 , 32'h0004B371 , 32'hFFFE2E9B , 32'hFFFB44F0 , 32'h00064B1E} , 
{32'hE1EC8620 , 32'h02F4BBAC , 32'hD7C82500 , 32'hF84945E0 , 32'h17B91AE0 , 32'h02BD246C , 32'hEF1EE720 , 32'hFC962F28 , 32'hE9F417A0 , 32'h1C822F60 , 32'hF42435E0 , 32'h0192D7AC , 32'hF2030B40 , 32'hF7A7B4F0 , 32'hEF028DA0 , 32'h0DEFD580 , 32'hE758D240 , 32'hF5EE01F0 , 32'hF862FE08 , 32'h21101FC0 , 32'h03DC8770 , 32'hEA194E20 , 32'hFF76AA7C , 32'h116A1600 , 32'h1721D220 , 32'h016C4450 , 32'hEA9132A0 , 32'hF016D2A0 , 32'hEA331480 , 32'hEBCC3900 , 32'h082A4B00 , 32'h00209494 , 32'hFD2DC208 , 32'hFDD3A950 , 32'h0374F588 , 32'hF346ACB0 , 32'h0A3D4F70 , 32'hF78A9500 , 32'h082B2340 , 32'h0AC0D520 , 32'h0BDB7600 , 32'hEDFC1700 , 32'h04718A50 , 32'hFB0A4AD0 , 32'h06437F58 , 32'hEF9197E0 , 32'h18690E80 , 32'hF2F520F0 , 32'hF763F840 , 32'h10DE67A0 , 32'h0241C414 , 32'hDF01AF40 , 32'hFECD501C , 32'hFB2ECEB8 , 32'hF81D5F60 , 32'hF94BB5B8 , 32'hF7EDE910 , 32'hF524A840 , 32'hFB48FE10 , 32'hF7E2B8C0 , 32'hF75EE400 , 32'h08327620 , 32'hF8F97250 , 32'h05766150 , 32'hF2DFB7F0 , 32'h052955C8 , 32'hFD34FF20 , 32'hFB159F78 , 32'hF5C79A40 , 32'hF7AF9530 , 32'hF48183D0 , 32'hFFF45643 , 32'hFD9735D8 , 32'hFE29589C , 32'h01D69208 , 32'hF6883540 , 32'hFE5C6958 , 32'h11EFB540 , 32'hFBD8EE68 , 32'h0642B8E0 , 32'h03CB52D8 , 32'hF7EB16D0 , 32'hF2A4CBA0 , 32'hF9640B10 , 32'hFA8F7368 , 32'hFFD33BF0 , 32'h03D6A698 , 32'hFCB62358 , 32'hFE8FC1A4 , 32'hFFF9C274 , 32'hFFFC6915 , 32'hFFFEB38D , 32'hFFFF9641 , 32'h00018156 , 32'h00041F1B , 32'hFFFF2992 , 32'h00052299 , 32'h0000D830 , 32'h00091DBD , 32'h00015CA4} , 
{32'hBEC02700 , 32'h50A72300 , 32'hF098F0E0 , 32'hE2C0F160 , 32'h21D7DD80 , 32'hBEB63500 , 32'h4F77DA80 , 32'h4B7FFE00 , 32'hCDEC1C00 , 32'hFA5A7ED0 , 32'hD995B680 , 32'h2BEBC5C0 , 32'h28261840 , 32'hE6877F40 , 32'h07368D28 , 32'h292D8980 , 32'h2156D740 , 32'h1E81F4A0 , 32'h0F661860 , 32'hD7DA7B80 , 32'h17FFC4A0 , 32'h127F0EE0 , 32'h06D717A8 , 32'h31A18740 , 32'h0F0B7F40 , 32'hEFCABF60 , 32'h0F3CE0F0 , 32'hD9BF2BC0 , 32'h00E763CD , 32'hECDD8480 , 32'hDDADA240 , 32'hFE91FBF0 , 32'h0261019C , 32'hF9DD3870 , 32'h043029F8 , 32'h08E0EAC0 , 32'hF8726B30 , 32'h021C2F44 , 32'h06CDFB68 , 32'h14E044E0 , 32'h178DB500 , 32'h00D89C1F , 32'h0024DE3D , 32'hF04834D0 , 32'hEE26A120 , 32'hFFECDFAC , 32'h15FDD9C0 , 32'h105AB440 , 32'hF15C34E0 , 32'h0EE68660 , 32'hFA887900 , 32'h0CEFA990 , 32'hF618CB00 , 32'hFF4C780B , 32'hF8CB8690 , 32'hFD23C670 , 32'hF0DA6910 , 32'h03C95410 , 32'hFEE0C73C , 32'hFF1CB549 , 32'h0F42DF40 , 32'hE8E00A20 , 32'hF5837530 , 32'h17788700 , 32'hFBB3D058 , 32'h009EEA62 , 32'h04389D90 , 32'hFB35B3E0 , 32'hFFCA0AA2 , 32'hF588A100 , 32'h0135707C , 32'hFDD2B43C , 32'hEE848C00 , 32'hFA5886D8 , 32'h02118148 , 32'hF9AF9760 , 32'h047D1300 , 32'h01543974 , 32'h0099E335 , 32'hFD20486C , 32'hF968B100 , 32'hFF8CABB8 , 32'hF88A1040 , 32'hFE5A6ACC , 32'h012F7494 , 32'hF998F248 , 32'hFE0C392C , 32'h03FB4E4C , 32'hFFECC7E3 , 32'h00E162B3 , 32'h00014312 , 32'hFFFFA3BF , 32'h0002C8CB , 32'hFFFF22A6 , 32'hFFFFA26E , 32'hFFFD65F9 , 32'hFFFF8E89 , 32'hFFFD7797 , 32'h000048C7 , 32'h00018FF8} , 
{32'hE96A6DE0 , 32'h008EF0AC , 32'hEA523AC0 , 32'h1E939180 , 32'h0A49D040 , 32'h1EB13740 , 32'hFA4D7660 , 32'hFB868B90 , 32'hED13A860 , 32'h0C39EAA0 , 32'h01EA2F34 , 32'h0CAEE900 , 32'hF6C16550 , 32'hF1E76950 , 32'hE18707E0 , 32'h06A23B18 , 32'hE96C6B40 , 32'hF82A2098 , 32'h026B3F8C , 32'h042B30E0 , 32'hF67255F0 , 32'h0AE39A80 , 32'hFCB853BC , 32'hFB17D948 , 32'h0EB70100 , 32'h02F5C678 , 32'hEF458880 , 32'hFF8F82FE , 32'hF1F11960 , 32'hE0707400 , 32'h14394C80 , 32'h15D41E40 , 32'hFF4FE734 , 32'hFD4B8408 , 32'hF7C947E0 , 32'hFF305DFB , 32'h0C40B770 , 32'h0564CCF8 , 32'hFEC116F8 , 32'h0AB51B60 , 32'h002B4242 , 32'h07574458 , 32'h0C7E49C0 , 32'hFC9035F8 , 32'hFD688B94 , 32'hF5E3BED0 , 32'hFB487238 , 32'h04D87448 , 32'h02C11378 , 32'hFBF3B2E8 , 32'hF2081E60 , 32'hEA859C80 , 32'hF3E52570 , 32'hF15F1680 , 32'hF99397E8 , 32'hF1653830 , 32'hFBC9B6C8 , 32'h0EC37AF0 , 32'h03A814CC , 32'hFC22ED60 , 32'h04FA1F78 , 32'hFC493A50 , 32'hFB0AB5D0 , 32'hFD217B34 , 32'hFF2BB1C7 , 32'hFF257BE8 , 32'h05A266C0 , 32'h0C514910 , 32'h0617A7A8 , 32'hF5263510 , 32'hF927D920 , 32'h0406D568 , 32'hF4B02270 , 32'h00271624 , 32'h00F3D549 , 32'h052CF4E0 , 32'h004AFC04 , 32'h002B98B8 , 32'hF8AE2B10 , 32'hFBCE3658 , 32'h0BB3CF30 , 32'hFCC395BC , 32'hFE9AA5E8 , 32'hFCABDEDC , 32'h01C42C8C , 32'h02D0344C , 32'h05A3A980 , 32'hFC91261C , 32'h0196DBF8 , 32'hFFB91952 , 32'hFFFBE3A1 , 32'h00076358 , 32'h0003CEA0 , 32'h0002A2A2 , 32'h0000C649 , 32'h00017C80 , 32'hFFFC2B99 , 32'h0000314F , 32'hFFFB8688 , 32'h00004997} , 
{32'hF5503DF0 , 32'h0937D120 , 32'h02AC9368 , 32'h0E99F610 , 32'h03152E8C , 32'hFEB29014 , 32'hF723DD80 , 32'h0720FD98 , 32'hFBCED8E8 , 32'hF7A88260 , 32'hF2DD67C0 , 32'hFE06FC58 , 32'h08DD8E00 , 32'hF55028E0 , 32'h0235E2F4 , 32'hFFC7BF32 , 32'hF01658A0 , 32'h0A354F90 , 32'hFE880360 , 32'h0216671C , 32'hF6352A90 , 32'hF3E005E0 , 32'hFFDDBE3F , 32'h0C64A200 , 32'h033D6268 , 32'hFC2741A0 , 32'h0A00C560 , 32'hFA6C4E80 , 32'hF35849B0 , 32'h09E22FA0 , 32'hF0DAF920 , 32'hF01604C0 , 32'hFA3006F0 , 32'h00504C45 , 32'hF342A910 , 32'h04F99750 , 32'h09070320 , 32'h10630F60 , 32'h0958C1D0 , 32'h002EDEFB , 32'h07161440 , 32'h06712678 , 32'hFD877F88 , 32'h0591D8E8 , 32'hF3637340 , 32'h0599D070 , 32'hF8B40078 , 32'h053DFAF8 , 32'hFBDDED18 , 32'hFED7CCFC , 32'hFE9B9D40 , 32'h047C3248 , 32'hF67FACA0 , 32'h0501B688 , 32'h06EE4318 , 32'h07C6DDB0 , 32'hFF6A1D2F , 32'hFAEE7CA8 , 32'h054707E8 , 32'h0B056440 , 32'h0942B710 , 32'hF7B672B0 , 32'h06186AD8 , 32'hFEEE3508 , 32'hFC5A9D90 , 32'hFAF2F348 , 32'h03340448 , 32'h008561DA , 32'hFC9501E8 , 32'h00D7D8AB , 32'hF9E860C8 , 32'hFEB176A0 , 32'h04940CC0 , 32'hFFDC8BAE , 32'h03E44738 , 32'hFE358A10 , 32'h10869520 , 32'hFD98C218 , 32'hFE15F058 , 32'hFF1CB6F1 , 32'h0020B010 , 32'h04CE8148 , 32'hFF857E05 , 32'hF951FA88 , 32'hF9D6C8F8 , 32'h023CBD94 , 32'h0192B1FC , 32'hFE46F314 , 32'h02015DC0 , 32'h008E73BA , 32'hFFFBDC5E , 32'hFFF75588 , 32'h0001A30D , 32'hFFFEA137 , 32'h00030EC1 , 32'h000485EA , 32'h00013598 , 32'h00027704 , 32'h00086794 , 32'h00000064} , 
{32'h0D1E2090 , 32'hE2F9F6E0 , 32'h0A8AA280 , 32'hE217EA20 , 32'h10A06BE0 , 32'hE146DD20 , 32'hE9E04960 , 32'hD34808C0 , 32'hCC13D800 , 32'h1A47E9E0 , 32'h24CCA900 , 32'hF55E8780 , 32'hE31D4FE0 , 32'hE460ECE0 , 32'hEAFA3F60 , 32'hD8A1E580 , 32'hF97A7928 , 32'h1F85C520 , 32'hE229C3A0 , 32'hEE6C49E0 , 32'hFF17E006 , 32'h0C09B9C0 , 32'hF62DD150 , 32'hF8CFDA90 , 32'h0BFD4410 , 32'hEDE12D40 , 32'hF9460818 , 32'h0D036E50 , 32'hDB534280 , 32'hDFCAECC0 , 32'h007139EA , 32'hF1971330 , 32'hFB20F030 , 32'hF74587C0 , 32'h049D3C78 , 32'hF91A4E00 , 32'hE597B960 , 32'h1FE62140 , 32'hFC0ED354 , 32'hE8CF3740 , 32'h1848F2C0 , 32'h01FB0784 , 32'h20202040 , 32'hFFA2AC91 , 32'hEA2FA4C0 , 32'h05398620 , 32'h04D783F8 , 32'hFADBEC10 , 32'h0BF21990 , 32'h125EF700 , 32'h06B5E400 , 32'h07A01038 , 32'h13925AC0 , 32'h053BF3D8 , 32'hFAE98A78 , 32'h067AAA38 , 32'hDEF9D600 , 32'hF8C4A610 , 32'hF614B500 , 32'h0A9D16F0 , 32'h0485C340 , 32'hFEF14040 , 32'hE7B2E620 , 32'hFF3610C8 , 32'hFBBE72C0 , 32'hFDF55800 , 32'hF3180D10 , 32'hFFA08E05 , 32'h05FE3BC8 , 32'h08FFF290 , 32'hFBD314C8 , 32'h05F7B1B8 , 32'h12252CA0 , 32'hF8520CA0 , 32'hFB9C44B8 , 32'h055F1388 , 32'h026E9970 , 32'hFE21DF94 , 32'h00C9632C , 32'h06679150 , 32'hF9B13580 , 32'h09492AD0 , 32'h02021CA4 , 32'hF5124250 , 32'h017181C0 , 32'hFDF4529C , 32'hFEB3AA54 , 32'h024E0124 , 32'hFD965D20 , 32'hFE936AF0 , 32'hFFFE0A1A , 32'hFFFF77BF , 32'h0002E37F , 32'hFFFD1560 , 32'h00020A01 , 32'h00001302 , 32'hFFF89A3C , 32'hFFFDD78C , 32'h00010939 , 32'hFFFDE0C5} , 
{32'h18B194C0 , 32'h068FE8F8 , 32'hFDA7F628 , 32'h0C04BDE0 , 32'h1DA5B420 , 32'h09D8E740 , 32'hE3665980 , 32'h12236840 , 32'h36898B80 , 32'hE3376F80 , 32'h0ABFE280 , 32'hFF0091FC , 32'hF87397E0 , 32'hE887C7A0 , 32'h06046188 , 32'hDFA01580 , 32'h0A51FA30 , 32'h0E252060 , 32'h1BF6A7A0 , 32'hF70AC310 , 32'h15BFAF80 , 32'hFF049ACD , 32'hFF09C1CF , 32'h06449940 , 32'hF38E3840 , 32'hFCBFBDA0 , 32'h28C01200 , 32'h0F1ADC60 , 32'h06BC10B0 , 32'h09D1C020 , 32'hFA568548 , 32'h0B712E60 , 32'hF9A598A8 , 32'h090F2D40 , 32'hEAD7E040 , 32'h141F6A60 , 32'hFC45C9B8 , 32'hFBA14068 , 32'h16EBCA40 , 32'h0AD187E0 , 32'hEC3F6780 , 32'h26395E00 , 32'hF9456C98 , 32'h048E8EB8 , 32'hE97EE920 , 32'h105DDB60 , 32'h0D5BC890 , 32'h05F11250 , 32'hFBAC6450 , 32'hECE8E000 , 32'hFE587E10 , 32'h1134DF60 , 32'hF0FBAB80 , 32'h031CB5C4 , 32'hF07365C0 , 32'hFBB3D818 , 32'hF7022ED0 , 32'hED6DB1C0 , 32'hFF7C16B5 , 32'hFF0B6D61 , 32'h045CD8F8 , 32'h0641B9F8 , 32'h00EFBA1E , 32'hF5BBCF50 , 32'h0156470C , 32'h03488224 , 32'hF83A3800 , 32'hF344C990 , 32'hF9FF3930 , 32'hFF72B9A4 , 32'h0138913C , 32'hF5035940 , 32'hF8228650 , 32'h04FDADD8 , 32'h0646BB08 , 32'h04B0BD28 , 32'h09E9DFD0 , 32'h0A643470 , 32'hFEC1AD78 , 32'h0536A5B0 , 32'hF7693EB0 , 32'h01B14260 , 32'hFD161A7C , 32'hFFF0D7B1 , 32'hFB7FAFC0 , 32'hFE863200 , 32'hFF920088 , 32'hF734CC90 , 32'hFEFBFE68 , 32'h007881C5 , 32'h0001C7BA , 32'hFFFD7226 , 32'h0000D149 , 32'h0005CA73 , 32'h00029B27 , 32'hFFFCC953 , 32'h00047CFA , 32'h00031917 , 32'hFFFF67F9 , 32'h00055DB2} , 
{32'hFFFB7877 , 32'h0004239F , 32'hFFFCC809 , 32'hFFF9B754 , 32'h0008619C , 32'h000E7CA9 , 32'hFFFB9033 , 32'hFFFB42E4 , 32'hFFFEAFAC , 32'hFFFC4DFB , 32'hFFFF4B69 , 32'hFFF35C95 , 32'hFFFFF921 , 32'hFFFF3298 , 32'h0006E90B , 32'h0000FB9D , 32'h0002ACE3 , 32'hFFFB0A81 , 32'h00048B78 , 32'hFFFADCE2 , 32'h0000C0BC , 32'hFFF8CBE7 , 32'h000C2A2C , 32'h0001FB73 , 32'hFFFFC515 , 32'h00013DAF , 32'hFFFE37F2 , 32'h0007DB6B , 32'h000C640B , 32'hFFFDD24B , 32'h00024386 , 32'hFFFE46F4 , 32'hFFFAAB66 , 32'hFFFA8172 , 32'h0008BE0F , 32'h0003CC65 , 32'hFFF8E6B6 , 32'h000D78F5 , 32'h0004F35E , 32'hFFFC64BA , 32'hFFF9C6AE , 32'h0000E792 , 32'h00083CF0 , 32'h00056003 , 32'hFFF7B382 , 32'hFFF8C872 , 32'h0003086C , 32'hFFF45366 , 32'h00054E3F , 32'hFFFF0D58 , 32'h00076C68 , 32'h0001E71E , 32'h0002313B , 32'hFFFE0C3C , 32'hFFFFD1F4 , 32'h000144D0 , 32'hFFF84A61 , 32'h0001409C , 32'hFFFFA208 , 32'h0004DE10 , 32'h0005626A , 32'hFFFF5E72 , 32'hFFFFA1A3 , 32'h00003F54 , 32'h00010644 , 32'hFFF8CDE9 , 32'h0006737F , 32'h0000BC52 , 32'h00048835 , 32'h000238DE , 32'h00006E76 , 32'hFFFE7D96 , 32'hFFFB74EE , 32'h00039BB1 , 32'hFFFF1C5A , 32'hFFFDA8A8 , 32'hFFF123F5 , 32'h00033FFD , 32'h000297DA , 32'h000800D0 , 32'hFFFB3714 , 32'h0006CC39 , 32'hFFFF773E , 32'hFFF97507 , 32'h0008A935 , 32'h000096C5 , 32'hFFF79CA2 , 32'h0004DB44 , 32'hFFFF64D1 , 32'h0008FEBF , 32'hFFFFB2DC , 32'h0008E462 , 32'h00076117 , 32'hFFF3B0E2 , 32'hFFFF6BBF , 32'hFFFD7841 , 32'hFFFB782F , 32'h0004E00A , 32'h000BFABA , 32'h000556CF} , 
{32'h1A202020 , 32'h587E7580 , 32'h2F1CBB00 , 32'h2302D400 , 32'h56C9A480 , 32'hEC851BE0 , 32'h0EF24710 , 32'h1A700960 , 32'hFAB2F738 , 32'h2CE20780 , 32'hC428D340 , 32'h153C3060 , 32'h119C4E40 , 32'hFA5F5C10 , 32'h0F9BEFC0 , 32'h2D6E6880 , 32'h0E349800 , 32'hFC4EF4E0 , 32'hE06C8A00 , 32'h01489E28 , 32'h10345100 , 32'h20551D40 , 32'h04E5B7C0 , 32'hDA70E940 , 32'h014002F4 , 32'h151D11C0 , 32'hF6534B70 , 32'h11314F20 , 32'hEE4C8C60 , 32'h06D0CAB8 , 32'hFCB94034 , 32'h0471ED38 , 32'hF66BDEB0 , 32'hF5B7C160 , 32'hE0E5A9C0 , 32'h042B0EB8 , 32'h139BF3E0 , 32'hE1144740 , 32'hFCF90D0C , 32'hEE63DE60 , 32'hF6F97A00 , 32'h07BCA6E8 , 32'h060A0FA0 , 32'hFA3738A0 , 32'h136FF840 , 32'h03BB9368 , 32'h064E2AB0 , 32'hF94D8100 , 32'hF1BB67B0 , 32'hF98F7648 , 32'h05A0D148 , 32'hFED86E2C , 32'hF96E3C78 , 32'h040F7668 , 32'hF9A8B868 , 32'h0D2DDEA0 , 32'hED8C3FC0 , 32'hFB05CC08 , 32'hF9D36698 , 32'hDF0AC540 , 32'h01ECA7EC , 32'h0AAB9D90 , 32'h04700B50 , 32'h0550AA88 , 32'h09420DA0 , 32'h05996200 , 32'hFD9CC714 , 32'hFFF45F19 , 32'h06931850 , 32'h10237680 , 32'hEEA38B00 , 32'hEFCA9420 , 32'h0073EC22 , 32'hECA843E0 , 32'h0487EEB0 , 32'h0D0434B0 , 32'h04B45670 , 32'h035C29F8 , 32'h01AC7EC4 , 32'h0673BB88 , 32'hFD152294 , 32'hF8B8DDB8 , 32'h06514A80 , 32'hFE6D2D80 , 32'h00ED1429 , 32'hFD77D784 , 32'h07560830 , 32'hFEAA9410 , 32'hFEC533E4 , 32'hFF9AF077 , 32'hFFFB3CC0 , 32'hFFFE0718 , 32'h0000C117 , 32'hFFFB7FC3 , 32'hFFFE4D9F , 32'h0002F1A8 , 32'hFFFE13C4 , 32'h00007EB6 , 32'hFFFEB874 , 32'h00004928} , 
{32'hF30299D0 , 32'hFEA59150 , 32'h21D1F940 , 32'hBB89B980 , 32'hD2512E80 , 32'hCE100240 , 32'hEB957C40 , 32'h04FBF798 , 32'h526C2980 , 32'h0C075590 , 32'hF9E2CD58 , 32'hFFF2D819 , 32'h0F347550 , 32'h106DF5C0 , 32'h079DA910 , 32'hF0C7F060 , 32'hFE0A9AC0 , 32'h3921FF80 , 32'h0ECD9180 , 32'h1BD335C0 , 32'hD4246E00 , 32'hF91F3A40 , 32'hFD5B72FC , 32'hEDEAE320 , 32'h0E5049E0 , 32'hF5DCD180 , 32'h0572F038 , 32'h100015C0 , 32'hF566B6D0 , 32'hEFD44240 , 32'h1CCA7C20 , 32'hEB0E1BC0 , 32'hDCFDBDC0 , 32'hDF150240 , 32'h07604AF8 , 32'hF86A0830 , 32'hF1D38650 , 32'hF6651410 , 32'hF6BBEFE0 , 32'h04DB62A0 , 32'h083F3900 , 32'h0AF4B560 , 32'hE3DA1540 , 32'h13EE9BE0 , 32'h0A57EF50 , 32'hF9E0D530 , 32'hEDB4CE20 , 32'h0026131D , 32'hFE2795E0 , 32'hF66564A0 , 32'h068251F0 , 32'hF0CFCF90 , 32'h07E5B050 , 32'hFA4058A8 , 32'h093E1B40 , 32'hEC12C440 , 32'h07E90B00 , 32'hFCE5CADC , 32'h076D6718 , 32'hF5BE0540 , 32'hF3323B00 , 32'hF9EFB7A0 , 32'h04822DD8 , 32'h18D153C0 , 32'h065A0F28 , 32'h00F2B9BC , 32'h03A79540 , 32'h01AB2E48 , 32'h08F594C0 , 32'hFE40FEC4 , 32'hF5870B80 , 32'h0F68D450 , 32'hF5160320 , 32'hFBFC4190 , 32'h0757B3A0 , 32'h00D97DE1 , 32'h022BA0DC , 32'hFFDD034C , 32'hFF6291F9 , 32'hFA4E36C0 , 32'hF6C4F910 , 32'hFE177C14 , 32'hF93423C0 , 32'hFC3E8418 , 32'h0206BE90 , 32'h060636A8 , 32'hFC3D2FAC , 32'h0A602690 , 32'h044B97C0 , 32'h004FFE7A , 32'hFFFE2825 , 32'hFFFBC46B , 32'hFFFF49BB , 32'hFFFEB145 , 32'hFFFF0FA8 , 32'h000019BC , 32'h00034CAE , 32'h00034352 , 32'h00008B63 , 32'h0004046A} , 
{32'h0003EFE6 , 32'h00019513 , 32'hFFFC19D0 , 32'h0006382C , 32'h0009DF38 , 32'h0004944B , 32'hFFFF7BE1 , 32'hFFFACDE3 , 32'hFFFD758C , 32'h00028D64 , 32'h00005E22 , 32'hFFFB309C , 32'hFFFDD5EE , 32'h00030B40 , 32'h000AE507 , 32'h00079983 , 32'h00033B82 , 32'hFFFF09CE , 32'h0003AB6B , 32'hFFFF3468 , 32'h00045B61 , 32'hFFFCF4B3 , 32'h00013613 , 32'hFFF71B94 , 32'hFFFC2CE9 , 32'h0007CCE5 , 32'h000065E8 , 32'h00065FE6 , 32'h0002E2F7 , 32'h0004EE6D , 32'hFFFD6840 , 32'hFFFB83D6 , 32'hFFFD0EC2 , 32'h000157EA , 32'hFFFB73A5 , 32'hFFFE76E7 , 32'hFFFDA91B , 32'hFFFF7A90 , 32'h0002DE23 , 32'h00015432 , 32'h00000FC8 , 32'hFFFC09F8 , 32'h00002B87 , 32'hFFFD79A3 , 32'h0002EC8F , 32'hFFF9612F , 32'h00052913 , 32'h0003BA18 , 32'hFFFEDE3B , 32'h0000B248 , 32'hFFFFBD90 , 32'hFFFF751B , 32'h0003C422 , 32'hFFFCC0DA , 32'h0001D639 , 32'h00034FF7 , 32'hFFF8CA05 , 32'hFFFFDB2D , 32'hFFFC5B9C , 32'hFFFF0252 , 32'h0003F7E9 , 32'h0002CD2B , 32'h0000BCFB , 32'hFFFA7592 , 32'h0000F7DC , 32'h00078777 , 32'h00062CFF , 32'hFFF2950A , 32'hFFFE779D , 32'hFFFAA362 , 32'hFFFA4344 , 32'hFFFEF830 , 32'hFFFE1A8D , 32'h0000CF8A , 32'h00061D38 , 32'hFFF83316 , 32'h000091DA , 32'h000285B3 , 32'h00030C79 , 32'hFFEFDAF1 , 32'hFFFFF163 , 32'hFFFAC00B , 32'hFFFEB1D2 , 32'h000213A7 , 32'h0001C68B , 32'hFFFF6531 , 32'h0008482C , 32'hFFF7A425 , 32'hFFF7AE9D , 32'h000D4337 , 32'hFFFC7A1C , 32'h0000389F , 32'h00020E67 , 32'h0004ADDA , 32'h0001B4E1 , 32'h00021BC6 , 32'h0005784F , 32'hFFFFA6F1 , 32'h0003AF56 , 32'hFFFEDCCC} , 
{32'h7FFFFFFF , 32'h37D91680 , 32'h4149AB00 , 32'hE22A4460 , 32'h09E379D0 , 32'h36910F80 , 32'hC2980900 , 32'h1AE13E80 , 32'hDAB36B80 , 32'h23AAD480 , 32'hD388BA00 , 32'hF93DC350 , 32'hE8045020 , 32'h02F08928 , 32'h14FFA740 , 32'h1C4DA320 , 32'hFFF03B9D , 32'h06A85CF8 , 32'hFDCFC6E0 , 32'hF64B36F0 , 32'h1009CFE0 , 32'hEB8E15A0 , 32'h07D2EF78 , 32'h18597A80 , 32'h07688470 , 32'h069543E8 , 32'hF48B4B30 , 32'hECBF4980 , 32'hFC5DDF30 , 32'h1F42D3C0 , 32'hF934F5A0 , 32'h30C760C0 , 32'hEFAFC600 , 32'h16E9C1A0 , 32'hFFB1CBD1 , 32'hD55817C0 , 32'hF9D944B8 , 32'hEB1B77E0 , 32'h1ADF3360 , 32'hFA2B3718 , 32'h1621F580 , 32'hD1B55F00 , 32'h04B44BC0 , 32'h11A1F900 , 32'h00DA8128 , 32'h053A5310 , 32'hF548DC40 , 32'hF7D49BC0 , 32'hEF8F4B40 , 32'h06F1F4D0 , 32'hE7E90F40 , 32'h0122D124 , 32'hF9928770 , 32'h00CA1C97 , 32'hF848C8B8 , 32'hF5BE0A30 , 32'h07A210C0 , 32'h0124C780 , 32'h0D885780 , 32'h0F31FCE0 , 32'hFF4BC765 , 32'h0472D908 , 32'h0645F4D0 , 32'h02581584 , 32'h0B7ACCF0 , 32'hF69E1050 , 32'hF89DF970 , 32'h09634C00 , 32'hFB8C6AE8 , 32'h0E7C9FB0 , 32'h09090ED0 , 32'hFF50C5C4 , 32'hFD9E7858 , 32'h0474E108 , 32'hFB8838F8 , 32'hFBE62DE0 , 32'h0A6061E0 , 32'h0B1A37A0 , 32'h007E69CD , 32'h0231F92C , 32'h03E78510 , 32'h05680B80 , 32'h003C682E , 32'hFE88CF18 , 32'h02C2EF68 , 32'h01988604 , 32'hFB2E9D18 , 32'hFD026E38 , 32'hFE3D2A40 , 32'hFFF9280F , 32'hFFFF5966 , 32'hFFFF903B , 32'h00048A62 , 32'hFFFE3C92 , 32'hFFFFD4F3 , 32'hFFFF20CB , 32'hFFFDA331 , 32'h00026F0A , 32'hFFFFCD08 , 32'hFFFFB85F} , 
{32'hFFFBB72B , 32'h00007C98 , 32'h0001655A , 32'hFFFE88DF , 32'h0003082E , 32'h0002CE0F , 32'hFFFD8EA2 , 32'hFFF869CB , 32'h000065A0 , 32'h0004B25A , 32'hFFFDBA57 , 32'hFFFC2167 , 32'h00010C58 , 32'h0005012D , 32'hFFFFCC77 , 32'h0008D049 , 32'h00031E02 , 32'h00035032 , 32'hFFFF91DE , 32'hFFFB582A , 32'h0004EA76 , 32'h00037F57 , 32'h00009EB6 , 32'h00097F56 , 32'hFFFCF6D1 , 32'h0003A868 , 32'h000143CD , 32'h00018355 , 32'hFFFFD83D , 32'h0006AE42 , 32'h0002A56C , 32'h0005FE6F , 32'h00032849 , 32'h0000E696 , 32'h0004C923 , 32'h00036F0C , 32'hFFF879CE , 32'hFFFAD616 , 32'h00003621 , 32'h0009466C , 32'h0001035A , 32'hFFFBE855 , 32'h0007F36F , 32'h00045743 , 32'hFFFE7AB3 , 32'h00057918 , 32'hFFFAEEA9 , 32'h0005CCD4 , 32'hFFFD608F , 32'h00038606 , 32'hFFF6B56D , 32'hFFFF5FE0 , 32'h0002627F , 32'h0002E2F8 , 32'hFFFECEA9 , 32'h0004907C , 32'h0000F9D3 , 32'h000A1A72 , 32'hFFFE5080 , 32'hFFFEC953 , 32'h0000555D , 32'hFFF96315 , 32'h0003D0F5 , 32'h00007D60 , 32'h00009212 , 32'h00026F54 , 32'h00067E72 , 32'hFFF8B16E , 32'hFFF9902B , 32'h00062A11 , 32'hFFFABE38 , 32'hFFFA8844 , 32'h00087A6B , 32'h00036C0A , 32'h0003D265 , 32'h00014739 , 32'h00031E44 , 32'h0003EC8C , 32'h0000AAE4 , 32'hFFF81044 , 32'h00044C6E , 32'h0002A0C2 , 32'hFFFA1644 , 32'hFFFC53B7 , 32'h00073A54 , 32'hFFFFC3FE , 32'hFFF97331 , 32'h0005C0D2 , 32'h0006DF41 , 32'h0003EA96 , 32'hFFFF7E13 , 32'h0005D5AF , 32'hFFFF7A13 , 32'hFFFC6977 , 32'hFFF9F288 , 32'hFFFF9B5A , 32'hFFFD8A51 , 32'h00067854 , 32'hFFFC0BCA , 32'hFFFDF482} , 
{32'h23AB0340 , 32'hE3524660 , 32'hD878B240 , 32'hB746B700 , 32'hF12768A0 , 32'hD05E1200 , 32'h119F3600 , 32'hF5BD3FF0 , 32'hEB84F620 , 32'h0D4693A0 , 32'h1459ACE0 , 32'h1EC17B80 , 32'hFFA237F3 , 32'hCF6C8000 , 32'h08FE8D10 , 32'h308F7A40 , 32'h048C0F48 , 32'hFE443FAC , 32'hFF336C31 , 32'hF8C415F0 , 32'hEA5F1620 , 32'h0CAB4740 , 32'hE8ACDCC0 , 32'h023E14BC , 32'hFDAA4078 , 32'h252BB580 , 32'hEA7A4120 , 32'hFC3285EC , 32'hE0192520 , 32'h0D24CE90 , 32'h11FBC6C0 , 32'hF9239D38 , 32'hFE6BDF5C , 32'h10A7A460 , 32'h1D7FE660 , 32'h01C61574 , 32'h15E9B0C0 , 32'hF48ED920 , 32'hEB6A15E0 , 32'h0A401F00 , 32'hF84A19F8 , 32'h17B2AB20 , 32'hF37BB8E0 , 32'h0C3EDD20 , 32'hFADAAAE8 , 32'h06C81090 , 32'hF33A95F0 , 32'hF29AE570 , 32'hEF9BDBA0 , 32'hEE7E8080 , 32'hF87A4258 , 32'h04B9D7A0 , 32'h0121C050 , 32'hF89E6B60 , 32'hF0C4E150 , 32'h0A714100 , 32'h04B50BD8 , 32'hFEAEB4B4 , 32'h104B79E0 , 32'hEF87DD00 , 32'h00378193 , 32'hFA62BFB8 , 32'h06E24CA0 , 32'hEB27B8C0 , 32'hEA2C5500 , 32'hFC1C9934 , 32'hFA2A1D40 , 32'h04EDAA30 , 32'hFCA50B88 , 32'hFFD67BB9 , 32'hFF002E88 , 32'hFFDC93F8 , 32'hF31606B0 , 32'h03A77AB4 , 32'hFC53AD44 , 32'h03608120 , 32'h00F29FF5 , 32'hFE8469C4 , 32'h0E6E73E0 , 32'h06E990A0 , 32'h00BC9352 , 32'h046CA850 , 32'h02325EA0 , 32'hF90FF280 , 32'hF8DF14F0 , 32'h01018970 , 32'h00EFC32A , 32'h04166520 , 32'h0267A144 , 32'hFFB88ECA , 32'hFFFF6874 , 32'h000168C9 , 32'hFFFC4B92 , 32'h0004EE43 , 32'h00017986 , 32'hFFFCC56C , 32'hFFFD2187 , 32'h0002EA5C , 32'hFFFF01B8 , 32'h00028093} , 
{32'h38BC6240 , 32'hB7AE3700 , 32'h060D48A8 , 32'h30C50640 , 32'hC193DA80 , 32'h53070700 , 32'h485ABA00 , 32'h099C3F50 , 32'hDD571080 , 32'hD0144F80 , 32'h1C2CD400 , 32'h2197BE00 , 32'hFFE52F7D , 32'h2E7B6740 , 32'hC4321380 , 32'h1E721820 , 32'h1658B300 , 32'h3BE98300 , 32'h10853020 , 32'hD0C133C0 , 32'hFE9537A4 , 32'hFEAE77C4 , 32'h12CFD740 , 32'hDC6D4500 , 32'hEC713FC0 , 32'h0EF74450 , 32'hEBFCA0E0 , 32'hDE765400 , 32'hFA58E540 , 32'hE2AE64C0 , 32'hFA486620 , 32'hE3B82420 , 32'hE7CC63C0 , 32'h001DC36E , 32'hF3E27630 , 32'hFF5A50C1 , 32'h08D492F0 , 32'hEE4A5F60 , 32'h06FA1170 , 32'h10A3A560 , 32'hEEC64FE0 , 32'hF002ADE0 , 32'h112084E0 , 32'h0C256F80 , 32'h2F2AF280 , 32'h018396D4 , 32'h00E0D6AB , 32'h07248C88 , 32'hF4852A50 , 32'hFD328B70 , 32'h06266A10 , 32'hF7545FE0 , 32'hFE319E80 , 32'hF4D77100 , 32'h01FC8EC8 , 32'h06B2F488 , 32'hF6022E20 , 32'hF18ED660 , 32'hFD26B290 , 32'hF9FB3A38 , 32'h08154400 , 32'hFBC1F9B0 , 32'hF24120D0 , 32'hF98AE690 , 32'h0D45CB70 , 32'hF63FF660 , 32'hFD240204 , 32'hF84D8898 , 32'h04B0BBF0 , 32'hFA4B84C8 , 32'h0D947C50 , 32'h081A87F0 , 32'hFF884287 , 32'h00C3D9EB , 32'h00764A85 , 32'hFDCEA204 , 32'h0556A9F0 , 32'h00E8C278 , 32'h03B78388 , 32'hFAAAC920 , 32'hF97042E8 , 32'hFC04E694 , 32'hFF6B55F6 , 32'hFD81A854 , 32'h0176FE78 , 32'h009D3FDC , 32'h04147B18 , 32'hFDFDF65C , 32'h030E3338 , 32'hFEE4E06C , 32'hFFFDD2AD , 32'h0003841D , 32'h00017683 , 32'h0002C38E , 32'hFFFF92A7 , 32'h0000CF8E , 32'h0001E137 , 32'h0003DE6B , 32'h0007F388 , 32'hFFFF6AC9} , 
{32'h0003C905 , 32'hFFFA7AF4 , 32'hFFFEB3BD , 32'hFFFF0BCC , 32'hFFFECFF1 , 32'h0000DFF1 , 32'hFFFAB353 , 32'hFFF8E7F0 , 32'hFFF9CA7C , 32'h000BB0F1 , 32'hFFF7790E , 32'h0002F206 , 32'h00050362 , 32'hFFFD3098 , 32'h000B7F08 , 32'h0000DAC6 , 32'h0000E4CD , 32'h0000C26A , 32'h0008C3D0 , 32'h00015C4D , 32'h000115C9 , 32'hFFF79B68 , 32'h0003946F , 32'h00085DC7 , 32'hFFFF6F3D , 32'hFFFDB652 , 32'hFFFFB11F , 32'hFFFE7B89 , 32'h000290A2 , 32'h00074264 , 32'hFFFFFF2C , 32'hFFF55D59 , 32'hFFFFFE9A , 32'hFFFC7A47 , 32'h00028A14 , 32'hFFFC9C9A , 32'h0002C2A6 , 32'h0001F3B7 , 32'h0001A20A , 32'h0004C9FA , 32'h000051C2 , 32'hFFFB73DE , 32'hFFF9324D , 32'hFFFB8FF9 , 32'h00056792 , 32'hFFF76D87 , 32'h000024BF , 32'hFFFFFFD9 , 32'h00065BF2 , 32'h0003465D , 32'h0005849F , 32'h000118D9 , 32'hFFF881EE , 32'h0005E1B5 , 32'hFFFB4AB4 , 32'hFFFCC7FF , 32'h00066168 , 32'h0002C366 , 32'hFFFF0FD1 , 32'h00020597 , 32'h00034D01 , 32'hFFFDAF97 , 32'h00024A80 , 32'hFFFE63C4 , 32'h00028100 , 32'h0001C4A2 , 32'h0001E5FD , 32'h0001E285 , 32'hFFFC9B15 , 32'hFFFC8EB2 , 32'h0004F8B9 , 32'h000248BA , 32'hFFFC9BFC , 32'h0003098E , 32'h000917EA , 32'h000206BA , 32'h000169E9 , 32'hFFF62C4A , 32'hFFFFD054 , 32'hFFFF12FB , 32'hFFF7E57D , 32'h0001C97F , 32'h00014280 , 32'h00028F0C , 32'hFFFF97DC , 32'hFFFCBC93 , 32'h0005D1E6 , 32'h00050A1E , 32'h0005B993 , 32'h0001D4D2 , 32'h0003BE88 , 32'h00022CA9 , 32'h0002663C , 32'h00041263 , 32'h00049277 , 32'h0003A536 , 32'hFFFC4CFB , 32'h00000B3D , 32'h00017406 , 32'hFFFFEAF0} , 
{32'hFFF6F364 , 32'h0000BF19 , 32'hFFFE71CE , 32'hFFFC48E9 , 32'h0002CBCB , 32'hFFFF54B0 , 32'h000024B7 , 32'h000432AA , 32'hFFF9AFE2 , 32'h00017B0A , 32'hFFFDD0CE , 32'h00001891 , 32'h0002F3FB , 32'hFFFD121F , 32'h0006B124 , 32'hFFFCE40E , 32'h000695A2 , 32'hFFFE156D , 32'h0003A53C , 32'hFFFAB811 , 32'h00050E3B , 32'h0005CA1F , 32'hFFFAFE16 , 32'h000228D9 , 32'h0001ED93 , 32'hFFF969EF , 32'hFFFDE370 , 32'hFFFA0A06 , 32'hFFFF4AA4 , 32'h0001CDE7 , 32'hFFFA92FD , 32'hFFF80DF7 , 32'h0000F5AC , 32'hFFFA1379 , 32'h000156CB , 32'hFFFEF5F1 , 32'h00036BEF , 32'hFFFB2BEA , 32'hFFFFFB36 , 32'hFFFE7654 , 32'h0007B8A8 , 32'hFFFAAFFE , 32'h000152A3 , 32'hFFFDC3B7 , 32'hFFFBE647 , 32'hFFFDF813 , 32'h0000A42B , 32'hFFF967EC , 32'h00076C0B , 32'hFFFC8D7D , 32'hFFF901D3 , 32'hFFFEF48C , 32'h00064FA8 , 32'h0006E3A2 , 32'h00014DA2 , 32'h00005253 , 32'h00069430 , 32'h000518DA , 32'hFFF8C0E7 , 32'h00025762 , 32'hFFF85184 , 32'hFFFDB85F , 32'hFFFF4065 , 32'h000119BD , 32'h0004D115 , 32'h00065E63 , 32'h0006D712 , 32'h0004BA46 , 32'hFFF8A0BA , 32'h00018FC7 , 32'h00082282 , 32'h00034DE5 , 32'h0000087C , 32'h00030121 , 32'hFFF90439 , 32'h0008F76B , 32'h00017935 , 32'h00055D9F , 32'h00020632 , 32'hFFFDD6D4 , 32'h00076BB7 , 32'hFFFC7C1D , 32'h00039033 , 32'hFFFF8EF0 , 32'hFFFBFB8A , 32'h00074741 , 32'hFFFAEB37 , 32'h0005F53F , 32'h000497F0 , 32'h0001A75E , 32'hFFFA4F7E , 32'hFFFDBB69 , 32'h000353E4 , 32'h0000DD68 , 32'h0004AC19 , 32'h0003C303 , 32'h0003BAE6 , 32'h000257B7 , 32'h00057C8E , 32'h000583F2} , 
{32'hFFFB86B9 , 32'h00018620 , 32'h000020F1 , 32'hFFFA57BD , 32'hFFFF53B9 , 32'h00049CC8 , 32'hFFFAC6FC , 32'h00084A05 , 32'hFFFF3CF4 , 32'h00007E60 , 32'h0001DAEA , 32'h000166FC , 32'h000621C5 , 32'h00074D62 , 32'h0002B86D , 32'h000342E3 , 32'hFFFFF13D , 32'h0000E999 , 32'h000471E6 , 32'hFFFE330B , 32'hFFFA9271 , 32'hFFFBB375 , 32'hFFFE7E1F , 32'hFFFF3546 , 32'hFFFC2F69 , 32'h00021FFB , 32'h0001FC47 , 32'h0002FDA9 , 32'h0000EC48 , 32'hFFFD46DF , 32'h00008AA8 , 32'hFFFC53DC , 32'h0008CAA8 , 32'hFFF639C0 , 32'hFFFF217B , 32'h0008F524 , 32'hFFFE4A53 , 32'h00042EA6 , 32'hFFFA6802 , 32'h000232EA , 32'h0006B05C , 32'hFFFF05BD , 32'hFFFE1C86 , 32'hFFFBE93B , 32'h00055508 , 32'h0004DE91 , 32'h0002473F , 32'hFFFF304E , 32'hFFFECF35 , 32'hFFFF9399 , 32'hFFFEE20E , 32'h0003F862 , 32'hFFFCBFD6 , 32'h0001F35A , 32'h00052CE7 , 32'h00008760 , 32'h000632EC , 32'h0000CF91 , 32'h0003E79D , 32'h000329D7 , 32'hFFF6E139 , 32'h0006AF38 , 32'h000219D6 , 32'h0002CF3A , 32'hFFF99F9D , 32'h000843D2 , 32'hFFFE7C0D , 32'h00009C8C , 32'h000123B9 , 32'h000514F5 , 32'hFFFE0F4F , 32'hFFFCC9E9 , 32'h0002C58A , 32'hFFFCFC26 , 32'hFFF55981 , 32'hFFFF4D29 , 32'h0000C54F , 32'h0000254E , 32'h0002E568 , 32'h00012531 , 32'hFFFFD455 , 32'hFFF9790B , 32'hFFFCFADE , 32'h00069009 , 32'hFFFEDBA1 , 32'h0007909C , 32'hFFF68104 , 32'hFFFDB087 , 32'h0003800B , 32'hFFFFE8F4 , 32'hFFFD3953 , 32'h0001DCAD , 32'hFFFED58B , 32'hFFFDF869 , 32'hFFFDE4D9 , 32'hFFEF317B , 32'h00058EF1 , 32'hFFFBEB1F , 32'hFFFC6E22 , 32'hFFFDAE09} , 
{32'hFFF86B19 , 32'hFFFF12AB , 32'h000048E1 , 32'h00001CD1 , 32'hFFFAEF17 , 32'h000404F3 , 32'hFFFED601 , 32'h0002F2CD , 32'hFFFD9BBB , 32'hFFFCCD9B , 32'h00004A6C , 32'h00016C5A , 32'h00061333 , 32'h00011345 , 32'hFFFF4FA5 , 32'hFFFFF989 , 32'hFFF72485 , 32'h000557D8 , 32'h000285F6 , 32'h0006BA51 , 32'hFFFC8AED , 32'hFFFCE00D , 32'hFFFB3AEA , 32'h000138C9 , 32'hFFFFA57D , 32'hFFFDB601 , 32'hFFFCB8A2 , 32'hFFFC2E74 , 32'hFFFCCD19 , 32'h0004C84A , 32'h00044055 , 32'hFFFC3DDD , 32'hFFFE2A3C , 32'h000B7B50 , 32'h000248C6 , 32'h00002FAC , 32'hFFFC9CAD , 32'hFFFD3C3F , 32'hFFF6229C , 32'hFFFFC9BF , 32'h00018B8D , 32'h00064D5C , 32'h00023955 , 32'h00045997 , 32'h0001075D , 32'h0009A693 , 32'hFFFB29E5 , 32'hFFFD6649 , 32'h0005FC43 , 32'h00020F94 , 32'hFFFB9E2D , 32'hFFFA5C77 , 32'hFFFC11C8 , 32'hFFFE9E71 , 32'hFFF5CB65 , 32'h0000A104 , 32'hFFFD08D7 , 32'h000C2040 , 32'hFFF9664D , 32'hFFFE4FED , 32'hFFF27DE4 , 32'h00006C8A , 32'hFFFBD1BE , 32'hFFFBBAC2 , 32'h000077AA , 32'hFFFD57DD , 32'h0004ECF1 , 32'hFFFA5038 , 32'hFFFF51D2 , 32'hFFF921AF , 32'hFFF8830F , 32'hFFFB8D85 , 32'h000511A3 , 32'h00046608 , 32'h00069D11 , 32'hFFFFF07B , 32'hFFF974C1 , 32'hFFFECE44 , 32'hFFFA3C92 , 32'h00022492 , 32'h00096042 , 32'hFFFA91C7 , 32'hFFFBA336 , 32'hFFFF7C84 , 32'hFFF171F2 , 32'h0004467A , 32'h00009ED8 , 32'h0007C116 , 32'h0002BE1B , 32'h000332CA , 32'hFFFD4CD0 , 32'h0007A0F8 , 32'hFFFD7A07 , 32'hFFFEDCB1 , 32'hFFFC20C8 , 32'h00026E14 , 32'h0002DC24 , 32'hFFFC7EA1 , 32'h00067940 , 32'h000258C3} , 
{32'hFFF83FA1 , 32'hFFFF702C , 32'h000255B8 , 32'hFFFDCF2A , 32'hFFFE373C , 32'h00027BCE , 32'hFFFDE14A , 32'hFFFD0E1E , 32'hFFFD7DBA , 32'h0000E0C0 , 32'hFFFD6DF1 , 32'h0000292B , 32'hFFF9993B , 32'h0002AEFF , 32'h000188BB , 32'hFFFD06C3 , 32'h00008176 , 32'hFFF79A78 , 32'hFFFB75F1 , 32'h000CB33A , 32'hFFFD8F7A , 32'hFFFABC5F , 32'hFFFC9B61 , 32'hFFFD5C58 , 32'h000054D9 , 32'h0001ACB8 , 32'hFFFEBBCF , 32'hFFFD7839 , 32'hFFF9DFE6 , 32'hFFF9D38F , 32'hFFFEAF04 , 32'h00000A2C , 32'h00008A82 , 32'h00019F6F , 32'h0003B812 , 32'h0000A79F , 32'h00002245 , 32'hFFF3F070 , 32'hFFF8984E , 32'h0002B318 , 32'hFFFB6676 , 32'hFFFF51E7 , 32'hFFFF538E , 32'h0000DC70 , 32'hFFFE8934 , 32'h0008BE2C , 32'h0002561B , 32'h000244EF , 32'h00013079 , 32'hFFFF1033 , 32'h0003E69D , 32'h0003D706 , 32'h00050D4F , 32'hFFFDED61 , 32'h0003F9D1 , 32'h00047305 , 32'hFFFDBB82 , 32'hFFFE046F , 32'hFFFC6D5F , 32'hFFFA886D , 32'hFFFF2F0D , 32'hFFFF132F , 32'hFFFDD6DA , 32'hFFFA1E1C , 32'h00044630 , 32'h0006A23A , 32'hFFFEC128 , 32'hFFFDF1CE , 32'h0004D057 , 32'hFFF98C2E , 32'hFFFD9B66 , 32'hFFFB1463 , 32'h0001B6D5 , 32'hFFFF8B95 , 32'h00037562 , 32'hFFFC737B , 32'h0001E8A8 , 32'h000340AC , 32'hFFFB7A0A , 32'hFFFB3EA6 , 32'hFFFC07D0 , 32'hFFFE6DE4 , 32'h00034565 , 32'h000A7539 , 32'h000182A5 , 32'h00011D7F , 32'hFFFF388F , 32'hFFFE03AE , 32'h000628CA , 32'hFFFF8A38 , 32'h0008CDFF , 32'h0002A2B8 , 32'h000437BF , 32'h0002A944 , 32'h0004C886 , 32'hFFFA7196 , 32'hFFFE1796 , 32'hFFF8E6A3 , 32'hFFFFA25B , 32'h000000FD} , 
{32'h00026A05 , 32'h0004FA00 , 32'h00048DA7 , 32'h000550F5 , 32'hFFFFA5E8 , 32'h0000CCB9 , 32'h0004B649 , 32'hFFFBDFB3 , 32'h0002CD51 , 32'h0002808A , 32'hFFF98F1D , 32'h00056340 , 32'hFFFFCA5F , 32'hFFFB1870 , 32'hFFF89536 , 32'h0002131D , 32'h00052E98 , 32'h0009856B , 32'h000107C8 , 32'hFFFDA626 , 32'hFFFAD542 , 32'h0002B06A , 32'h0002BE4A , 32'hFFFAEF96 , 32'hFFF4CAA2 , 32'hFFFD8C12 , 32'h0001E478 , 32'h000555B5 , 32'h00066EB6 , 32'h0005460A , 32'hFFFD259F , 32'hFFF59D72 , 32'h00039D0E , 32'h0002C7F4 , 32'hFFF90729 , 32'hFFFEF9C7 , 32'hFFFCF67A , 32'hFFFEB9C9 , 32'h0004DFD7 , 32'hFFFD9E7B , 32'hFFFE5898 , 32'h000434FA , 32'h0001BE17 , 32'h0006254F , 32'hFFFBB274 , 32'h0006BFE7 , 32'hFFF76516 , 32'h0000ABE6 , 32'h000143E1 , 32'hFFFA8127 , 32'hFFFF7E8E , 32'hFFF93D30 , 32'h00025469 , 32'hFFF6FE52 , 32'hFFF9E68B , 32'h0002D45F , 32'hFFFE1C0E , 32'hFFFFAB71 , 32'h00020E1B , 32'h0004675C , 32'h0002DD16 , 32'h0001D369 , 32'h00026643 , 32'h00024EEB , 32'h0003463A , 32'hFFFD2EB0 , 32'h0006A0A9 , 32'hFFFE03A0 , 32'h00024F19 , 32'h0003909E , 32'hFFF8F96F , 32'hFFFDED95 , 32'h00004864 , 32'hFFFEEA9C , 32'h000271F5 , 32'h00031AE7 , 32'h00056C5B , 32'hFFFF2122 , 32'hFFFD24F3 , 32'hFFF9775C , 32'hFFFC0D66 , 32'h00008979 , 32'hFFFAABF9 , 32'hFFFF57E0 , 32'hFFFE2C0F , 32'h000425E9 , 32'h00076464 , 32'h00015691 , 32'h0008334B , 32'hFFF9BC70 , 32'hFFFF9E63 , 32'h00072268 , 32'h0001108B , 32'h0003CD00 , 32'hFFFDB7BA , 32'hFFFACB18 , 32'hFFFB302B , 32'hFFFD7CA7 , 32'hFFF922DB , 32'h00005698} , 
{32'h05983B68 , 32'hCAE5A340 , 32'h01749624 , 32'h209A3F00 , 32'hF18EBEC0 , 32'hFBCD8618 , 32'h138EA700 , 32'hDE7270C0 , 32'hE3EE3940 , 32'hF2181E20 , 32'h0D497C30 , 32'h120843C0 , 32'h17789960 , 32'h0DEA5B20 , 32'h1BD2A2C0 , 32'hE52D0180 , 32'h022977D8 , 32'h21EE52C0 , 32'hE5FA52A0 , 32'h1AA318E0 , 32'h1A67AA20 , 32'hF7AEF8E0 , 32'hF862E010 , 32'hEA949EA0 , 32'h14549CC0 , 32'h0290EDD8 , 32'h051A24A8 , 32'h0D3CCAD0 , 32'h05F954F0 , 32'hFAE3FA80 , 32'hFC3FBB80 , 32'hEF2435E0 , 32'hF443B550 , 32'h0912D5F0 , 32'h002782D4 , 32'h05CCF858 , 32'h03B2A9EC , 32'hF9A20038 , 32'hF9EC3580 , 32'h063C8830 , 32'h02EBEB5C , 32'h0ED84DA0 , 32'hF579B0E0 , 32'hFCD57958 , 32'hEE68C300 , 32'hFAA56818 , 32'h0592EAF8 , 32'hFB486B28 , 32'hF28212A0 , 32'h0D1AB440 , 32'hF367F9D0 , 32'hEC987420 , 32'hFCCD5FFC , 32'hF200BF50 , 32'hEC7E03E0 , 32'h0ED995C0 , 32'h078B2910 , 32'h006453BD , 32'hF95BF030 , 32'h087CE540 , 32'hFF2B32F2 , 32'h019F13BC , 32'hF5EEF520 , 32'hFEE8F70C , 32'hF36A5F80 , 32'h052F3090 , 32'hF6D623C0 , 32'h11879280 , 32'hFA1C0F80 , 32'hFE365120 , 32'h06A0B3B0 , 32'hF7ED00B0 , 32'h05A9EE28 , 32'h05C5F2A0 , 32'hFBE777D0 , 32'h0367C258 , 32'h076884C8 , 32'hF8A63E08 , 32'hF71C7490 , 32'hFC4AF300 , 32'h0371EA70 , 32'h04BBC2E0 , 32'hFE9494AC , 32'hFE14AB70 , 32'h067FDC68 , 32'hFB70E0B0 , 32'hFD7471A4 , 32'h05198180 , 32'h0575B3F0 , 32'hFFD67F89 , 32'hFFF972E5 , 32'hFFFFBD02 , 32'h0003D80E , 32'hFFF93240 , 32'hFFFDE12F , 32'hFFFFE753 , 32'h00005D56 , 32'h00016BFE , 32'hFFFECAF1 , 32'h0003CF2C} , 
{32'hE4F8EF40 , 32'h7FFFFFFF , 32'h1D650640 , 32'h121F6440 , 32'hFD3257F8 , 32'hF555B9C0 , 32'h3CB44880 , 32'h387C6480 , 32'hF9821AE0 , 32'hCEA008C0 , 32'hDCD38580 , 32'h0B1D30A0 , 32'hF02C5C70 , 32'hF2D29CC0 , 32'h2402D3C0 , 32'hF74F6D70 , 32'hFE76D91C , 32'h0624CA30 , 32'h03A85238 , 32'h0CB65110 , 32'h027BFA04 , 32'hFABD7EB0 , 32'hEB941400 , 32'h107E0480 , 32'hEA254340 , 32'hFFCDC871 , 32'hFC6CEC68 , 32'h0535A240 , 32'hF57AA6C0 , 32'h06625000 , 32'hE3A7A580 , 32'hF6470FD0 , 32'h18FA15E0 , 32'hF95710C8 , 32'hF4D22CA0 , 32'hFF686FA8 , 32'hE216C560 , 32'h2C0813C0 , 32'hDE720D80 , 32'hFD0B1394 , 32'hF055C830 , 32'hFBD9C1A8 , 32'h18596C60 , 32'hF3AEA220 , 32'h00D25DE7 , 32'hFB108E68 , 32'hF97BD978 , 32'hE5A98240 , 32'h00158C1D , 32'hF5EEACE0 , 32'hF23DF6A0 , 32'h09AAF4F0 , 32'h029B7708 , 32'hE53924E0 , 32'h12C92EE0 , 32'hF7183AB0 , 32'h1396C060 , 32'hF201C730 , 32'hFC0DD25C , 32'hED38EEA0 , 32'h138C0300 , 32'h02609A88 , 32'hFEFB4600 , 32'h08777B90 , 32'hFF202C6F , 32'h03B575D8 , 32'h0BD618B0 , 32'hFB2B89A0 , 32'h120F57C0 , 32'hF90ABEF0 , 32'hF9CA7928 , 32'h0651C2A8 , 32'h09FD6230 , 32'hFEA881EC , 32'h0D025790 , 32'h08690800 , 32'h080B49D0 , 32'hFAF25DB8 , 32'hFDC54AEC , 32'h013A65D8 , 32'h04FF91A0 , 32'hFDA5F218 , 32'hFE6F010C , 32'h029FBAC0 , 32'hFFAF4B95 , 32'h03DCA9E4 , 32'h095D46D0 , 32'h01C63A90 , 32'hFC40BB6C , 32'hFE97D7E4 , 32'h0003A8B4 , 32'h000108CC , 32'h00043967 , 32'hFFFC678C , 32'hFFFC5663 , 32'hFFF91C11 , 32'h0001E3E1 , 32'h0001D9BF , 32'hFFFECE0C , 32'h0000C8EA} , 
{32'h5F6B7380 , 32'hF5C85000 , 32'hA6C21900 , 32'h566AB100 , 32'hD6CE7EC0 , 32'hEC634340 , 32'hF3E82710 , 32'h2D796B00 , 32'h4B16DF80 , 32'hD92B6F00 , 32'hE3E095C0 , 32'h0221AA28 , 32'hB6E57C80 , 32'h16591360 , 32'h09A175A0 , 32'hFFC703BE , 32'h19931C80 , 32'h3412B640 , 32'h07845810 , 32'h1B826A80 , 32'h01D33900 , 32'hE164D480 , 32'hEBCA07C0 , 32'h2496F480 , 32'h2529DEC0 , 32'hF9F49148 , 32'h06EC5D90 , 32'hF4CBF460 , 32'h04846A68 , 32'hFB74EBE8 , 32'h0FB88D30 , 32'h0E04F270 , 32'h0F6478A0 , 32'hF242C510 , 32'hF66DCBD0 , 32'hFD6F76DC , 32'h01664B8C , 32'h060C7110 , 32'hDAF3DD00 , 32'h16871FA0 , 32'hF5472C20 , 32'h0373B7A8 , 32'h0FE5E910 , 32'hE81E1F20 , 32'hF39E3430 , 32'h04403FF8 , 32'h11B2BFE0 , 32'hF32D7F20 , 32'h07817C00 , 32'h1AB1D580 , 32'hD4600B40 , 32'h0B22EB70 , 32'h06D0E5B8 , 32'h005EC7FA , 32'h0DFC3800 , 32'h16F9A840 , 32'h063E7388 , 32'hEEA04AC0 , 32'hF967B2C8 , 32'h04441768 , 32'hFC2958C0 , 32'h0AE61460 , 32'hFDDA3F38 , 32'h00577671 , 32'hF650AEB0 , 32'h0A7A12C0 , 32'h01700A80 , 32'hFD66B2CC , 32'hFDB20E54 , 32'hFFD996A3 , 32'h01F99D84 , 32'h017E66D8 , 32'h0688C5A8 , 32'h00FD22CE , 32'h061D6B20 , 32'h062E4D90 , 32'hF81044A0 , 32'h0B8F2960 , 32'h054E68A0 , 32'hF7388BD0 , 32'hFD0C093C , 32'hFB6EC090 , 32'h0272ACD4 , 32'hFC190C38 , 32'h025D2530 , 32'hFF74D0D7 , 32'h01C718A4 , 32'h002198C8 , 32'hFBF256A0 , 32'h015956C4 , 32'hFFFE48B2 , 32'hFFFDD7C3 , 32'hFFFBFC03 , 32'h0004D051 , 32'h00017409 , 32'h00061B90 , 32'hFFFEB17E , 32'hFFFDEE89 , 32'h0000EAFF , 32'h0000A49C} , 
{32'h1B53D640 , 32'hF9D85C18 , 32'hFE2AD268 , 32'h0C4A06C0 , 32'hC6AD0B80 , 32'hE35EC2E0 , 32'hE2FC4F40 , 32'h0B1CAAB0 , 32'h230D68C0 , 32'hD18D47C0 , 32'hFE09B234 , 32'hFE585E44 , 32'h00B0DADC , 32'hE6CDBCA0 , 32'h1293C9E0 , 32'h234BCEC0 , 32'h16037B20 , 32'h0B34C040 , 32'hEDD80A60 , 32'hF1EFF100 , 32'hF5A98AF0 , 32'hE66BC7C0 , 32'hF2EF5640 , 32'h0D9FC390 , 32'h07063A38 , 32'hE67CAF00 , 32'h1E763FC0 , 32'h028EFC48 , 32'hF43CBFF0 , 32'h1EF177A0 , 32'hD51DCB00 , 32'h03AEC534 , 32'hEBD85EC0 , 32'h1C4EFBC0 , 32'hF8CCF900 , 32'hF371EB10 , 32'hFCEFFFBC , 32'hE92638E0 , 32'h07542948 , 32'h19545220 , 32'h081CA780 , 32'h043A3B98 , 32'h0B614640 , 32'h0342A100 , 32'hFF404669 , 32'h165AB8E0 , 32'hFCEF9798 , 32'hEBE6BF00 , 32'h20394D80 , 32'hFE4261A0 , 32'h09FB5900 , 32'hE0E0A860 , 32'hF72112E0 , 32'h0A76DE30 , 32'h02F4A2C4 , 32'h0878A970 , 32'hF349C730 , 32'h09237AF0 , 32'hF6C0FDB0 , 32'h074FC3C0 , 32'hFD57B7C0 , 32'hF2868910 , 32'hFA2CB280 , 32'hF7C70630 , 32'h0B43CC00 , 32'hFDA73E64 , 32'hF31BE240 , 32'hFF642EFF , 32'h0942D400 , 32'h056EF720 , 32'hF13CF120 , 32'h0B9BA410 , 32'h071372C0 , 32'h07341088 , 32'hFD1979F8 , 32'hFCF1957C , 32'h073A6620 , 32'h0054E360 , 32'hFCC06BBC , 32'hFE578CDC , 32'hFB026F18 , 32'h01A52BC8 , 32'h01EE054C , 32'h05DDFB70 , 32'hFF191180 , 32'hFC304B04 , 32'hFFF1E984 , 32'hFF2321A7 , 32'hFEFED960 , 32'hFFBDA958 , 32'h000196C2 , 32'hFFFE2E7A , 32'hFFFCC3AA , 32'hFFFCF348 , 32'hFFFB9D27 , 32'hFFFF7EF7 , 32'h00038B32 , 32'hFFFD02E3 , 32'hFFFDCE7F , 32'h0000CB54} , 
{32'h22527A80 , 32'hD57C9600 , 32'hFDAC8F2C , 32'h0C146B40 , 32'hC046ED80 , 32'hD6310840 , 32'hF0053510 , 32'h102C5FE0 , 32'h25E67340 , 32'hD5BE48C0 , 32'h084F57A0 , 32'hF3540A90 , 32'h10EBA340 , 32'hF43E73D0 , 32'hEC06B500 , 32'h25FDD200 , 32'h1C60DDC0 , 32'hEFE3BD40 , 32'hFC807E2C , 32'h0FD1FEF0 , 32'h0069438A , 32'hE920C3E0 , 32'h0FC64810 , 32'h18001C60 , 32'h0E6DF340 , 32'h03BE82EC , 32'hFB2B1220 , 32'hFB2745B0 , 32'hF17DB670 , 32'hE3B5E8C0 , 32'hF41D1C00 , 32'h02CC8F70 , 32'hE8A4C180 , 32'h0E62B1D0 , 32'hFFB04C69 , 32'h0619D038 , 32'hE6A08C20 , 32'hFE8CC84C , 32'h0CDD57B0 , 32'hEC08EFC0 , 32'hFF3DE73A , 32'h044714B8 , 32'h05C70258 , 32'hF2FB0CF0 , 32'h046436B8 , 32'hFB9C4050 , 32'hE7D74720 , 32'hE2301340 , 32'hE9883B00 , 32'h1CB86D80 , 32'hFBB4F548 , 32'hFAD7A9B8 , 32'hDB39A4C0 , 32'h09CF8FF0 , 32'hFB5DD228 , 32'h06DDFB00 , 32'hFC263140 , 32'h07BF75B0 , 32'h0105A7E8 , 32'h027A2360 , 32'hEB2A54C0 , 32'h0B407E90 , 32'h042E65F8 , 32'h06F1C130 , 32'h026867F4 , 32'h01915DE4 , 32'h014E4AFC , 32'h0951F6D0 , 32'h0A247650 , 32'hEBE0ADA0 , 32'h0259025C , 32'h02DBBD04 , 32'h00D177AE , 32'hFD771D94 , 32'hFE3879EC , 32'hFF9679F8 , 32'hFF0AC08F , 32'hFD7C6B84 , 32'h01152820 , 32'h08352E70 , 32'hFD7CDF64 , 32'h021C3754 , 32'h0A43BD40 , 32'hFBBA95E8 , 32'hFE156AD4 , 32'h03FB2B98 , 32'hFF51B9DF , 32'h026822B4 , 32'h088152E0 , 32'h00455D13 , 32'h0007CC26 , 32'hFFFD81E6 , 32'hFFFD4EF1 , 32'h000039CC , 32'h00013121 , 32'hFFFF7E3B , 32'hFFFEE496 , 32'h00034CCF , 32'h0000392F , 32'hFFFC6A2D} , 
{32'h04F37AE8 , 32'hFBD4B5A8 , 32'hD7B24780 , 32'h226A5A80 , 32'h13B56A00 , 32'hC8F07600 , 32'hC6BDCBC0 , 32'hD95EC5C0 , 32'hE6246200 , 32'h0838D2D0 , 32'h023D41F4 , 32'h0DDB4200 , 32'h0F6B9D40 , 32'h03AA31B8 , 32'hE8A6B3A0 , 32'h2C9C5C00 , 32'h090F4330 , 32'h114F46E0 , 32'hF71B71E0 , 32'hE93877E0 , 32'hEB0FB3A0 , 32'hFB6D3370 , 32'h24EEBFC0 , 32'h1DF268A0 , 32'h02534FBC , 32'h16589300 , 32'h0BE7A120 , 32'hF54CB450 , 32'hE60E5A60 , 32'hDF029180 , 32'hFC3F562C , 32'h11724820 , 32'h04EDA578 , 32'hFA62C870 , 32'h0075B061 , 32'hFF188943 , 32'hDC2EB480 , 32'h0B06DA80 , 32'hF9A42058 , 32'hF475B3A0 , 32'hFBAD5160 , 32'h030D651C , 32'h17339CA0 , 32'hE2AA9F60 , 32'h0E3526A0 , 32'h04B4ED28 , 32'hFE8B5328 , 32'h0B382780 , 32'h00094612 , 32'hEC59E900 , 32'hF9AC03A0 , 32'h160336A0 , 32'h0A33B760 , 32'hFE61EB18 , 32'hDEAE4BC0 , 32'hE9263F40 , 32'hFF0D86C1 , 32'hF9EA0618 , 32'hF998BA08 , 32'h001A425E , 32'hFC316AAC , 32'hFBD10030 , 32'hF9D14D20 , 32'h070FCAB8 , 32'hFBF64B58 , 32'h077FA4E0 , 32'hEC009340 , 32'hFD7F20A8 , 32'hF20F7DD0 , 32'hF981EED8 , 32'hFEE88918 , 32'hFC46742C , 32'h014F9568 , 32'h05473CC8 , 32'hFAF38188 , 32'h042FAF60 , 32'hFEDA7154 , 32'hFF794257 , 32'h04D077F8 , 32'hFC10466C , 32'h00A21258 , 32'hFC51DCC4 , 32'h059ADC98 , 32'h04AFE840 , 32'h070EE198 , 32'h06DC5680 , 32'hFEC9D400 , 32'hFF1557EC , 32'hFED5CC5C , 32'hFF590583 , 32'hFFFDF046 , 32'hFFFD1A09 , 32'hFFFF76DD , 32'hFFFD1AA2 , 32'h0001E463 , 32'hFFFDCC19 , 32'h0001B830 , 32'h00021DE9 , 32'h00001281 , 32'h00002FA7} , 
{32'h00086F1F , 32'h00030681 , 32'hFFFFDD06 , 32'h0001500D , 32'h00078F78 , 32'h0000155D , 32'h0001DFFD , 32'hFFFFB589 , 32'hFFF9B3F1 , 32'hFFFC3F66 , 32'hFFF95FD8 , 32'h0005C097 , 32'h00025F77 , 32'h000535A6 , 32'h0002E9E3 , 32'hFFFC79FD , 32'hFFF87A24 , 32'hFFFC646D , 32'hFFF770AB , 32'hFFFE2082 , 32'hFFFF8FB2 , 32'hFFFF342D , 32'hFFFB9CE7 , 32'h00032544 , 32'h00071A3E , 32'h000394D1 , 32'h00015326 , 32'h000225C6 , 32'hFFFEA3E2 , 32'h0001B891 , 32'hFFFC5C23 , 32'h0002381C , 32'hFFFB5AF1 , 32'hFFFF33B1 , 32'h00082F77 , 32'hFFFAB498 , 32'hFFFE56F8 , 32'h00094E09 , 32'h000259B8 , 32'hFFFCC5AA , 32'h0008922A , 32'hFFF3590E , 32'h00012D00 , 32'h0001AF43 , 32'h00085EDB , 32'hFFFB9165 , 32'h0001F7A6 , 32'hFFFC131F , 32'hFFFF6B9F , 32'hFFFA58F4 , 32'h0006D7A0 , 32'h0002EDFD , 32'hFFFCE1B5 , 32'hFFF90657 , 32'hFFF997BA , 32'hFFFC4853 , 32'hFFFFF025 , 32'hFFFE4C5A , 32'h0001988C , 32'h00023E17 , 32'h00040E64 , 32'h000262EF , 32'h00039AA7 , 32'h00017E95 , 32'hFFF45437 , 32'h0008358A , 32'hFFFEA4D5 , 32'h000148BF , 32'h000AE692 , 32'h000218EA , 32'h0008491A , 32'h00015A59 , 32'hFFFCA19A , 32'hFFFA886F , 32'h0003A606 , 32'h0006677C , 32'hFFFFDA16 , 32'hFFFD5968 , 32'hFFFF2D3C , 32'hFFFB242F , 32'h00036804 , 32'h0006935D , 32'h000274D8 , 32'hFFFECDE2 , 32'h0001CD40 , 32'hFFFCF6F2 , 32'h0003E33D , 32'hFFFE3CD2 , 32'h0000CA33 , 32'h0004141E , 32'hFFFEDACF , 32'h0008C971 , 32'hFFFDA571 , 32'hFFFC7236 , 32'hFFF9E9B1 , 32'hFFF9DEAC , 32'h0005B466 , 32'h00002DEF , 32'h000411F7 , 32'h00003BA2} , 
{32'h00033955 , 32'h000CDE45 , 32'hFFFE0EC0 , 32'h000232EA , 32'h0000E80C , 32'h00035792 , 32'hFFFCE735 , 32'h00010759 , 32'h0003F367 , 32'hFFFB6F3A , 32'hFFFD2F01 , 32'hFFF8D1E0 , 32'hFFF8EA6D , 32'hFFFD676D , 32'h0006452A , 32'h00033FE8 , 32'h0009880E , 32'h0003B506 , 32'hFFF75D23 , 32'h0008388E , 32'h00026538 , 32'hFFFDD1D9 , 32'h0000E784 , 32'hFFF9C6D9 , 32'hFFFC5DAE , 32'hFFFC427E , 32'h0003405D , 32'h0002F814 , 32'h00045A6E , 32'hFFFF4C2D , 32'hFFF6E3AE , 32'h000576FA , 32'h000649AA , 32'hFFF9CF93 , 32'hFFFFA78B , 32'hFFF9302A , 32'h00073CC8 , 32'h00051814 , 32'h00002B24 , 32'h00048468 , 32'hFFFB89F8 , 32'h000492C9 , 32'hFFFB4C75 , 32'hFFFDA8A5 , 32'hFFFE45BB , 32'h000AD4D4 , 32'h0001DDED , 32'hFFFC402F , 32'hFFF94C8B , 32'hFFFF556D , 32'h0002306C , 32'hFFFF2F41 , 32'hFFFE17F1 , 32'h000E0149 , 32'h00059E23 , 32'h0003AA79 , 32'h00007651 , 32'h00019571 , 32'h0008121D , 32'hFFFBF014 , 32'hFFFA9C8A , 32'hFFFE363C , 32'hFFFA0F6E , 32'hFFFB8817 , 32'h0004F09C , 32'hFFFB248E , 32'h00067707 , 32'hFFFDCE0F , 32'hFFFD531B , 32'hFFFDB932 , 32'hFFFC9BB5 , 32'hFFFE0AE6 , 32'h00034F14 , 32'hFFFBD05E , 32'hFFFDD9E8 , 32'h0002F57E , 32'h0005AD11 , 32'h000717CD , 32'hFFFDC7EB , 32'h00036296 , 32'h0000C829 , 32'h000161C7 , 32'h00027E77 , 32'h0003DF20 , 32'hFFFEBA38 , 32'h0005EE6A , 32'hFFFD73C4 , 32'h000823DC , 32'hFFFE3FB6 , 32'h00057EF6 , 32'h0003BD15 , 32'hFFF9F2F2 , 32'hFFFC7297 , 32'hFFF8C7DE , 32'hFFFB23D5 , 32'hFFFDAA80 , 32'h00021BC1 , 32'h0000BC05 , 32'h0004078C , 32'hFFFD3B27} , 
{32'hFFFDB3A4 , 32'hFFF87AB6 , 32'hFFFC916C , 32'h0001DEBE , 32'hFFFE2669 , 32'hFFFC46C6 , 32'h0003821F , 32'hFFFACC24 , 32'h0003BE5C , 32'hFFFA7DEF , 32'h0001E634 , 32'hFFF887DB , 32'hFFFE34DD , 32'hFFFF7BC7 , 32'h0003336B , 32'h0009FAF6 , 32'h00071399 , 32'hFFFF7328 , 32'hFFFA82DD , 32'hFFFCCF70 , 32'hFFFE7B6E , 32'h00039F06 , 32'hFFFC5D12 , 32'h0002951F , 32'hFFFE9FA9 , 32'hFFFE53E3 , 32'hFFFBAFBE , 32'h00010EE2 , 32'hFFFD5882 , 32'h0005E3D0 , 32'h0002DCE5 , 32'h0004E65B , 32'h00047B63 , 32'hFFFE9304 , 32'hFFF93312 , 32'hFFFBC7E6 , 32'hFFFC352E , 32'hFFFF12F8 , 32'hFFF8F2D6 , 32'h000791B0 , 32'h000077E1 , 32'h0000E019 , 32'h00032DE2 , 32'h0001B4A8 , 32'h00014989 , 32'hFFFD5117 , 32'hFFFE137B , 32'hFFFD4182 , 32'h000351B7 , 32'h00002DCF , 32'h00014C49 , 32'h0002FC86 , 32'h000BC2D0 , 32'h00018239 , 32'h000625A4 , 32'hFFFB0C53 , 32'hFFFCE589 , 32'h00013F03 , 32'h0005A742 , 32'hFFFE2795 , 32'h00047E3C , 32'h000413A1 , 32'hFFFDC364 , 32'hFFFFCDFE , 32'h000376A0 , 32'h000383B4 , 32'hFFFC3CA6 , 32'hFFFFABAA , 32'hFFFC1533 , 32'hFFFF7ED7 , 32'hFFFB5A31 , 32'h0003014F , 32'h00032A8E , 32'h0001261C , 32'h00002876 , 32'hFFFDB96B , 32'h0003903A , 32'h00007572 , 32'hFFFBB165 , 32'h0000D1DC , 32'hFFFFB48E , 32'h00021FDA , 32'h00006983 , 32'hFFFC908E , 32'hFFFEF54B , 32'h000306D8 , 32'h00056D1A , 32'h0001AA34 , 32'h000460A1 , 32'hFFFFC092 , 32'hFFFE7A09 , 32'hFFFEC031 , 32'h000812F1 , 32'h000300E4 , 32'hFFFED242 , 32'hFFFF395D , 32'h0002EC39 , 32'h0003060A , 32'hFFFF353F , 32'hFFFFF3F8} , 
{32'hFFFA5870 , 32'h000695B2 , 32'h00015514 , 32'hFFFC2F06 , 32'hFFFDCEEA , 32'hFFFA1A8A , 32'hFFFDEAF9 , 32'h0002AF6D , 32'hFFFD2913 , 32'hFFFE9524 , 32'hFFFAEE41 , 32'h0003F9DF , 32'hFFFDC420 , 32'hFFFB8761 , 32'h000B34E6 , 32'h00001117 , 32'hFFFCE95C , 32'hFFF87B82 , 32'hFFFDB5F0 , 32'h0006A21F , 32'hFFF78759 , 32'hFFFD9500 , 32'h00007956 , 32'hFFFB262D , 32'hFFF8B1A4 , 32'hFFFABD67 , 32'h0001B6F8 , 32'hFFFF4B7C , 32'hFFF810A8 , 32'hFFF8DD6E , 32'h0005B1A1 , 32'h000355A6 , 32'hFFFCD24B , 32'hFFFEB629 , 32'h0001467A , 32'hFFFFA9CE , 32'h0001DFA1 , 32'hFFFA14AA , 32'hFFFBEE23 , 32'hFFFC2173 , 32'h000458D3 , 32'hFFF9572B , 32'hFFFA69A3 , 32'hFFFF787D , 32'hFFFE9E7D , 32'hFFFDCBCD , 32'h000229F5 , 32'hFFFB7DEE , 32'hFFFD7EEE , 32'hFFFDB8E3 , 32'h00074DAD , 32'hFFFDE43A , 32'h00090C1E , 32'hFFFCEE6E , 32'hFFFEB954 , 32'hFFF8D8C6 , 32'h0003A995 , 32'hFFFC887C , 32'h00039C9E , 32'hFFFF97D3 , 32'h00018590 , 32'h000B4A76 , 32'hFFFF9DFE , 32'hFFF91EF6 , 32'hFFF88624 , 32'hFFFFA18E , 32'h0002457E , 32'h0009A867 , 32'h0008FD2E , 32'hFFFDEF48 , 32'h00004E48 , 32'hFFFCA0BB , 32'hFFFEDC79 , 32'hFFFD49F7 , 32'hFFFB02F8 , 32'hFFFB67B6 , 32'h00052CCD , 32'hFFFC3E0B , 32'hFFFEE78D , 32'hFFFC966A , 32'h00003FE5 , 32'h0003D979 , 32'hFFF8DB8C , 32'hFFFAA8E7 , 32'h0001E9E5 , 32'h000710C5 , 32'hFFFC9914 , 32'hFFFE7E15 , 32'hFFFFB78E , 32'hFFF8D501 , 32'hFFFBC87D , 32'hFFFDE9E5 , 32'h00095840 , 32'hFFFD4D0F , 32'h0001F4F8 , 32'hFFFBC1B4 , 32'hFFFCC750 , 32'h000C550B , 32'hFFFDC3DA , 32'hFFFE1D83} , 
{32'hFFFE7761 , 32'hFFFEFA8E , 32'hFFFC6C41 , 32'hFFFFB292 , 32'h000CB1C7 , 32'h000105C8 , 32'h0002230C , 32'h00047513 , 32'h00013B57 , 32'h0005F2AE , 32'hFFF7EDAF , 32'h00063F15 , 32'h000173F7 , 32'hFFFA2A29 , 32'h0003D7DD , 32'h0004D60E , 32'hFFF9B098 , 32'h00039684 , 32'hFFFE4390 , 32'hFFFAECE6 , 32'hFFFFD647 , 32'h000789C0 , 32'h0001D73D , 32'h000F205E , 32'hFFFD5789 , 32'hFFF3BB8A , 32'hFFF93805 , 32'hFFFAF325 , 32'hFFFB7B15 , 32'h00083A30 , 32'hFFFFA677 , 32'hFFF0828F , 32'h000B086F , 32'h0003D2BA , 32'h00039777 , 32'h00021C85 , 32'hFFFD872C , 32'hFFFBE645 , 32'hFFF6F28A , 32'hFFFED8E4 , 32'h000136E9 , 32'hFFFFD56D , 32'hFFFAF9F9 , 32'h0006CBBA , 32'hFFFCA82A , 32'h0002BCBC , 32'hFFFD87AA , 32'h0008ED4D , 32'hFFFC0935 , 32'hFFF17815 , 32'h00065D4E , 32'hFFF5AC0F , 32'h0003FE4D , 32'hFFFC12D2 , 32'h0001C2D7 , 32'hFFFA9CCF , 32'hFFFFBA2C , 32'hFFF5F508 , 32'h00006D99 , 32'hFFFD7E24 , 32'hFFFD5110 , 32'hFFF92E94 , 32'h00014244 , 32'h000076F8 , 32'hFFFE78B6 , 32'h00043238 , 32'h0000FAB1 , 32'h0004C937 , 32'h000967DF , 32'hFFFDAFA9 , 32'hFFFE4400 , 32'h00007FAD , 32'h00035F17 , 32'hFFF72034 , 32'h00003D63 , 32'h00032AA0 , 32'hFFFF6512 , 32'h00082EE3 , 32'h00040E5C , 32'h0009C781 , 32'hFFFC9CA8 , 32'h0006FDD8 , 32'h00039240 , 32'h0001BD15 , 32'h000330BE , 32'hFFF87121 , 32'h0000EC26 , 32'hFFFEAF4E , 32'hFFF9F691 , 32'h00000442 , 32'h00018025 , 32'h000469A2 , 32'hFFFA50BE , 32'h000310A4 , 32'hFFFE4663 , 32'hFFFA5761 , 32'hFFFBC3FF , 32'h0002408B , 32'h0007949D , 32'hFFFCED57} , 
{32'h0A2DA860 , 32'h11E3D100 , 32'h08943370 , 32'hF2063830 , 32'h06506AA0 , 32'h0BFCD720 , 32'hF548A4E0 , 32'h0BA6C080 , 32'h2D28AB80 , 32'hEE9CADC0 , 32'hF2E68470 , 32'hF825CC80 , 32'h1084F7A0 , 32'h0A5C68B0 , 32'hFAE8C020 , 32'hF254EBD0 , 32'hF7BEBDB0 , 32'hF25FB6D0 , 32'h25663880 , 32'hFDE0D494 , 32'h0AC218D0 , 32'hFAD789A0 , 32'hCED12F40 , 32'hF941CCA8 , 32'h26EF8740 , 32'hF1EDF710 , 32'hFA297F78 , 32'h03BE1AE0 , 32'hED717EE0 , 32'hFD82026C , 32'hEC36C7A0 , 32'hE5B8C2A0 , 32'h0660A818 , 32'hFA692900 , 32'hFDACB75C , 32'hFEBCDD7C , 32'h1913EB20 , 32'hED294320 , 32'hE7A8DF20 , 32'hFADC26F8 , 32'hF0019E00 , 32'hFA950420 , 32'hEC75BD80 , 32'h0A218A50 , 32'h0660D438 , 32'hF8E6A5C0 , 32'h27D79440 , 32'hEC90D760 , 32'h04D67298 , 32'hFF5BDA6C , 32'h19D153C0 , 32'hF738EDF0 , 32'hFEC4F690 , 32'h10768960 , 32'h073A1BC8 , 32'h0323C7A4 , 32'hFBD79448 , 32'h05D79BB0 , 32'h0D78C7E0 , 32'h023CE150 , 32'h00C1F1BA , 32'h0B2DA620 , 32'hF5556500 , 32'h05AAF9C0 , 32'h01EAD414 , 32'h02CDB8F4 , 32'hF87F2DC8 , 32'hF8AF6DA8 , 32'hFDB519B8 , 32'hEEC49500 , 32'hFF8549E8 , 32'hF5174900 , 32'hFA842DF0 , 32'h070F7F00 , 32'hFA176AA8 , 32'h0179761C , 32'hFC8CFC68 , 32'hF9875238 , 32'hF4C0E7C0 , 32'hFDEA98D8 , 32'hF54ADC40 , 32'hFCDC2F94 , 32'h00A9E08D , 32'hFCD109FC , 32'hFDCCC094 , 32'h034DC17C , 32'hFB4E9190 , 32'h019E93B8 , 32'hF6FCABC0 , 32'hFF1618A3 , 32'h00011FD1 , 32'h0001917B , 32'h000123E6 , 32'hFFFD4D8A , 32'h00020FB0 , 32'hFFFB7B7B , 32'hFFFAA514 , 32'h0001E318 , 32'h00004D9E , 32'hFFFDAF90} , 
{32'h00AB9A1C , 32'h538ECF00 , 32'hF9FE1238 , 32'hF07C17C0 , 32'hF01E4580 , 32'hFD301288 , 32'hFE89B8CC , 32'h0A676A80 , 32'hEF272F80 , 32'hD86AB7C0 , 32'hF390F340 , 32'h1FFD39A0 , 32'hE88DE6A0 , 32'h0EDBED70 , 32'hE5616CA0 , 32'h1F2D0DA0 , 32'h16212260 , 32'h065F1B20 , 32'h0E534DE0 , 32'h07AB4BF0 , 32'hEB272F60 , 32'h12BEEAC0 , 32'h089B6BF0 , 32'h04331AC0 , 32'hEA4056C0 , 32'h03A993A8 , 32'h0FEBD080 , 32'hDB211540 , 32'h27AB7C00 , 32'hF3EA37B0 , 32'h049A7870 , 32'hF6995F90 , 32'h1854CF00 , 32'h0CE27350 , 32'h04F94760 , 32'hCFDC26C0 , 32'h04BDA378 , 32'h1C324CA0 , 32'h09656940 , 32'hEBDED820 , 32'hFBF20678 , 32'h102C39C0 , 32'hFCA64298 , 32'h06FE0CC0 , 32'h1C3C95C0 , 32'h07A220A8 , 32'h09B14410 , 32'hF443FC30 , 32'h00CD7FF3 , 32'hFF30BB13 , 32'h191BA320 , 32'hEB2A21C0 , 32'h0863CB10 , 32'h0F315550 , 32'hE927E1C0 , 32'hFD5B8128 , 32'hF94BB8A0 , 32'hF0F4B8E0 , 32'h10E2E640 , 32'h047E5FF0 , 32'h0830F910 , 32'h06187240 , 32'h096F2A50 , 32'hF8B4E270 , 32'hFE204398 , 32'hF66A7EF0 , 32'h102BAA80 , 32'hFE55854C , 32'hFF764AD2 , 32'h001E8180 , 32'hF40BBC70 , 32'hFD99639C , 32'h0563B2C8 , 32'h0A7E1BE0 , 32'hFE4CCC50 , 32'h0C2AF210 , 32'hFF8F1F6F , 32'hFB6599B8 , 32'hF6F59E20 , 32'hFB35FC98 , 32'h074A7AE8 , 32'h09B4EC60 , 32'hFA8EE068 , 32'hFF7D73C6 , 32'hFB148338 , 32'h086AA9A0 , 32'h02FC57F4 , 32'h011F649C , 32'hF9C379A0 , 32'h00141DA8 , 32'hFFFFB74D , 32'hFFFFF0A0 , 32'hFFFF7FB3 , 32'hFFFF723F , 32'hFFFE3733 , 32'h0000C9C6 , 32'hFFFF2204 , 32'hFFFDB35A , 32'h00006554 , 32'h000191EC} , 
{32'h2A110B40 , 32'hFB35F3E0 , 32'hF92F3BE0 , 32'h1F9B3700 , 32'hB5131800 , 32'hE91483E0 , 32'hB76B8B80 , 32'hE2E33EA0 , 32'h22129E40 , 32'hE7AE6C40 , 32'hAEEE4180 , 32'h14109E00 , 32'h44272600 , 32'hF9C7F6B8 , 32'h0870CD00 , 32'h0DBD0880 , 32'h0BCA70C0 , 32'hF57F6050 , 32'hE63C3A80 , 32'h1D1231C0 , 32'h2F2D9C80 , 32'h16A44AC0 , 32'h05D3E698 , 32'hDB0DD940 , 32'h108862E0 , 32'hECE5C500 , 32'h04A3E780 , 32'hFEFCA8F8 , 32'h00F9CF7F , 32'hF4288140 , 32'h19163360 , 32'h061FE848 , 32'h0E96E030 , 32'hFCE59B94 , 32'hF43A9650 , 32'hFDE002E8 , 32'hF3BC9DE0 , 32'h08D54DD0 , 32'h276F6F80 , 32'h291B0A00 , 32'hF0F89B80 , 32'hF5D0F090 , 32'h1899F120 , 32'hF1DD0E20 , 32'h04938AA0 , 32'h15C08260 , 32'hEE768BE0 , 32'hED016EE0 , 32'h03A6B6B4 , 32'hFA3247E0 , 32'h054C6550 , 32'h0CC258D0 , 32'hFD676784 , 32'hE3160AE0 , 32'hFFDABDB3 , 32'hF4EE4890 , 32'h08C65180 , 32'h0B3E9D50 , 32'h133DBAA0 , 32'h03D15324 , 32'hF39F4870 , 32'hFD8C14A0 , 32'hEF0B3660 , 32'hFAE0AF70 , 32'hFE0B8EC0 , 32'hF8B67FF8 , 32'h05502190 , 32'h02A98714 , 32'hFCA57A20 , 32'hFA962660 , 32'hF3351880 , 32'hF37383C0 , 32'h03E3B238 , 32'h0268C370 , 32'hFC2C8590 , 32'h04E8B658 , 32'hF8D4E350 , 32'hF8DD6218 , 32'h08261A20 , 32'h0BD6FC10 , 32'hF7AE22F0 , 32'h0578F0A8 , 32'hFC88D52C , 32'hFB5E21D0 , 32'h01B3E058 , 32'hFA6D0B40 , 32'h016EBA40 , 32'h07CBEA60 , 32'hFAFC7958 , 32'h01B92644 , 32'hFFFE64BC , 32'hFFFFCECC , 32'h00025479 , 32'h0003A1EC , 32'h0001DCF3 , 32'hFFFE5FDB , 32'hFFFD3E56 , 32'hFFFE8969 , 32'h0001F237 , 32'h0002BB14} , 
{32'h0004E9CA , 32'hFFFF7706 , 32'hFFFDF372 , 32'hFFF869FB , 32'hFFFECEA0 , 32'hFFFC4D57 , 32'h00065B87 , 32'h0004C0EC , 32'hFFFF6F62 , 32'hFFFEB381 , 32'h0006B6D7 , 32'h000295F5 , 32'h0005632E , 32'h000A279B , 32'h00069476 , 32'hFFFECBC0 , 32'h0001AEA3 , 32'h00073C13 , 32'hFFFE3E85 , 32'hFFF9890F , 32'h000890B9 , 32'hFFFAB8E7 , 32'hFFFA850A , 32'hFFFCD0C9 , 32'hFFFDAEE9 , 32'h00044CAE , 32'hFFFCB9FF , 32'h00023A25 , 32'h000864CB , 32'h00038319 , 32'h0002D1DB , 32'hFFFB0E59 , 32'hFFFAAC5A , 32'hFFF87655 , 32'hFFF8E722 , 32'h0004BDFB , 32'hFFFE4646 , 32'h00036F98 , 32'h0002D59E , 32'h0000BA17 , 32'hFFFE47B2 , 32'h000622D3 , 32'h0004FF91 , 32'h0001D56C , 32'h000187D1 , 32'hFFFB81E5 , 32'hFFFC29EC , 32'h0000310F , 32'hFFFD225A , 32'h000562A4 , 32'hFFFEBC1E , 32'hFFFF5526 , 32'h00021E5B , 32'h0000043F , 32'h0008B9CA , 32'h0000F1D6 , 32'hFFFE6E51 , 32'h00008AFE , 32'hFFFD011D , 32'hFFFF5EFA , 32'hFFFCA1D3 , 32'hFFFC11A8 , 32'h0005AEBC , 32'h0002DB0F , 32'hFFFDD3E1 , 32'hFFFB11EE , 32'h000206ED , 32'hFFFFC74F , 32'hFFF95335 , 32'hFFFEC708 , 32'hFFFCDC57 , 32'hFFF70647 , 32'hFFFCDF83 , 32'h00027CAC , 32'hFFFDEB78 , 32'h0000EBE3 , 32'hFFFA6929 , 32'hFFFBA124 , 32'hFFF736F0 , 32'h00058004 , 32'h00014030 , 32'hFFFE5522 , 32'h0003839D , 32'h0004E39E , 32'hFFF97D7B , 32'hFFFC0ABD , 32'hFFFAA3D4 , 32'h000005E7 , 32'h000B80CC , 32'h000633D7 , 32'h000FC0E7 , 32'hFFF501F8 , 32'hFFFB17FC , 32'h00068D5D , 32'hFFFC8439 , 32'h0000F512 , 32'h00021488 , 32'h0003ED6D , 32'hFFF9B545 , 32'hFFFE41D8} , 
{32'hFFFC7BD7 , 32'hFFFAE6BE , 32'hFFF7B15F , 32'hFFFBF9E1 , 32'h0002B4CF , 32'h00044980 , 32'h00018B2B , 32'h000077F3 , 32'hFFFB76AE , 32'h00008122 , 32'h00089B41 , 32'hFFFB117E , 32'h00012810 , 32'hFFFD0A07 , 32'hFFFD6519 , 32'h00001E50 , 32'hFFEFB6A9 , 32'h00076B7E , 32'h0007D747 , 32'h00027D2B , 32'hFFFFF5E2 , 32'h0005CD8C , 32'hFFFF5299 , 32'hFFFAD322 , 32'h0002C7E0 , 32'hFFFE3299 , 32'hFFFC52EF , 32'h0004A2C2 , 32'h00085805 , 32'h00029B86 , 32'h0004629F , 32'h00000E77 , 32'hFFFF5961 , 32'hFFFBCBBC , 32'hFFFC5C89 , 32'h00029DCC , 32'hFFFBCB79 , 32'h0006FC9F , 32'hFFF63370 , 32'h00061B48 , 32'h000696DA , 32'hFFFAB6B1 , 32'hFFFF4E0B , 32'h0006FF5F , 32'h0003963E , 32'h00065663 , 32'h0001E4E4 , 32'h0004F479 , 32'hFFFA5655 , 32'h00024DF9 , 32'hFFFD3D10 , 32'hFFFE471C , 32'h00011674 , 32'hFFFFAEE1 , 32'hFFFC6226 , 32'hFFFF63D5 , 32'hFFFDD762 , 32'h0007A0D4 , 32'hFFF8B89E , 32'h000493C2 , 32'hFFFCB272 , 32'h00014EF2 , 32'h0001A492 , 32'hFFFE3E6F , 32'hFFFB324F , 32'hFFFDDA00 , 32'hFFFFC167 , 32'h0005CB6A , 32'h00070CC4 , 32'h0000794C , 32'h0008F1EA , 32'h00084266 , 32'h0002DD71 , 32'hFFFC9254 , 32'hFFFAFCE8 , 32'hFFF2CD68 , 32'hFFFBD758 , 32'h000030E6 , 32'h0007CA5A , 32'h0004CB8B , 32'h0000AB71 , 32'h0006A54C , 32'hFFFE91B1 , 32'hFFFC54C2 , 32'h0003BBFF , 32'h00032A0D , 32'hFFFFA3EF , 32'h00023855 , 32'hFFFD183C , 32'h00018F92 , 32'h000D8D4D , 32'h00057DDB , 32'hFFFD8AA6 , 32'h000235A7 , 32'hFFFB1EC3 , 32'h0003CAB7 , 32'hFFFE4171 , 32'hFFF8734A , 32'h000AAF6B , 32'hFFF86F41} , 
{32'hFFFEAA4F , 32'h00024FFF , 32'hFFFF14E5 , 32'h00020EF4 , 32'h00003BAC , 32'hFFFCC354 , 32'hFFFC11CF , 32'hFFFCA181 , 32'h00015815 , 32'hFFFD4F77 , 32'h0000907F , 32'hFFFE059E , 32'hFFFAD38D , 32'hFFFB5F39 , 32'hFFFF3369 , 32'hFFF7DEB5 , 32'h00019F16 , 32'hFFFADC84 , 32'h0000F1C1 , 32'h0008F995 , 32'h00039010 , 32'h0003E409 , 32'hFFFEE921 , 32'h0000B9B8 , 32'h0003F5CC , 32'h00034B5C , 32'hFFFCE740 , 32'h0001F719 , 32'h0006BC21 , 32'hFFFD3577 , 32'hFFFEDF8E , 32'hFFFB43B4 , 32'hFFFEC34F , 32'hFFFA5FEE , 32'hFFF70EA7 , 32'hFFFF87EE , 32'hFFFB5249 , 32'h000210BE , 32'hFFFB5C65 , 32'h0006916A , 32'h00039B2D , 32'h000228ED , 32'h0000B8A0 , 32'hFFFB208F , 32'hFFFEC920 , 32'hFFFAA3A4 , 32'h000B571A , 32'h0001EECA , 32'h0000ABB6 , 32'hFFFBFD7E , 32'hFFFC735C , 32'hFFFC55A7 , 32'h0001DDCB , 32'hFFFAAE74 , 32'hFFFC74BB , 32'hFFFD04F1 , 32'hFFFCB5B7 , 32'hFFF9BCDF , 32'hFFFAED03 , 32'h00012252 , 32'hFFF636E2 , 32'h0000A7F8 , 32'hFFF63119 , 32'hFFF93948 , 32'hFFFDCAF6 , 32'h00033C55 , 32'h000711E1 , 32'hFFFEBA32 , 32'hFFFCC6A0 , 32'hFFFF6C1C , 32'h00049F7B , 32'hFFFE32B4 , 32'hFFF98036 , 32'h00013450 , 32'hFFF97749 , 32'h0003225C , 32'hFFFCDDF6 , 32'h0005591F , 32'h0004A4E3 , 32'h00029129 , 32'h000543A4 , 32'hFFFC5DCF , 32'hFFFC7801 , 32'h00038728 , 32'h0002CA24 , 32'h000259CD , 32'hFFFD3CD6 , 32'h0002EE1F , 32'h0000E15A , 32'h000768DE , 32'h000764F4 , 32'h0002C59D , 32'h00042C26 , 32'h000389EB , 32'h0003A018 , 32'hFFF9EC85 , 32'hFFFD7BDB , 32'hFFFB195B , 32'h00034DE4 , 32'h000185BE} , 
{32'h0008D28B , 32'hFFF94C61 , 32'hFFFD75F5 , 32'h00022C8D , 32'hFFF2B0F2 , 32'hFFFBC264 , 32'hFFFFEE18 , 32'hFFFDEA1D , 32'hFFFBF24D , 32'hFFFC9508 , 32'hFFFFBF7C , 32'hFFFEF5C6 , 32'hFFFA94DA , 32'hFFFA13EA , 32'h00002414 , 32'h0007D71F , 32'h00032B57 , 32'hFFFC0FAB , 32'hFFFE221B , 32'h0001F309 , 32'hFFFFB1EB , 32'h0005E2AE , 32'hFFFD6126 , 32'hFFFDBE4A , 32'h00020275 , 32'h00043C9C , 32'h000192B1 , 32'h0006BFB8 , 32'hFFFCED47 , 32'hFFFDB4D3 , 32'h00010B7A , 32'h00062738 , 32'hFFFE074D , 32'hFFFFDC4C , 32'hFFFFCF33 , 32'hFFFE8EA7 , 32'hFFFA59D8 , 32'hFFFE11B9 , 32'hFFF42B02 , 32'h0008BBF9 , 32'hFFFF55C6 , 32'h00036917 , 32'h000880C8 , 32'h0003CFA3 , 32'hFFF90F62 , 32'hFFFD9B2F , 32'h0006268F , 32'hFFFAD2A9 , 32'hFFFCEA87 , 32'hFFF95BF0 , 32'h000C1EF8 , 32'h000B3EE0 , 32'hFFFBDD2D , 32'hFFFEE25A , 32'hFFF610C5 , 32'hFFFE6C33 , 32'hFFFCDCF1 , 32'hFFFC6139 , 32'h0005D54D , 32'h0005759F , 32'hFFF82C03 , 32'hFFFD0824 , 32'h00053544 , 32'h00010AC2 , 32'hFFFCAE09 , 32'hFFFDBA97 , 32'hFFFB202E , 32'h000CDAAF , 32'h0000024E , 32'hFFFC2B37 , 32'h00046351 , 32'hFFFC2FC2 , 32'hFFF85B74 , 32'h0001BF03 , 32'h00019798 , 32'h000116F8 , 32'hFFFBA258 , 32'h000635E1 , 32'h00003B7D , 32'hFFFE5BE8 , 32'h00020C92 , 32'h00078483 , 32'h00047D95 , 32'h0000B37B , 32'h00026C30 , 32'h0001EAFB , 32'hFFFD9F11 , 32'hFFFC4D9A , 32'hFFF72372 , 32'h00016628 , 32'h00029165 , 32'h000527CD , 32'hFFF72B9E , 32'hFFFE1461 , 32'h00095455 , 32'h00069423 , 32'h0005DB86 , 32'hFFFA71A9 , 32'h0005B3AB , 32'hFFFF28B0} , 
{32'hE96E9160 , 32'hF7B2FDC0 , 32'hE7AD4660 , 32'h0BE2CC80 , 32'h24464440 , 32'h2B9C4A00 , 32'h11CFC000 , 32'h03120048 , 32'h07547420 , 32'h0B252ED0 , 32'h1187C320 , 32'h091F8850 , 32'hE48C8960 , 32'hF184A920 , 32'h03B3226C , 32'hF80D0A48 , 32'hFEABF484 , 32'h0C209500 , 32'h085ED790 , 32'h1F5BA020 , 32'hE66DBEE0 , 32'h0EC25BF0 , 32'h0710FD50 , 32'hE97A3EA0 , 32'h12B26CE0 , 32'hE0147FA0 , 32'hF27DD690 , 32'h06C03CA0 , 32'hFC1A9DB0 , 32'hF82F7FB8 , 32'h0AE76C50 , 32'h0CC7B280 , 32'hF9083970 , 32'hFD826A2C , 32'h07D7B778 , 32'hEF662340 , 32'h0CF69D50 , 32'h102EF920 , 32'h01B6BF18 , 32'h173A8320 , 32'h09B918D0 , 32'hFD2CE40C , 32'h085A6280 , 32'h185F4020 , 32'hFD1606A8 , 32'h096D3EF0 , 32'h052D76F8 , 32'h0132A00C , 32'hF7E955A0 , 32'h013176DC , 32'hEF1001E0 , 32'hFF7C116B , 32'hFC747330 , 32'h002256A7 , 32'hF011EBA0 , 32'h181557C0 , 32'hFBF9F3B8 , 32'h070DEA00 , 32'h07C90EE0 , 32'h021559C4 , 32'h0BB3F9C0 , 32'hF1E27370 , 32'hF9E7FA18 , 32'h0236C2AC , 32'h0062B21C , 32'h0E50F260 , 32'h023DF060 , 32'hFFC925CD , 32'hFDCC9084 , 32'h00CA8EDC , 32'h0231E868 , 32'h0EAF10F0 , 32'hF65945B0 , 32'h096F70A0 , 32'h0307C6CC , 32'h045C10A8 , 32'hF7C79A30 , 32'hF4FE0240 , 32'hFE718D20 , 32'h040ED088 , 32'h0B4F1470 , 32'hF079C4A0 , 32'hFFA5F37E , 32'hF9F448B0 , 32'hFADEF6F8 , 32'hFEF0BCEC , 32'h04370DF8 , 32'h01A8D3CC , 32'hFC975818 , 32'h00B43BCF , 32'h00010AAF , 32'hFFFB5675 , 32'hFFFE645C , 32'hFFFA1981 , 32'hFFFD123D , 32'hFFF99FB4 , 32'h00067767 , 32'h00029169 , 32'hFFFC71B5 , 32'hFFFDBF99} , 
{32'h822EAC00 , 32'h8FF36780 , 32'hF1AB5260 , 32'hE19B59A0 , 32'h1C0881E0 , 32'hCB6D3580 , 32'h45F5F500 , 32'h25038CC0 , 32'h35108A00 , 32'hD2660C80 , 32'h25A1A700 , 32'hD312CCC0 , 32'hD4A8BC00 , 32'hE042AC40 , 32'h5248BF80 , 32'h06CC9790 , 32'h57A0D380 , 32'hF71D8F00 , 32'hEC5DD880 , 32'h0BC032B0 , 32'h037AC024 , 32'h1162AD80 , 32'h22CF1580 , 32'hEC4020C0 , 32'h16B6C480 , 32'hEDEF1BA0 , 32'hCBADCD80 , 32'hEF5A9320 , 32'hF78129F0 , 32'hF9427FB8 , 32'h00310333 , 32'h01173904 , 32'h3386F180 , 32'hFD3EFAC0 , 32'hD4FAEB80 , 32'hF77BDE00 , 32'h101056A0 , 32'hFB8CD568 , 32'h147DCB80 , 32'hE5EC8160 , 32'hEF380680 , 32'h081516D0 , 32'h07B97220 , 32'h184AA620 , 32'h080C53D0 , 32'h01A57C04 , 32'hE97DE6A0 , 32'h0C9751A0 , 32'hF2E0C7A0 , 32'hF0D8B940 , 32'hFB7F3F10 , 32'hFC2D97E8 , 32'h0B5A3180 , 32'h0647AED0 , 32'h04E7B460 , 32'h02DC4A48 , 32'hF50352F0 , 32'h12DC6C60 , 32'h046C6CC0 , 32'h05C97608 , 32'h0A627200 , 32'h0CB92EE0 , 32'h03402CF8 , 32'hFC83588C , 32'hF8BBFA20 , 32'h058898C8 , 32'hF7B51510 , 32'h029F3DF0 , 32'hF6B2C030 , 32'hFB904FF0 , 32'hF8EDFBA8 , 32'h073FEE38 , 32'h03C8D218 , 32'h09822A90 , 32'h015A5080 , 32'h06ED2BA8 , 32'h059CDD38 , 32'h002CFB7A , 32'hFA8B2EF0 , 32'hFDEEBCA0 , 32'hFC1B8D18 , 32'hFC6D4B9C , 32'hFFED63F8 , 32'hFD0BCA4C , 32'h0590CC70 , 32'h053C6960 , 32'hFBF95048 , 32'h009D0595 , 32'h03BD5DB8 , 32'h00C951C8 , 32'hFFFF942A , 32'h000220FB , 32'h00040A58 , 32'h0000DF53 , 32'h0002321D , 32'h00024640 , 32'hFFFD8AB1 , 32'h00010D8D , 32'h0004239F , 32'h000035F8} , 
{32'h00021BE4 , 32'h00078AD6 , 32'h000004E1 , 32'h00005F62 , 32'hFFFA975E , 32'h00012080 , 32'h0006D638 , 32'hFFFEA3C1 , 32'h0003FCF6 , 32'hFFF800E8 , 32'h00005412 , 32'h0003EC93 , 32'h000793CA , 32'h00020392 , 32'hFFFEFB60 , 32'hFFFBAB5B , 32'h0008214A , 32'h00038CDE , 32'h00026776 , 32'hFFFDCD3C , 32'hFFFF95F1 , 32'hFFFFA979 , 32'h0002C061 , 32'hFFFD566B , 32'hFFFEF39C , 32'h0001909F , 32'h0004E4A1 , 32'h0000B669 , 32'hFFFF9E98 , 32'h000173F5 , 32'h00037138 , 32'hFFF6A9C9 , 32'h0001464D , 32'h000278BA , 32'hFFFEA9AC , 32'hFFFFC3FD , 32'h000272B4 , 32'h0000C359 , 32'hFFFD81EA , 32'hFFFA6836 , 32'hFFFFCCB9 , 32'h00013DF8 , 32'h0001E05C , 32'h0005A7BB , 32'h00003FD7 , 32'hFFFF1ED2 , 32'hFFF9CCE7 , 32'h0000C312 , 32'h0007120A , 32'hFFFC91A4 , 32'h000077D1 , 32'h000792E4 , 32'hFFFFB3FF , 32'hFFFF8D42 , 32'hFFF76609 , 32'hFFFC51B3 , 32'h00043EAE , 32'h00069BEC , 32'h000392D3 , 32'hFFFE56BE , 32'hFFF89E49 , 32'h000081DC , 32'hFFFD7EA6 , 32'h0002B13B , 32'hFFFF1C96 , 32'hFFFC9B21 , 32'hFFFE5FB2 , 32'hFFFBC1F0 , 32'h0009660B , 32'hFFF94688 , 32'h00011ED4 , 32'h0008C1F1 , 32'h0002980B , 32'hFFFB1478 , 32'hFFFDC838 , 32'h000192F8 , 32'hFFFC7A81 , 32'hFFFEC392 , 32'hFFFBA471 , 32'hFFF9149B , 32'h00084413 , 32'hFFFAC13C , 32'hFFFD325A , 32'hFFFDC5B9 , 32'h000548FE , 32'h0000EE4C , 32'h0003A078 , 32'h00004154 , 32'h00069A90 , 32'hFFFE3E3A , 32'h0002E11C , 32'hFFF67230 , 32'hFFF7B27E , 32'hFFFB2695 , 32'hFFFBC1EA , 32'hFFFF7EC5 , 32'hFFF87554 , 32'h00028F27 , 32'h00031543 , 32'h0002F61C} , 
{32'h00097E63 , 32'h0005C0A1 , 32'h00026309 , 32'hFFFCE0CD , 32'hFFFB41AD , 32'h00049651 , 32'hFFF6AB7D , 32'h00022EBF , 32'hFFF6DA07 , 32'hFFFE1DA1 , 32'h00025A1D , 32'hFFF68C71 , 32'hFFFD7120 , 32'hFFFB4D24 , 32'h00038980 , 32'hFFFF4BD5 , 32'hFFFBC676 , 32'hFFFE45DA , 32'hFFFF77E5 , 32'hFFFA7523 , 32'hFFFD48B9 , 32'h00033380 , 32'h0000CE12 , 32'hFFFE1F16 , 32'h00032647 , 32'hFFFE30A8 , 32'h000308F3 , 32'hFFF74B14 , 32'h000683FE , 32'h0001BE82 , 32'h0002D506 , 32'hFFFEDD54 , 32'h00036BDF , 32'hFFFF03F2 , 32'h000365B1 , 32'hFFFF745D , 32'hFFFC191B , 32'hFFFEFDF5 , 32'h0004128E , 32'h0001F75C , 32'hFFFBF213 , 32'h00047192 , 32'hFFFEF2D1 , 32'hFFFEB367 , 32'h000349DB , 32'h000225D2 , 32'hFFFE0C76 , 32'hFFFF2E5E , 32'h00017295 , 32'h00022A84 , 32'h0001ACEE , 32'hFFFBCBEB , 32'h00075D90 , 32'h000159DA , 32'h00006141 , 32'hFFFDC79A , 32'h000447F3 , 32'h00025954 , 32'h00029403 , 32'hFFF874F9 , 32'hFFFD269D , 32'hFFF9F1F4 , 32'hFFFAF883 , 32'h00028523 , 32'hFFFD6E58 , 32'hFFF9B7B0 , 32'hFFFF9706 , 32'hFFFB8C65 , 32'hFFFA929C , 32'h00095B5D , 32'h0002ECB3 , 32'hFFFAF29A , 32'hFFFF3BCF , 32'hFFFEFAF3 , 32'hFFFBB330 , 32'h0000887D , 32'h00062DBB , 32'h00045154 , 32'h0000BAF1 , 32'h00041A8F , 32'hFFFCF4D7 , 32'h0001B75E , 32'hFFFEA369 , 32'hFFFBB337 , 32'h00038387 , 32'hFFFDF08A , 32'hFFFF5B65 , 32'h00088DFC , 32'hFFFB6F7B , 32'h0005530D , 32'hFFFE1069 , 32'hFFF2F78F , 32'h0000D4E9 , 32'hFFFFCE7A , 32'h0004412A , 32'hFFFA1D7B , 32'h0000AADB , 32'hFFFAEB3F , 32'hFFFF85D8 , 32'hFFFFEFAE} , 
{32'h00003556 , 32'hFFF8EEE5 , 32'hFFFAF00F , 32'hFFFEFEE5 , 32'hFFFE5C5B , 32'h0008A884 , 32'hFFFFF2B7 , 32'hFFFFC12D , 32'h0007F0C6 , 32'hFFFA702B , 32'h0004F6FB , 32'h00069505 , 32'hFFFC81B6 , 32'h0003217D , 32'hFFFB1640 , 32'h00005D2D , 32'h00043B12 , 32'h0002CCDD , 32'hFFFC356E , 32'hFFFC2D27 , 32'h0002CCAD , 32'h000199DC , 32'h000254C3 , 32'h0004E3A0 , 32'hFFFD056B , 32'h0002C1B6 , 32'hFFF6A57E , 32'h000115FB , 32'h00032CCD , 32'hFFFCEB61 , 32'h0000693E , 32'h00007554 , 32'h00018054 , 32'hFFFE4FF2 , 32'h0003B6B3 , 32'hFFFFA6DD , 32'h0000D167 , 32'hFFFB1E90 , 32'hFFFBAE58 , 32'hFFF9937D , 32'h00056C39 , 32'hFFFA6F76 , 32'hFFF8E9E3 , 32'h0002228C , 32'h000EDADD , 32'h00015C5B , 32'hFFFEAAE2 , 32'hFFFC554E , 32'h000D3FD6 , 32'hFFFC18B6 , 32'h00065FF4 , 32'hFFFE9D02 , 32'h00020D4D , 32'hFFF41748 , 32'hFFFC4002 , 32'h0003438B , 32'h0003D67C , 32'h0003214E , 32'hFFF9118B , 32'hFFF86EF5 , 32'h000499C4 , 32'hFFFC7A1A , 32'hFFFD1834 , 32'hFFFCA573 , 32'hFFFE2C8A , 32'hFFFB8DF3 , 32'hFFFE19AA , 32'hFFF93167 , 32'h00025673 , 32'hFFFD619C , 32'h00049A6B , 32'h0000C80E , 32'hFFFDDEA5 , 32'hFFFDD462 , 32'hFFFC5BE5 , 32'h0008A183 , 32'h000663E9 , 32'h0009668E , 32'h00012707 , 32'h00025425 , 32'hFFF5410E , 32'hFFFED27A , 32'hFFFB9356 , 32'hFFFD7A7E , 32'hFFF717E7 , 32'h00005C51 , 32'h00091704 , 32'hFFFD019F , 32'hFFFF4F1D , 32'hFFFE7408 , 32'hFFFBFEE1 , 32'hFFFFE1F7 , 32'hFFFC842D , 32'hFFFE6499 , 32'hFFFD251D , 32'hFFFD105D , 32'h0000BC8C , 32'hFFFBDA73 , 32'h00001D3C , 32'h00021D36} , 
{32'h41228C00 , 32'hB1E14B80 , 32'h24862500 , 32'h9F42E380 , 32'hA4092180 , 32'hFEDC87DC , 32'h4A312800 , 32'hEAF37520 , 32'hACE14900 , 32'hFF0DF3F8 , 32'h18B37EC0 , 32'hEE6FCCE0 , 32'hEECE2420 , 32'h1F5D49A0 , 32'hFD6C69A0 , 32'hB98B2D00 , 32'h0D9AA560 , 32'h1D9C1820 , 32'h07D64670 , 32'h1A500D00 , 32'h15299D60 , 32'h11974DE0 , 32'hEF2DB540 , 32'h1959D800 , 32'h33BC2B40 , 32'h14B6F840 , 32'hFE450A78 , 32'hEF733760 , 32'h0E3484D0 , 32'hF2D94BC0 , 32'h1B475520 , 32'h08097810 , 32'hF0262BD0 , 32'hF2450EC0 , 32'hEE265B80 , 32'hF3485770 , 32'h0A6151A0 , 32'hFC9824FC , 32'h13826B20 , 32'hF7C87F40 , 32'hF4990640 , 32'h067D18F0 , 32'hF1FAEF10 , 32'hEFC92A40 , 32'hFDF3BE8C , 32'h229F5F40 , 32'hD5C15D40 , 32'hFC097274 , 32'h0B07C5E0 , 32'h06178480 , 32'h0F28FF00 , 32'hFA94E368 , 32'hEF9B3DE0 , 32'h053A6C20 , 32'hFCB55858 , 32'h0157CF68 , 32'hF56F6200 , 32'h017611B0 , 32'h03E23A50 , 32'hF2AEC1E0 , 32'hFF746662 , 32'hFE40ED14 , 32'hF1387B90 , 32'h05431D30 , 32'hEE0286C0 , 32'hF5661AC0 , 32'h04D07FD0 , 32'h06019D78 , 32'hFF46E391 , 32'h0948DBC0 , 32'h02EA6AEC , 32'hF3DC4B90 , 32'h021EAC04 , 32'h06EAAA50 , 32'h08CC6D80 , 32'hF79F16F0 , 32'h052002D8 , 32'hFB97EDD8 , 32'hFD5E5458 , 32'hFEC122E8 , 32'h07D7D8F0 , 32'hFD44335C , 32'hFF23D902 , 32'hFF6E23F1 , 32'hFCE7E608 , 32'h05E3B7C0 , 32'hFC7777C4 , 32'hFCA635F8 , 32'hF8BDDDC0 , 32'hFFD741A7 , 32'hFFFBAA86 , 32'hFFFFD8AE , 32'h00010A98 , 32'hFFFECED2 , 32'hFFFDAB6C , 32'hFFFD5892 , 32'h0003643F , 32'hFFFDECEE , 32'hFFFCDA0F , 32'hFFFF99DB} , 
{32'h09A302A0 , 32'hB4632200 , 32'h1381E660 , 32'h17775B00 , 32'hE87B5360 , 32'h7FFFFFFF , 32'hC2BF1100 , 32'h0BDC3DE0 , 32'h41948880 , 32'hC17A2BC0 , 32'h1D21C360 , 32'h421C2000 , 32'h04311670 , 32'hDF64FB40 , 32'h0C7A9330 , 32'h3F07B3C0 , 32'h085014A0 , 32'h1D4DC980 , 32'hE387B120 , 32'hFE9237A8 , 32'h0965FE20 , 32'h1FD2AAE0 , 32'hF13B7D80 , 32'hE9318200 , 32'h1CD3AD60 , 32'h19204660 , 32'hEBB8C3A0 , 32'h047BE400 , 32'h14E1AB80 , 32'h0056A7EA , 32'h03E4D5D4 , 32'h1BA1B5A0 , 32'h0386778C , 32'hF91486C0 , 32'h0982ADB0 , 32'h17936B60 , 32'hEB971C00 , 32'h0C0FD2E0 , 32'hE86A9480 , 32'hFE3F12FC , 32'h16B9EFA0 , 32'h101EDCE0 , 32'h08B59030 , 32'h0B2CF880 , 32'hFF42DBBD , 32'h02E88DC8 , 32'h0E90FD30 , 32'h055F23D0 , 32'hF5E3D290 , 32'hFB3D0508 , 32'h048545E0 , 32'hF8D49EE0 , 32'hFF8ADA07 , 32'h09A7E020 , 32'h0CE733C0 , 32'hFF67957B , 32'hE3508F40 , 32'h097FCF80 , 32'h0018FFCD , 32'hFE4F4828 , 32'hFA9F1868 , 32'hECD7FCA0 , 32'h03FB5B0C , 32'hFCC99378 , 32'h00D6A241 , 32'hED105FC0 , 32'h03A10220 , 32'hFE8C7F74 , 32'h02162718 , 32'h07D7CF20 , 32'hFFBF944F , 32'hFB110408 , 32'h031EA024 , 32'hF8279628 , 32'hFD9E0528 , 32'hFFAD400F , 32'h0566CF20 , 32'h06DD2558 , 32'hFDB33C8C , 32'h009800B1 , 32'h05123F18 , 32'hFD62CBF8 , 32'hFF104E10 , 32'h0235DF10 , 32'h020E369C , 32'h074B7600 , 32'hFCD65344 , 32'h044D7C08 , 32'hFFDA2733 , 32'hFF34C400 , 32'h0006B7D7 , 32'hFFFFF443 , 32'hFFFFBB74 , 32'hFFFDC3D2 , 32'h0000AE86 , 32'hFFF98B27 , 32'h00027B35 , 32'hFFFCAF67 , 32'hFFFEECA0 , 32'h00005DF1} , 
{32'hA2D5F700 , 32'h9D009380 , 32'h0FF1F7D0 , 32'h156C1180 , 32'hCAEB3600 , 32'hA0C96A80 , 32'hD0B2BF00 , 32'h0EFAE9E0 , 32'h1B445C60 , 32'h271A3A00 , 32'h1C83A600 , 32'h263EED40 , 32'h20F8E940 , 32'hF2715C10 , 32'hC316C500 , 32'h0F517370 , 32'h0066EE99 , 32'h07388E80 , 32'hDE629DC0 , 32'h01900908 , 32'h02E25974 , 32'h15AC1500 , 32'h148FEEE0 , 32'h1CB60100 , 32'hD8C99500 , 32'hC6A45600 , 32'hFF054D31 , 32'hFE1F1124 , 32'h33FA4000 , 32'hF7EEE690 , 32'h0C740120 , 32'h01B424D4 , 32'h1773C1E0 , 32'hF8E81D78 , 32'h0EEAD0E0 , 32'h0797A400 , 32'hFFC19F6F , 32'hF5A3A1C0 , 32'h079E5A28 , 32'h09F13400 , 32'hEFDA4AE0 , 32'hF764DC10 , 32'hF25CF0F0 , 32'h1050A240 , 32'h0073892C , 32'hF6AFFB60 , 32'hF2FE7D40 , 32'h025107AC , 32'h179B1C80 , 32'hF84355F8 , 32'hEF0A3E20 , 32'hF4246F90 , 32'hF4E82E50 , 32'h08BB2170 , 32'h16581A60 , 32'h0615D970 , 32'hF57DD530 , 32'hE9FF2C00 , 32'h0B174B40 , 32'hFDE2E69C , 32'h0E67C530 , 32'h08B3F2D0 , 32'h0238DC78 , 32'h09F17680 , 32'hED147E00 , 32'h0E0B4390 , 32'h00FFE475 , 32'h0FAFF070 , 32'hF6EFCA20 , 32'h076948F8 , 32'hFCB51DB8 , 32'hFAB7E960 , 32'hFE6D6398 , 32'hFC055DFC , 32'hF4C28AB0 , 32'hFE0D90CC , 32'h058731D8 , 32'h0891D140 , 32'h049B8658 , 32'h008286F1 , 32'hF9AC08E8 , 32'hFDF7C490 , 32'h02871B24 , 32'hFFB69986 , 32'h027437B0 , 32'hFD27C390 , 32'h037FC16C , 32'h0228CF98 , 32'hFDCF0B18 , 32'hFA34E540 , 32'h0002A258 , 32'hFFFEC17C , 32'hFFFE0CD4 , 32'hFFFFE64D , 32'h0002AC3A , 32'h00008BD2 , 32'h00003B10 , 32'h0001B057 , 32'hFFFEF7B7 , 32'hFFFEAC9E} , 
{32'hFFF90B9E , 32'hFFFEE503 , 32'hFFFE16E6 , 32'h0002C716 , 32'h00029D25 , 32'h00011B2F , 32'hFFFC916B , 32'hFFFF19E3 , 32'hFFFA0ED3 , 32'hFFFEBF8F , 32'hFFFFD689 , 32'h0000029E , 32'hFFFE59AD , 32'hFFFE08B5 , 32'hFFFB4A2E , 32'h0001BFB9 , 32'hFFFB20FA , 32'hFFFDC79E , 32'h000510C7 , 32'h0001D117 , 32'h00023D3C , 32'h000B585C , 32'hFFFA8D36 , 32'h00078717 , 32'hFFFC92A0 , 32'hFFFC6F95 , 32'h0000EE49 , 32'hFFFE7B32 , 32'h000F27A7 , 32'hFFFE2030 , 32'hFFFE940B , 32'hFFF9EFD7 , 32'h00027F9C , 32'h0004D0D9 , 32'hFFFC2F90 , 32'hFFFB2A1A , 32'hFFFE1F74 , 32'hFFFE4C94 , 32'h0000DB20 , 32'hFFFD0B66 , 32'h000427C7 , 32'h00006B24 , 32'h00049E5F , 32'h00024770 , 32'hFFFBF2FB , 32'h000540F8 , 32'hFFFDA3AB , 32'h00060547 , 32'h000BAF3D , 32'h00037B2B , 32'hFFFE88B7 , 32'h00041861 , 32'hFFFF0AD5 , 32'h000198A5 , 32'h0003F30D , 32'h00058179 , 32'h0001558D , 32'h000243E6 , 32'hFFFE954F , 32'h0002B65D , 32'hFFFD0FDF , 32'h00014F55 , 32'h00004DAA , 32'h000A0201 , 32'h0004B119 , 32'h0003FB7E , 32'hFFFE35F2 , 32'hFFF6F345 , 32'h000087FF , 32'h0001A9E0 , 32'h00099F8A , 32'h00005164 , 32'hFFFD9E68 , 32'h00032CE8 , 32'hFFF8750E , 32'hFFFFE252 , 32'hFFFF98A0 , 32'hFFF928E6 , 32'hFFFD4664 , 32'hFFFE8F9C , 32'hFFFD7C05 , 32'hFFF852EE , 32'hFFFC342D , 32'hFFFCFDCA , 32'h00032972 , 32'h0003E349 , 32'h000221A0 , 32'hFFFA4A69 , 32'hFFFB6689 , 32'h00041A58 , 32'hFFFE0755 , 32'hFFF57965 , 32'h0001C01F , 32'h00046BBE , 32'hFFFB71A2 , 32'h000E38C6 , 32'hFFFE8E3A , 32'hFFFDF961 , 32'hFFFFA4E9 , 32'h00028465} , 
{32'h00032B16 , 32'h0002FC1F , 32'hFFFA5F4F , 32'hFFFF050F , 32'hFFFB96D5 , 32'h00039ABC , 32'hFFF73972 , 32'hFFFA7D8B , 32'hFFFD60B6 , 32'h00011C42 , 32'hFFF0D4EB , 32'h0003A7EE , 32'h000191A5 , 32'h000127BD , 32'hFFF7D771 , 32'h0008B6DF , 32'h0001FBE5 , 32'hFFFAB819 , 32'hFFF941D8 , 32'hFFFE8206 , 32'h00073BE3 , 32'h0001A0F5 , 32'h0000B653 , 32'h00063336 , 32'h000C4145 , 32'h00050064 , 32'h0000AB36 , 32'hFFFD05B7 , 32'h00076369 , 32'hFFFB9441 , 32'h00040EB7 , 32'h000099C3 , 32'h00093ABD , 32'h00069F62 , 32'h0000EDAC , 32'h000597F5 , 32'hFFF67BE8 , 32'h00084BEC , 32'h0000EE8E , 32'hFFFB0869 , 32'h0000E81E , 32'hFFFDA95D , 32'h0008A911 , 32'h00012B85 , 32'h0000C782 , 32'h0007899E , 32'h000ADACA , 32'h000BE115 , 32'hFFF8A393 , 32'h00022144 , 32'h00001CD3 , 32'h0001A635 , 32'hFFFBCCC5 , 32'h0006F6D3 , 32'hFFFFCD9D , 32'hFFFF7E09 , 32'h0001AC20 , 32'h0006958B , 32'h0008C7CC , 32'hFFFB205F , 32'hFFF9AA85 , 32'h00019848 , 32'hFFFCC67D , 32'hFFF8F694 , 32'hFFFDB039 , 32'hFFFCC46D , 32'hFFF811D3 , 32'hFFFBF969 , 32'hFFFEDDEA , 32'h00001E0E , 32'hFFFC8299 , 32'h00028F02 , 32'h0009AD60 , 32'h000665CF , 32'hFFFAFD93 , 32'hFFF9D59A , 32'h00047D81 , 32'h0007D891 , 32'h0003E490 , 32'hFFFD4A4C , 32'hFFFD59CB , 32'h0007A996 , 32'h00012F1E , 32'h0001E894 , 32'hFFF9D55A , 32'h00039E35 , 32'hFFF88E84 , 32'hFFFF0B50 , 32'h000B7D44 , 32'hFFFA9167 , 32'hFFF20527 , 32'hFFFA4B2B , 32'h000A0F4F , 32'h00058B1A , 32'hFFFDA4DE , 32'hFFFADA6B , 32'h0002B63E , 32'h00023765 , 32'hFFFBFD1B , 32'hFFFB37FF} , 
{32'h0006D198 , 32'hFFFDC520 , 32'hFFFE156D , 32'h00056BD7 , 32'h0002D3F9 , 32'hFFFFA4B5 , 32'h00046ED5 , 32'hFFFC8E44 , 32'h00034228 , 32'hFFF7A415 , 32'h00021D0E , 32'hFFFC9104 , 32'h000399B5 , 32'h0002888B , 32'h0001423F , 32'hFFFB3A9D , 32'h000904E1 , 32'h000828F7 , 32'hFFFC3629 , 32'hFFFF1558 , 32'h00036631 , 32'hFFFB8C3A , 32'h0006346B , 32'hFFFD9470 , 32'hFFFFFA2B , 32'hFFFEAAB3 , 32'h00060A63 , 32'hFFF7A58E , 32'hFFFE1A1F , 32'hFFFF0C09 , 32'h000720AE , 32'hFFFFA293 , 32'h0000B5C0 , 32'h0001FD4B , 32'h00068D37 , 32'hFFFDF557 , 32'hFFFDFCAA , 32'h0000559C , 32'h00002D6F , 32'h0003B13A , 32'h00034052 , 32'h00022744 , 32'hFFF9200B , 32'hFFFFFCB9 , 32'h00088A15 , 32'hFFFC9E11 , 32'hFFFDFCF8 , 32'h00058FAE , 32'h0002AEBE , 32'hFFF9EBEF , 32'hFFFDF9C4 , 32'h0005D214 , 32'hFFFD532D , 32'hFFFCF0F7 , 32'h000073F6 , 32'h0000CEBE , 32'h00004228 , 32'hFFFDFB74 , 32'h00080998 , 32'hFFFB2E2C , 32'hFFFFCBDE , 32'h00005700 , 32'h0003D2AF , 32'h000539CF , 32'h0001D566 , 32'h0006C345 , 32'hFFFE3D45 , 32'h00007730 , 32'h00024FA9 , 32'h0001B899 , 32'h0001115C , 32'h000D7882 , 32'hFFFE9FC1 , 32'h00072BA5 , 32'h0001C45D , 32'h000D2C12 , 32'h0000678B , 32'h0003C496 , 32'h00039477 , 32'hFFF76284 , 32'h00018B0D , 32'h00038F3C , 32'h0005127D , 32'hFFFBD14F , 32'hFFFEB6DC , 32'hFFF9E42E , 32'hFFFF4E05 , 32'h0000B324 , 32'hFFFFA7BB , 32'h00013485 , 32'h0008AD0C , 32'hFFFDB5FE , 32'hFFFCA5D7 , 32'hFFFE6B1A , 32'h0005F822 , 32'hFFF98DF0 , 32'hFFFD380E , 32'hFFFDE225 , 32'hFFF63E7D , 32'h0002F037} , 
{32'h0A8224B0 , 32'hF1C49800 , 32'h0F7C3810 , 32'hE24BDD60 , 32'h01BC9C18 , 32'hE54064C0 , 32'h13F86100 , 32'hEA0137C0 , 32'hFBBBF138 , 32'hFDF1F890 , 32'h1148D1E0 , 32'h00FBE286 , 32'h0A64ECB0 , 32'hF5D0F6C0 , 32'hE6BCAB80 , 32'hE48C6BE0 , 32'h1A296880 , 32'hFE1B0F24 , 32'hF9244090 , 32'h1AA9FA80 , 32'h1AD13640 , 32'hF0BDBF40 , 32'h0AF08260 , 32'h09BFF5A0 , 32'h117CC6E0 , 32'hF41F8BD0 , 32'hF9BE3EA8 , 32'hFBD31ED0 , 32'hFC358F34 , 32'hFF299FF1 , 32'hF5A93870 , 32'hF09B7C20 , 32'hFE910DD4 , 32'h055D1298 , 32'h07946080 , 32'h023517CC , 32'hF76E83E0 , 32'h0A1A0E70 , 32'h046BBB38 , 32'hF2D38470 , 32'h13DA8020 , 32'h0A219150 , 32'hF8803828 , 32'hEE8EB500 , 32'h116C8700 , 32'h0FCB07E0 , 32'h13E80A40 , 32'hF359BB60 , 32'hF3ED9E70 , 32'h036577B0 , 32'hFC2ACD48 , 32'h0459A2B8 , 32'h0EE3E470 , 32'h040865C0 , 32'hF795F520 , 32'h0407AF18 , 32'h1165D2E0 , 32'hF28A8260 , 32'hFBEF56B8 , 32'hF8CAF1C8 , 32'h05F441F8 , 32'h0820D780 , 32'h0B7462F0 , 32'hF8FEF6C0 , 32'h017EA03C , 32'h022E4F3C , 32'hFD8F7BDC , 32'h08ABDAC0 , 32'hFEF4D394 , 32'h12AEA160 , 32'hFF88DD43 , 32'h0FC27140 , 32'hF79D2CF0 , 32'h0239B494 , 32'hFD0C0974 , 32'hFBAC94E8 , 32'h0A372810 , 32'hF8306FF8 , 32'hFABFE118 , 32'hFD8FC2EC , 32'hF3728040 , 32'h06D97F50 , 32'hFF93834A , 32'hFDD7FBD8 , 32'h017C1940 , 32'h00E396EF , 32'h03E047BC , 32'h00096DEA , 32'hFEB55EEC , 32'h00A26610 , 32'hFFFF7B1A , 32'h000659EB , 32'h0001A19B , 32'hFFF4E897 , 32'h0002CC67 , 32'hFFFF30C6 , 32'h0000D823 , 32'h0000D587 , 32'hFFFE6535 , 32'hFFFD3FC3} , 
{32'h06869DA0 , 32'h06548338 , 32'h1816B660 , 32'hF8A54000 , 32'h0E8F89C0 , 32'h1B78B000 , 32'hFB381380 , 32'hEB2A6500 , 32'hFCDD50C4 , 32'hEDB05BA0 , 32'hF4326310 , 32'hF3662FB0 , 32'hEFFC47A0 , 32'hEF4D0E40 , 32'h110F4F00 , 32'h1217D6A0 , 32'hE6AEFC80 , 32'hEE316D00 , 32'hFB497C10 , 32'h0A857240 , 32'hF24A9D20 , 32'hF08648E0 , 32'hF8870C18 , 32'hF33803C0 , 32'hFF019380 , 32'h04351160 , 32'h0330AA9C , 32'h10DA9560 , 32'hFA494480 , 32'hFF6E31F2 , 32'hFBA32B48 , 32'hEC7C46E0 , 32'h129BAA80 , 32'hEEF4D500 , 32'h008BA06F , 32'hE772BBC0 , 32'hFCA7BDA4 , 32'hECD1EB40 , 32'h01C41E10 , 32'hF6185500 , 32'hF27E75B0 , 32'h03D9A7B0 , 32'h1105DC80 , 32'hE8F9FC80 , 32'hF560DD10 , 32'h0217C14C , 32'hFBE9EE20 , 32'h10A511A0 , 32'hF8C57610 , 32'hFC821BF4 , 32'h023D74B8 , 32'hFC24D4D8 , 32'hFFE03E05 , 32'h0593DCD8 , 32'h0CC012D0 , 32'h02C61504 , 32'hF6B49DA0 , 32'hF1A8ED10 , 32'hF9D189E0 , 32'hFDE0DF50 , 32'hF9BE1448 , 32'hF238E1B0 , 32'h0708EE50 , 32'h004F3A83 , 32'h0312BFD4 , 32'hFD017474 , 32'hFFDE5740 , 32'h0606DD08 , 32'hFA1D0268 , 32'hEDDDB560 , 32'h0BB02C50 , 32'h0F06E1D0 , 32'hF709ECF0 , 32'h00482BFA , 32'hFC866AE4 , 32'h013A8F18 , 32'h06627778 , 32'h008E17B1 , 32'h0A54CED0 , 32'h03000158 , 32'hFCADB02C , 32'hFC96C2CC , 32'h03650E98 , 32'hF9C4D610 , 32'hFA29D678 , 32'hFB4DF178 , 32'hFC57BED4 , 32'hFB6B09F8 , 32'hFFA02682 , 32'hFFA1CA1E , 32'hFFFC86F3 , 32'h000390B2 , 32'hFFFDDF55 , 32'h00010C07 , 32'h0001A635 , 32'hFFFAB7C2 , 32'hFFFDFEFC , 32'hFFFEDC11 , 32'hFFFCC895 , 32'h0001D644} , 
{32'h5D274700 , 32'hC92A7B00 , 32'hC5CB1580 , 32'h2ABDFD80 , 32'hCB13E480 , 32'h85280E80 , 32'h308B3780 , 32'hC3A163C0 , 32'hFEB03B4C , 32'h5F386800 , 32'hE66DD0E0 , 32'h03717E04 , 32'hD9043400 , 32'h23E11900 , 32'h3AF50600 , 32'h24EADBC0 , 32'h20B13B80 , 32'hFE794034 , 32'h0D646D70 , 32'h017F3230 , 32'h2160C580 , 32'hD368DF80 , 32'hF0F6DC30 , 32'hF6EF39C0 , 32'h00D8A8A2 , 32'h0B8283E0 , 32'hF2B37FF0 , 32'h0B74C640 , 32'h0554C4A8 , 32'hF6107EB0 , 32'h04123690 , 32'hE54CF600 , 32'hF8086A30 , 32'h162B2660 , 32'hF70D8880 , 32'hFCC7E4F4 , 32'hFD9F8094 , 32'h116DC140 , 32'h0A9E8E80 , 32'h0C66CD10 , 32'h135F0E00 , 32'h03345160 , 32'h0609F6C0 , 32'h0CADEAA0 , 32'h0F46E380 , 32'hC5A69180 , 32'h072BB038 , 32'h0FB5C7D0 , 32'h0D6C24E0 , 32'hFA564C30 , 32'hFCCAF94C , 32'hF840A270 , 32'h14C90860 , 32'hF642DD70 , 32'h015728B8 , 32'h00803616 , 32'h0024F4C1 , 32'h03BE1CDC , 32'h0136E7A4 , 32'hF9413218 , 32'h04A7BD90 , 32'hFC7632C0 , 32'h09C39350 , 32'hFD3C059C , 32'h00BD1DA1 , 32'hF6FFCF10 , 32'h08D44470 , 32'h0435BC78 , 32'h03E72AE8 , 32'hF8E2AD60 , 32'h0DA44FF0 , 32'hFBF7EF50 , 32'h06FE05E8 , 32'hFAFFD348 , 32'hFCA8E320 , 32'h03CA4170 , 32'h07357060 , 32'h02584B04 , 32'h041F32F0 , 32'h04CE63C0 , 32'h00A59EB1 , 32'h06A4A7F8 , 32'hFD47E390 , 32'h049318F0 , 32'hFB9CEB18 , 32'h0296EEF0 , 32'hF91224B0 , 32'hFA9AC378 , 32'hFE7243B8 , 32'hFEC7D570 , 32'h00002C37 , 32'hFFFF0104 , 32'hFFFF6F75 , 32'h00020B05 , 32'hFFFE2F40 , 32'h0000E230 , 32'h00026944 , 32'hFFFC9C0D , 32'hFFFD7D03 , 32'h00004CE8} , 
{32'h00028219 , 32'hFFFB8877 , 32'hFFFD5CBC , 32'hFFFD39A5 , 32'hFFFBC849 , 32'h0003223E , 32'h0001166A , 32'hFFFD1675 , 32'h0003C87A , 32'h00031689 , 32'h00068EC0 , 32'hFFFFF415 , 32'h00078FA0 , 32'h0001B031 , 32'hFFFF5482 , 32'h0001C05D , 32'h00024999 , 32'hFFF6069B , 32'hFFFC5863 , 32'hFFFEB038 , 32'h000600E9 , 32'hFFFF08EF , 32'hFFFB13C7 , 32'hFFFA53F9 , 32'hFFFEC644 , 32'hFFFD565C , 32'hFFFE9A4B , 32'hFFFF9C78 , 32'h00028860 , 32'h0009321B , 32'h0004BA17 , 32'hFFFAD495 , 32'h00016FF2 , 32'hFFFDB7F7 , 32'h00006E62 , 32'hFFF363E4 , 32'h0003EAA2 , 32'h0002D754 , 32'hFFFDE2BB , 32'hFFFE0571 , 32'h00038545 , 32'h0004DC5D , 32'hFFFAEE8B , 32'hFFFDE56E , 32'h00088320 , 32'h0000BDB4 , 32'h000099BF , 32'h0004DEDD , 32'hFFFF17CA , 32'h000184A6 , 32'h00000242 , 32'h00019BC5 , 32'h00025467 , 32'hFFF9ACB1 , 32'hFFFE8470 , 32'hFFFF06C6 , 32'hFFFF30FF , 32'hFFF7E908 , 32'hFFFA4159 , 32'hFFFE19F7 , 32'h00006050 , 32'h0001B6F6 , 32'hFFFF6077 , 32'h000B18BF , 32'hFFFE71BE , 32'hFFFD1D46 , 32'hFFF613A6 , 32'hFFFEE395 , 32'hFFFFC4E6 , 32'hFFFFDCCC , 32'h00017CCC , 32'h0001443A , 32'hFFF7887C , 32'hFFFD1880 , 32'hFFF68EF8 , 32'h0003797E , 32'hFFFD42DB , 32'h00027C29 , 32'hFFFDA3A5 , 32'h0005A502 , 32'hFFFC32E5 , 32'hFFFE75FE , 32'h000A06EF , 32'hFFF7190E , 32'h0004AE8E , 32'hFFFC8A4D , 32'hFFF95159 , 32'h00065541 , 32'h000329DD , 32'h00034C18 , 32'h000543A0 , 32'hFFFBC264 , 32'hFFF4C223 , 32'hFFF85CFA , 32'h00068A0D , 32'hFFF85BC6 , 32'hFFFEE45F , 32'h00001356 , 32'h00072681 , 32'h000090E6} , 
{32'h00EE50A6 , 32'h061497D8 , 32'hF9DA67E0 , 32'hF97D1478 , 32'hFB9B2220 , 32'h021C7C50 , 32'hF4522F30 , 32'h00322160 , 32'h019A3FE0 , 32'hFACA53D0 , 32'h01AE69E0 , 32'hFE98FB70 , 32'h0197BE48 , 32'h02CAD924 , 32'h040A6A20 , 32'h072CFAB0 , 32'hFBAF0B18 , 32'hFDDC78E0 , 32'hFF2E4469 , 32'hFD849DE4 , 32'hF5F2DCD0 , 32'hFD3BA9A8 , 32'hF6D8D2E0 , 32'hF6439080 , 32'hFFDB4888 , 32'h0442D1D8 , 32'hFABE4410 , 32'h07BD9360 , 32'hFA231668 , 32'h01BC12D8 , 32'h04FBFD50 , 32'hFE84A1B4 , 32'hFA141160 , 32'hFC1B05D8 , 32'h02E4B398 , 32'hFFF8B44D , 32'hFCC874D4 , 32'hFDC957B4 , 32'h0065CEFD , 32'hF753D720 , 32'hFFD1A39C , 32'h04030B50 , 32'hFEDE94B8 , 32'h04FF85F0 , 32'hFE6180E4 , 32'hFB1C46E8 , 32'h0147DCA4 , 32'h0269FF90 , 32'hF977CD20 , 32'hF85852E8 , 32'hFBE2F8D8 , 32'h039B5934 , 32'h00E347D4 , 32'hFE61A02C , 32'hFFAD30E1 , 32'h0128F730 , 32'hFE298D0C , 32'hFC7816B8 , 32'h040405D0 , 32'hFD6B8C60 , 32'h02E4147C , 32'hFF0E758C , 32'hFE6BB8D4 , 32'h0007C3A2 , 32'h02354248 , 32'h0512AF28 , 32'hFCCBBBEC , 32'hFC60B064 , 32'h001BDCB3 , 32'hFF4B94BB , 32'h00A66C23 , 32'h026B3634 , 32'h013371C8 , 32'h047FC818 , 32'hFD790A64 , 32'hFDC915A4 , 32'hFEAB2BAC , 32'h03AB976C , 32'hFCC3B10C , 32'hFD08209C , 32'hFF0EEE0A , 32'h003A8446 , 32'hFD7D1404 , 32'hFF41A2CF , 32'h009EB0B1 , 32'hFFB69BFC , 32'hFC534B34 , 32'h067D40B0 , 32'h013D597C , 32'hFFE70A2D , 32'hFFFDDFF1 , 32'h0007BFFA , 32'hFFF54DD5 , 32'h0002E776 , 32'hFFF8CFA1 , 32'h0003FAC2 , 32'h000C8DC9 , 32'hFFFCC7CB , 32'hFFFF1E49 , 32'h00009F2F} , 
{32'hFFFA7815 , 32'hFFF6F53A , 32'hFFFE949C , 32'hFFF7443B , 32'h0003B58D , 32'hFFF56356 , 32'hFFFB2FE6 , 32'hFFFA652F , 32'h000A38AA , 32'h0001C82F , 32'h0001F05D , 32'h000502AA , 32'hFFFA9DC3 , 32'h0000B42E , 32'h001060CB , 32'h0008890B , 32'hFFFA7207 , 32'h0006458F , 32'h0001445E , 32'h000657D1 , 32'hFFF292A4 , 32'hFFF16BCC , 32'hFFFBDD74 , 32'h0008C424 , 32'hFFF78CF1 , 32'hFFFADCA3 , 32'h00047D88 , 32'hFFFEABAE , 32'h000564FF , 32'h0002768E , 32'hFFF80EF4 , 32'hFFFDE113 , 32'h00058F3C , 32'h0004526A , 32'h0002F3AA , 32'h0000C9DA , 32'hFFFBEA3B , 32'hFFF75560 , 32'h0000CE97 , 32'hFFFF5DA3 , 32'hFFFACAC0 , 32'h00040FD0 , 32'hFFFA509B , 32'hFFFBC2C6 , 32'h0007D56F , 32'hFFF24AAC , 32'h0000DAAD , 32'h00020894 , 32'hFFFE0064 , 32'h0004018E , 32'h000658ED , 32'hFFFFA6BB , 32'hFFFDD713 , 32'hFFF317D7 , 32'hFFFB9078 , 32'h0003FD74 , 32'h00023E60 , 32'h00003319 , 32'hFFFF62BE , 32'h0007FE68 , 32'h000682F7 , 32'h00028F34 , 32'hFFFE59B8 , 32'hFFFE3036 , 32'hFFF7D0BF , 32'hFFFF64A6 , 32'hFFFEAA29 , 32'hFFFFFDDA , 32'hFFFE45A2 , 32'hFFFBA288 , 32'hFFFC1D91 , 32'h000D34BB , 32'h000329EE , 32'h00061DEF , 32'hFFF3D3DD , 32'h00003C43 , 32'h00026FCB , 32'h0007F8E1 , 32'hFFF9BBBC , 32'hFFFA70C9 , 32'h0000AC41 , 32'hFFFEA05C , 32'hFFF9D561 , 32'hFFF27270 , 32'hFFFA6D9B , 32'h0003072B , 32'h000226C8 , 32'hFFF9642A , 32'hFFFFD94A , 32'hFFFF44F1 , 32'hFFFD2A39 , 32'h000321E3 , 32'h00033E2F , 32'h0001B4C9 , 32'h0001C704 , 32'h00006BF0 , 32'hFFFF6D9B , 32'h0002C86F , 32'hFFFE21A0 , 32'hFFF79589} , 
{32'hF6AE08F0 , 32'hF0017150 , 32'h21B30600 , 32'hE12953C0 , 32'h224FA6C0 , 32'h27AF1D00 , 32'h52B7C080 , 32'hF1E26750 , 32'hDD400980 , 32'h6069D400 , 32'h09B96390 , 32'h069EE250 , 32'hECB36320 , 32'hF1DDB3E0 , 32'hD151C780 , 32'hD41BEFC0 , 32'h058D0DA0 , 32'h01B0B720 , 32'h09165580 , 32'h046A1620 , 32'h2884E940 , 32'h0BB24E20 , 32'h32207740 , 32'hEC91F220 , 32'hF052CF80 , 32'hE8196C20 , 32'hFA6FD5F0 , 32'h1DEDC820 , 32'hF7CAEE20 , 32'h06A0E2F8 , 32'h0465FA58 , 32'h127BEC60 , 32'h1D23A2C0 , 32'h011C15A0 , 32'h14983720 , 32'h13A2F1C0 , 32'hFB9DE2F0 , 32'h01501330 , 32'hD12B91C0 , 32'h15B99260 , 32'hF52A5700 , 32'h03A6A0EC , 32'h12851940 , 32'hE72623A0 , 32'hFDAB9674 , 32'hFAAB2058 , 32'h0041E105 , 32'h0140E028 , 32'hF0434370 , 32'h0DC60400 , 32'h01478DD0 , 32'hFDF68924 , 32'hF642E4F0 , 32'hF371DF30 , 32'hFDB722C0 , 32'h13531B20 , 32'h0539BBF8 , 32'h0D905A50 , 32'h038CBBBC , 32'h0315D1D8 , 32'hFB68DD20 , 32'h01BF5148 , 32'hF9677580 , 32'hFC7BBF80 , 32'h07561178 , 32'hFD364DA8 , 32'h03F5BFF4 , 32'hF973AC90 , 32'hFC900F18 , 32'h08C03600 , 32'hF559D730 , 32'h01296A04 , 32'hFEDEEB5C , 32'h038641A8 , 32'h0D911570 , 32'hFD2C54A4 , 32'h01C02E68 , 32'hFBD69D40 , 32'h0343C2C4 , 32'h02AF4B1C , 32'hF631D9A0 , 32'h02BEA3A8 , 32'hFC2B33C0 , 32'hFC236BCC , 32'hFAAE4AC0 , 32'h03211748 , 32'hFA5B0930 , 32'hFBAE1FA0 , 32'h039023A4 , 32'hFFBB0A2D , 32'h000538F5 , 32'h000280B6 , 32'h00000626 , 32'hFFFF8371 , 32'h000164A0 , 32'h000087A4 , 32'h000305A9 , 32'hFFFEE207 , 32'h00016BEC , 32'hFFFF81A8} , 
{32'h0004BB8D , 32'hFFF0235A , 32'h000E21DA , 32'hFFFF02FF , 32'h00067D7F , 32'hFFFA430A , 32'hFFFF9BFA , 32'hFFFCBF4C , 32'h00000DDE , 32'h0006447D , 32'hFFFBA36B , 32'hFFFF9CB5 , 32'h0001C87F , 32'h0006574F , 32'hFFFD735C , 32'hFFF5D6AB , 32'h00001156 , 32'h000357BC , 32'hFFFBEC24 , 32'hFFF8A87B , 32'h0002B8B8 , 32'h0008A7C6 , 32'hFFF522E6 , 32'hFFF7CE7F , 32'h000C9D44 , 32'h00044B37 , 32'hFFFF2133 , 32'h0000BFA8 , 32'hFFFC4BE2 , 32'hFFFFB6F7 , 32'hFFF89B70 , 32'h00066E5C , 32'h0002C94E , 32'hFFF87CE3 , 32'hFFFE3BA3 , 32'hFFFC50A0 , 32'h00035340 , 32'h0004534E , 32'h0002B79F , 32'hFFFC1751 , 32'h00028EC1 , 32'hFFF96F44 , 32'hFFF7A715 , 32'hFFF746C5 , 32'hFFF29E12 , 32'h0000BE67 , 32'h000137EA , 32'hFFF90DEF , 32'h0009D9CB , 32'h00045CCC , 32'hFFFEF034 , 32'hFFFE29FF , 32'h00067CB9 , 32'h0007F0BB , 32'h000BEF93 , 32'hFFFC81E1 , 32'hFFFE9B17 , 32'h00089483 , 32'h00053A8E , 32'h0006EE61 , 32'hFFFD129B , 32'hFFF6593B , 32'h00042640 , 32'h000316F9 , 32'hFFFF9663 , 32'hFFFBBC92 , 32'hFFF98FD2 , 32'h000B1F0E , 32'hFFFD845E , 32'hFFFD5A88 , 32'h0008FAC8 , 32'hFFF49867 , 32'h0002E5EC , 32'h00062417 , 32'h0009FE1D , 32'h00027E09 , 32'h0001A3DB , 32'h00035959 , 32'hFFFC1B4D , 32'hFFF841BF , 32'h0002A942 , 32'hFFFF5EB1 , 32'h00063D63 , 32'h000662FC , 32'hFFF63667 , 32'h000C876B , 32'hFFFDB22B , 32'hFFFAD8E9 , 32'h00037BE2 , 32'hFFFE9FD5 , 32'h0000AF43 , 32'h0001ADD4 , 32'h000441B9 , 32'h000611E6 , 32'hFFFF100B , 32'h0002A603 , 32'hFFFA664A , 32'hFFFE3DE8 , 32'hFFFE6042 , 32'h0001F009} , 
{32'h29485A80 , 32'hA8946F00 , 32'h4E7E6E80 , 32'h031526B4 , 32'h69EF1D80 , 32'h7FFFFFFF , 32'hB9FFB380 , 32'hEBECB6C0 , 32'hDCE848C0 , 32'h38BA9140 , 32'h1538CAE0 , 32'hD9A7CD80 , 32'h2C4A0FC0 , 32'h0F106520 , 32'hE52A2960 , 32'hFA4878C8 , 32'h3B4A9B80 , 32'h0EFB5380 , 32'hCFD14B00 , 32'h3EC1F380 , 32'hFEB16574 , 32'h05E40148 , 32'h18091840 , 32'h1D9A3C00 , 32'h19611340 , 32'hD952B240 , 32'hFC615AE0 , 32'h0131D514 , 32'hE980BF60 , 32'h198E16A0 , 32'hFEF26BA8 , 32'hDEB07640 , 32'hFFD5C953 , 32'h08CBB970 , 32'h16B23140 , 32'hF8C9B350 , 32'h000ADDFB , 32'h36C9B9C0 , 32'h14E00FC0 , 32'h05236FF8 , 32'hF974B958 , 32'hFE496370 , 32'hF6C2FDA0 , 32'h077B7EA0 , 32'hF68D5940 , 32'hF759CCB0 , 32'hF51FA390 , 32'h0816F290 , 32'h07075420 , 32'hE998F1A0 , 32'h0D88F580 , 32'h0D6CF4A0 , 32'h09680690 , 32'hEC9B1BE0 , 32'hF94C4698 , 32'hF78DEAD0 , 32'hEBBE6980 , 32'h06DFE5E8 , 32'hF8D67A28 , 32'h01BA4BB4 , 32'h00A12315 , 32'h07421B70 , 32'h0573E5D0 , 32'hFDF51C84 , 32'h0BDD6810 , 32'hFD7EEB90 , 32'h072DBBC0 , 32'hFCECD638 , 32'h0680C5A8 , 32'hF3046F70 , 32'h03B79F24 , 32'hFC953E44 , 32'hF95BE958 , 32'h0542F2F8 , 32'hFF813F96 , 32'h00381567 , 32'hF6259070 , 32'h07BF8528 , 32'hFF896F47 , 32'hF6406F50 , 32'h00669397 , 32'hFC6124CC , 32'h0926B130 , 32'h00092E1E , 32'hFD5A9D60 , 32'hFD44E238 , 32'h008A06D9 , 32'hFE094E4C , 32'hFEAF9C78 , 32'hFF12DA9A , 32'h000064A0 , 32'hFFFD4B5D , 32'hFFFBE881 , 32'h000224E3 , 32'hFFFDB7AE , 32'h0000B1C4 , 32'h0001D0A5 , 32'h00022326 , 32'h0002E9A4 , 32'hFFFFD912} , 
{32'hFFFCD550 , 32'h0001DD16 , 32'h000431B6 , 32'hFFFEB85A , 32'h0000868D , 32'hFFFCA287 , 32'h00030AAD , 32'h00057839 , 32'hFFFC0AA1 , 32'hFFFC36AC , 32'h0003F9A7 , 32'h000526F7 , 32'h00001654 , 32'hFFFA6611 , 32'h0002F8CB , 32'hFFFB305C , 32'hFFFF15E2 , 32'h00039176 , 32'h00003263 , 32'hFFFC57C1 , 32'hFFFD1C43 , 32'h0005B0F1 , 32'h0004305E , 32'hFFF8BA6C , 32'hFFFDBD49 , 32'h00012AE7 , 32'hFFFA919C , 32'h00087288 , 32'hFFF975BF , 32'h0004D733 , 32'h00017482 , 32'hFFFB29AC , 32'hFFFBCABC , 32'hFFFF061C , 32'h0000709D , 32'h0000AC56 , 32'h00075072 , 32'h000C605E , 32'hFFF8F000 , 32'h00002005 , 32'hFFF92C1A , 32'h0001415F , 32'hFFFA814B , 32'h0006B6C4 , 32'h00037255 , 32'hFFFAFD6D , 32'hFFFCBA02 , 32'hFFFFD589 , 32'h00002940 , 32'h000E8487 , 32'hFFFC53E4 , 32'hFFFDEC89 , 32'hFFFB5744 , 32'hFFF8A753 , 32'h0001605F , 32'h0003686F , 32'h0001D4E8 , 32'h0002C16B , 32'h00090F5B , 32'hFFFC1A6F , 32'hFFF7358C , 32'h00002ECB , 32'hFFFF59D9 , 32'h000293F3 , 32'h0000A996 , 32'h0004CCBB , 32'hFFF98856 , 32'h0008AAAA , 32'h0007874A , 32'hFFFEE56B , 32'h00074D9B , 32'h0004FDBC , 32'hFFF7327E , 32'hFFFEACE7 , 32'h0009E592 , 32'hFFF99AFF , 32'hFFF68165 , 32'hFFF94319 , 32'hFFFD4FCD , 32'hFFF909E8 , 32'h0002393D , 32'h00042CFE , 32'hFFFED05D , 32'hFFFE0163 , 32'hFFFEBF57 , 32'h000489B5 , 32'hFFFC43BB , 32'hFFFD0CD8 , 32'hFFF86AFF , 32'hFFFA5F2A , 32'h000868C4 , 32'hFFF89AB2 , 32'hFFFEF0EA , 32'h000311E5 , 32'hFFFF1A52 , 32'hFFFB9736 , 32'h000171CE , 32'hFFFBA3B9 , 32'h0000A5BA , 32'h00045F2C} , 
{32'h0C270770 , 32'h7FFFFFFF , 32'h3B746E40 , 32'h2EDD0AC0 , 32'h37AA6980 , 32'h145BB0C0 , 32'h6DBB1480 , 32'h5DF61500 , 32'h2C480640 , 32'h33F0F500 , 32'hDE638840 , 32'h0ACA8CC0 , 32'h0BF97C40 , 32'h09D04CF0 , 32'hF1313F20 , 32'hFA0B55C8 , 32'h2FDC3700 , 32'hE6AB0960 , 32'hDF7DF6C0 , 32'hFECC7820 , 32'hE9992A40 , 32'hF0CA8C60 , 32'hECCD1080 , 32'h1E7CAFE0 , 32'hEB3B9DA0 , 32'hF1FEEE00 , 32'hF2BB3A40 , 32'h1EC743A0 , 32'h06FBA0E0 , 32'hE0241C80 , 32'hEF01BB20 , 32'hCB25D980 , 32'hFE16EB64 , 32'hEAA150A0 , 32'h01122BCC , 32'hF3BB1360 , 32'hFB589CA0 , 32'h08455720 , 32'h1B50F400 , 32'hF9715F00 , 32'hD018FA00 , 32'hF6E689D0 , 32'h0F237F80 , 32'hF40E4C10 , 32'hEB9E7680 , 32'h1824CB40 , 32'h08C4DF20 , 32'h014AF2B0 , 32'h1223D0C0 , 32'h037C42F4 , 32'hF349DB40 , 32'hF48CBA70 , 32'h02FF5540 , 32'hFC6CD9E0 , 32'h09860B70 , 32'hFA33E438 , 32'hF63F2DA0 , 32'h01C0D8B4 , 32'h06880458 , 32'h00CC0654 , 32'hF38DA680 , 32'hEF965B00 , 32'h047CB920 , 32'hF7BC0960 , 32'hF9395580 , 32'h0749C348 , 32'hFCF8FEC0 , 32'h073041A8 , 32'h03F8EE48 , 32'h0BBEA460 , 32'h04C527C0 , 32'h01C3BD0C , 32'h05F62918 , 32'hFA175308 , 32'hF54C42C0 , 32'hF8D4B520 , 32'hF76F0DF0 , 32'hFC7D6610 , 32'hFD515164 , 32'h00D49438 , 32'h0B9773D0 , 32'h00ADE67D , 32'hFBE41BD0 , 32'h00A9D976 , 32'hFF9EA79B , 32'h054BAC88 , 32'hFCAF42A4 , 32'h004002E4 , 32'h04A40BE8 , 32'h01077070 , 32'h00005C55 , 32'hFFFF980A , 32'h0000B297 , 32'h000308F1 , 32'h00026136 , 32'hFFFE62AF , 32'h0000F9B0 , 32'h00028E9C , 32'h0000A4A7 , 32'hFFFF5014} , 
{32'h3D0A2680 , 32'hF242AE00 , 32'hEEE858A0 , 32'h3FF50E00 , 32'hFEE220C4 , 32'hE296E6E0 , 32'hF0978130 , 32'hF6FA65D0 , 32'hF6F72C50 , 32'hBB8A8980 , 32'hF04502F0 , 32'h2B8BFD40 , 32'hEB3C0180 , 32'h17AA0F60 , 32'hD2990380 , 32'hDF20E6C0 , 32'h20A2F780 , 32'h021F46D4 , 32'h0ABE1B00 , 32'hF6DD5430 , 32'hE72664C0 , 32'hE936B720 , 32'h1916A0A0 , 32'h031DA850 , 32'hF55F77B0 , 32'h05C1BEC0 , 32'h0A667420 , 32'hF2BCC7A0 , 32'hB5B03480 , 32'hF7D424D0 , 32'hECE19700 , 32'hE3B3DCE0 , 32'hF73ECF40 , 32'h015DD60C , 32'h0CA0D0B0 , 32'hEF29CDE0 , 32'h0ECF6700 , 32'hFA02D2A0 , 32'h07FD3C08 , 32'hEF11D200 , 32'h04D1D118 , 32'hF5A85270 , 32'hFA001760 , 32'h07752340 , 32'hE2835B00 , 32'h089E1340 , 32'hF482B310 , 32'hFDED8F20 , 32'h039F9298 , 32'hFB59AD30 , 32'hFF035C6B , 32'h13FC5780 , 32'hF7462250 , 32'h014AD4C4 , 32'hFBA1B988 , 32'h0804BB20 , 32'hFF33F03A , 32'hF25FFB10 , 32'h08F927B0 , 32'h04B28AF0 , 32'hFBEE9900 , 32'h0C968FB0 , 32'hFE7815EC , 32'hFA2E6938 , 32'h093DAE10 , 32'hF8579610 , 32'hFF0052D1 , 32'h0CC35260 , 32'h0A240180 , 32'hF8368838 , 32'hF552A7E0 , 32'hFCA9B0AC , 32'hFD0F3D3C , 32'hFECF8BE4 , 32'hFC49D3A8 , 32'h00C419E7 , 32'h03C7BA34 , 32'hFFB5B880 , 32'hF963E3A0 , 32'h03BF8268 , 32'hFE517C90 , 32'hF65446F0 , 32'hF61897C0 , 32'h10555820 , 32'h0663D7D0 , 32'hFCDEC9C4 , 32'hF9005030 , 32'hFCF608D4 , 32'hFFCC009A , 32'hFE93233C , 32'h00029791 , 32'hFFFEB038 , 32'h0001383D , 32'h00016F2A , 32'hFFFE373B , 32'hFFF8C624 , 32'hFFFF6C70 , 32'hFFFF0602 , 32'hFFFD2C08 , 32'h00028F65} , 
{32'h7FFFFFFF , 32'h28DDAC40 , 32'h73A28080 , 32'h9CC80800 , 32'hB65B9080 , 32'h0C198FA0 , 32'h080E8470 , 32'hE77B0C00 , 32'h04A759A8 , 32'hE74C6420 , 32'hC016FC40 , 32'h0CDC0E90 , 32'h0E3AC330 , 32'h3156C1C0 , 32'hE46E0600 , 32'h0A0A8A10 , 32'h316D8980 , 32'hFE495F04 , 32'h18683E60 , 32'h190050C0 , 32'hF40F01C0 , 32'hD2E862C0 , 32'h1DC8D720 , 32'hFECC05EC , 32'hFCAC8504 , 32'h348124C0 , 32'h2B255540 , 32'h081C71B0 , 32'h00D05033 , 32'h0E2DF500 , 32'h1854DDA0 , 32'hD7578C00 , 32'h1D2B0620 , 32'h0478F7F0 , 32'hFD540024 , 32'h0F4A2BE0 , 32'hF3C3A260 , 32'hF63714D0 , 32'h017DB8B0 , 32'h071D44A8 , 32'h01EC89C4 , 32'h1A058AC0 , 32'hF2C7CB30 , 32'hFFF08ACC , 32'h0414EE00 , 32'hF84E4900 , 32'h03A263B4 , 32'h11A817A0 , 32'hF28AF140 , 32'hFA42AFE0 , 32'hF2FBB180 , 32'h04E6F210 , 32'hF3AF94C0 , 32'hF0F87350 , 32'h0D88AF70 , 32'h0210686C , 32'hECDEE820 , 32'h0D3B4B20 , 32'hE9A634C0 , 32'h09AB1360 , 32'h0285F438 , 32'h08CBE6A0 , 32'hF2E735D0 , 32'hF1092F50 , 32'hFCD0F364 , 32'h092BF060 , 32'hFB787DA0 , 32'hF7691370 , 32'hFEC04D2C , 32'h00647D46 , 32'hF8A9DED0 , 32'hFA891548 , 32'h04E20CF8 , 32'hF5F50F00 , 32'hFE98FF9C , 32'hFFFA51B3 , 32'hF803BD58 , 32'hFA08E130 , 32'h0108C02C , 32'hFF9E799C , 32'h0B25BD10 , 32'h047D1938 , 32'hFB94C520 , 32'h030D3E98 , 32'hFD69AE48 , 32'hFC1B6D94 , 32'h02C06C04 , 32'h02223430 , 32'hFAE54D50 , 32'hFFDE4A19 , 32'h000550CD , 32'h0000741D , 32'hFFFE4B94 , 32'hFFFC9075 , 32'h0001B2FB , 32'hFFFEA88B , 32'h00009076 , 32'h0000FDA6 , 32'hFFFF5607 , 32'hFFFD2F0B} , 
{32'h19446420 , 32'hB3F70600 , 32'hF2477160 , 32'h7FFFFFFF , 32'h10E8F340 , 32'h4436D200 , 32'h18840C40 , 32'h97393600 , 32'h4D933E80 , 32'h0E598DB0 , 32'h154A9740 , 32'h381F6D00 , 32'hDD548EC0 , 32'h3695D680 , 32'hDB69BA00 , 32'h06E13550 , 32'h23A2A480 , 32'hD86518C0 , 32'h1FE4BCC0 , 32'h0DCB86A0 , 32'hEC9F2C00 , 32'h27AD4AC0 , 32'hF89B5BC8 , 32'h2522DFC0 , 32'hF0C5BEB0 , 32'h05E34F08 , 32'h25C10900 , 32'h2C6BFF40 , 32'h041D0EC8 , 32'hE3B04A80 , 32'hE15AFF00 , 32'hEB0412E0 , 32'h0067EF87 , 32'h11FF6220 , 32'hEE4742C0 , 32'hE6766000 , 32'hEBD0D740 , 32'hEB993680 , 32'h0ED5DAA0 , 32'hF9D67E30 , 32'h1F44B860 , 32'hF4F5F070 , 32'hF4BC4F60 , 32'h06D63438 , 32'h02BCD308 , 32'hF508ADE0 , 32'hF462A490 , 32'h04E9D110 , 32'hE9170760 , 32'h0FA386B0 , 32'h07999118 , 32'h0BC01D60 , 32'hFB866070 , 32'h00134970 , 32'hF3CF5170 , 32'h08577A90 , 32'h13927F60 , 32'h12F25200 , 32'h0720DA38 , 32'h09796D90 , 32'hFDD748D0 , 32'hFE832614 , 32'hFFE5E23E , 32'h05CBD028 , 32'hEEBC0C60 , 32'h07402238 , 32'h05A2D678 , 32'hF5B30E50 , 32'hFDD65CA4 , 32'h09BE5000 , 32'hFFF2685A , 32'h013292F0 , 32'hFF8EB94C , 32'hFBDBF7D0 , 32'h00E490BE , 32'h01CCCAF4 , 32'h05062FA8 , 32'h093F2530 , 32'hFCBF9B80 , 32'h032EC7AC , 32'hFFA43C89 , 32'h020394D4 , 32'hFFF71BE4 , 32'hFA666BF0 , 32'hFD055CE8 , 32'h02EA1E5C , 32'h04AE4E50 , 32'h018ECE94 , 32'hFFB907B7 , 32'h00BA2BED , 32'h0000C454 , 32'h00042B1F , 32'hFFFFF957 , 32'h00006217 , 32'h00014A43 , 32'hFFFE780E , 32'hFFFF784A , 32'hFFFEB487 , 32'hFFFF784B , 32'h00001335} , 
{32'h00040693 , 32'h00021588 , 32'hFFFAFC6C , 32'h00077C8C , 32'h00031016 , 32'hFFF80F45 , 32'h0001F7A1 , 32'hFFFD2790 , 32'h0006464F , 32'h000431B1 , 32'hFFF690A7 , 32'hFFF6D3FA , 32'hFFF5E4FD , 32'h0001FB69 , 32'h0004C6C2 , 32'hFFFEA531 , 32'hFFFFA2B9 , 32'h00024912 , 32'hFFFEF046 , 32'hFFFD687A , 32'hFFF96A8F , 32'h00032F1B , 32'hFFFAC3E8 , 32'h0002BF16 , 32'hFFFFD14D , 32'h0000E5BE , 32'h0005D13D , 32'hFFFBEE76 , 32'hFFF72543 , 32'h00028E14 , 32'h00011079 , 32'hFFFDEC8B , 32'hFFF704D7 , 32'h00070495 , 32'h0007558C , 32'hFFFB2E1A , 32'h00015C84 , 32'h00040529 , 32'h0000A1F9 , 32'hFFFB817C , 32'hFFFE8A5B , 32'hFFFB71E9 , 32'h00004059 , 32'h00000B97 , 32'hFFFEEBF6 , 32'h000316C0 , 32'hFFFD76B6 , 32'hFFFFC17D , 32'hFFF841F8 , 32'h0000B06F , 32'hFFFE7E16 , 32'h00020306 , 32'hFFFDE4F6 , 32'hFFFA4F7E , 32'h000050B9 , 32'h0002CC16 , 32'h0000B725 , 32'hFFFD6C2C , 32'h00002BCD , 32'h000667C3 , 32'h0002E4F4 , 32'h00039D2A , 32'hFFFF135C , 32'h00035AC8 , 32'h00028573 , 32'h0007590D , 32'hFFFED357 , 32'hFFFD6AF5 , 32'hFFFB67A6 , 32'h00056758 , 32'hFFFBC1F1 , 32'h0004E153 , 32'h00037CBF , 32'h0004E6EF , 32'h0002F3AF , 32'hFFFA45CF , 32'h00038D40 , 32'hFFF9AD5A , 32'hFFF99224 , 32'h000621D9 , 32'hFFFDEE77 , 32'h00062AC4 , 32'hFFFEB60B , 32'h0000EA96 , 32'hFFF54E27 , 32'h00019AEB , 32'hFFFB27AF , 32'hFFFB3FE0 , 32'h00092F21 , 32'hFFFA8964 , 32'h0007ABC3 , 32'h00014524 , 32'hFFFFF08D , 32'h0000F71B , 32'h0000B26A , 32'h0001577B , 32'h0001B2FB , 32'hFFFD5D8A , 32'h0000C449 , 32'h00014A3D} , 
{32'h08C4B860 , 32'h04F388C8 , 32'h3224C680 , 32'hDB2E6780 , 32'hFA8BB408 , 32'hC2F48040 , 32'h0BDF5D50 , 32'hE3608DA0 , 32'hEB930D80 , 32'hF3C1E1A0 , 32'hE75FB260 , 32'hD8818540 , 32'h0093047C , 32'h019CB730 , 32'h05B35480 , 32'h086B2140 , 32'hF52AD3E0 , 32'h0322DD9C , 32'hFA2F3B00 , 32'hF7D21E40 , 32'h1139DB80 , 32'hE3E86740 , 32'hF2A47D60 , 32'h14F2D180 , 32'hD5C15500 , 32'h1E817680 , 32'hE0B26540 , 32'h0EB6EFE0 , 32'h0A29BE50 , 32'h09957690 , 32'hF4110240 , 32'hD0945080 , 32'h06516390 , 32'hF2FBE2C0 , 32'h0EF4B3B0 , 32'h2159B440 , 32'hF8BF2760 , 32'hF84D6A48 , 32'hEE018D80 , 32'hF71F2CC0 , 32'h063630E8 , 32'hF1BD3DF0 , 32'h068CD2D8 , 32'hFE770330 , 32'hFABACAB8 , 32'h0BB39280 , 32'hF1DD3BE0 , 32'hF1E2B760 , 32'hF13CA640 , 32'h14198000 , 32'h1F717720 , 32'h000037E5 , 32'h09A277C0 , 32'h0FC315E0 , 32'h0675EE48 , 32'hFA9CA718 , 32'hF6816050 , 32'hF24E8B20 , 32'hF44413F0 , 32'h08B38390 , 32'hFF0CC688 , 32'hFD524480 , 32'hFF3422DE , 32'hFD7C8504 , 32'hFD27F1E8 , 32'h0C300130 , 32'h0912D170 , 32'h05C969B0 , 32'hF9E9DE80 , 32'hFFC3B9D0 , 32'hFF018C36 , 32'hF6B73E30 , 32'hF669CF70 , 32'h0E0347E0 , 32'h0311F500 , 32'h01AB2FB8 , 32'h00D13D03 , 32'h0621A780 , 32'h08590330 , 32'h021CAF1C , 32'h00CF947E , 32'hFF735C79 , 32'hFEEEE264 , 32'hFA860608 , 32'h072DC3C8 , 32'hFD06469C , 32'hFDF72674 , 32'h00B32F39 , 32'h0178DF20 , 32'hFE9B4BF0 , 32'h0002A399 , 32'h0003B5C3 , 32'h00026A10 , 32'h0000C78C , 32'hFFFBB61A , 32'hFFFDBAA3 , 32'hFFFF155C , 32'h000278FE , 32'hFFFC3A39 , 32'hFFFFB2CF} , 
{32'hF4128CE0 , 32'hFE742F50 , 32'h0716A8B8 , 32'hFC286C7C , 32'hFEF99E04 , 32'hFA4CA098 , 32'h001D53E5 , 32'h02046E5C , 32'h093EC430 , 32'h0246EB5C , 32'hF7F78EE0 , 32'h0B6E19D0 , 32'h09C20370 , 32'hF6D1DF60 , 32'hFFD877AB , 32'hF9DEC1C8 , 32'hF76375A0 , 32'h1D2760C0 , 32'hF685F550 , 32'h0A844D10 , 32'hF6E77F50 , 32'hFDAEDF98 , 32'hFDBF6EC4 , 32'hFBC7A1E0 , 32'hFF85CC3A , 32'h05383058 , 32'h06B75AC0 , 32'h0019489A , 32'h030462B8 , 32'hFB3BC540 , 32'h089D1400 , 32'hFD34ACBC , 32'h04F827C0 , 32'hFD53D334 , 32'h04B045C8 , 32'h011318DC , 32'hFE09A67C , 32'hFFD278D3 , 32'hF6D78D80 , 32'hFE27EC50 , 32'hFA29C740 , 32'h0958B930 , 32'hF2A2A170 , 32'hF94701D8 , 32'hFEA42F64 , 32'h073C04B0 , 32'hF7E3C0E0 , 32'hF41B1650 , 32'h075C4B48 , 32'hFBE0B998 , 32'hFA132A38 , 32'hFBA55C50 , 32'h0071B68F , 32'h03FD1578 , 32'h0F2DB830 , 32'hFB5C2708 , 32'hFCA41758 , 32'h01FAA2D8 , 32'h068939A0 , 32'h04D00888 , 32'hF9F8B058 , 32'hFE3597F8 , 32'h0DF839C0 , 32'hFE625A48 , 32'hF9E038C0 , 32'hFF2D3016 , 32'hFB46E220 , 32'hF4AC83E0 , 32'h08922170 , 32'h029B2D38 , 32'hFF657CAB , 32'hFBD16FC0 , 32'hFE77F844 , 32'h01FDAB6C , 32'hF7EF6110 , 32'hFFF076BC , 32'h06331D40 , 32'hFFFDA335 , 32'hFE266EF8 , 32'hFBE46A70 , 32'h01B66900 , 32'hFBE318B8 , 32'h03DE3C70 , 32'h020CC8E4 , 32'hFB4ED520 , 32'h015AE750 , 32'hFC12D260 , 32'hFC61B0BC , 32'hFEF83A10 , 32'h009F9BC3 , 32'hFFFBA5C0 , 32'hFFFF0C6F , 32'h0004FAF6 , 32'hFFFAAD49 , 32'h0007D122 , 32'h0001DDF5 , 32'hFFFD5FA0 , 32'hFFFC1897 , 32'h00047DB5 , 32'hFFF98A80} , 
{32'hFFFE6683 , 32'h0005C7CA , 32'hFFF8F5BE , 32'hFFFE4E0B , 32'hFFFBF957 , 32'hFFFFB271 , 32'h00009490 , 32'h0008CF2B , 32'h000332F9 , 32'hFFFA18D1 , 32'h0001E7F6 , 32'hFFFBA8A9 , 32'hFFF93B58 , 32'h0001FB49 , 32'h00023978 , 32'hFFFC423A , 32'h00010C4C , 32'hFFF934DE , 32'h0000E7DB , 32'hFFFC39D0 , 32'hFFF7F226 , 32'hFFFC8C74 , 32'h00065027 , 32'h0001E1C3 , 32'hFFF6BAA9 , 32'hFFFD623E , 32'h00005732 , 32'hFFFCDF77 , 32'hFFFB8FEA , 32'h0005491B , 32'h0000A62A , 32'h000251B8 , 32'h00068002 , 32'hFFFC8E31 , 32'hFFFE4E65 , 32'hFFFCCBC4 , 32'hFFFE1DF9 , 32'hFFFC6727 , 32'hFFFD0503 , 32'h00033F3D , 32'h00064B58 , 32'h00010718 , 32'hFFFDE4FE , 32'hFFFE8A98 , 32'h000809E3 , 32'h00041F02 , 32'h000003E5 , 32'hFFF95B12 , 32'h00005872 , 32'h000507ED , 32'hFFFE3587 , 32'h00025A64 , 32'h0002D913 , 32'hFFF47F6B , 32'hFFFAB988 , 32'h0001922B , 32'hFFFEA2CE , 32'h0000215C , 32'h00007C99 , 32'hFFF90951 , 32'h0007F726 , 32'hFFF8A4BB , 32'hFFFB4036 , 32'hFFFF84BB , 32'h000A7383 , 32'h000246FD , 32'h000225F8 , 32'h000093A1 , 32'hFFFF8F6C , 32'hFFFBE32E , 32'hFFF9FEB9 , 32'h000280C5 , 32'hFFFAF06E , 32'h0003A71C , 32'hFFFFECF3 , 32'h0003F25E , 32'h00019F85 , 32'hFFF8A9C5 , 32'h00038DE8 , 32'h0002094A , 32'h0005E11A , 32'hFFF88F3E , 32'hFFFED7D9 , 32'hFFFC35E8 , 32'h00033AE5 , 32'hFFFD5065 , 32'h00019147 , 32'hFFF4CC66 , 32'hFFFD8D5C , 32'h0008EB4F , 32'h00050038 , 32'hFFFECBD8 , 32'hFFFC0B70 , 32'hFFFE8D6A , 32'hFFFE69A2 , 32'h00003B06 , 32'h0000B230 , 32'h0003C2D9 , 32'hFFFC2A8B , 32'hFFFEE485} , 
{32'h136EC3A0 , 32'hE7E87000 , 32'h14BC7000 , 32'hF144F710 , 32'h3336F040 , 32'h05A7F9A0 , 32'hE37C43C0 , 32'h32FBD6C0 , 32'hF87E3848 , 32'hFC0D793C , 32'h088831A0 , 32'hEA5D1780 , 32'hFEFC5944 , 32'h0AAEEB50 , 32'hF9654990 , 32'hE0D9CC80 , 32'h04E83248 , 32'h1C7E4BE0 , 32'h03DCAFD0 , 32'h03E027C4 , 32'h09E97FE0 , 32'hE3DD0E40 , 32'h0BB6DE20 , 32'hFD9FB27C , 32'hFA252CB8 , 32'hE7631840 , 32'hE08C36E0 , 32'h34CF3640 , 32'h03FC2580 , 32'hE25786A0 , 32'h053AEF18 , 32'h006554E5 , 32'h0297C048 , 32'h12AC8FC0 , 32'hFEF60784 , 32'h0FFAE9A0 , 32'h19325020 , 32'h09960360 , 32'h07DC3788 , 32'hF7F8EEE0 , 32'h000D4E94 , 32'hFAFA8668 , 32'hFEBF5D14 , 32'h05E4CAA0 , 32'h038DE884 , 32'h03FECCB0 , 32'hFCA39E7C , 32'hF2C7C1A0 , 32'h0402CA18 , 32'hEC53F320 , 32'hFA09C060 , 32'hEE8B9520 , 32'h0D960870 , 32'h0D3EB900 , 32'h061E1DE0 , 32'hEF897C80 , 32'h0C3AE240 , 32'hF778ACD0 , 32'h03556C6C , 32'hF9FCE590 , 32'h0111E74C , 32'hE3187B40 , 32'hF8A70448 , 32'hFFD7A54F , 32'h123669C0 , 32'hFF2DFF34 , 32'h02AF6F08 , 32'hFEDD29AC , 32'hF8056848 , 32'hF5343B90 , 32'h0745CFA8 , 32'hFE5C6744 , 32'hF9D8B780 , 32'hFC196E44 , 32'h0D1FD290 , 32'hF9D3A7E0 , 32'h055F2780 , 32'hFE984444 , 32'h07535D88 , 32'h03CF804C , 32'hFBD1AC30 , 32'h0AFFACB0 , 32'hFAA98AE0 , 32'h096EB230 , 32'hFCFC3280 , 32'h00325F97 , 32'h01D958BC , 32'h0376DA38 , 32'h0060B475 , 32'h00E21A45 , 32'hFFFD71EF , 32'h0001F6FE , 32'h0000AEDB , 32'h00029023 , 32'h0000EFA9 , 32'hFFFCD131 , 32'hFFFD5285 , 32'hFFFD97D7 , 32'hFFFFB7B8 , 32'hFFFDE197} , 
{32'hFFFEEA62 , 32'h00021E37 , 32'hFFFB8D0C , 32'h0002C485 , 32'h00018993 , 32'hFFFFAD68 , 32'h00008860 , 32'hFFFA4B12 , 32'hFFF54260 , 32'h0000795B , 32'hFFFDE6C7 , 32'hFFFA98FF , 32'h00000519 , 32'hFFF8E5F4 , 32'h0002DDA7 , 32'h0002AA83 , 32'h00044795 , 32'hFFFC1EB8 , 32'h00021201 , 32'hFFFFD2D7 , 32'h000237A7 , 32'hFFFF72F3 , 32'hFFFD9532 , 32'hFFFF0FE5 , 32'hFFF9F379 , 32'hFFFC2F6C , 32'hFFFEB703 , 32'hFFFFA14D , 32'hFFFC3894 , 32'hFFFB7748 , 32'h000A43FF , 32'hFFFF08E3 , 32'h0005331C , 32'hFFFD7184 , 32'hFFFC5DC6 , 32'hFFFB5910 , 32'h000246CB , 32'h000130F2 , 32'hFFFE0FDC , 32'h00045244 , 32'h0003CBFC , 32'hFFFCE67A , 32'h00016ED8 , 32'hFFFD89B5 , 32'hFFFEC025 , 32'hFFFD056E , 32'h0006035E , 32'h0001391F , 32'hFFFE957F , 32'hFFF43359 , 32'h00006F57 , 32'hFFFF7177 , 32'hFFF885F9 , 32'hFFFF89A1 , 32'h000266DD , 32'hFFF5A664 , 32'hFFF65407 , 32'hFFFF1ACA , 32'h0001A631 , 32'hFFFDDE32 , 32'h000532F9 , 32'h000D41D8 , 32'h000667AC , 32'h0004FCC5 , 32'hFFFCFC74 , 32'h0002E1FB , 32'h0001B715 , 32'hFFF8B431 , 32'h000147E7 , 32'hFFFEA756 , 32'hFFFE870F , 32'h0006519F , 32'hFFFF30EF , 32'h0001F452 , 32'h00034689 , 32'h00018A64 , 32'hFFFE733F , 32'hFFFB793E , 32'hFFF3DC7D , 32'hFFFF7619 , 32'hFFFEC4CD , 32'h0001A640 , 32'hFFF6EAA9 , 32'hFFFEBF74 , 32'h00046E24 , 32'hFFF95F49 , 32'h0006B1B7 , 32'h0009FF4A , 32'h00032003 , 32'hFFFBD749 , 32'h0001AE05 , 32'hFFFDE1E5 , 32'hFFF8D325 , 32'h00015280 , 32'hFFFBBD62 , 32'hFFFFB986 , 32'hFFFCFA15 , 32'hFFF70068 , 32'h00026F50 , 32'hFFFF8E94} , 
{32'h03733D94 , 32'hF9337868 , 32'h0DC59EA0 , 32'hF858AD70 , 32'hFE229DE8 , 32'h0E8234F0 , 32'h020DFB74 , 32'hFDE7D218 , 32'h03E6A188 , 32'hFECE490C , 32'hECC601C0 , 32'h03002030 , 32'hF645DD70 , 32'hF15A7230 , 32'hEF70FB60 , 32'h019851B8 , 32'hFF863330 , 32'hFE428A34 , 32'hFA10CDF8 , 32'hFE388BE0 , 32'hF87561D0 , 32'hF71F6E60 , 32'hFBF5D358 , 32'h0813A5E0 , 32'hF4F7F310 , 32'h04647668 , 32'hFB67BA20 , 32'hF4469D10 , 32'h044410F0 , 32'hF67DCA60 , 32'h0317B3A8 , 32'h04ADDC70 , 32'h040BF548 , 32'h0338BFEC , 32'h0E0F4770 , 32'hF62A5FC0 , 32'hF92FB8E8 , 32'h0410CEC0 , 32'hFC7AF884 , 32'hFD4E6C9C , 32'hFE0100B0 , 32'h05929B18 , 32'h071005A8 , 32'h108C1620 , 32'hFDCA5F74 , 32'h01CDC7EC , 32'h03AAF864 , 32'h006428A0 , 32'h02DCD28C , 32'hFD79D254 , 32'hFE1B2238 , 32'h0A6307D0 , 32'hFFEEA503 , 32'hFE56E8AC , 32'hFD9E0F00 , 32'hFA78F0D0 , 32'h0F287CB0 , 32'hF5EDE980 , 32'hFAD79CD8 , 32'h0978D2B0 , 32'h0836DFA0 , 32'h043D1B70 , 32'hFA21AD18 , 32'h0DF17BE0 , 32'h03E7DD80 , 32'hF37AA8C0 , 32'hFCD0A39C , 32'hF3EAE530 , 32'hF64383F0 , 32'hFE4D663C , 32'h021047C8 , 32'hF6D40B80 , 32'h020FADBC , 32'hF84B04D8 , 32'hFD89CA34 , 32'hFC49AA0C , 32'hFB8A2880 , 32'hFCEEF2EC , 32'hFC07D80C , 32'h012EAF2C , 32'hF78E7A70 , 32'hFAA6F0C8 , 32'h00E4D87B , 32'hF9959930 , 32'hFE357414 , 32'h075C30B8 , 32'h00820DD0 , 32'h072DBD68 , 32'hFF020A96 , 32'h00FBC741 , 32'hFFFBDF04 , 32'hFFFB0452 , 32'hFFFDD3AF , 32'h0006D48C , 32'h00011935 , 32'hFFFD0754 , 32'h0000BD36 , 32'hFFFCF1C5 , 32'hFFFD119E , 32'hFFFFF77D} , 
{32'h4FF53400 , 32'hD9D3BD40 , 32'h6DA85880 , 32'h04C81B80 , 32'h26527300 , 32'h42446180 , 32'h26307F00 , 32'h026BB2C8 , 32'h1531EAE0 , 32'h1C271940 , 32'hA4BCF680 , 32'h24A1A640 , 32'hFBC0EAE8 , 32'h1E225960 , 32'h21D2E900 , 32'h1048E8E0 , 32'hE709F480 , 32'hE171BB00 , 32'hDC486A00 , 32'h1A5BF180 , 32'hF0AA3330 , 32'hF091C500 , 32'h0BD12CE0 , 32'hEAC9ED40 , 32'h2EEEB900 , 32'hF0922C00 , 32'h0A597820 , 32'hEA1BA8A0 , 32'hD49C7EC0 , 32'hF83C4830 , 32'hE8EBE0E0 , 32'hFB2360A0 , 32'h16822340 , 32'h0E002A60 , 32'h0EB822A0 , 32'h17DB35E0 , 32'h06DEB210 , 32'hE1D27DA0 , 32'hFB41A9E0 , 32'h02620AC8 , 32'hF8DC1200 , 32'h0E346B20 , 32'h095F7F60 , 32'h0373F2C0 , 32'hF050B590 , 32'h013B21E8 , 32'hF55C9130 , 32'h14EC0F00 , 32'h0F9FBB40 , 32'h0F923FA0 , 32'hF36C5270 , 32'hFF2B094A , 32'h064BEF40 , 32'h0DC80270 , 32'hF40A19C0 , 32'hEAA9E260 , 32'h162892A0 , 32'hE52B18A0 , 32'hFB0348C8 , 32'hFF565F8C , 32'h024010D8 , 32'hF5567690 , 32'h16A994E0 , 32'h06A628A8 , 32'hFBF02728 , 32'hFAC9DBA8 , 32'hF8985E60 , 32'hF9309E60 , 32'h02792C68 , 32'h04CC87C0 , 32'hFF222E6C , 32'hF90701C0 , 32'h03037710 , 32'h0A22EC90 , 32'hFE264640 , 32'hF9158CA0 , 32'h011B789C , 32'hFCA7A398 , 32'hFA7CE078 , 32'h076C52F0 , 32'hFF170526 , 32'hF8E262B8 , 32'h041DF388 , 32'hF82CD3B8 , 32'h03899E10 , 32'h05504F68 , 32'hFDD0F598 , 32'hFD34E82C , 32'hFD33628C , 32'hFF48B06D , 32'h00021FED , 32'h000143C9 , 32'h00017647 , 32'hFFFC7252 , 32'h00005446 , 32'h0001A080 , 32'h0002378B , 32'hFFFD2A64 , 32'hFFFFB871 , 32'hFFFF2B53} , 
{32'h73917E80 , 32'h276F4B40 , 32'h1BB00BE0 , 32'h0E7292A0 , 32'h0CAF5E60 , 32'h3735F880 , 32'hD5E57180 , 32'hEF373D40 , 32'h19552600 , 32'h0B54D0D0 , 32'h04BECBB0 , 32'hECC66180 , 32'hFAA43B40 , 32'hEBF4DD00 , 32'h08E068B0 , 32'h10923820 , 32'h19B13F40 , 32'hFD5A85AC , 32'h2DE7E780 , 32'h094E6440 , 32'h189D7D00 , 32'h0642F9F0 , 32'h034FBEE8 , 32'h0EEBF010 , 32'h0B27CB80 , 32'hE5E036E0 , 32'h12BB7BC0 , 32'hDEC198C0 , 32'h0D4C74A0 , 32'h0C111C90 , 32'hE0BE8740 , 32'hE7537F00 , 32'hF359CB10 , 32'hF1848110 , 32'hE14F2960 , 32'hFBEFEFF0 , 32'hF9C2BC98 , 32'h06B64498 , 32'hEF4D6B00 , 32'hE9620660 , 32'hFEA45BCC , 32'hF9D7B9A0 , 32'h06295690 , 32'hEEF15F20 , 32'hF86ECB60 , 32'h04AAF8A8 , 32'hF93782D0 , 32'h172DEF00 , 32'hEB73FEA0 , 32'hF7456D40 , 32'h045388A8 , 32'hF9518250 , 32'hF09B1DF0 , 32'hF05FDF50 , 32'h020EF23C , 32'h138C9AC0 , 32'h0AF04340 , 32'hFF526171 , 32'h0D564880 , 32'hF0EC77E0 , 32'h17B4AA60 , 32'hF330F670 , 32'h04A54040 , 32'h00308901 , 32'h0D0C0EE0 , 32'hFE55CA64 , 32'hFDF015E8 , 32'h06611FD8 , 32'hF918A090 , 32'h039E20AC , 32'h059F50D0 , 32'h0303EA64 , 32'h07557F98 , 32'h0600B230 , 32'h058219F0 , 32'h0B4C7950 , 32'hFCC6A59C , 32'h05E2FE08 , 32'h035E6CC0 , 32'h0629B0B0 , 32'hFBA65760 , 32'h00E935AA , 32'hFE7A0E08 , 32'hFF74D67D , 32'hFAF81A48 , 32'hFC70F210 , 32'hF6125B20 , 32'h057FD468 , 32'hFEF5C118 , 32'hFE930D10 , 32'hFFFD92E2 , 32'hFFFED2BF , 32'h000216F1 , 32'hFFFFE6CC , 32'hFFFD9D20 , 32'h0001161D , 32'hFFFEA72F , 32'hFFFCDD6D , 32'h0002ED86 , 32'hFFFDB2FF} , 
{32'hFFFA2572 , 32'h00047633 , 32'hFFFC27F1 , 32'h000261B1 , 32'hFFFAC783 , 32'hFFFF4E21 , 32'h0000369C , 32'h000327E4 , 32'h00046212 , 32'h0008834D , 32'h000012C3 , 32'h0003F017 , 32'hFFFDA625 , 32'h0008C73F , 32'h0006154E , 32'hFFFF5888 , 32'h0000D549 , 32'hFFFB6174 , 32'hFFFE1E69 , 32'h000851F4 , 32'hFFFE036B , 32'h000580EC , 32'hFFFDC53C , 32'hFFFBF461 , 32'h00007503 , 32'hFFF858F1 , 32'hFFFA493E , 32'hFFF928B3 , 32'hFFFA963A , 32'h0003D34D , 32'hFFF8B32A , 32'hFFFEF5C1 , 32'hFFF74076 , 32'h0002640D , 32'hFFFBDDE9 , 32'h0000FBD0 , 32'hFFFDDA2F , 32'h0000FF34 , 32'hFFFC058E , 32'h00008BC4 , 32'h0003F0D9 , 32'h0000D421 , 32'hFFFA3CD9 , 32'h00051B80 , 32'hFFFD60A3 , 32'hFFFC4822 , 32'h0002BEF6 , 32'h000732C8 , 32'h0001A625 , 32'h000A1411 , 32'h0004C2D7 , 32'hFFF19CBA , 32'hFFFE920F , 32'hFFF4229C , 32'hFFFB452B , 32'h0008FF82 , 32'hFFFE7DC7 , 32'h0003FEC1 , 32'hFFF9C59F , 32'h000232FB , 32'hFFFEDDA9 , 32'hFFFC607D , 32'h00063262 , 32'hFFFE571F , 32'hFFFCEAB1 , 32'hFFFB8440 , 32'hFFF8E739 , 32'h000389A1 , 32'hFFFF5FEB , 32'h0004BF7C , 32'h000505D6 , 32'h000801A8 , 32'h00015C6D , 32'hFFFC2E20 , 32'hFFFD614B , 32'hFFF79DCF , 32'h0002CEA5 , 32'hFFFFC60F , 32'hFFFC21B9 , 32'hFFFB3173 , 32'hFFF97DFD , 32'h00058905 , 32'h00097C4F , 32'hFFFEC994 , 32'h000220D2 , 32'hFFFE7699 , 32'hFFFB7736 , 32'hFFFFC6B5 , 32'hFFFB0A25 , 32'hFFF90341 , 32'hFFFD2AF4 , 32'h0005F2F7 , 32'hFFF61C49 , 32'hFFFB2787 , 32'h0002B483 , 32'h00021C30 , 32'h0002C114 , 32'h0001FCFD , 32'h0000534D , 32'hFFFA4BFF} , 
{32'h0004DD42 , 32'h000462EF , 32'hFFF9037C , 32'hFFFD293F , 32'hFFF5B323 , 32'hFFFF3F39 , 32'h00022351 , 32'hFFF7635F , 32'h0002C4D9 , 32'h000548CD , 32'hFFFC3EF6 , 32'h000A0DE3 , 32'h00062906 , 32'hFFFE4442 , 32'hFFFB894E , 32'hFFFC4210 , 32'h00035190 , 32'hFFFE2215 , 32'h00035388 , 32'h000317B9 , 32'hFFFC79C9 , 32'hFFFE0B9D , 32'hFFFE700B , 32'hFFF477D1 , 32'hFFFE6436 , 32'hFFFD1542 , 32'hFFF88DC5 , 32'hFFFF5718 , 32'h000678FD , 32'hFFFF1992 , 32'h0004BB86 , 32'h00060F4C , 32'hFFFBE1EC , 32'h00085D0F , 32'hFFF9FBFE , 32'hFFF7CC07 , 32'h00012504 , 32'hFFFF5C4C , 32'h000507B6 , 32'h00048152 , 32'h0000A304 , 32'h0003D0E8 , 32'hFFFFDA9D , 32'h00096B61 , 32'h000468B7 , 32'h0002A3AE , 32'h0000F0CA , 32'h000196E8 , 32'hFFF678EE , 32'h000153C4 , 32'hFFFAC67F , 32'h0003B194 , 32'h00025782 , 32'hFFF9885E , 32'hFFFCC10F , 32'h0003FE6F , 32'h00051FAC , 32'h0001EA5F , 32'h00073FD2 , 32'hFFFAF1AC , 32'hFFFB2620 , 32'hFFFFCFB3 , 32'h0000DA6F , 32'hFFFD7611 , 32'hFFFEC706 , 32'hFFFF6ACE , 32'hFFFBBFFE , 32'hFFFDCBE6 , 32'h0001CB61 , 32'hFFFF88DB , 32'hFFFAE981 , 32'hFFFF853B , 32'h000D217C , 32'h0000EABD , 32'h0004FDAA , 32'h00002156 , 32'hFFFC5848 , 32'hFFFA35C3 , 32'hFFFE0C63 , 32'hFFFCC237 , 32'h0002BAAF , 32'h0004E2EC , 32'h0004C986 , 32'h00040E05 , 32'hFFFA118F , 32'h00024BC7 , 32'hFFFFBF69 , 32'h00023CFE , 32'hFFFF7C8F , 32'hFFFA6F0E , 32'hFFFE3DBE , 32'h0000EE91 , 32'hFFFB7792 , 32'h00017317 , 32'hFFFDC42A , 32'hFFFBDEA9 , 32'hFFF9F7D8 , 32'h00000F52 , 32'h000159F5 , 32'hFFFC0FDC} , 
{32'hA8645580 , 32'h22BD5540 , 32'h2CDB63C0 , 32'hFEEC2FF8 , 32'h0B0B0070 , 32'h21CBDA80 , 32'hF244E180 , 32'hED11A4E0 , 32'hC38D3240 , 32'h0450D1C0 , 32'hE1376FC0 , 32'hD59169C0 , 32'h0C9EB990 , 32'h3D69E380 , 32'h01A8E768 , 32'h06A692D0 , 32'hF4AE4300 , 32'hFC5A40A4 , 32'hF58AE360 , 32'h1BF1CD20 , 32'h15D7B520 , 32'h09081BC0 , 32'hFE5D7174 , 32'h12371A20 , 32'h06905988 , 32'hD8766980 , 32'hE3D4B980 , 32'hEC144540 , 32'h043E1680 , 32'h053575C0 , 32'hF5B3CF90 , 32'hE53BD5A0 , 32'hE1387AA0 , 32'h077A2C50 , 32'hE67D71A0 , 32'h126EE5E0 , 32'h1419FEC0 , 32'hE3DB2100 , 32'hF0F7F770 , 32'hE8465640 , 32'h0B853C70 , 32'h1A663700 , 32'h0D911DE0 , 32'h0B3C6BD0 , 32'h0BD23B60 , 32'hF08842D0 , 32'h043E3908 , 32'hE4CC48A0 , 32'h07BAB708 , 32'h0F15F4F0 , 32'h01404CE8 , 32'h1BB17000 , 32'hFD96B588 , 32'h053874B8 , 32'h044695A8 , 32'hFC626DE8 , 32'hFFE62E48 , 32'h02674FD4 , 32'h0D09B8A0 , 32'hFA321690 , 32'hFA2F5060 , 32'hFA20DCB8 , 32'hF244AA30 , 32'hF531E730 , 32'hF4A7B670 , 32'h063FF160 , 32'h007A2855 , 32'hFC9E3EA8 , 32'hF5744280 , 32'h06511790 , 32'hF0918720 , 32'h087B3DD0 , 32'h0DCC2790 , 32'hFEC7C22C , 32'hFBE70750 , 32'h0885B7D0 , 32'h0B411630 , 32'h09013BA0 , 32'h0ADE2E50 , 32'hFECD3CAC , 32'h02373CF4 , 32'hF3A70990 , 32'h0120ADB0 , 32'h0581B208 , 32'hF8C1A3D0 , 32'h011AF658 , 32'h00519AC6 , 32'h06678DF0 , 32'h00A1DB48 , 32'h0190E700 , 32'h0002E030 , 32'hFFFF4632 , 32'hFFFEC77B , 32'h0005F28E , 32'hFFFFFA44 , 32'hFFFF5EF8 , 32'h0001C257 , 32'h00037059 , 32'hFFFC3B34 , 32'h00009909} , 
{32'h0005DD36 , 32'h00032C57 , 32'h000128B2 , 32'hFFFCC811 , 32'hFFFACB19 , 32'h000718CC , 32'h000354CF , 32'h00035E8F , 32'hFFFCD9E2 , 32'hFFFACDF4 , 32'h0006318F , 32'hFFFF29A5 , 32'hFFFF6042 , 32'h00025FB0 , 32'hFFFF0739 , 32'h0006EB99 , 32'h000412B2 , 32'hFFFF80A3 , 32'hFFFC71D1 , 32'hFFFA5E4C , 32'h00023CA3 , 32'h0001F633 , 32'h00042F7B , 32'h000270C0 , 32'h0000778C , 32'h000903AA , 32'h0006F0A9 , 32'h00076649 , 32'hFFFB27AB , 32'h0007FD76 , 32'hFFF3BB13 , 32'h000348F5 , 32'h0001B4C9 , 32'hFFFEB2AD , 32'hFFFD6BD0 , 32'h00078E21 , 32'hFFFCC23E , 32'hFFFB826C , 32'hFFFE8B0A , 32'h0002394B , 32'hFFFDC14A , 32'hFFFA768C , 32'h0001063E , 32'h0006AF3A , 32'hFFFD3FB8 , 32'hFFFDE0A6 , 32'hFFFE0CBE , 32'hFFFB33A0 , 32'h0002B3EC , 32'hFFFFDA06 , 32'h0005B8BD , 32'h00034C7B , 32'h000889D5 , 32'h0003718E , 32'h000218F3 , 32'hFFFB05E5 , 32'hFFFAFC72 , 32'h000A4E1C , 32'hFFFD561C , 32'hFFFD939C , 32'h000216EC , 32'hFFFCCFE8 , 32'h0004887E , 32'hFFF976BD , 32'hFFFBD558 , 32'hFFFBCB2C , 32'hFFFA4A5B , 32'hFFFC51F1 , 32'h000514B1 , 32'h0009E03A , 32'hFFFE6A76 , 32'h0001F816 , 32'h0000909E , 32'h0000795A , 32'hFFFEB239 , 32'hFFFD11FF , 32'hFFF9F249 , 32'h000000D0 , 32'h00037862 , 32'h0001FD46 , 32'h00076E62 , 32'hFFFE0080 , 32'h0000B987 , 32'h00022585 , 32'h000904F2 , 32'hFFFD3ECB , 32'hFFF9584D , 32'hFFFA56EA , 32'h000559EC , 32'hFFFA7409 , 32'h000112C4 , 32'h00055E2A , 32'h0007A019 , 32'hFFFFAE81 , 32'hFFFCC827 , 32'h000145CC , 32'hFFF9385E , 32'hFFFB0FA0 , 32'h000589DA , 32'h00050C6C} , 
{32'h5B7E8A80 , 32'h076889B0 , 32'hF0D270A0 , 32'h32122040 , 32'h2C97C300 , 32'h104DD720 , 32'hF2250900 , 32'hE004A5A0 , 32'hDD10C340 , 32'h0B968720 , 32'hE4D18D40 , 32'h24095480 , 32'h2F16B300 , 32'h1102AC60 , 32'h1F4806E0 , 32'hFDB2BEF8 , 32'h0AB66750 , 32'hFF2EFDEC , 32'hE5B0DDE0 , 32'h13CC4B80 , 32'hFF43C3F7 , 32'hEC3F0100 , 32'hDBB93180 , 32'hDBC6E680 , 32'hF4EF4CC0 , 32'hE411C760 , 32'hFC831A98 , 32'hDAE9C740 , 32'h36B93840 , 32'hF8CCEAB0 , 32'h2F671FC0 , 32'h13B43B80 , 32'h15398080 , 32'hFE37E51C , 32'hD4F53840 , 32'hE4586140 , 32'hDD891380 , 32'hF796C140 , 32'hEA5D9180 , 32'h02A72E28 , 32'h007D8F3E , 32'hF9CE0068 , 32'hEB35DA20 , 32'hF8F42FF0 , 32'hDD22A7C0 , 32'h0983F410 , 32'h0576CAF0 , 32'hEF9AA820 , 32'hEF568940 , 32'h00496C33 , 32'h08A886A0 , 32'h03B4128C , 32'h0E3F3A30 , 32'h0D17C330 , 32'hF57C2C70 , 32'h0A831890 , 32'hF29431E0 , 32'h07818490 , 32'hFF0C0E76 , 32'hFDB8E804 , 32'hEF742840 , 32'hFAE2E5E0 , 32'hF9FE08C0 , 32'h0D5AF710 , 32'h0E50F530 , 32'h0D2AAD20 , 32'hFFC95993 , 32'h0D7B90A0 , 32'h03409A98 , 32'h04247898 , 32'h0F1583D0 , 32'h0E8C95D0 , 32'hFE14E0F4 , 32'hFB3D8D00 , 32'h000934F2 , 32'hFF5FF773 , 32'hFFE49EE3 , 32'h01240090 , 32'h00CC2B27 , 32'h05B28208 , 32'hF8A329E0 , 32'hFFF99AE6 , 32'hF9EF9018 , 32'h08300E80 , 32'h022C5E78 , 32'h01319678 , 32'hFDB7BA4C , 32'hFCA22F5C , 32'hFCC69E80 , 32'hFFFC7319 , 32'h00058D61 , 32'hFFFE47AC , 32'hFFFEC129 , 32'h0002D353 , 32'h0001C325 , 32'h00009A63 , 32'h0000F777 , 32'h0004AC65 , 32'h00007D3B , 32'hFFFF4798} , 
{32'h000574ED , 32'hFFFCF5E0 , 32'h000094A7 , 32'hFFFF1752 , 32'h00004E80 , 32'hFFFB4183 , 32'h00015D9C , 32'hFFFF1967 , 32'h00001FA2 , 32'h0001F2CD , 32'hFFFEDFDB , 32'h0001A516 , 32'hFFFC708E , 32'h00079D0F , 32'h00033016 , 32'h00090B6F , 32'hFFFC4F7E , 32'h00058835 , 32'h00058753 , 32'hFFFEBDA6 , 32'h00020AB2 , 32'hFFFDE757 , 32'h0002AB1B , 32'h0005FB2D , 32'hFFF6804C , 32'h000137CC , 32'h00004442 , 32'h00064F6F , 32'h0001D4B2 , 32'hFFF93803 , 32'h00024B8D , 32'hFFF6141E , 32'h000601FB , 32'h000238D5 , 32'h0000D4FA , 32'h000DC4E0 , 32'h0002CEB8 , 32'h00058318 , 32'hFFF91545 , 32'hFFFCD051 , 32'h0005A1F4 , 32'hFFFEDF43 , 32'h000009CD , 32'hFFFA7E9B , 32'hFFFAFD46 , 32'h00087F67 , 32'h00060288 , 32'h000227F3 , 32'hFFFA047B , 32'h0000AF6E , 32'h00003EFD , 32'hFFF7DD4D , 32'h00005922 , 32'hFFFFA3C7 , 32'hFFFA4A7C , 32'hFFFFBCC2 , 32'h0007520D , 32'hFFFF0620 , 32'h00046C93 , 32'hFFF7874D , 32'hFFF6CBDE , 32'h00033ACB , 32'hFFFB0FF4 , 32'hFFFAC631 , 32'h000190A0 , 32'h00083946 , 32'h0002EBD8 , 32'hFFF159CE , 32'h000762C4 , 32'h000709BF , 32'h0002926E , 32'h00005DBC , 32'hFFFDAF0B , 32'hFFFC1DDF , 32'hFFFDE5F7 , 32'h00002F48 , 32'h000632E8 , 32'hFFFFA4DA , 32'hFFFDEF80 , 32'hFFF38B1F , 32'h0004312A , 32'h00015D7E , 32'hFFFEEC87 , 32'h0002FF35 , 32'h000698E8 , 32'hFFFBCADF , 32'h0009486A , 32'h0000AE08 , 32'h0001395B , 32'hFFFF32C2 , 32'h0000F1FE , 32'h0002AD9F , 32'hFFFB2FFE , 32'h00015EFC , 32'hFFFDC283 , 32'h00089C45 , 32'h000725ED , 32'h00009419 , 32'h000A2867 , 32'h000099D4} , 
{32'hFF0C5781 , 32'h05767DD0 , 32'hFFBA4057 , 32'h042EA0C8 , 32'hFCD65AE0 , 32'h0AEA7DD0 , 32'hFD883F14 , 32'h085BB030 , 32'h0182A55C , 32'hFBD2C158 , 32'h0A4F5B60 , 32'h05518D08 , 32'h0B5BDA20 , 32'h06587518 , 32'hFF6E9041 , 32'h068D3B88 , 32'h0500B890 , 32'hFC875E34 , 32'hFB6075B8 , 32'h06E126F0 , 32'hFD047E54 , 32'h03DF21D4 , 32'h065CB200 , 32'h033BAF9C , 32'h0A6A9F70 , 32'hFA8BDD58 , 32'h04FBDD40 , 32'h08D5FD50 , 32'hFF1BBF73 , 32'hFCAB78E4 , 32'hFA3613A0 , 32'h033A71A0 , 32'h027B17F8 , 32'hF388F6F0 , 32'hFDE5A7C0 , 32'h024E2FB4 , 32'h05338220 , 32'h017FE2A0 , 32'h06865E18 , 32'h046AECD0 , 32'h01AA9C9C , 32'hFDA314E0 , 32'hFE7C0770 , 32'hFA0165D0 , 32'h00A2FA36 , 32'h0474FC98 , 32'hFFC8446D , 32'h04A7ACF8 , 32'hFF54D7FD , 32'h03F19F0C , 32'hFAB43058 , 32'hFD7C6528 , 32'h048A4270 , 32'h034388F0 , 32'hFCAB1E24 , 32'h07711B90 , 32'hFE2E4AEC , 32'h014996DC , 32'h00E28715 , 32'hF8B8D5D8 , 32'hF8C8F828 , 32'h03B6ACCC , 32'h036AB788 , 32'h05354EC0 , 32'h067DB3D8 , 32'h03554A24 , 32'hFF065B43 , 32'hFB35E1A0 , 32'h068B95E0 , 32'h02995190 , 32'hFD896ECC , 32'h02846B4C , 32'hFEF9A6DC , 32'hF762D380 , 32'hFCE92938 , 32'hFF95008F , 32'h02E2E46C , 32'h0043DEBD , 32'hFED80008 , 32'hFE85CBF8 , 32'h041930D0 , 32'hF9AA3018 , 32'h04749928 , 32'h004D555E , 32'h0604EA78 , 32'hFE6777B0 , 32'hFFA99F76 , 32'hFE5CED54 , 32'h0091411D , 32'h0089D977 , 32'hFFFBDCAA , 32'hFFFE3123 , 32'hFFFEF82D , 32'hFFFDA88E , 32'h0001526E , 32'h00060638 , 32'hFFFA8DE2 , 32'h0004F668 , 32'hFFFFCEEA , 32'hFFFC6A8C} , 
{32'h0000D5DD , 32'hFFF8DAF1 , 32'hFFF87C3B , 32'h0005ACEC , 32'h0003268C , 32'hFFFCA0A5 , 32'h0007A82B , 32'h000061A2 , 32'h0001195B , 32'hFFFC6CCA , 32'h00007236 , 32'h00094310 , 32'hFFFF08AB , 32'h0002171D , 32'hFFFE9E79 , 32'h0001BEA8 , 32'h000527A1 , 32'hFFFE4C89 , 32'hFFFBB73F , 32'h00026130 , 32'h00007FE4 , 32'h0001E5B5 , 32'h00030571 , 32'hFFFF4A1C , 32'h00048380 , 32'hFFFC472C , 32'hFFFF455B , 32'h0006300C , 32'h00059EAE , 32'h0003E619 , 32'h000202F5 , 32'hFFF9B47E , 32'hFFF9015E , 32'h00055293 , 32'hFFF7F99E , 32'h0002C205 , 32'hFFFF1ED9 , 32'hFFF91702 , 32'hFFFFD206 , 32'h0002EDC1 , 32'hFFF650EC , 32'h00041873 , 32'hFFFC0409 , 32'h0007198C , 32'hFFFD01E5 , 32'hFFFC64A1 , 32'hFFFA3E3B , 32'hFFFBFB81 , 32'hFFFC414F , 32'h00014FDC , 32'hFFFF8436 , 32'h00077036 , 32'hFFFFD497 , 32'h000AE9EC , 32'hFFFDC05B , 32'hFFFD9D91 , 32'h00045B74 , 32'hFFFF1A27 , 32'hFFFD7C61 , 32'hFFFFA9CD , 32'hFFFF52C0 , 32'h0005E84F , 32'hFFFE6040 , 32'hFFFF9AA5 , 32'h0005A2E9 , 32'hFFFE08A9 , 32'hFFFF195B , 32'hFFFE9CA3 , 32'hFFFCE1EC , 32'h0004FFBC , 32'h00000FFC , 32'hFFFA60F6 , 32'h00019A4C , 32'hFFFFB7B1 , 32'hFFFA17FF , 32'h0002D64A , 32'hFFFA04DC , 32'h00021B73 , 32'h00041795 , 32'h000A36D8 , 32'hFFF74CF9 , 32'h0002F930 , 32'h00033BC9 , 32'hFFFF376A , 32'h000A4191 , 32'h000492D4 , 32'h00013925 , 32'hFFF50F5C , 32'hFFF50B99 , 32'hFFFA4BB0 , 32'hFFFEB0C3 , 32'h0009B4A3 , 32'hFFFCC259 , 32'h0001F97C , 32'h00034700 , 32'hFFFE4FBD , 32'h00003A88 , 32'h00031517 , 32'h00039F8A , 32'hFFFDC0A7} , 
{32'h3B75CC40 , 32'h5CAAC900 , 32'hD09A1100 , 32'hDEAFDB00 , 32'hFBE14F40 , 32'hFB508530 , 32'hFE82706C , 32'h13B18EA0 , 32'h23808000 , 32'hF890B880 , 32'hF0B31630 , 32'h0EFE4910 , 32'hE133B320 , 32'hDED11000 , 32'hD0756500 , 32'hE6D8E8A0 , 32'h065DB258 , 32'hE8F91C20 , 32'h0A327580 , 32'hF4983620 , 32'h0C577690 , 32'h1DB06D20 , 32'hED3D1DA0 , 32'h0983FA90 , 32'hF44A8F00 , 32'h0AE2AF90 , 32'hDD2D4AC0 , 32'hFDCD7614 , 32'h0177B8C4 , 32'hF88F6FC8 , 32'h097242A0 , 32'hEA4D7220 , 32'h008046D4 , 32'hE7CEACA0 , 32'h01A7DC44 , 32'hF5C4D520 , 32'hE8970800 , 32'hE3D63960 , 32'h0E81B640 , 32'hF8C734D0 , 32'hF034E770 , 32'h0D8815C0 , 32'hFFF09A58 , 32'h24670080 , 32'h04E02888 , 32'h0AD57B20 , 32'hFAF4B8A0 , 32'h08C97AD0 , 32'hFBEB7088 , 32'h09D49820 , 32'hF52004C0 , 32'h1504EFA0 , 32'h01BBA7F4 , 32'hF16D3F40 , 32'h09855030 , 32'hFCD67F34 , 32'hF85B75F8 , 32'hF8E85218 , 32'hFD938540 , 32'hFF7CDED2 , 32'hFCC7100C , 32'hF0915EC0 , 32'h043058F0 , 32'h145AF9E0 , 32'h08299A20 , 32'h02F340FC , 32'hF3C62F40 , 32'h0384A998 , 32'hFD755DB4 , 32'hFDBB6B44 , 32'hFF1F00C2 , 32'hFB3ABC90 , 32'hF82589D8 , 32'h020B24BC , 32'h040224E0 , 32'h0D7BE630 , 32'h036DAA64 , 32'h00FAFD44 , 32'h05318628 , 32'hF7FB2260 , 32'hFF625B0B , 32'h0902E900 , 32'h028C2D94 , 32'h062AFF00 , 32'hFC21D34C , 32'h03DAD40C , 32'h08059250 , 32'hFD468EF0 , 32'h01CC4EEC , 32'h001C016B , 32'hFFFDB828 , 32'hFFFFDCA5 , 32'h0001D42E , 32'hFFFABDB4 , 32'hFFFEAE68 , 32'h00028E63 , 32'hFFFF685B , 32'hFFFA63F0 , 32'h000274F0 , 32'hFFFE358A} , 
{32'h000049BC , 32'h0000C650 , 32'h00050A12 , 32'h00027543 , 32'hFFFB0B93 , 32'h00037DCB , 32'hFFFE5EDE , 32'hFFFD7316 , 32'h0003F665 , 32'h0008C342 , 32'hFFFD9F06 , 32'hFFFB2000 , 32'hFFFDCDD0 , 32'hFFFC4889 , 32'hFFFF7552 , 32'h000052A8 , 32'h0006D015 , 32'hFFFE84B2 , 32'hFFFFB44A , 32'h00035497 , 32'hFFFEEA45 , 32'h00002F39 , 32'hFFFE5A62 , 32'h0006CA01 , 32'hFFFB51DE , 32'hFFFF25A0 , 32'hFFF4AC55 , 32'h000450B8 , 32'hFFFE7E93 , 32'h000462FF , 32'h0002D03D , 32'hFFFD3742 , 32'h000539BE , 32'h0006E11C , 32'h00075683 , 32'hFFFDAA23 , 32'h00081CE8 , 32'h000609D5 , 32'hFFFB93BA , 32'h00015557 , 32'hFFFC0673 , 32'hFFFE443D , 32'hFFFA78D0 , 32'hFFFF0CA3 , 32'h0000467D , 32'h0002FDE3 , 32'h00058A98 , 32'hFFFDDF41 , 32'hFFFD1E10 , 32'h00081580 , 32'hFFFE517D , 32'h0003E4BF , 32'hFFFCE423 , 32'hFFFE1F7C , 32'h00029445 , 32'hFFF8FD85 , 32'h00070F59 , 32'hFFFAB5C4 , 32'h0008A0AA , 32'hFFFF2682 , 32'hFFFF8EDD , 32'hFFFBCBA2 , 32'h0006405C , 32'hFFF78757 , 32'h0000F694 , 32'hFFFBC210 , 32'hFFFED98B , 32'h000074EC , 32'hFFFFBDD5 , 32'h00078691 , 32'hFFFD9B22 , 32'h000298EE , 32'h0000D701 , 32'hFFFA7237 , 32'h00072D26 , 32'hFFF7723E , 32'hFFFCD95E , 32'h00012C2F , 32'h000089C2 , 32'h00027395 , 32'hFFF77144 , 32'hFFFCB6FF , 32'h000921B5 , 32'hFFF8022A , 32'h00056AD8 , 32'hFFF99B89 , 32'h0007D770 , 32'h0001B3D4 , 32'h0000F125 , 32'h00017916 , 32'hFFFCAEB8 , 32'hFFFCBDE3 , 32'h0004019D , 32'hFFFE3FF6 , 32'h00016C82 , 32'h0008EB02 , 32'hFFFBFF06 , 32'hFFFBFD3E , 32'h0000AC53 , 32'hFFF9A48A} , 
{32'h00030AF0 , 32'hFFFC6469 , 32'hFFFD0231 , 32'hFFF7C473 , 32'hFFFB7EB5 , 32'h00034C30 , 32'h00031C95 , 32'hFFF9888F , 32'hFFFB78C9 , 32'hFFFBF02D , 32'hFFF7E410 , 32'hFFFC251C , 32'hFFFFDD92 , 32'h0000E40C , 32'hFFFB8185 , 32'h00019F8C , 32'h0000AAB7 , 32'hFFFDDDAE , 32'hFFF1894B , 32'h0001EC98 , 32'h00079621 , 32'h00029062 , 32'h0004BA99 , 32'hFFF930EE , 32'hFFFD892E , 32'h00018D87 , 32'hFFF8F0B0 , 32'h0000AA00 , 32'hFFF9894D , 32'h0007AAF1 , 32'h00069205 , 32'hFFFB1A67 , 32'h0001F386 , 32'hFFFFE189 , 32'hFFF9B448 , 32'h0002922A , 32'h0007CBC4 , 32'h000320CF , 32'h00033D12 , 32'hFFFF800B , 32'hFFFE370D , 32'hFFFC430D , 32'h0004A610 , 32'h0003E9C5 , 32'hFFFDE786 , 32'hFFFEDE16 , 32'hFFFDE38E , 32'hFFFB9747 , 32'h00002273 , 32'hFFFDFB76 , 32'hFFFA5941 , 32'hFFFE5EC8 , 32'hFFFD100E , 32'hFFF9F819 , 32'h00048EBC , 32'h00033D36 , 32'hFFFD2742 , 32'h0008F71B , 32'hFFFE0C48 , 32'hFFFB4ECD , 32'hFFF7A7FB , 32'h00043C46 , 32'hFFFF0BF0 , 32'h0001A07B , 32'hFFFB952A , 32'hFFFD3F26 , 32'h0002C746 , 32'h0003C36C , 32'h0005EBA3 , 32'hFFF69CDE , 32'hFFFE8AC7 , 32'h00002C87 , 32'hFFF77B58 , 32'hFFF512A5 , 32'h00047E3B , 32'h000230EA , 32'h0005FD2B , 32'hFFF5EE59 , 32'hFFFE49C6 , 32'h00037630 , 32'h00058E00 , 32'hFFFFA49F , 32'h000362AA , 32'hFFFD0F31 , 32'hFFFA7AF0 , 32'hFFFE0044 , 32'hFFFD120E , 32'h00036F2C , 32'hFFFD2ADA , 32'hFFF94001 , 32'h0004FA1F , 32'h000650A1 , 32'hFFF6B564 , 32'hFFFE0091 , 32'h000B5D5D , 32'hFFFDA8F4 , 32'h0004E01A , 32'hFFFB8417 , 32'h00008343 , 32'h00028857} , 
{32'hFFFAFA99 , 32'hFFFFB6FC , 32'h0002A9D4 , 32'hFFFE866E , 32'h00035F31 , 32'hFFFC9DD1 , 32'h0000A291 , 32'h00021CC8 , 32'hFFFD15C8 , 32'h0000B523 , 32'h0003A3BB , 32'hFFFFF3C9 , 32'h0005B884 , 32'h00027C43 , 32'h00010741 , 32'h0003FD69 , 32'h0001E450 , 32'hFFFC837E , 32'h000A5BA0 , 32'hFFFF196C , 32'h000009C4 , 32'hFFFC95A4 , 32'h0000B8D0 , 32'hFFFFF1E5 , 32'hFFFB6D2D , 32'h000158FD , 32'hFFFD25E2 , 32'hFFFAA5B6 , 32'h000AF26E , 32'h0003038F , 32'hFFFC69B9 , 32'h0006862E , 32'h00008F1E , 32'hFFFDE0DC , 32'h0003935D , 32'h0003FB61 , 32'h0009E3B8 , 32'hFFF8D9C2 , 32'h000A38BF , 32'hFFFE8865 , 32'hFFFC37EF , 32'hFFFD18E0 , 32'h0003A87A , 32'h0008C0DF , 32'h0003E73E , 32'hFFFE2DD6 , 32'h0002D99A , 32'h00030A75 , 32'h0003D154 , 32'hFFF78F6A , 32'h0004136D , 32'hFFFC97AD , 32'hFFFEE55B , 32'hFFF4F118 , 32'h00055828 , 32'h00058EB4 , 32'h00010846 , 32'hFFF80A88 , 32'hFFF8AC39 , 32'hFFFA5071 , 32'h000333F5 , 32'hFFFB1B29 , 32'hFFFF7587 , 32'h000843D7 , 32'hFFFE1ABB , 32'h000423AF , 32'hFFFBA0F7 , 32'h00006BCF , 32'h00012299 , 32'hFFFF24FF , 32'hFFF807D0 , 32'h00007146 , 32'h0003499B , 32'hFFFFF22A , 32'h000086C7 , 32'hFFFFB698 , 32'h0004F006 , 32'h00016D6F , 32'h0004D7AA , 32'h0002C5B1 , 32'h00063424 , 32'hFFFFC526 , 32'h000288C6 , 32'h0006E0CC , 32'h000334F3 , 32'hFFFC6D7D , 32'hFFFB707F , 32'hFFFE4A60 , 32'h00011C5D , 32'h0001A106 , 32'hFFF72B1E , 32'hFFF820FA , 32'hFFFAFD81 , 32'hFFF870CA , 32'hFFFF7A5E , 32'h0006EF20 , 32'h00000EC0 , 32'h0003B6E0 , 32'hFFFA72FA , 32'h0001EDD9} , 
{32'hF3C9E290 , 32'hFBE041F8 , 32'hC8E9EA80 , 32'hCFB247C0 , 32'hAE565C80 , 32'hE6C19640 , 32'h0FFE6310 , 32'h008EFF4E , 32'hCD46F580 , 32'h2BE330C0 , 32'h0D968B70 , 32'h0BDD0650 , 32'h0BB79DE0 , 32'hF3579430 , 32'hE8E51900 , 32'h3CE9DD80 , 32'h14CF65A0 , 32'h114C4300 , 32'hD2A51D40 , 32'h2CA27A40 , 32'hD9F64AC0 , 32'hFB892580 , 32'h0A597390 , 32'hE79CBC00 , 32'hF0172A20 , 32'hF533F910 , 32'hE5ED1A80 , 32'h0DEC6BE0 , 32'hFC13A8E8 , 32'h03AAEEC4 , 32'hE0EEB760 , 32'h03E73BA0 , 32'h046D3498 , 32'h156DABC0 , 32'h0B292BB0 , 32'hD3F02B80 , 32'hF021A960 , 32'hF8E0C5B0 , 32'h026D4034 , 32'hF7C6B330 , 32'h061B0288 , 32'h20E1DE40 , 32'hFD0B93D4 , 32'hEDD9F320 , 32'hFF8FFE7D , 32'hFDCB49B4 , 32'h13AFAB20 , 32'hF3A6EA60 , 32'h03907C44 , 32'h029602D4 , 32'hEF369FC0 , 32'hFEC5DA5C , 32'h00164E14 , 32'h0DB249A0 , 32'h047CEA38 , 32'hFCED99F0 , 32'h07C1BBE8 , 32'hF8953000 , 32'h000F28AE , 32'hFE4C2E98 , 32'hF7931360 , 32'hF6D68460 , 32'h06D37268 , 32'h024F67E4 , 32'h0862B4E0 , 32'hFB8EED20 , 32'hFED79200 , 32'h004D9CC7 , 32'hFA365188 , 32'hFB62EEC0 , 32'hF9FDFCA8 , 32'hF842F730 , 32'hFF912917 , 32'hF652F650 , 32'h0A2D1CB0 , 32'h0AD70000 , 32'hFD022828 , 32'hF596CB00 , 32'h0524B820 , 32'hF845A3D0 , 32'hFD060174 , 32'h00696045 , 32'hF8AB0D00 , 32'h026B6378 , 32'hF5024930 , 32'hFE20DDB8 , 32'hF8761598 , 32'hFC0D1E34 , 32'hFB5765E0 , 32'h015966F0 , 32'h00007B2C , 32'hFFFF0377 , 32'h00024BD7 , 32'hFFFCB2AE , 32'h00003139 , 32'hFFFF1205 , 32'hFFFCBC0E , 32'h0002B154 , 32'hFFFE9B6C , 32'hFFFFEB25} , 
{32'hC6C0CB80 , 32'h0E370820 , 32'hEF3BA600 , 32'h49C50B80 , 32'h2DAB9280 , 32'hD1279780 , 32'h2343CAC0 , 32'hA6EA5B00 , 32'h0D5008A0 , 32'hF759D330 , 32'h0083330C , 32'hD4574B00 , 32'hB48DB080 , 32'hFD7E3600 , 32'h0D848F60 , 32'h163C0920 , 32'h03CB0BD0 , 32'h493EAD00 , 32'hFB724A88 , 32'h38D23F80 , 32'hFF739F25 , 32'h3AF802C0 , 32'hFECF9B5C , 32'hDFA3E500 , 32'hEC072980 , 32'hEA50E200 , 32'hED26B540 , 32'h02C58DEC , 32'h160B9740 , 32'hF61914C0 , 32'hDF137E80 , 32'h001322AC , 32'h02244F64 , 32'hF743C500 , 32'h0F592CD0 , 32'hFEF89244 , 32'hF45076F0 , 32'hF81D9F60 , 32'h02921084 , 32'h107CE6A0 , 32'h005715BA , 32'h01459D70 , 32'hF1D6AEB0 , 32'h082CC040 , 32'hF8895ED0 , 32'h0482C000 , 32'h0F317C10 , 32'hF99B1680 , 32'hF55EF640 , 32'h06AA76C8 , 32'hFABF4430 , 32'h13A79A40 , 32'hEEE7F3C0 , 32'h07722D58 , 32'h03A0C304 , 32'hF40DC450 , 32'hF8B79238 , 32'hF51CB240 , 32'hFC253718 , 32'h02E61178 , 32'h05F73068 , 32'hF6DECCB0 , 32'h07CA7FE8 , 32'hF63F8F80 , 32'hFA2433C8 , 32'hF840CB90 , 32'h06FAB380 , 32'hF3B3D710 , 32'h0ACB48D0 , 32'h0AE5C3E0 , 32'hFF4FC605 , 32'hF43E53F0 , 32'hF9424108 , 32'h09E10530 , 32'hF1B16DE0 , 32'hF5BC5840 , 32'hF86C74A8 , 32'hF5940F30 , 32'hFFD61488 , 32'h04680148 , 32'hF9490108 , 32'h02C4AC04 , 32'hFE5066B8 , 32'h0955F210 , 32'h00FAA0CE , 32'hFD3CB2FC , 32'h014F30F8 , 32'hFD4AA4EC , 32'h025D7F64 , 32'h0009281D , 32'h0000275A , 32'hFFFF780C , 32'hFFFBBE4F , 32'h0001670C , 32'hFFFA4264 , 32'h0000D097 , 32'h000092E3 , 32'h00022B75 , 32'h00036BB9 , 32'h00038691} , 
{32'hFFFE5B96 , 32'h0008CBF6 , 32'h00003128 , 32'h0000EDAE , 32'h000D89AF , 32'h0003C8C4 , 32'h000013BE , 32'h0002402F , 32'h00016B50 , 32'h00042FFA , 32'h00038BA7 , 32'hFFFCD569 , 32'hFFFEC1F4 , 32'hFFFF9DBF , 32'h0006F896 , 32'h0000F99A , 32'h00065B39 , 32'h000586D1 , 32'h00067CD9 , 32'hFFF77E67 , 32'h0001D256 , 32'hFFF02DA7 , 32'hFFFAD080 , 32'h00048911 , 32'hFFFE390D , 32'hFFF86AE3 , 32'h0005A0C9 , 32'h0001B8E7 , 32'hFFF91B6E , 32'hFFFD1E89 , 32'hFFF8CFA6 , 32'h000D2BC0 , 32'h0008F474 , 32'hFFFF6B9E , 32'hFFF8DE57 , 32'hFFFFEFFD , 32'h0003CDAB , 32'h00038995 , 32'hFFFF2B2C , 32'h0004049C , 32'hFFFFD2D1 , 32'hFFFC46E0 , 32'hFFFEF282 , 32'hFFFF90DE , 32'h00042DE6 , 32'h00023DE9 , 32'hFFFCAE48 , 32'h00015AD5 , 32'hFFFE05DA , 32'h00072F3C , 32'hFFF7048F , 32'h00019036 , 32'hFFFDD1E2 , 32'hFFFD38EC , 32'h0009446D , 32'h000098AB , 32'h00009C37 , 32'hFFFBAEBE , 32'h0001555F , 32'hFFFA1ACF , 32'hFFFD9B8E , 32'h00054C9D , 32'hFFF8F5B8 , 32'h00037BBA , 32'hFFFDA445 , 32'hFFF43FC2 , 32'hFFFECFCF , 32'h0003C8C1 , 32'h00023FEE , 32'h00070218 , 32'hFFFB6A1F , 32'h00031B5C , 32'hFFFB6C2F , 32'h0002019D , 32'h00014D1E , 32'hFFFEE3E1 , 32'h00090047 , 32'h0009D953 , 32'hFFFEF6F4 , 32'hFFF6AA22 , 32'hFFFC0F07 , 32'h0005FE9C , 32'h0000C61C , 32'h000507B6 , 32'hFFFDFABE , 32'h00047ECF , 32'hFFFFE476 , 32'h0007879E , 32'h000399D4 , 32'h00069737 , 32'h0000D1FB , 32'h00002E2D , 32'h0000CFEC , 32'hFFFD3629 , 32'hFFF71927 , 32'hFFFC9FE6 , 32'hFFFBA83F , 32'h00032BD0 , 32'hFFFA314B , 32'hFFFA4032} , 
{32'hFFF93D3A , 32'hFFF721B4 , 32'h0000CC00 , 32'hFFFFD683 , 32'h00026221 , 32'hFFFF7E9F , 32'hFFFF2325 , 32'h0001CC1B , 32'hFFFD830F , 32'hFFF9737B , 32'hFFFAD839 , 32'h00096D16 , 32'hFFFC500C , 32'h0000CE5E , 32'hFFFDA1A4 , 32'h0005D73D , 32'hFFFFFF80 , 32'h000418D6 , 32'hFFFC2718 , 32'h0002C5C9 , 32'hFFFEABA9 , 32'hFFF7A4E1 , 32'h0000257F , 32'hFFFE9742 , 32'h000FDED0 , 32'hFFFCDC1B , 32'h00001BFB , 32'hFFFFF885 , 32'h000292BE , 32'h000185EB , 32'h00028C8E , 32'h0003B4E8 , 32'h0001CC3C , 32'hFFFF1157 , 32'hFFF93AAD , 32'h0002BDA1 , 32'h000550F7 , 32'hFFFCDBC4 , 32'hFFFC4B63 , 32'hFFFA2BF6 , 32'hFFFE2AA0 , 32'hFFF849DD , 32'h0000EC9F , 32'h0006B8A5 , 32'h000CA5B5 , 32'h0001F5A8 , 32'hFFFE1448 , 32'h0000A04A , 32'hFFF67BA6 , 32'hFFF902A7 , 32'hFFF58DE7 , 32'h0000269F , 32'hFFFEED24 , 32'h00085AC4 , 32'hFFF9A798 , 32'hFFF989B7 , 32'h00016EB8 , 32'hFFF94BA4 , 32'h000A0D0B , 32'hFFFAACF6 , 32'hFFFB7D07 , 32'hFFFF607E , 32'hFFFF8ACD , 32'h00027E40 , 32'hFFFBE3FC , 32'hFFF9C067 , 32'hFFF8C2B2 , 32'hFFFD968C , 32'h0004F059 , 32'h00029383 , 32'h00010478 , 32'hFFFF8EFC , 32'h00040521 , 32'hFFFE3D80 , 32'h00053C58 , 32'hFFFD5AE8 , 32'hFFFB9A84 , 32'hFFF0178B , 32'h0003C51F , 32'h00023D2B , 32'h000304A7 , 32'hFFFD60B4 , 32'hFFF6382F , 32'h00072AC5 , 32'hFFFCA44D , 32'hFFFB0064 , 32'h00036D1F , 32'hFFF75533 , 32'hFFFCD87A , 32'hFFFEA912 , 32'hFFFACE42 , 32'hFFF6AC0F , 32'hFFF7AC28 , 32'hFFFAD6EC , 32'hFFFD8F5D , 32'h00009D7F , 32'hFFFAEA1E , 32'h00035AEA , 32'hFFFE2C7F , 32'hFFFE64FA} , 
{32'h00034817 , 32'hFFFEE1C9 , 32'h00097C55 , 32'h00008DC6 , 32'hFFF8C01D , 32'h00038EE0 , 32'h000066D9 , 32'h00031370 , 32'hFFFD4C01 , 32'hFFFF52BA , 32'h0004AAFF , 32'h0006F906 , 32'h00029D79 , 32'h00081E62 , 32'h00071BFF , 32'hFFF5D21C , 32'hFFFB6D1A , 32'hFFF9C8D1 , 32'h0000B284 , 32'hFFFF2C90 , 32'h00004AB8 , 32'hFFFFFEB3 , 32'h00076522 , 32'hFFFF2B39 , 32'hFFFE36C3 , 32'hFFFDD707 , 32'h0009E5CC , 32'h000065A8 , 32'h00004BB4 , 32'h000468E0 , 32'hFFFEBCCA , 32'hFFFDE258 , 32'hFFFE507B , 32'h0004609B , 32'h000A53CC , 32'hFFF838A2 , 32'hFFF7165C , 32'h00032165 , 32'hFFFAF8F6 , 32'hFFFC306F , 32'hFFFC21F2 , 32'h0001905F , 32'h000145CD , 32'hFFFE4E6E , 32'hFFFEAF1D , 32'h0005A02F , 32'h00039DE7 , 32'hFFF67B0D , 32'hFFFAADC5 , 32'h00051B7C , 32'hFFF5B3B8 , 32'hFFFC8A71 , 32'h0004E328 , 32'hFFFD5049 , 32'h000496A8 , 32'h000AFD23 , 32'h0001C821 , 32'hFFFF5585 , 32'h00019D57 , 32'h0003A33F , 32'hFFFC7582 , 32'hFFFF3308 , 32'h0004AF14 , 32'hFFFF5C2E , 32'h0009F1C3 , 32'hFFFF7963 , 32'h0003882B , 32'hFFFA2A10 , 32'h000033E7 , 32'h000AB781 , 32'hFFFF5F78 , 32'hFFF73F55 , 32'h00013514 , 32'h0002E9E9 , 32'hFFFE87DA , 32'hFFFF0A1A , 32'hFFFE69DA , 32'h000305E7 , 32'h0001B7A2 , 32'hFFFBDEB3 , 32'hFFFB2015 , 32'hFFF5BBCF , 32'hFFFE2EB9 , 32'hFFFEC530 , 32'hFFFC3DA7 , 32'h00045028 , 32'hFFFEF5E3 , 32'h000421FC , 32'hFFFFA17D , 32'hFFFBC9D3 , 32'hFFFB22BD , 32'h000A49E6 , 32'hFFFB1784 , 32'h00073968 , 32'h0000C9CC , 32'h0006C9DA , 32'hFFFBC213 , 32'h00021AF1 , 32'hFFFE885B , 32'h0005A674} , 
{32'hFFFEE6AC , 32'hFFFF9BC9 , 32'h0002F404 , 32'hFFFD485A , 32'hFFFE03EA , 32'hFFFEBFAE , 32'h0007DFF1 , 32'h000531D0 , 32'h000143B6 , 32'h00003070 , 32'h0000154E , 32'h00017F9D , 32'h00010B13 , 32'h00005C6F , 32'h000076A0 , 32'h0007A043 , 32'hFFFB1AFA , 32'h0003C403 , 32'hFFFD5A4D , 32'h00023FFD , 32'hFFFA8ED1 , 32'hFFFBDEBE , 32'hFFFC893F , 32'h0001C391 , 32'hFFFAF07D , 32'h00090062 , 32'h00021574 , 32'h0002F63E , 32'hFFFD652B , 32'h000406BA , 32'hFFFE6530 , 32'h00048646 , 32'h0003C0C6 , 32'hFFFC3168 , 32'hFFFB27B0 , 32'hFFFB23A2 , 32'h0000BCBE , 32'h0000C487 , 32'h00021FDB , 32'hFFF64E9A , 32'h0002F1B1 , 32'h00006276 , 32'hFFFE24CA , 32'h000C056F , 32'h0003744F , 32'hFFFC478F , 32'h00000E65 , 32'hFFFC08E7 , 32'h0001B477 , 32'hFFFF5A30 , 32'h0000FA03 , 32'h00031E36 , 32'h000777B7 , 32'h00001F2A , 32'hFFFCDE11 , 32'h00039675 , 32'h0003DE14 , 32'h0006DF14 , 32'h0001732A , 32'h0000DE24 , 32'hFFFDFA64 , 32'hFFF9F927 , 32'h0001E100 , 32'hFFFF0D5B , 32'hFFF852A5 , 32'hFFFE6C43 , 32'hFFFB2E1D , 32'h0000A674 , 32'hFFFF07BB , 32'h000309D4 , 32'h0001A2D9 , 32'h0002682F , 32'hFFFEF1E3 , 32'hFFFD8003 , 32'hFFFF59C2 , 32'hFFF6221F , 32'h000070A3 , 32'h0001D534 , 32'h0000AD9B , 32'h0007A2DA , 32'hFFFE97B4 , 32'h0002EB49 , 32'hFFFDC021 , 32'hFFFFFEEC , 32'h0003AA47 , 32'hFFFD9ABA , 32'h0006AEF7 , 32'h00072BDD , 32'h00051F8E , 32'h00032C41 , 32'hFFFF940B , 32'hFFFE67DF , 32'h000104F7 , 32'hFFFD49EB , 32'h0004140B , 32'hFFFA89B4 , 32'h0005802D , 32'hFFF98EF8 , 32'h0001910A , 32'h0000007B} , 
{32'hDA2F2B80 , 32'hDF2932C0 , 32'h3CB00F40 , 32'h34E69A40 , 32'h4022EB80 , 32'h40F72F80 , 32'h2E5F1900 , 32'hED291840 , 32'h132FB020 , 32'h16928DC0 , 32'hB6DBAA80 , 32'hFD27EA10 , 32'hF9A58A68 , 32'hFBB62730 , 32'hD27BE300 , 32'h098EABC0 , 32'hD0FB7800 , 32'hE6801880 , 32'hF22D8070 , 32'h20DD1FC0 , 32'hFBB64EB8 , 32'h0CB7C9B0 , 32'hCFBD90C0 , 32'hEBFBAB20 , 32'hEE210560 , 32'hFCA938CC , 32'hFEFEA128 , 32'hDA521B80 , 32'hFAB253E0 , 32'h07C1F668 , 32'h00419756 , 32'hF6530B40 , 32'hF7F1A240 , 32'h09E35190 , 32'h15053CE0 , 32'h17A036A0 , 32'hF414D310 , 32'h135D3F20 , 32'h0476B8D0 , 32'h1EB7B2A0 , 32'h18E0B9C0 , 32'hF5310640 , 32'h04210BE8 , 32'h0FF7E380 , 32'h23D9B100 , 32'h04C20208 , 32'h0090C542 , 32'hF88B8ED8 , 32'hFC30E8EC , 32'hEB506B80 , 32'hF20AB080 , 32'h006BBA07 , 32'hF77684E0 , 32'h185F19E0 , 32'h0619E7E8 , 32'h00889A31 , 32'hF425EDF0 , 32'hF68D1B60 , 32'h08264490 , 32'hF1506E10 , 32'hF43246A0 , 32'h151E2160 , 32'hFC0DB820 , 32'h075E3818 , 32'hF74BDF00 , 32'h09CD7110 , 32'hFD24C198 , 32'h0B302C80 , 32'hFCF74280 , 32'hF7D5B600 , 32'h0AC64560 , 32'hFF694673 , 32'h0E875980 , 32'h07057DB8 , 32'h0E81EA20 , 32'h077E3118 , 32'hFE3A2000 , 32'hFB178B28 , 32'hF7EBCD60 , 32'h00D9CF62 , 32'hFE778B10 , 32'h070B9A18 , 32'hFC18D1EC , 32'h035B2994 , 32'h07313460 , 32'h037AE4EC , 32'hFC307028 , 32'hFC26CC80 , 32'h02854FBC , 32'h0085E501 , 32'hFFFB66CF , 32'hFFFE83BF , 32'h000271EB , 32'h0000FACC , 32'h00010572 , 32'hFFFF2A70 , 32'hFFFB7F77 , 32'hFFFE4278 , 32'h0002B599 , 32'h00015FA1} , 
{32'h1EC4B8C0 , 32'h18D0AC80 , 32'h41168E00 , 32'h223D7240 , 32'hD209D040 , 32'hDF886700 , 32'hF5FC5EF0 , 32'hE4C89D60 , 32'hDA6FA740 , 32'h0DE0A000 , 32'h0F8284C0 , 32'h219EC280 , 32'hDD765440 , 32'hF7EE67F0 , 32'hE73B4F20 , 32'hF65C3A10 , 32'hFBBFB658 , 32'hF8A705E8 , 32'hDC84F8C0 , 32'hF53F6A90 , 32'h0B602D70 , 32'hFB3C1448 , 32'h0A997070 , 32'hF8189FB0 , 32'h2C0EC580 , 32'hFF602C39 , 32'h08FA0480 , 32'h0F50C600 , 32'hF7CE6D20 , 32'h21A87C80 , 32'h13DA10A0 , 32'h109C7840 , 32'hF1477010 , 32'h06F034D8 , 32'hF26A6700 , 32'h11FC0EA0 , 32'hFF617810 , 32'hF0CA4E10 , 32'h0F41BC00 , 32'h0410D2A0 , 32'hD11F09C0 , 32'hFF178F65 , 32'hFFF8AA22 , 32'hF63CDAD0 , 32'h03F3ED24 , 32'hF3D24170 , 32'h05976888 , 32'hF2E122E0 , 32'hF770D800 , 32'hF0FE7820 , 32'h0A685180 , 32'h15A5B520 , 32'h086F7E80 , 32'h20653440 , 32'hFADBF6E0 , 32'h00C20E2E , 32'h06999888 , 32'hFD93300C , 32'hFABEB680 , 32'h04D229A0 , 32'h204B0480 , 32'hFAE15798 , 32'h00556F28 , 32'h0B101410 , 32'hFC240A30 , 32'h04DF1210 , 32'hF6E1B3E0 , 32'hFB29BF20 , 32'h1F5DBC20 , 32'h07E4DC10 , 32'h0B285DA0 , 32'h00292AFB , 32'hFA39F688 , 32'hFEBDA60C , 32'hF8C9D280 , 32'h07695858 , 32'hFD4E357C , 32'hFBF289F8 , 32'h04C4BE20 , 32'hFAFF1BF8 , 32'h04F339C8 , 32'h077013B0 , 32'hFAA701B0 , 32'hFCE544C4 , 32'h02B6011C , 32'h07F41678 , 32'h037234EC , 32'h059209C8 , 32'h02ED24B0 , 32'h000B2494 , 32'h000081C8 , 32'hFFFC385D , 32'hFFFFCE67 , 32'h0007ACB9 , 32'h0004FA79 , 32'hFFFD5E16 , 32'h0000BBEB , 32'h0001E8C3 , 32'h0000F49F , 32'hFFFFCFB2} , 
{32'h3EECBB00 , 32'h1351D640 , 32'h53648F80 , 32'hE052E260 , 32'h0FB8F520 , 32'hB6D1E300 , 32'hB8C7FF80 , 32'h06517EC0 , 32'hC7013900 , 32'hF1F6C5A0 , 32'h02C45830 , 32'hEDCECC60 , 32'h0B27BF40 , 32'h29C2D980 , 32'hFF2C970B , 32'h11CDFAE0 , 32'hE9DB85E0 , 32'h0424C388 , 32'h08A7C390 , 32'h093EDDD0 , 32'hFD02B054 , 32'hFC36F0CC , 32'hDE18A280 , 32'h04034268 , 32'h0890C340 , 32'hE34B31C0 , 32'h124D7B60 , 32'h1A1CC7E0 , 32'hD4057F40 , 32'hF25F4360 , 32'hEFDE5600 , 32'h192E1220 , 32'h272E3FC0 , 32'hFB69A8B0 , 32'h03D4FB7C , 32'hF4D56C30 , 32'hDF24D900 , 32'h02CDDFF8 , 32'hF4F16D00 , 32'h062DBD98 , 32'hFA3E9CA0 , 32'h0B121610 , 32'hE73A9960 , 32'h25F0A800 , 32'hFDDFE3D8 , 32'hF3AFC020 , 32'h07B33C30 , 32'h037F7910 , 32'hF3BF7EA0 , 32'hF871E568 , 32'h02C4F818 , 32'h15649D60 , 32'hFF46BBBB , 32'hF8747620 , 32'hF1CB4F10 , 32'h0C79BDA0 , 32'hFCA4DE64 , 32'h0A1A7490 , 32'h0C3D3400 , 32'h05115688 , 32'h148F8F60 , 32'hFD165898 , 32'h03023414 , 32'hFE91CFB0 , 32'hFCAE53DC , 32'h03EB7434 , 32'hF8EF1418 , 32'hFF92B6A0 , 32'h01BBF8E0 , 32'hFA2D6A08 , 32'hFE4221BC , 32'hFD12DF1C , 32'h045DF658 , 32'hF684DEE0 , 32'h0BB99B00 , 32'hFBE2E660 , 32'h028EF90C , 32'hFCDCCDC4 , 32'hFA704BC8 , 32'hFCC1C9AC , 32'h03234E48 , 32'h04D68560 , 32'hFD05DEE0 , 32'h05056878 , 32'h01F87458 , 32'h014B89F0 , 32'hFEB539AC , 32'hFEFFBC98 , 32'h05111410 , 32'hFFC5AEDB , 32'hFFFE91EE , 32'h00067BD4 , 32'hFFFFD116 , 32'hFFFF1836 , 32'h0005E3FF , 32'h0003A5E7 , 32'hFFFE0C06 , 32'hFFFE34FD , 32'h000026AF , 32'hFFFD44B8} , 
{32'hE7B187A0 , 32'hE1D13240 , 32'hC44D1A40 , 32'hFD956BAC , 32'h8C9C8180 , 32'hE83F0140 , 32'hD2C26000 , 32'hDFFF3D00 , 32'hD0B53400 , 32'hFE10BBFC , 32'hD7E01800 , 32'h34C51880 , 32'hE2A28360 , 32'hE1A80660 , 32'h00B3B0A3 , 32'h14709120 , 32'h1C6D3120 , 32'hEA7D4BA0 , 32'h1865DAE0 , 32'hD94C5240 , 32'hED5561A0 , 32'hD60A0980 , 32'h031425F8 , 32'hCA44A940 , 32'h100EA200 , 32'hC260DCC0 , 32'hDFCD6C40 , 32'h0573BFB8 , 32'hEB1499E0 , 32'hF8738AD8 , 32'h07294020 , 32'hD6EED080 , 32'hFBA2D3D0 , 32'h10AB62A0 , 32'hF904D078 , 32'hF1B54810 , 32'hF55D3180 , 32'hFEB205E8 , 32'hD887DC40 , 32'hE9DCA100 , 32'hFA6443A8 , 32'hF6000A10 , 32'hE2BBD4E0 , 32'hFA573780 , 32'hFAEE69D0 , 32'h136C17E0 , 32'hFAA04EE0 , 32'h06424D68 , 32'h05C72EA8 , 32'hEBE09180 , 32'hF8DB4070 , 32'h025FE68C , 32'hFF941A2F , 32'hFBDD3D30 , 32'h01322DB8 , 32'hFD0272A4 , 32'h08E7E960 , 32'h0785A370 , 32'h017451B8 , 32'hF74DAD10 , 32'hFEC78884 , 32'hFF45BE0A , 32'hECD860E0 , 32'h0703FAB0 , 32'hFB140C18 , 32'h0062C725 , 32'h06BA5C10 , 32'hF85542D0 , 32'hEF1C5E80 , 32'h0ED8A4C0 , 32'hFB3A58D0 , 32'hF268F0E0 , 32'hFE8BE240 , 32'hFE9720DC , 32'h061444A8 , 32'hF4B25C70 , 32'hF7D3DE20 , 32'h05A34498 , 32'hFA3F6860 , 32'h0061EBD8 , 32'h08B358E0 , 32'h04B183E0 , 32'h0A631A60 , 32'hFC1C40C4 , 32'h0585E618 , 32'hFE7A527C , 32'h043FAB48 , 32'hF6C8B620 , 32'h04FEC678 , 32'h014B167C , 32'hFFFECA9C , 32'hFFF95814 , 32'h00023761 , 32'h000245C7 , 32'hFFFE4CFA , 32'hFFFEE40B , 32'h0000011E , 32'hFFFFD3B4 , 32'h00049DA2 , 32'h0001295D} , 
{32'hD40E9A00 , 32'hC475BF80 , 32'h2D8C2400 , 32'h0A1E84C0 , 32'hCE437800 , 32'hE328F3C0 , 32'h101EBD60 , 32'h1B210040 , 32'h1FB99F00 , 32'hE8BCB3C0 , 32'h0A046560 , 32'hEF452EC0 , 32'h04C3AC38 , 32'hE0A2AD00 , 32'hDA6D0AC0 , 32'h1E330860 , 32'hF74878C0 , 32'h1A32C1A0 , 32'hFD5AB828 , 32'h2B59E040 , 32'h28390380 , 32'h0EC9F910 , 32'h05BD0EF8 , 32'hFD7E7A8C , 32'hF02BF120 , 32'hEDB4FC40 , 32'h0A540720 , 32'hE4435840 , 32'hF3166780 , 32'hEDDFB4E0 , 32'h0C5AD1A0 , 32'hF944CF40 , 32'h009B16F2 , 32'hFE1E3F1C , 32'h112DC620 , 32'hF9674FA0 , 32'h19B54F20 , 32'hF354B3C0 , 32'hF0E64AC0 , 32'h005E4C0D , 32'hF9577DD8 , 32'h008B56DF , 32'hF30555C0 , 32'hF4984540 , 32'hE3C7A3A0 , 32'hE380B4A0 , 32'hEB8BD5C0 , 32'hE5C6FE00 , 32'hFDC7E214 , 32'hF8823730 , 32'h0D375A30 , 32'h0E0D4F80 , 32'hFAA12280 , 32'hFFA7C2E7 , 32'hFBE42BC0 , 32'hF6708AA0 , 32'h09F6A300 , 32'h14828FA0 , 32'hF0C8BB00 , 32'hF969D610 , 32'hFD90EED0 , 32'h0862E1B0 , 32'h06ED7850 , 32'h033E81D0 , 32'h17FF82A0 , 32'h02A3FEAC , 32'h0F74F9E0 , 32'hF82C8F08 , 32'h08E8A970 , 32'h01DB57A0 , 32'hF7DCE6F0 , 32'h06C5ABB0 , 32'h032F0A84 , 32'hF5DA85C0 , 32'hF21BA100 , 32'h003C59A8 , 32'hFE8811F0 , 32'h0BF60010 , 32'hFD8D4118 , 32'hFD47786C , 32'h0385AB98 , 32'h0A4AA150 , 32'h005F8253 , 32'h016BEE1C , 32'h068BDCF8 , 32'hFEEF145C , 32'hFF70EFC6 , 32'hFC996310 , 32'hFCD89744 , 32'h024AC0C0 , 32'hFFF59DD2 , 32'h0002A60F , 32'h0005BCBE , 32'hFFFE15DA , 32'h000103C4 , 32'h0000E139 , 32'h0005191B , 32'hFFFAD110 , 32'hFFFF1483 , 32'h0000A42B} , 
{32'hFFFD610D , 32'hFFFB406D , 32'h0007727F , 32'hFFFE4CE4 , 32'hFFFD7471 , 32'h0001AF46 , 32'h00009F6B , 32'hFFFCC2C7 , 32'hFFFC5F29 , 32'hFFFE08A8 , 32'h0005A947 , 32'hFFF8F117 , 32'hFFFB0D05 , 32'hFFFB80F9 , 32'hFFF91E30 , 32'h0005E5DC , 32'hFFFEE12D , 32'h00064D0A , 32'h0000646E , 32'hFFFF637B , 32'hFFFD73F2 , 32'h0005B70C , 32'h00079D37 , 32'hFFFED80B , 32'hFFF9983B , 32'h00047D4B , 32'hFFF9AB7E , 32'hFFF7BC54 , 32'h0000EBC6 , 32'hFFFEC1A5 , 32'hFFFC6558 , 32'hFFFD24A6 , 32'hFFFAB561 , 32'h0000C241 , 32'hFFFD50F7 , 32'hFFFEEA99 , 32'hFFFF61C7 , 32'hFFFE615B , 32'hFFFCB2BA , 32'h000A4972 , 32'hFFFE8422 , 32'hFFFF7397 , 32'h000161C7 , 32'h000383E2 , 32'hFFFD24A5 , 32'hFFFC163B , 32'h00003B55 , 32'h0004B448 , 32'hFFFA5FCF , 32'hFFFBA3E4 , 32'hFFFE9338 , 32'hFFFBB5D5 , 32'h0002433F , 32'hFFFD0B7F , 32'hFFFD818A , 32'hFFFD9FA2 , 32'hFFFFF0A1 , 32'h00027245 , 32'hFFFB7B5A , 32'h0003488A , 32'hFFFA6F13 , 32'h0004CF3F , 32'hFFFCCFF6 , 32'hFFFF6EAB , 32'hFFFA55C0 , 32'hFFFDEA3C , 32'hFFFC7585 , 32'hFFF9298B , 32'h00010EDE , 32'h000B2582 , 32'hFFFAB667 , 32'h0000C4C8 , 32'hFFFF5D6E , 32'hFFFB7D31 , 32'hFFFE30BF , 32'hFFFDC4DA , 32'h0001248B , 32'h00002A90 , 32'h000107F2 , 32'hFFFF71A9 , 32'hFFFF1F77 , 32'h0005DF0B , 32'h00005CE3 , 32'hFFFF7243 , 32'h0004568D , 32'h000097D2 , 32'hFFFB4834 , 32'hFFFECE25 , 32'h0003EAD9 , 32'h00079C8E , 32'h00006027 , 32'hFFFCC770 , 32'hFFF9A507 , 32'h0008D53F , 32'h0002D403 , 32'hFFFFCB57 , 32'hFFFC983D , 32'h00071D30 , 32'h00022249 , 32'hFFFF7F03} , 
{32'h00030B1B , 32'hFFFBFC05 , 32'h0004BED1 , 32'hFFFDEF41 , 32'hFFFDCDC1 , 32'hFFFD4E5F , 32'hFFF9D13E , 32'h0003355B , 32'h0006A0B0 , 32'h0000DBD4 , 32'h0004CA0C , 32'hFFFE1740 , 32'h00028745 , 32'hFFFA54AC , 32'h0005A498 , 32'hFFFE5084 , 32'h0007FDF5 , 32'hFFFB086C , 32'h00041E12 , 32'h00003FCF , 32'h00011CBD , 32'h0005520E , 32'h0003B9CC , 32'hFFFA4CF1 , 32'hFFFB9A23 , 32'hFFFD02FC , 32'hFFF39433 , 32'h00055E75 , 32'h000047B0 , 32'h0002B2BD , 32'h000A7D14 , 32'hFFFB7B94 , 32'hFFF9C50D , 32'hFFFF7EDE , 32'h0000A0B4 , 32'hFFF97306 , 32'h0001E7FC , 32'h00029C6E , 32'h00028E3A , 32'hFFFD7800 , 32'h00062048 , 32'hFFFCAEE1 , 32'hFFFF7D06 , 32'hFFFE9BC9 , 32'h0006AB75 , 32'h000ECED7 , 32'h000945F2 , 32'hFFF7B811 , 32'hFFF18CE0 , 32'hFFFAB6B6 , 32'h00028298 , 32'hFFFC483B , 32'h000088CC , 32'hFFF60ACB , 32'h00016451 , 32'hFFF9594B , 32'hFFFCF569 , 32'hFFFEAB00 , 32'h00059D02 , 32'h0003C3EF , 32'h0004E724 , 32'hFFFE980E , 32'hFFFF309A , 32'hFFFFB779 , 32'hFFFE2A83 , 32'hFFFF667C , 32'h00026477 , 32'hFFFEF5DC , 32'hFFFDA32C , 32'hFFF999DD , 32'h00072D8D , 32'hFFFB20A9 , 32'hFFF95871 , 32'hFFF9CC43 , 32'h0000D4AB , 32'h0005ECFE , 32'h00014265 , 32'hFFFBADCB , 32'h0003B6EE , 32'h00031639 , 32'hFFFEAB4F , 32'h0000CE41 , 32'h00040932 , 32'hFFFAB7BB , 32'h0000F69A , 32'h000A170D , 32'h0001F771 , 32'h000A0AA3 , 32'h000A45DC , 32'hFFFC04FE , 32'hFFFD0EAC , 32'hFFFFA966 , 32'h0001B2EC , 32'hFFFD4A82 , 32'h00005922 , 32'h0002E807 , 32'h0006A9AA , 32'hFFFFD397 , 32'hFFFF863C , 32'hFFF938E7} , 
{32'h000136CE , 32'h0005D19E , 32'h000337CE , 32'h000308AD , 32'h00086B0C , 32'hFFFFE2A0 , 32'h00061364 , 32'hFFFF1001 , 32'h00048061 , 32'hFFFFED9A , 32'h000553B7 , 32'hFFFF5855 , 32'h000270FC , 32'hFFFC9AB1 , 32'h000431E3 , 32'hFFFEA272 , 32'h000948F1 , 32'hFFFC5464 , 32'hFFFEF339 , 32'h00060793 , 32'h0000DC02 , 32'hFFFF9D7D , 32'h0005FC19 , 32'hFFFAFCAB , 32'h00042D24 , 32'h0001B6E1 , 32'hFFF6BC2B , 32'h0000EF95 , 32'h00016B22 , 32'h0003F789 , 32'h00004A33 , 32'hFFFDD038 , 32'h00075095 , 32'h00021EB5 , 32'h00030B45 , 32'hFFF84343 , 32'h00088890 , 32'h00037CB0 , 32'h0005C8A5 , 32'h0003EE48 , 32'hFFFDAFA8 , 32'h0002A63B , 32'hFFFEF3C5 , 32'h000920F1 , 32'hFFFF7101 , 32'h0004F74D , 32'hFFFDE4E3 , 32'h0001574E , 32'h000460EC , 32'hFFFD6D6E , 32'hFFFD956D , 32'h0000A6FD , 32'h00069299 , 32'hFFF97A44 , 32'h0003F64B , 32'hFFFEE654 , 32'h000835B5 , 32'hFFFB9F67 , 32'hFFFE1F5C , 32'h0000BD16 , 32'hFFFD9C98 , 32'h0004ADFF , 32'hFFF78727 , 32'hFFF7ACC9 , 32'h0001990D , 32'hFFFDB4DC , 32'h0004F4D8 , 32'h00040AD5 , 32'h000444D1 , 32'hFFFFBE1F , 32'h00011715 , 32'h00041C2F , 32'hFFFB151F , 32'hFFFFDDED , 32'h0005F7F4 , 32'hFFFDDD7E , 32'h00042BD6 , 32'h00083FF4 , 32'hFFF70685 , 32'hFFFD48EE , 32'h0003F11B , 32'h000A89DA , 32'hFFF6A020 , 32'h00051F7A , 32'hFFF65EBA , 32'h000791FC , 32'hFFFAF9D3 , 32'hFFFDEA9E , 32'h00002BF2 , 32'hFFFF453E , 32'h0004A294 , 32'hFFFD8942 , 32'hFFFB9210 , 32'h0000D5AE , 32'h000154FF , 32'hFFFEC622 , 32'hFFFFD273 , 32'hFFFD556B , 32'h0000F5AF , 32'hFFFD3650} , 
{32'h076B1240 , 32'h08C3C420 , 32'hEA8EE040 , 32'h08AE7050 , 32'h025A39EC , 32'h059E2900 , 32'hEFBD63E0 , 32'h0F6F9AD0 , 32'h05484620 , 32'h0ED462F0 , 32'h169BF640 , 32'h014D8C00 , 32'h13853AA0 , 32'hFEF0FF10 , 32'h049609B0 , 32'hFC440D2C , 32'hFF910761 , 32'h0B0A7170 , 32'h0A879530 , 32'h0D1FC990 , 32'h0F202A20 , 32'hFD328884 , 32'hFD0CFEB8 , 32'h03EA20C8 , 32'h009578AE , 32'h07A0ADB8 , 32'h0A178F50 , 32'h03013F70 , 32'hF1AF1EA0 , 32'h04F5DC18 , 32'hFAFE2A88 , 32'hF59BF340 , 32'h01AC84E4 , 32'hDF0F5380 , 32'hF677D2D0 , 32'h00349169 , 32'h0B64AA70 , 32'h0CD570D0 , 32'hFACF1A80 , 32'hFEA51038 , 32'hF8E7E760 , 32'hFC5D2F14 , 32'hF57FEE50 , 32'hE903B520 , 32'hFF6A1FDE , 32'hFE635188 , 32'h0B8CC2F0 , 32'hFCD4C4DC , 32'hFE4D3D1C , 32'h0A4417E0 , 32'h0A3A9360 , 32'hFC36D0FC , 32'h014FC8CC , 32'hFD267278 , 32'h03A6D390 , 32'h0EFCFE20 , 32'hF30438C0 , 32'h09838640 , 32'h07103FD8 , 32'h0113CCD0 , 32'hEE93A5E0 , 32'hFBF3A8C0 , 32'h01356050 , 32'h0034ECA8 , 32'h065B59F8 , 32'hF8DC0A38 , 32'hFC952EE0 , 32'hFD35B498 , 32'hFEDDC2EC , 32'h09C358F0 , 32'hFFF762FF , 32'h03051318 , 32'h03F39B1C , 32'h02E631EC , 32'hFBFB1B68 , 32'h041A8490 , 32'h0653BDB8 , 32'h01430140 , 32'hFB8D1DA0 , 32'hFC26DF70 , 32'hFF83E8F0 , 32'hFAF4E2E0 , 32'hF75E9DA0 , 32'h00748B75 , 32'h07C42CC8 , 32'h07513348 , 32'h0857F190 , 32'hFBF92328 , 32'h05A97960 , 32'hFE9E2688 , 32'hFFFDC1A0 , 32'h00048D1F , 32'hFFFBBFB8 , 32'h00008612 , 32'h00029C82 , 32'hFFFEC0B2 , 32'h00024674 , 32'hFFFC3626 , 32'h0001563D , 32'hFFFF311C} , 
{32'h00076405 , 32'hFFF9DCA0 , 32'h00006A59 , 32'h0008025A , 32'hFFF9B66B , 32'h0000A148 , 32'hFFFCB115 , 32'h0002BC50 , 32'hFFF71655 , 32'hFFF85C64 , 32'hFFFE31F9 , 32'h0001B304 , 32'h000A02E2 , 32'h0001BAC9 , 32'h0004AE9F , 32'h0007C2CA , 32'hFFFD4F39 , 32'hFFFFA3B6 , 32'hFFFF32CE , 32'hFFFFC919 , 32'hFFFE88D5 , 32'hFFFCD6AE , 32'h00040929 , 32'h0000DA53 , 32'h000556AB , 32'hFFF96A97 , 32'h000467A4 , 32'h00000350 , 32'h000482BE , 32'h0006E60D , 32'hFFFCD2A6 , 32'h0003FA91 , 32'hFFFDC41A , 32'hFFFDBC23 , 32'h00008E7D , 32'h000598EE , 32'hFFFFA853 , 32'h00032948 , 32'h00021F0D , 32'h0005861D , 32'h0003A379 , 32'hFFF97E26 , 32'h0000DA9E , 32'h00041357 , 32'h00015DF1 , 32'hFFFD7113 , 32'h000901F8 , 32'hFFF9289E , 32'hFFFFB607 , 32'hFFFE41C0 , 32'hFFFB59A4 , 32'h0000B40F , 32'h0005A964 , 32'hFFFABAC2 , 32'h0003D323 , 32'hFFFF17AC , 32'hFFF378B8 , 32'hFFF83ADB , 32'hFFFFC334 , 32'hFFF00B88 , 32'h0000007B , 32'h00041BC8 , 32'h000882C2 , 32'h0001F600 , 32'h0003A21E , 32'h0000CC4F , 32'hFFFE3626 , 32'hFFFD6DD2 , 32'h00010ED6 , 32'hFFFD4DC1 , 32'hFFFB306A , 32'h00048D41 , 32'h0000AC84 , 32'h00021653 , 32'h00001484 , 32'hFFF95549 , 32'hFFF61B3F , 32'hFFFD6443 , 32'hFFFD7F64 , 32'h0003E328 , 32'hFFFA98AA , 32'h000200A8 , 32'h000654EB , 32'h0003868D , 32'h00018171 , 32'h0003EFDA , 32'hFFFEFB56 , 32'hFFF898ED , 32'h0000DA12 , 32'hFFFDD611 , 32'hFFFA1855 , 32'h000662B9 , 32'hFFFFCC8F , 32'h00062A60 , 32'hFFFA0E79 , 32'hFFFDAF8F , 32'hFFFF13F2 , 32'h0002E3CF , 32'h000445DA , 32'hFFF7D3ED} , 
{32'h00011E3D , 32'hFFF6DF5D , 32'hFFFAF951 , 32'hFFFEB400 , 32'h00045EFC , 32'hFFFCB1B4 , 32'h0000CDB0 , 32'h0003047C , 32'h000541FE , 32'hFFFC9E61 , 32'hFFFFBE23 , 32'hFFFE382B , 32'hFFFC17DD , 32'hFFF8AEFD , 32'h00027EF0 , 32'h00007201 , 32'hFFF97D58 , 32'h00041A2A , 32'h0000BC70 , 32'h0006D145 , 32'h00005708 , 32'h00035E29 , 32'h0001701E , 32'hFFF4D854 , 32'hFFFE6F5C , 32'h00054DC4 , 32'h000571AB , 32'hFFFAEEBC , 32'hFFFB2537 , 32'h00009FAA , 32'h00034EFC , 32'h000AEA37 , 32'h00044E2D , 32'hFFFEB2C2 , 32'h0004B0CA , 32'h00009ECA , 32'hFFFFF543 , 32'hFFFAFA29 , 32'h0004C840 , 32'h000BE311 , 32'hFFFE0D40 , 32'h0001686C , 32'hFFFF70D5 , 32'h00009813 , 32'hFFFE9A84 , 32'hFFFD0621 , 32'h0003855A , 32'hFFFD61D5 , 32'hFFF6B145 , 32'hFFFFCAF5 , 32'hFFF74FB5 , 32'h00056604 , 32'hFFFAD6C5 , 32'hFFF555A8 , 32'hFFF744E9 , 32'hFFFC889A , 32'h00007516 , 32'hFFFD2D43 , 32'h00007D86 , 32'h000733A1 , 32'h0005ECC2 , 32'hFFFCCE16 , 32'hFFFE4861 , 32'h0003BDE6 , 32'h0003276F , 32'hFFFAECED , 32'hFFFB2B0D , 32'hFFFE683E , 32'hFFF5A39D , 32'hFFF9B320 , 32'hFFF57312 , 32'hFFFE158F , 32'h000119EA , 32'hFFF97F98 , 32'h0001B209 , 32'h000073CA , 32'h0007BA6F , 32'hFFFB49CA , 32'h000A30EE , 32'h0007EDCC , 32'h000222D2 , 32'hFFFF8944 , 32'h00000976 , 32'hFFFF9D6D , 32'hFFFF7317 , 32'h00066CB1 , 32'hFFFB701D , 32'h000039B8 , 32'hFFFE53E0 , 32'h00021807 , 32'h000AE75C , 32'hFFFC3CF2 , 32'h000883D7 , 32'hFFFCDAFF , 32'hFFF6DE7F , 32'hFFFFE73F , 32'h0009F0DA , 32'h00087260 , 32'hFFFE3185 , 32'h00037844} , 
{32'h0FF343D0 , 32'hEA4D15A0 , 32'hF2D6C2A0 , 32'h1612CE20 , 32'h09FAE110 , 32'hDE512400 , 32'hE254B5A0 , 32'hF9E22CD8 , 32'h0CAEB970 , 32'hE5FBB8E0 , 32'h08F28990 , 32'hF2A50D00 , 32'h1B5DB380 , 32'hF4417A00 , 32'h11D804E0 , 32'h0D23CB30 , 32'hFC24C914 , 32'hFE6E09D8 , 32'h002E72D0 , 32'h051A5F38 , 32'hF057CA00 , 32'hFD1F4D00 , 32'hF9583B10 , 32'h0EADD3E0 , 32'hFF5189E1 , 32'hFF5A3D11 , 32'h0A9AA9B0 , 32'hE7734FE0 , 32'hFD21A5FC , 32'hE06EE8E0 , 32'h03A3857C , 32'h0F967980 , 32'hF815D010 , 32'h0151F41C , 32'hE39F04A0 , 32'hFAF8B028 , 32'h04CEABB8 , 32'h0A1DAC90 , 32'h0B462C70 , 32'h00762C36 , 32'h10169E80 , 32'hFF36D676 , 32'hFB765090 , 32'h04DC9C18 , 32'hF5B09B00 , 32'hFE997E04 , 32'hFE55B630 , 32'hFAE980F8 , 32'h0FB80D90 , 32'hFB660158 , 32'h12EE5CE0 , 32'h123DCE40 , 32'h070E3790 , 32'h066BF268 , 32'hFB908FC8 , 32'hF0C89000 , 32'hFE7A3EBC , 32'hF5EF91A0 , 32'hF8CCDAE8 , 32'hF322D6A0 , 32'h02F0BB2C , 32'h0A35F120 , 32'h00A6000C , 32'h02502F18 , 32'hFE0337C4 , 32'hF3AA41B0 , 32'hFF030B0B , 32'hFBF92E98 , 32'h023C4E28 , 32'h030F4D38 , 32'h048C2398 , 32'hFD547344 , 32'h0B6F67C0 , 32'hF7C3FB40 , 32'h0AEEB430 , 32'hFD63DAE4 , 32'hFA98D3B0 , 32'hF73F4000 , 32'h0C20AA70 , 32'hF29AEE30 , 32'h00155177 , 32'hFD36A6AC , 32'h016C6320 , 32'hF23CBDE0 , 32'hF5447EE0 , 32'hFF17D355 , 32'hFFC0E0AE , 32'hF979EEB0 , 32'h0689FD50 , 32'hFF41454B , 32'h0002B35C , 32'h00048214 , 32'hFFFE1BFB , 32'h0001CB4F , 32'h0000EEF3 , 32'hFFFF3428 , 32'h00032D30 , 32'hFFFFC45F , 32'hFFFE093F , 32'hFFFF89B0} , 
{32'hFE3C2B3C , 32'hD3401800 , 32'h87F62E80 , 32'hB3DC4400 , 32'h32FCCE80 , 32'hFD2C451C , 32'hF7232AE0 , 32'hE6DF7820 , 32'hECB5DCE0 , 32'hF3ABEE40 , 32'hCA996580 , 32'hF1361880 , 32'h1AB345C0 , 32'h079EF7A8 , 32'hF82C0C40 , 32'hF24B23A0 , 32'h01C6D85C , 32'h11059600 , 32'h2DC1EF40 , 32'h18F3C0E0 , 32'hD396C100 , 32'h09EA9F50 , 32'h1292A080 , 32'h07F984B8 , 32'hE5BD8D80 , 32'h040E2260 , 32'hEB1C2820 , 32'hFB564C30 , 32'hC582BE00 , 32'hF5BC74C0 , 32'hF09C4CB0 , 32'h00A109A6 , 32'h0B2B4270 , 32'hDC4E9F00 , 32'hF60B5680 , 32'h25C27240 , 32'hFEADB600 , 32'hE7F77A80 , 32'h19F48EE0 , 32'hFD96EB94 , 32'h17AD8B60 , 32'hE582F6C0 , 32'h00753B03 , 32'hF9B9C478 , 32'h01F8FCEC , 32'hF8ABDEA8 , 32'h0765F1D8 , 32'hF20F2CC0 , 32'h1E72F640 , 32'hF4ED7B50 , 32'hFA31E368 , 32'hF71C4FD0 , 32'h0591AF30 , 32'h0ED015B0 , 32'h0FDA2370 , 32'h2523C6C0 , 32'hFD51323C , 32'h142A8780 , 32'hF66CBEE0 , 32'hFAECE938 , 32'h08B5F030 , 32'hFFFA55F6 , 32'h076A4BB8 , 32'h0867B860 , 32'h0CB826B0 , 32'hF2B85690 , 32'h0154B3A0 , 32'h0461D910 , 32'h0177EC6C , 32'h11D0E560 , 32'h0E199570 , 32'hFAE0EE50 , 32'hFDE780F4 , 32'hF9F90958 , 32'hFC7C1978 , 32'h024AC974 , 32'hFE634068 , 32'h00515367 , 32'h012DF450 , 32'h011FBF04 , 32'h014D7B54 , 32'hFD831038 , 32'h0655CD38 , 32'h02078294 , 32'hFA7C2448 , 32'h0023E46E , 32'h05398B88 , 32'h043A2B08 , 32'hFC92C210 , 32'h0160EC80 , 32'hFFFF3CA8 , 32'hFFFE8901 , 32'h00012DB7 , 32'h0002588F , 32'h0003AC20 , 32'hFFFDBF28 , 32'h000320BF , 32'hFFFF13A5 , 32'h000017B3 , 32'h0002793F} , 
{32'h0002EBE2 , 32'hFFFC3741 , 32'h00060CB4 , 32'h0000C467 , 32'h0004A793 , 32'h000B21DA , 32'hFFF8DAE8 , 32'h0000E0F4 , 32'h000198F7 , 32'h00088438 , 32'h00005188 , 32'hFFFAC60E , 32'hFFFD8ED0 , 32'hFFFD7951 , 32'hFFFD0F59 , 32'h0006C745 , 32'h0000A1ED , 32'hFFFA1848 , 32'hFFF70107 , 32'hFFFF4198 , 32'h00081A64 , 32'hFFFFDBA9 , 32'hFFFF8AF2 , 32'h00018A46 , 32'h0003A0D3 , 32'hFFFE8308 , 32'hFFF6FBEA , 32'hFFF89B2F , 32'h0001BBA0 , 32'h0000B4F2 , 32'hFFF7A9A2 , 32'hFFFB434A , 32'h0005569A , 32'hFFFD8090 , 32'h000169C9 , 32'h000004D0 , 32'h000149AA , 32'h000169B0 , 32'hFFFC68F3 , 32'h00078121 , 32'hFFFD3128 , 32'hFFFBC700 , 32'h0000323B , 32'h0006D45A , 32'h00029DEB , 32'hFFFC21FB , 32'h00043ADC , 32'h0001FA0A , 32'hFFFB4496 , 32'hFFFED11B , 32'h00028E2B , 32'hFFFD0EA0 , 32'h000210A0 , 32'h0002B377 , 32'hFFFEB80F , 32'h0003A57E , 32'h00031F88 , 32'h00027304 , 32'h00033910 , 32'hFFFF3001 , 32'h00006340 , 32'hFFFFD893 , 32'hFFF6FF9A , 32'hFFFE0564 , 32'hFFFDF2DC , 32'hFFFE4361 , 32'h0001D013 , 32'hFFFA1F1F , 32'h0000EF24 , 32'h000BD6E2 , 32'hFFFCE2BC , 32'h0002E6E6 , 32'h00053491 , 32'hFFFC9740 , 32'hFFFF65A3 , 32'h00044CB9 , 32'hFFFD3D3B , 32'hFFFA28E1 , 32'hFFFB4FAC , 32'h00002BF4 , 32'hFFFFC7C6 , 32'h0004514F , 32'hFFFB844F , 32'hFFFBF818 , 32'h0003C6CA , 32'h00037620 , 32'hFFFF52F8 , 32'hFFFC8F29 , 32'h00004E5B , 32'h000494F8 , 32'hFFFD4B8E , 32'h0006B51F , 32'h000753CD , 32'hFFFCF82F , 32'hFFFD6970 , 32'h0004BE99 , 32'hFFF3DF89 , 32'hFFFB0830 , 32'hFFFBC2F4 , 32'hFFFEE438} , 
{32'h9E98AB80 , 32'h7FFFFFFF , 32'h0DCA3050 , 32'h07B335E8 , 32'h019CE444 , 32'hF71740B0 , 32'h3F7A5400 , 32'hF34A2A00 , 32'h1EB05AC0 , 32'hD7261D00 , 32'hD096C900 , 32'hE52E0280 , 32'hDB133600 , 32'h33F01600 , 32'h2677A0C0 , 32'h03B8D51C , 32'hC502A080 , 32'hFA8ACED0 , 32'h0961B250 , 32'hD0B27440 , 32'hF6107190 , 32'h09A17FF0 , 32'h16DC4F20 , 32'h212826C0 , 32'h35357840 , 32'h06F01220 , 32'hF7156850 , 32'hF7B2FA70 , 32'hE9A18C80 , 32'h10EB1A60 , 32'h026DC78C , 32'hF9A041E8 , 32'h080B39A0 , 32'h012AC2DC , 32'h1B2A42E0 , 32'hEC415AA0 , 32'hF8226CF0 , 32'h187B0FA0 , 32'h04254158 , 32'h0A9AB850 , 32'hF42B9DC0 , 32'h07A257E0 , 32'h07140810 , 32'hFCF22AC0 , 32'h04B72B88 , 32'h15FF94A0 , 32'h0516FD88 , 32'hF824D318 , 32'hF708BF50 , 32'hFC207004 , 32'h07604DF0 , 32'h07FFA780 , 32'h02BE9A98 , 32'h015CC480 , 32'hF0C561A0 , 32'h0EB03AD0 , 32'hF0A2FB10 , 32'hFD84C38C , 32'h046DC400 , 32'hE90476C0 , 32'hEBACF5E0 , 32'hF911EB70 , 32'h018EC4A8 , 32'hF8118838 , 32'h085DCFE0 , 32'h09F1C9B0 , 32'h03793AE0 , 32'h00EF7C5B , 32'h02ECE994 , 32'h07A71940 , 32'h083C0050 , 32'hF97D6568 , 32'hF42FB1B0 , 32'hF4E92770 , 32'hF852CFF0 , 32'h01C26B7C , 32'hFFEEEE0F , 32'h09E206D0 , 32'h029A1D98 , 32'hFFA426FB , 32'hF8868AC0 , 32'h0BBC6C40 , 32'hFC48BA90 , 32'h01F9A728 , 32'h0007E47B , 32'h01172D10 , 32'hFF3083E1 , 32'h011FF5AC , 32'hFE97AC40 , 32'h00F48F6C , 32'hFFFD2649 , 32'h00003152 , 32'hFFFD2863 , 32'hFFFFA8DB , 32'h00003222 , 32'h0002F3EF , 32'hFFFE1711 , 32'h0001A8AF , 32'hFFFF6601 , 32'hFFFC10A1} , 
{32'hF0E148A0 , 32'h224EA840 , 32'hF89E21B0 , 32'h09569A00 , 32'h0ED242B0 , 32'h0E138050 , 32'h0CF27A40 , 32'hF5F8F720 , 32'hFB1E6B28 , 32'h0AF5AEA0 , 32'hFC3B7E40 , 32'h0000ED0D , 32'hD5306D00 , 32'h007B151F , 32'h0835E340 , 32'h0B49B960 , 32'hFDD98C94 , 32'h12ED9E80 , 32'h0CD2A5C0 , 32'hF0A68030 , 32'hF423B9E0 , 32'h058014A0 , 32'h11DAF9A0 , 32'hF2063750 , 32'hFBC9E150 , 32'hEEC42BE0 , 32'hF8398818 , 32'h0D571D80 , 32'hFD58DDFC , 32'h102079C0 , 32'h0F418420 , 32'hFAB1B150 , 32'hFD8B8CC0 , 32'hF3D5B360 , 32'hFD3AAD24 , 32'h1608A780 , 32'h08FD88B0 , 32'h09672780 , 32'hFC9125F4 , 32'h1288B1A0 , 32'h02269110 , 32'hFBCC0B30 , 32'h026475D8 , 32'h07F3D920 , 32'hFC51DFC0 , 32'h003F05B0 , 32'hF3F33A90 , 32'h04A27B88 , 32'h00C83A05 , 32'h06A1B908 , 32'hFC72A12C , 32'hF086D150 , 32'hFCFFB484 , 32'hEBA635A0 , 32'hF5CE5530 , 32'h045F4C40 , 32'h006AB1A6 , 32'h08AA78E0 , 32'hFCCBEB24 , 32'hF5EF0C80 , 32'hEE5EE380 , 32'h022F42C8 , 32'hEE8D6300 , 32'hF7845780 , 32'h0E935C80 , 32'h05F75728 , 32'hF535FD90 , 32'hF247FB10 , 32'h06F86768 , 32'h037DD428 , 32'hFA1B3478 , 32'hF5BC8F00 , 32'hF7683ED0 , 32'h031213FC , 32'hF96B6CE8 , 32'h02C5CC0C , 32'h0D471830 , 32'h02383E80 , 32'h0583D048 , 32'h019820F8 , 32'h05D28C20 , 32'h034549E8 , 32'hFECFED98 , 32'h07517370 , 32'hFA5EC048 , 32'h0872BD40 , 32'hF6BC3AC0 , 32'h020882C8 , 32'hFE786F08 , 32'hFEC5C1D4 , 32'h00042B35 , 32'hFFFB4BBA , 32'h00022F95 , 32'hFFFF5974 , 32'h000612B1 , 32'h00030C05 , 32'hFFF9EB77 , 32'hFFFF4E19 , 32'h0000EB48 , 32'h000152BF} , 
{32'h08C61DF0 , 32'hFD83A200 , 32'hDDF41100 , 32'hE64C7240 , 32'h022E0384 , 32'h0457DED0 , 32'h20F66BC0 , 32'hDDA45840 , 32'hEA088CA0 , 32'hF3A5ADB0 , 32'h128385A0 , 32'h195B81A0 , 32'hE472C500 , 32'h12E74EA0 , 32'hF9397A70 , 32'hFB950FC0 , 32'h191BDDA0 , 32'hE9377860 , 32'h042FDAB8 , 32'hFD656930 , 32'h23DC91C0 , 32'h0FE750B0 , 32'hFD88A7C8 , 32'h1A385100 , 32'h1AD76A80 , 32'h03833C10 , 32'h05B14900 , 32'h30584D40 , 32'h0FD69420 , 32'h02D55C74 , 32'hFB56BBD0 , 32'hFD40941C , 32'hFAE29790 , 32'hFD9AF8E4 , 32'h0D8982E0 , 32'h01CFEB28 , 32'h03C8E100 , 32'hDE3CEF80 , 32'hF5A78670 , 32'hF82A0EB8 , 32'hFCA7A738 , 32'h018AB44C , 32'h0A3C18B0 , 32'h2D8D63C0 , 32'hEB431F20 , 32'h05356540 , 32'hFD146BE4 , 32'hF8D6D510 , 32'h0E548710 , 32'hF1AEC4B0 , 32'hF396A690 , 32'h04DFEE00 , 32'hF8FFB9D8 , 32'hFED1F9F0 , 32'hF4D691D0 , 32'hEC276780 , 32'hFECD8C3C , 32'hF6CFB450 , 32'h04558CF0 , 32'hFA9BCFD0 , 32'h0322E7E8 , 32'hFD176B8C , 32'hF7E02780 , 32'h071F2940 , 32'h06600D20 , 32'hFD1B5AC4 , 32'h07EC5BC8 , 32'h068DD570 , 32'hFEFA397C , 32'hF47B40E0 , 32'h0DD46360 , 32'hFE35A7D8 , 32'h131F5B20 , 32'hFD5F603C , 32'hFD0638C8 , 32'hFFB5B97A , 32'h036CAB30 , 32'h0A7EF8F0 , 32'h066C70D0 , 32'h0137E158 , 32'hFEAAB5C8 , 32'hFC6E5D94 , 32'h01B848D4 , 32'hFD127ABC , 32'h010DF22C , 32'hFBCCD208 , 32'hFF5DE2B3 , 32'h019D864C , 32'hFBC624A8 , 32'h0165A20C , 32'hFFFC63EF , 32'h000218A2 , 32'hFFFFB6C6 , 32'hFFFC10F6 , 32'hFFFDB1F9 , 32'h000310E3 , 32'h0000573B , 32'hFFFF8850 , 32'h0003A3AF , 32'hFFFEC19F} , 
{32'hD672B8C0 , 32'h014A6A64 , 32'hC0AFA680 , 32'h283BE0C0 , 32'hB4F6E880 , 32'h29718500 , 32'hFB356298 , 32'h2A3B1A00 , 32'hF7C17C60 , 32'h0A0C8A40 , 32'hFD33108C , 32'hFE15BE8C , 32'hF67E7300 , 32'h1F38A540 , 32'hFB25A2E8 , 32'hF04C8D60 , 32'hDBFF2EC0 , 32'hDF946280 , 32'hFA4B5BE0 , 32'h1D10B4A0 , 32'hE21D7BC0 , 32'hEAD94B40 , 32'h0767C0C0 , 32'hE6680D40 , 32'hF4870DF0 , 32'h00F3A195 , 32'hFDE6A3E0 , 32'hF579F7B0 , 32'hF5082E20 , 32'h02D0A9E0 , 32'hF213B0C0 , 32'h1C12D020 , 32'h06B3B1B0 , 32'h056E8CE0 , 32'h01DE53E0 , 32'h136BA160 , 32'hE5BA0D20 , 32'h01D6CCA0 , 32'h037F1B8C , 32'hF0F18280 , 32'hDAE40B00 , 32'hFD048224 , 32'h05A8CD60 , 32'h20196940 , 32'hEAEA5EA0 , 32'h0A2F3D30 , 32'h17896180 , 32'h0D2283C0 , 32'hF46F8D70 , 32'h09DB7A70 , 32'h0787C740 , 32'hFEABEDA0 , 32'hE5538960 , 32'hF81C5190 , 32'h100A0580 , 32'hFAEC4C10 , 32'hF39EDBC0 , 32'h014E5504 , 32'h02A7EA7C , 32'hFBFA1F50 , 32'h00C3DD3E , 32'hFFA14041 , 32'hF2606600 , 32'hFC9E6460 , 32'hF8B7F370 , 32'hEFC374C0 , 32'h1330FD00 , 32'h0E142310 , 32'hFD86A71C , 32'hFBCC7518 , 32'h02C33358 , 32'h026EB6EC , 32'h011AF950 , 32'hF6F50860 , 32'hF7D1F8D0 , 32'h0033A3B6 , 32'h057E39D8 , 32'hF6F741B0 , 32'h0770FAF0 , 32'hFB0DC0A8 , 32'hFA054758 , 32'hFFAAFF0F , 32'h035B7440 , 32'hFF45F84C , 32'hFD610040 , 32'h01E9C6E8 , 32'hFD5CC220 , 32'hFE83B448 , 32'hFD243A48 , 32'h0149FA28 , 32'h0000697D , 32'h0004C7E4 , 32'h0000CEF0 , 32'hFFFDEAE3 , 32'hFFFFF8F1 , 32'h00021105 , 32'h0002C75C , 32'hFFFC8658 , 32'h0001036C , 32'hFFFF2032} , 
{32'hFFFC2787 , 32'hFFF96E71 , 32'hFFFC34D8 , 32'h00048FFF , 32'h0002A3B4 , 32'hFFF9B23A , 32'hFFFE7402 , 32'h0002D32F , 32'h000353C2 , 32'h00056C89 , 32'h0005B1EB , 32'hFFF551A8 , 32'hFFF88A7B , 32'h0003B6EA , 32'h00044BF8 , 32'h00059222 , 32'hFFFC68F8 , 32'hFFF8E675 , 32'hFFFE7237 , 32'h0000E8F2 , 32'hFFFA9050 , 32'h00062523 , 32'hFFFA90F2 , 32'h00038FAA , 32'h0004AB9C , 32'h000185BB , 32'h0004EB5E , 32'hFFFF8B6C , 32'h00010B0D , 32'h00049C68 , 32'h0004370F , 32'h0000D4E9 , 32'hFFFD662B , 32'h0002DB95 , 32'h000242BD , 32'h0001D101 , 32'h000031C5 , 32'h00022926 , 32'hFFFB7BB1 , 32'hFFFDFC51 , 32'h0004B23B , 32'hFFFECF6B , 32'h0000DBC5 , 32'hFFFEAA15 , 32'hFFFC3EA5 , 32'h0001BEE8 , 32'h0000DCC4 , 32'h000211A0 , 32'h000635CF , 32'h00098935 , 32'h00025964 , 32'h0005E540 , 32'h00013A3E , 32'h0007C4BF , 32'hFFFA0479 , 32'hFFFBAD8E , 32'hFFFB36AA , 32'h00098A04 , 32'hFFFECB2E , 32'h0000D351 , 32'h000406B0 , 32'hFFFEB921 , 32'hFFFB8C1B , 32'hFFF81B2F , 32'hFFFECC36 , 32'h0002F580 , 32'h00020C13 , 32'hFFFA0A96 , 32'hFFFDED44 , 32'hFFFEBB70 , 32'hFFFF6889 , 32'hFFFCDEA7 , 32'h00037D6D , 32'h0004F40E , 32'h0008714D , 32'hFFFA64FB , 32'h0000D542 , 32'h0001B4C6 , 32'hFFFCFF0A , 32'h00029965 , 32'h000053B3 , 32'h00049B87 , 32'hFFF8EA8D , 32'hFFFE5B26 , 32'h00023094 , 32'hFFFFC917 , 32'hFFFCA6AD , 32'h0000ED72 , 32'h0006CD88 , 32'h000077A9 , 32'h0001CE7B , 32'h00075989 , 32'h0003598A , 32'h0005A98D , 32'hFFFE392A , 32'h0000E0F9 , 32'hFFFCC45D , 32'h0006F92A , 32'h0002F0B7 , 32'hFFFFDC09} , 
{32'h13810CA0 , 32'hF3895ED0 , 32'hF3168B30 , 32'h1944A740 , 32'hCBCB0E80 , 32'h1A9A7920 , 32'h10CF8500 , 32'h0C660B60 , 32'hFB6B51F0 , 32'hF802B860 , 32'h09E862D0 , 32'hF4D93BB0 , 32'h0A93C4E0 , 32'hFF14B160 , 32'h0DA1C630 , 32'h1D05EF60 , 32'h0E3CB0E0 , 32'hD62727C0 , 32'h0DC7E960 , 32'h15338780 , 32'h14459620 , 32'hF5B181B0 , 32'hFEFC73C4 , 32'h048B6E10 , 32'hF1FAB0E0 , 32'h05EF67E8 , 32'hF2F9C220 , 32'hFBC95770 , 32'h00310099 , 32'hE2595F00 , 32'hFCEB1450 , 32'hFFCC05D2 , 32'h10ACD500 , 32'hF2AFA2B0 , 32'h0C6C0CC0 , 32'hFC90C42C , 32'h0751B848 , 32'h1F3FCAA0 , 32'h1BEA2520 , 32'h07574140 , 32'h2679AF40 , 32'hFC3695D8 , 32'h0499C5D0 , 32'h06CD6290 , 32'hFCB0EF14 , 32'h06217148 , 32'hF0DBC4E0 , 32'hF6439590 , 32'hF5C2AEE0 , 32'hE8C50300 , 32'hFD50A5A4 , 32'hEF574EC0 , 32'hFED664DC , 32'h179196A0 , 32'hFA2BFD68 , 32'h11A1FEE0 , 32'h002AFD0E , 32'hF77EA6B0 , 32'h0427B848 , 32'hF94AA390 , 32'hFD3217AC , 32'hF694E920 , 32'h04255F40 , 32'h06DAFCD8 , 32'hF9D47200 , 32'h1DB55CA0 , 32'hF8E7D268 , 32'hF5F398B0 , 32'h068EB590 , 32'h07AB8C98 , 32'hFAC4B9A8 , 32'hF95DF590 , 32'hF1E639D0 , 32'h02EC1660 , 32'hFFE3319A , 32'hF6ABC650 , 32'h04C42A90 , 32'hF24335A0 , 32'h0A9ECAF0 , 32'hFE925DDC , 32'h0306D9A8 , 32'hFD64B6AC , 32'h0582C7C0 , 32'hFBF4DCD8 , 32'h0187F8EC , 32'hF6D20420 , 32'h0184C7A8 , 32'hFFBEBF88 , 32'hFCB66DD0 , 32'h013B8B90 , 32'h000228F0 , 32'h0006695A , 32'h00010EEA , 32'h0004303B , 32'hFFFF45F3 , 32'h0001BAC6 , 32'h0002CC93 , 32'hFFF9B3BB , 32'h00013C57 , 32'hFFFDF235} , 
{32'h282C65C0 , 32'h16850AA0 , 32'h395C8200 , 32'h186E08E0 , 32'h21F02C00 , 32'hC005B880 , 32'h1D3731A0 , 32'h2B1191C0 , 32'hD349FB00 , 32'hD47E1C40 , 32'hF20C1150 , 32'h2088A040 , 32'hE9A4A940 , 32'hF11C46A0 , 32'h0E4D13D0 , 32'hE4A7D360 , 32'hF9E09648 , 32'h16AEA280 , 32'hFC15CAF8 , 32'h087275B0 , 32'hE5CCE360 , 32'h2EEAB380 , 32'h05897AF8 , 32'hE60E6200 , 32'h114E9D20 , 32'hF0183CF0 , 32'h01B08F94 , 32'h2D2FCC00 , 32'hEDF715E0 , 32'h14A15920 , 32'hEC93DFA0 , 32'h19D0F720 , 32'hFBE94E70 , 32'h1A6FB4A0 , 32'h1450A960 , 32'h143B6DE0 , 32'hFE14D178 , 32'h04945000 , 32'h2501C5C0 , 32'hE23AF200 , 32'h0CB3B4A0 , 32'h066FE940 , 32'hDFFF8EC0 , 32'hF61BA9C0 , 32'h0AF8D000 , 32'hE9C49DA0 , 32'hF5633F80 , 32'h07583690 , 32'hEF39B000 , 32'h032BDB04 , 32'hFEFD8F1C , 32'hEFE9FE80 , 32'hF4720B00 , 32'hF10E4F40 , 32'h09C89300 , 32'hFC4FF28C , 32'h0A0FE490 , 32'h00EF232A , 32'hEB08E600 , 32'hFC6A9DAC , 32'hE5A2C940 , 32'hF2FCF9F0 , 32'hFBA3C958 , 32'h045D0770 , 32'hFCACD87C , 32'h0B34FD80 , 32'hFA1038B0 , 32'hFBFA9518 , 32'hEF6FC260 , 32'hFB314028 , 32'h061C6DF8 , 32'h0D072220 , 32'h09F9ADB0 , 32'h0B5FE250 , 32'hF3BD3670 , 32'h0D8B1820 , 32'hF675A340 , 32'hFF377BD6 , 32'h00BC39B9 , 32'hFA244F40 , 32'hF8453CF0 , 32'hFF4B4537 , 32'h0185972C , 32'hFFDD051A , 32'h02324D70 , 32'hFFADA7F9 , 32'h023EF684 , 32'hFE0E1D18 , 32'hFC50A434 , 32'hFF7666B4 , 32'h000210FC , 32'hFFFCD658 , 32'hFFFFB124 , 32'h00064A67 , 32'h0001220C , 32'hFFFE4430 , 32'h00024506 , 32'hFFFE4BD9 , 32'h00017DDD , 32'h00014DE6} , 
{32'hF67D4230 , 32'hFC20EDC0 , 32'hF3D7D8A0 , 32'h1A0C89C0 , 32'hF9612398 , 32'h02B12910 , 32'hF5391A60 , 32'hEE3FCA40 , 32'hF131E7E0 , 32'h05B79088 , 32'hEC09BC60 , 32'hFC048A08 , 32'h0F34DED0 , 32'h003E0CDC , 32'hF31DD9F0 , 32'hF6ED1330 , 32'h07E8EBD0 , 32'h12F559A0 , 32'hF0B07BA0 , 32'hFCB936B0 , 32'hF4A0D540 , 32'h00174E88 , 32'hFF50825F , 32'h0FC83D00 , 32'h049A88E8 , 32'hFABA26B8 , 32'hF4E42460 , 32'h0A56B420 , 32'h00EC3A27 , 32'h01141904 , 32'hFB462AB0 , 32'h032EA830 , 32'hFC0F956C , 32'hF710AF80 , 32'hEDC058A0 , 32'h03996800 , 32'hF9A41078 , 32'h18343DE0 , 32'hF600BB80 , 32'hDFF734C0 , 32'h0FBFB140 , 32'hFAE461E8 , 32'h0743B960 , 32'hF92D6BD8 , 32'hFDF46B64 , 32'hFB1027B0 , 32'hFE99DD74 , 32'hFBC39E20 , 32'h0509FA78 , 32'h0239A388 , 32'h0B354450 , 32'hF81F17F0 , 32'hFF768187 , 32'hFE0CE1AC , 32'hFD0837C8 , 32'h01D34A94 , 32'h09FE6480 , 32'hFDF7567C , 32'h0C262050 , 32'h0400EC88 , 32'h0AF5ADE0 , 32'hF6A13BC0 , 32'hFE6C206C , 32'hFA8ECAD8 , 32'hFA5FDBF8 , 32'hFF0E0778 , 32'hFEB94C94 , 32'hF7773650 , 32'hFCEC6664 , 32'hFA7759F0 , 32'hFA2603D8 , 32'hFD948190 , 32'hFA9C84F8 , 32'hF80647F8 , 32'hF44F7E50 , 32'h0BD1F950 , 32'h00CFCEFC , 32'h07B02C58 , 32'hFD911AA0 , 32'h02F59F0C , 32'h00AB8DF8 , 32'hFA7A30A8 , 32'hF9CEC978 , 32'h0346B1A4 , 32'hFF88D008 , 32'h013A51D4 , 32'h010B1438 , 32'hF9086DA8 , 32'hFD296590 , 32'h004B2B83 , 32'h00014BE9 , 32'h00081F25 , 32'hFFFFA311 , 32'h0000D6AE , 32'hFFFE3218 , 32'h00028A48 , 32'hFFFD54D0 , 32'h000073A9 , 32'h00004196 , 32'h000156E5} , 
{32'hFFFFBB89 , 32'hFFFA339F , 32'h0001650A , 32'hFFFBD1EA , 32'hFFFF64AC , 32'hFFFF294D , 32'h00015A2B , 32'hFFF4F540 , 32'h00043DA1 , 32'hFFFBC876 , 32'hFFFEE334 , 32'hFFFECA83 , 32'hFFFB3E0E , 32'hFFFFA2AE , 32'hFFFD6760 , 32'h00010F7F , 32'hFFFCD9AC , 32'hFFFBDEFC , 32'hFFFB3A65 , 32'h0002BE4B , 32'hFFFBEAA3 , 32'h00036A56 , 32'h00026288 , 32'h0002414C , 32'hFFFC5439 , 32'hFFFC2039 , 32'h00031BA0 , 32'h0006B0A1 , 32'hFFFA1033 , 32'h0004BECB , 32'h000241D5 , 32'hFFFA2C0C , 32'hFFFF6EC0 , 32'hFFFF08D9 , 32'h0001C884 , 32'hFFFCC136 , 32'h00008D88 , 32'hFFF54974 , 32'hFFF8DC2E , 32'hFFF9064F , 32'h0003164C , 32'h00047702 , 32'h0006BF4E , 32'h0001EE6A , 32'hFFF99330 , 32'h00025377 , 32'hFFFF3125 , 32'hFFF88761 , 32'hFFFC50B5 , 32'hFFFBD665 , 32'h000110C5 , 32'hFFFEBAE9 , 32'h0000383F , 32'hFFFD43B1 , 32'h00080633 , 32'h00038630 , 32'h0001179C , 32'hFFF84A75 , 32'hFFFDDC05 , 32'hFFF596E9 , 32'hFFFC9EFB , 32'hFFFFBEA8 , 32'h000AEFDD , 32'h0000C678 , 32'hFFFD1F49 , 32'hFFF7CE14 , 32'h0000F599 , 32'hFFFDE5BA , 32'h000960C0 , 32'h0001030F , 32'hFFFEADD5 , 32'hFFF7F377 , 32'hFFFC1E8F , 32'hFFFE7EFF , 32'hFFFD2546 , 32'h0001B1EC , 32'hFFFFB4DF , 32'hFFFACCBA , 32'hFFFD7577 , 32'h0001576F , 32'hFFF425D7 , 32'h000861B1 , 32'hFFFF7CE7 , 32'h0003924B , 32'hFFFB79D0 , 32'h0000EB55 , 32'hFFFF5C83 , 32'hFFFE2711 , 32'h00032F2A , 32'h000850A7 , 32'h0002F080 , 32'hFFFE5E2D , 32'h0000D208 , 32'h0007804A , 32'h0003D5EE , 32'h0004F5E4 , 32'hFFFEA592 , 32'hFFFE40A2 , 32'hFFFE0A4F , 32'hFFFE0EBC} , 
{32'h49875500 , 32'h083CFD70 , 32'hD8466FC0 , 32'h8A7F8000 , 32'h141723A0 , 32'hD6BC1DC0 , 32'h98E5C480 , 32'hE9E7B100 , 32'hDF88D080 , 32'h060AA1B8 , 32'hF883D830 , 32'h2CBCA880 , 32'hDC2915C0 , 32'h0254742C , 32'h0A81D0F0 , 32'h154D3060 , 32'hD63898C0 , 32'hD57A2440 , 32'h112C2B20 , 32'h3BB5DF80 , 32'hF9D0C508 , 32'h241AB3C0 , 32'h0321C494 , 32'hF2D6ECC0 , 32'hF8C83A70 , 32'hEE022BC0 , 32'h0FA3D7A0 , 32'hFF45D7D3 , 32'hFAE27218 , 32'h045D5BF8 , 32'h125712A0 , 32'hF74D1DE0 , 32'h098FF940 , 32'h097C8A40 , 32'hFEE8B548 , 32'hFDD0159C , 32'h109EF1A0 , 32'hFD6F1114 , 32'h09325F10 , 32'hFB240E28 , 32'hF4A9E330 , 32'hFAE680B8 , 32'h27DBC740 , 32'hFF000A80 , 32'hFC296518 , 32'h192DAFA0 , 32'hE783C520 , 32'hFDBE9F64 , 32'hEC71EBA0 , 32'h15C9D380 , 32'h0A7A5C10 , 32'hE896F000 , 32'hFC9580E8 , 32'hF527E080 , 32'h1EB39000 , 32'h047386C0 , 32'h053F3778 , 32'hEA0344A0 , 32'hFE2E10B8 , 32'h0B021BC0 , 32'h017AAB88 , 32'h113CEC60 , 32'hFA702908 , 32'h09276310 , 32'h09104250 , 32'hFF013C47 , 32'hF5317E30 , 32'hEAAC5080 , 32'h082F2A20 , 32'hFBA0A2C8 , 32'h08F5C060 , 32'h02C8AACC , 32'h016A9E3C , 32'hFB091A20 , 32'hF90A5860 , 32'hFD26CDAC , 32'h07EBA9D8 , 32'h0309324C , 32'hFABF2FF0 , 32'hFD2F29A8 , 32'h02C7E520 , 32'h06E26090 , 32'hFC56B62C , 32'h01A86118 , 32'hFCA29140 , 32'h0190A810 , 32'h0213B030 , 32'hFD944AE4 , 32'h02D50910 , 32'hFFBBC248 , 32'h00022BE1 , 32'h00001C67 , 32'h0000F863 , 32'hFFFE9F3A , 32'hFFFCE4B4 , 32'h0001CC58 , 32'hFFFFB48E , 32'h0000E5A8 , 32'hFFFF2758 , 32'hFFFEE5E5} , 
{32'hC0E80780 , 32'h681B8500 , 32'hF6F85DB0 , 32'h7FFFFFFF , 32'h41C55000 , 32'hC8538400 , 32'h44D07600 , 32'h81403480 , 32'h0F2D4560 , 32'hA1067580 , 32'h018650C8 , 32'hDD485180 , 32'h3238B240 , 32'hD2273900 , 32'hE0BDB0A0 , 32'h0A6F5800 , 32'hF3BC3C10 , 32'h09B7D950 , 32'h32A4E200 , 32'hE9FD4C40 , 32'hE9B4DD80 , 32'h1C030EC0 , 32'h01E97358 , 32'hDEE7FF80 , 32'h26BA7740 , 32'hD86D4080 , 32'h00EEF842 , 32'h136380C0 , 32'hF8D673C0 , 32'h18C80040 , 32'h1E7400E0 , 32'hFA3EE0D8 , 32'hFDB68700 , 32'hE2FA4700 , 32'h030342F8 , 32'hFE4BB138 , 32'hEB534FE0 , 32'hFD315E74 , 32'h133B83C0 , 32'hFFF81CD6 , 32'hFD9374CC , 32'hF9288018 , 32'h18127CA0 , 32'hF8091E90 , 32'h048F37C8 , 32'hF0EF4670 , 32'hF8D0D7D8 , 32'hF3B73D70 , 32'hFCEA50AC , 32'hF463EF00 , 32'hFA50F7D0 , 32'hF594FD80 , 32'h0638AFC0 , 32'hFD37FE18 , 32'h0A371DE0 , 32'hEB1313A0 , 32'h01F8E1BC , 32'hF8AAC9C8 , 32'hF920EC80 , 32'h00A34548 , 32'h0D79D5B0 , 32'h033504C0 , 32'h002B0D7D , 32'hFDED8D68 , 32'h0076D31C , 32'h05698A10 , 32'h006D41FC , 32'h08032240 , 32'hFC40E754 , 32'h083789C0 , 32'h0219B6DC , 32'hFB615818 , 32'h06BCB9C8 , 32'hFD3E56AC , 32'h0385DED8 , 32'hF7DF7700 , 32'hFF8C5520 , 32'h041BB550 , 32'hFD0A98AC , 32'h02B69F08 , 32'h08BA9620 , 32'hFD318BCC , 32'hFA188050 , 32'hFD129DBC , 32'hFDD1E09C , 32'h01C6DE20 , 32'hFB208980 , 32'hFDE8D620 , 32'hFF6F3A09 , 32'h00B55D3E , 32'h0004ECD3 , 32'h0001CA1E , 32'hFFFCFA67 , 32'hFFFBE969 , 32'hFFFEC061 , 32'hFFFF54C9 , 32'hFFFE0EF8 , 32'hFFFEB79E , 32'hFFFB0D2C , 32'hFFFBE7B6} , 
{32'h52799080 , 32'h141CA080 , 32'h2029D540 , 32'hDE82DEC0 , 32'h326460C0 , 32'hE0327E60 , 32'hF4EE2500 , 32'hE6BA07C0 , 32'h078E2710 , 32'h04F14AE8 , 32'h2D9544C0 , 32'h52013A00 , 32'hF364FC10 , 32'h0F77AE70 , 32'hEFA2D9A0 , 32'h036DDC9C , 32'hEFF2CC40 , 32'hE6405BE0 , 32'h082DD450 , 32'h044A6858 , 32'h04DD1448 , 32'hF8FA2408 , 32'h09DE8760 , 32'h04D04320 , 32'h060CD308 , 32'h10EE0AC0 , 32'hE53DB600 , 32'hF6DF60F0 , 32'hF8FF5418 , 32'h11B8A1C0 , 32'h069FEDB0 , 32'hFF910D80 , 32'h0458B8E8 , 32'h19277040 , 32'hF80E1EF8 , 32'hE4ED38A0 , 32'hFC2B59D8 , 32'hF38D3CD0 , 32'h0ABB9B30 , 32'h0A9405E0 , 32'h08CD0060 , 32'h024CCE58 , 32'hFE07ADD0 , 32'h0CAB0FD0 , 32'hFCCA42E8 , 32'h0577ED30 , 32'h013EDC54 , 32'hFEFC6A28 , 32'h1595A6C0 , 32'h0CD226C0 , 32'hEE371CA0 , 32'h04707940 , 32'hFD861910 , 32'hF502C420 , 32'h008D6F5C , 32'hF10E6080 , 32'hE74E1D40 , 32'h15AD91C0 , 32'hE86AEA20 , 32'hEA5CC760 , 32'hFFD1FAAD , 32'h03D4F9CC , 32'h07B79730 , 32'h0616DA98 , 32'h0BCD9C70 , 32'h136AF280 , 32'h0AC1BF10 , 32'hF3F8F6B0 , 32'hF3A4EED0 , 32'h0ADE4150 , 32'hFEBD1AD0 , 32'hFF4C842E , 32'h12CBEF40 , 32'h0AF7FA20 , 32'h055B7AC8 , 32'hFEEB2C4C , 32'h06D34048 , 32'hF4B8BA50 , 32'h05DFB738 , 32'hF60EBE30 , 32'hF431B710 , 32'hF8AC5950 , 32'hFCFCD3E4 , 32'h0336C8D8 , 32'h04CE4B08 , 32'h000E4F95 , 32'h001405B8 , 32'h05AC9D58 , 32'h0023B854 , 32'hFFD2C7E5 , 32'hFFFDE505 , 32'h000697AC , 32'h00044DB8 , 32'h0001E194 , 32'hFFFFCF26 , 32'hFFFE76B6 , 32'hFFFEED5D , 32'h0000C050 , 32'h0000DACB , 32'hFFFDA92B}
};

logic signed [31:0] US_3 [100][10] ='{
{32'hEFD23C60 , 32'hBE4A8D00 , 32'hA4565E80 , 32'hEF8CC1A0 , 32'h64630800 , 32'h217EDB00 , 32'h0B1AA330 , 32'hE3898D00 , 32'h21C5DF00 , 32'hD6568AC0} , 
{32'h60C0C800 , 32'hC1ACA4C0 , 32'h297FDA40 , 32'hF49E9AA0 , 32'hB9EF0700 , 32'hF5CCB770 , 32'hFE49A470 , 32'h04106470 , 32'h2046FBC0 , 32'h02BF85A4} , 
{32'h2B24CF00 , 32'h00BA751D , 32'hC5E9D000 , 32'h4A910D80 , 32'h0196F3D4 , 32'hC48614C0 , 32'h66C48880 , 32'hDFF28200 , 32'h0C6FAE50 , 32'h01FB7934} , 
{32'h0002103F , 32'hFFFF2038 , 32'h00021300 , 32'h0006E369 , 32'h000780D7 , 32'hFFF73533 , 32'h00054E80 , 32'hFFFFCCD5 , 32'hFFFCF104 , 32'h00083741} , 
{32'hFFFA04CA , 32'h00080627 , 32'hFFFDAB59 , 32'hFFFF4EAF , 32'hFFFFC34F , 32'hFFFE757B , 32'hFFF96838 , 32'hFFFCEAE0 , 32'h000255C9 , 32'hFFFF0CC8} , 
{32'h035FA5C0 , 32'h69952E80 , 32'hA1D3C080 , 32'hF314D780 , 32'h223E3440 , 32'h28650F80 , 32'hC7A2B500 , 32'hE0E73480 , 32'hD97B1CC0 , 32'hEEAD7700} , 
{32'h4FB5EC00 , 32'h3591CC40 , 32'h1045A480 , 32'hF56341F0 , 32'h0A749820 , 32'h02C0814C , 32'hF8D7C3E8 , 32'h2FD0DA00 , 32'hF4B20470 , 32'hF1BA6DF0} , 
{32'hF8315D48 , 32'h558C2D00 , 32'h341850C0 , 32'hF8E5D2E8 , 32'h8EE1F300 , 32'h2BF2BB00 , 32'h1D9FB7A0 , 32'h31B75040 , 32'h1FA031A0 , 32'hD542B800} , 
{32'hFFFFC4FB , 32'h000B9D9A , 32'hFFFEBE76 , 32'hFFFB6DAD , 32'hFFFA6F3B , 32'h00018FFE , 32'hFFFA52A9 , 32'hFFFAF7A2 , 32'hFFFB4D6E , 32'h0007D29B} , 
{32'hFFE3C2B0 , 32'hE7776DA0 , 32'h7E6D2D00 , 32'h77E88880 , 32'hD8B42D00 , 32'h339A5E00 , 32'h092E8390 , 32'hF65132B0 , 32'h01851614 , 32'hD9BB4540} , 
{32'h165B4300 , 32'h2E681700 , 32'hBEBEF380 , 32'hC529BA40 , 32'h10968C20 , 32'h07AD4010 , 32'h1C0EF1C0 , 32'hB77EFD00 , 32'hF14B9B50 , 32'hFAE47A70} , 
{32'hC2BEF240 , 32'h5E60BD00 , 32'hBB46C000 , 32'hDDE51580 , 32'hE7511D40 , 32'hE0A305E0 , 32'h5EBDE100 , 32'h0F26C670 , 32'hEDC92C20 , 32'hF2D74D20} , 
{32'h029156D0 , 32'h911F8400 , 32'h4E005600 , 32'h712E1680 , 32'h53232480 , 32'hDE878C00 , 32'h4BE2D200 , 32'hE42296E0 , 32'hF14D6620 , 32'hE5FC42E0} , 
{32'h19E67A40 , 32'h3B383700 , 32'h45C52680 , 32'h05DB91A8 , 32'hCABEBCC0 , 32'hFB388B88 , 32'h0334AB44 , 32'hFB34EA68 , 32'hE5E59DA0 , 32'hCD235E40} , 
{32'hE38B2660 , 32'hABCB3F80 , 32'hD64BF500 , 32'hF1A4B5E0 , 32'h0902E940 , 32'hCBF6B4C0 , 32'hE2C19AC0 , 32'h22E61D40 , 32'h3FA7FD40 , 32'hD1A866C0} , 
{32'h096F2CB0 , 32'hDEC39400 , 32'h1D236E20 , 32'h8BE5FB00 , 32'hCE63FE80 , 32'h06D5A900 , 32'hDE093880 , 32'h4CBBD480 , 32'h15F2F540 , 32'hF1AC5FE0} , 
{32'h7FFFFFFF , 32'hF9CECD38 , 32'h0DDC6220 , 32'hD4B46240 , 32'hC9650B80 , 32'hF64F6FF0 , 32'h39928140 , 32'h38D22DC0 , 32'h08BCDC80 , 32'hE88F6D80} , 
{32'h42D10900 , 32'hF434BCD0 , 32'hD5A9C300 , 32'h45191100 , 32'hD889EF40 , 32'hC043D900 , 32'h17AFE880 , 32'h47C37900 , 32'hFEC82B88 , 32'hE08D6840} , 
{32'h59D7BA00 , 32'hC3AED700 , 32'hFCE81B00 , 32'hFAB3CD50 , 32'hE12C2CA0 , 32'hB74C1800 , 32'hAE972F80 , 32'h137A5F80 , 32'hD4D2E9C0 , 32'hD54365C0} , 
{32'h0000F019 , 32'h0002CE43 , 32'h0002FABE , 32'h000104E4 , 32'h000330C9 , 32'hFFFD5C55 , 32'h00029109 , 32'h0004CB0F , 32'h000028AB , 32'hFFFE22FD} , 
{32'h583E1480 , 32'h64034500 , 32'h48C46B00 , 32'h212DB000 , 32'h1AB00A40 , 32'hEE69ADA0 , 32'hF78C7B90 , 32'hA5035D00 , 32'h16652EA0 , 32'hC2AB98C0} , 
{32'hDC21E600 , 32'h145D6B60 , 32'h4B68FE00 , 32'hC373D1C0 , 32'hF893F478 , 32'h9C0EB800 , 32'hEBB4DF60 , 32'hECA881A0 , 32'h16302AE0 , 32'hE0FF0A00} , 
{32'h32EBF6C0 , 32'hA0C15A00 , 32'h18C9A300 , 32'hA2B7C080 , 32'hF28F6AC0 , 32'h2286DAC0 , 32'hFE43CB2C , 32'hFA1AD078 , 32'h02558C30 , 32'hFC04E1B8} , 
{32'h000376D6 , 32'h00011037 , 32'h000164DD , 32'h000277A3 , 32'hFFFD767F , 32'hFFF97BFB , 32'h0006CE03 , 32'h00017C35 , 32'h0005FD3D , 32'hFFFDA3B9} , 
{32'h7FFFFFFF , 32'h1DB2C5A0 , 32'hC32997C0 , 32'hF5E02420 , 32'h0AFFD330 , 32'h2BF35600 , 32'hEED84880 , 32'hF0E88620 , 32'h4381BD80 , 32'hDE8422C0} , 
{32'h34863EC0 , 32'h6F53D180 , 32'hF50A8CA0 , 32'h144C6160 , 32'h4255C400 , 32'h23EDE9C0 , 32'hF3F51020 , 32'hFECA9AF4 , 32'h087CB3B0 , 32'hF099DA30} , 
{32'h21B041C0 , 32'h28898DC0 , 32'hFC8D9E10 , 32'h07A198F8 , 32'h3DA6B700 , 32'hE0681140 , 32'h122136C0 , 32'h0F0BCC90 , 32'h348EAB80 , 32'hEBA7D680} , 
{32'h27302A00 , 32'h2023F0C0 , 32'h1B4393E0 , 32'hE7119D40 , 32'h01A0D618 , 32'hF2D26FC0 , 32'hDC550040 , 32'hE2DB2680 , 32'hD9478200 , 32'hF2C2F870} , 
{32'hF69FE160 , 32'hDE5CBF40 , 32'hE84AC920 , 32'hCCDB88C0 , 32'hF51F2A10 , 32'h24447240 , 32'hD79EA4C0 , 32'h403F4D80 , 32'hD017A400 , 32'h15E620E0} , 
{32'hC0E8B680 , 32'hE7E41960 , 32'h9B26C880 , 32'hF35D80F0 , 32'h1D8B5480 , 32'hFCE5479C , 32'h2BA7FC80 , 32'hB953DD80 , 32'hBCE44A80 , 32'hD56EE100} , 
{32'h7BBD8580 , 32'h303EEC40 , 32'h5B915880 , 32'hE6968C20 , 32'hEA33BE40 , 32'hE7F393A0 , 32'h3FFFC380 , 32'h143F1960 , 32'hA276CC00 , 32'hC4739700} , 
{32'h4C07B780 , 32'hA610DA80 , 32'h4C2DF380 , 32'hF4FC3FF0 , 32'hE8300440 , 32'h34DE46C0 , 32'h143E82E0 , 32'hD4FBDC00 , 32'hB5296F80 , 32'h010DC890} , 
{32'h7FFFFFFF , 32'h292DE480 , 32'h2AB27340 , 32'h2DAEAFC0 , 32'h1ED71040 , 32'hDAF61800 , 32'h358A8F80 , 32'h28A69B40 , 32'h20961F00 , 32'hE8F6B840} , 
{32'h915B6F00 , 32'hFDA5F9C0 , 32'h4E496880 , 32'hC2C73540 , 32'h4C560980 , 32'hAB5D3B00 , 32'h7296B100 , 32'h5337B880 , 32'h04821ED8 , 32'hEA104DA0} , 
{32'hFFFC0F51 , 32'h000301F1 , 32'h0006055E , 32'hFFF79637 , 32'h0006E45D , 32'hFFFFE2E8 , 32'hFFFD4B7D , 32'hFFF7ED8E , 32'h0006DA08 , 32'h0002D1CF} , 
{32'hF86B2E10 , 32'hB0223E00 , 32'hE7348900 , 32'h1D25E4C0 , 32'h319E4A40 , 32'h9AE21A80 , 32'h024FF088 , 32'hFFA54132 , 32'hF576A360 , 32'hF01BD340} , 
{32'hEABC0860 , 32'hE5CA9D20 , 32'hBA0B4580 , 32'h0F445FA0 , 32'h2C63A680 , 32'h1A938820 , 32'h2A6D9A80 , 32'hE3D2F520 , 32'h0796AB60 , 32'hFF4618A2} , 
{32'h041491E8 , 32'hABEE4600 , 32'h65A98180 , 32'hA93DA880 , 32'hF05E5A30 , 32'h45262D80 , 32'hF1DDC200 , 32'hE7358480 , 32'h16B55180 , 32'hE8D84360} , 
{32'h374F80C0 , 32'hC0F8C600 , 32'h0D672E50 , 32'hBD0C2A00 , 32'h1F5199C0 , 32'hF4D4F2B0 , 32'hD22EBD40 , 32'h10B8CC60 , 32'h3DD6F380 , 32'hEB9A5D80} , 
{32'h41727800 , 32'hB96D6200 , 32'hFCF4A550 , 32'hC7E7B140 , 32'h1F214FA0 , 32'h4242F380 , 32'hF6953C00 , 32'h1BAC9420 , 32'hDAA397C0 , 32'hF55CCD80} , 
{32'hC67DEC40 , 32'h3022D880 , 32'h5CC5AC00 , 32'h049ACD80 , 32'hCE48C980 , 32'h25201540 , 32'h18E0C8E0 , 32'hA9A93780 , 32'h340DA200 , 32'hF43FF760} , 
{32'h019AEBD0 , 32'hFCFBAEF0 , 32'hF8DB01F8 , 32'h074D20D8 , 32'h00B9761A , 32'hF8B77918 , 32'hFF7DD676 , 32'h03813060 , 32'hF675E560 , 32'hF9E79008} , 
{32'hF6B36E60 , 32'h15006400 , 32'h0D8AD760 , 32'h1D21B300 , 32'hFA315E08 , 32'h07555C30 , 32'hF3A44530 , 32'h10EE6B00 , 32'hD6310740 , 32'h02681440} , 
{32'hD5AB5E40 , 32'hE54F14E0 , 32'h50C8CF80 , 32'hEF33E0E0 , 32'h52F20280 , 32'hCCD3DC40 , 32'hD85A04C0 , 32'hE142B400 , 32'h20F2A880 , 32'hE7069500} , 
{32'hF3924860 , 32'h1074EDA0 , 32'h7FFFFFFF , 32'hF98FE948 , 32'h98223300 , 32'hF0A39F00 , 32'h01AEFC70 , 32'h2F50A140 , 32'h3A91F8C0 , 32'hEEDB8C40} , 
{32'hDD17B9C0 , 32'h20877DC0 , 32'hACEE3800 , 32'hD480ED40 , 32'hCC286400 , 32'h2A1B4C40 , 32'h509BDB80 , 32'h010E78BC , 32'h1BB1BDA0 , 32'h0095FE93} , 
{32'h04A027E0 , 32'h7FFFFFFF , 32'hF7320630 , 32'h13E47420 , 32'h255F23C0 , 32'hF2F85650 , 32'h35339740 , 32'hE7A37640 , 32'hB08A2600 , 32'hEA1D2940} , 
{32'h4CD1D280 , 32'hF1332760 , 32'hE60838E0 , 32'h669D3280 , 32'hCBDEAE80 , 32'hD9D07EC0 , 32'hE0120EC0 , 32'h16FCA460 , 32'hC6B96180 , 32'hE6CA4CA0} , 
{32'hF706ABC0 , 32'h7FFFFFFF , 32'h0B3CCDF0 , 32'hEAF27CA0 , 32'h14A83F00 , 32'h27DB0F40 , 32'h3F09C640 , 32'h415D0A80 , 32'hF32EBC70 , 32'hE558FDA0} , 
{32'hB09AE580 , 32'h552C5880 , 32'hEDF0E8E0 , 32'hC8DE8100 , 32'hB87FA880 , 32'h16C01860 , 32'h2768F1C0 , 32'hAF73E780 , 32'h24B39A80 , 32'hEB436740} , 
{32'hFC33ECD4 , 32'h34371900 , 32'h2BE748C0 , 32'h05B7C990 , 32'h74C77680 , 32'hF3D12810 , 32'hF3E9A860 , 32'hB1ED5A80 , 32'h1373BBA0 , 32'hDB812BC0} , 
{32'hF00DF5B0 , 32'hD965A700 , 32'hCC040B80 , 32'hE1EEDA20 , 32'h584CA000 , 32'h51626800 , 32'h5666F200 , 32'hF3F0F9A0 , 32'h317165C0 , 32'hED4083E0} , 
{32'h47E2C580 , 32'hC69AAE00 , 32'hC9B9D080 , 32'h7303A280 , 32'hBCB4ED80 , 32'h00546B60 , 32'h1DAB5340 , 32'h1C0DD9E0 , 32'h2342CFC0 , 32'hFA600CF8} , 
{32'hC9BE9200 , 32'h12D2C700 , 32'h01151910 , 32'h395788C0 , 32'hFE2A3AD4 , 32'h2E07AFC0 , 32'hE98A1520 , 32'h4E116580 , 32'hCD229980 , 32'hFADA3660} , 
{32'hEC635620 , 32'h0D433CF0 , 32'h092458F0 , 32'hE6D5CEC0 , 32'h3DB97B00 , 32'hCEA33840 , 32'hCE2664C0 , 32'h362DCBC0 , 32'hF5E23620 , 32'hF438B710} , 
{32'hE1B19120 , 32'h1685EFC0 , 32'hC8B89FC0 , 32'hF1B87450 , 32'hF994B828 , 32'h0BA2DB80 , 32'hB0D97C80 , 32'hF5DF0B40 , 32'h0A8BAD20 , 32'hF7B2B460} , 
{32'hB8855E80 , 32'hE54D7340 , 32'hACD3C780 , 32'hAE929A00 , 32'hE2FCF4E0 , 32'hB6A2BC00 , 32'hA92C7800 , 32'hF42F1E50 , 32'hDA87C6C0 , 32'hC905B440} , 
{32'h1C6DD180 , 32'h03B14FE4 , 32'h90A69180 , 32'h55A79F00 , 32'hA5846080 , 32'h07800828 , 32'hF78C4990 , 32'h09FD4910 , 32'hF4FE92A0 , 32'hEB075F60} , 
{32'hC96561C0 , 32'h24971C40 , 32'h37002D00 , 32'h3BA69300 , 32'hC5DE0400 , 32'h1167B600 , 32'h045FCF78 , 32'hF0C7B0F0 , 32'h12D5E3C0 , 32'hEC8A4420} , 
{32'hA6F9B280 , 32'h4B5AFD80 , 32'hCF00D800 , 32'hFEA009B8 , 32'hBDF46500 , 32'hB6AC1F80 , 32'h278D22C0 , 32'hDBC0BDC0 , 32'hC7062BC0 , 32'hE05BA9C0} , 
{32'hEA5C2D20 , 32'h91DF0300 , 32'h952FE200 , 32'hD03CBD40 , 32'h18A18A40 , 32'h19ACCCA0 , 32'hF9E8AEC8 , 32'h30AFDA80 , 32'hF6C5C9E0 , 32'hED60B020} , 
{32'h071F22C8 , 32'hE87B11A0 , 32'hDA3CB980 , 32'h0385BB80 , 32'h4F077600 , 32'h31C1C940 , 32'hEBDB1820 , 32'hCA089D00 , 32'hECB9FD60 , 32'h06968DC8} , 
{32'hF7DBCD20 , 32'hF740F110 , 32'hFF98E0F4 , 32'hAF90A380 , 32'h058E8990 , 32'hF72D8D00 , 32'h7FFFFFFF , 32'h0E26B360 , 32'h0AC92D30 , 32'hEAD5FA80} , 
{32'hCEB7B640 , 32'hDB4279C0 , 32'hD441F880 , 32'hDCA311C0 , 32'h106E5000 , 32'hEACA6360 , 32'h087CC500 , 32'hE4726440 , 32'hFA1154F0 , 32'hEE37D0E0} , 
{32'h3F4F2800 , 32'hE6DA6840 , 32'hB1470B00 , 32'h00B72533 , 32'h10D9CA40 , 32'h492FDA80 , 32'hDF99F600 , 32'hE9A2A600 , 32'h121AAE60 , 32'hEF689F80} , 
{32'hA4AD0080 , 32'hBACB4C80 , 32'h07958510 , 32'h00E5B147 , 32'h9D785E80 , 32'h4A8E5B00 , 32'hEFE96540 , 32'hEACA7200 , 32'hF1BBDE50 , 32'hD93E9680} , 
{32'hFFFC4E97 , 32'hFFFC5756 , 32'h0004755F , 32'h0000775C , 32'hFFF9FD84 , 32'h0002F897 , 32'hFFFA9312 , 32'hFFFC857D , 32'h0005E465 , 32'hFFF75254} , 
{32'h2F9B73C0 , 32'hF90EBCC8 , 32'hE38E5F80 , 32'h3AD70180 , 32'h13EF0660 , 32'hE25271C0 , 32'h2ACAFA00 , 32'h0F99E9C0 , 32'hC5CFF400 , 32'hDCF7F9C0} , 
{32'h0397E144 , 32'hE36E00E0 , 32'h09B377E0 , 32'hE5330DE0 , 32'hE6521200 , 32'h1318AEE0 , 32'h2E786A40 , 32'hF42399C0 , 32'hEE86AE60 , 32'hF6007CC0} , 
{32'h0D4AE880 , 32'hD151FCC0 , 32'hB10B1E00 , 32'h382B3880 , 32'h04C3F338 , 32'h277D0580 , 32'h234BE000 , 32'h1B51CE80 , 32'hF37EDE50 , 32'hE3B5C180} , 
{32'hDF6F5080 , 32'hFF9EE128 , 32'h26A50340 , 32'h0A65C340 , 32'h3ADA0BC0 , 32'h252C2E00 , 32'h054F4AD0 , 32'h4A0C0600 , 32'h00BBF486 , 32'hE1FA5380} , 
{32'h0F341AE0 , 32'h19E27E80 , 32'hEFAF16A0 , 32'h4E4CBA80 , 32'hE3EBBAE0 , 32'h121BFE40 , 32'h1E686240 , 32'h28175DC0 , 32'h142E9780 , 32'hEE6710C0} , 
{32'h1221C900 , 32'h48CDF900 , 32'h03F89004 , 32'hFA794C30 , 32'h47664880 , 32'h4A2CE800 , 32'hE71258C0 , 32'hED001840 , 32'hE9571E60 , 32'hE07AB9C0} , 
{32'h0940D030 , 32'hE87D5640 , 32'h071BB1D0 , 32'hCF997E00 , 32'hE9ACDEC0 , 32'hC0CF58C0 , 32'h17716BA0 , 32'hE2591960 , 32'hF30BC6F0 , 32'hFABC8640} , 
{32'h2065DCC0 , 32'hFE6EDEB0 , 32'h07500AE0 , 32'h3DE61600 , 32'h16BA71E0 , 32'h34E42980 , 32'h31F1D900 , 32'h4F320F80 , 32'h284FE740 , 32'hD205A0C0} , 
{32'h18F26CC0 , 32'hF2E8DBC0 , 32'h502B8900 , 32'hD6952CC0 , 32'h1122DAE0 , 32'hDE9E3F40 , 32'hDBDDE8C0 , 32'h11E17020 , 32'hE6FDF380 , 32'hF8E48030} , 
{32'hCCFE8940 , 32'h2D4020C0 , 32'h5615D380 , 32'h0A9085C0 , 32'h0513B4B8 , 32'h1DAEB020 , 32'h1528DB80 , 32'hFD96F530 , 32'h0B48B2D0 , 32'hFF4695F8} , 
{32'h3067C0C0 , 32'h50623480 , 32'hCD8A2780 , 32'h35CF2740 , 32'h206113C0 , 32'h49ACF000 , 32'hB0414C00 , 32'h068B2FD8 , 32'h0DADF880 , 32'hCD9E0100} , 
{32'h7FFFFFFF , 32'hBFF23D80 , 32'hEF1E9700 , 32'hECF61100 , 32'hD2CB8BC0 , 32'hF5D1E560 , 32'hC9667DC0 , 32'hE21813E0 , 32'h0D6CCEC0 , 32'hB92EB600} , 
{32'h426AB580 , 32'hB247A680 , 32'h5B861F80 , 32'h147BEEC0 , 32'hF6216C70 , 32'hEEF039C0 , 32'h0BE79650 , 32'hBBEE0E00 , 32'h46FD8A80 , 32'hF1F50D10} , 
{32'h98124E00 , 32'h033673C0 , 32'h1C113C80 , 32'h49365300 , 32'hE7E94A80 , 32'h136E80A0 , 32'hB6FC3200 , 32'hF83A15D8 , 32'h0E3C3A10 , 32'hD70FED80} , 
{32'hFFB3EEB3 , 32'h40E6AE00 , 32'h18E1B2A0 , 32'h7FFFFFFF , 32'hB4A2D100 , 32'hD08426C0 , 32'hEC8693E0 , 32'hB3A7C780 , 32'h18DB0BC0 , 32'h08BCF070} , 
{32'hE26196E0 , 32'h32830240 , 32'h4AB9E100 , 32'hC3B19C80 , 32'hDFACAAC0 , 32'h32DB4200 , 32'hD3EC5C00 , 32'h0AFBF8E0 , 32'hF94BC718 , 32'hE110B600} , 
{32'hFFFE0E9D , 32'h0006A5E7 , 32'hFFFE5C94 , 32'hFFFCAF7E , 32'h0005213C , 32'hFFFE4D92 , 32'hFFFB7A9A , 32'hFFFB414D , 32'h00020925 , 32'h00077D07} , 
{32'h0AFC45C0 , 32'h6931CA00 , 32'h038EB2C4 , 32'h07FE1050 , 32'h488E6C00 , 32'h40DB7900 , 32'h055A92A0 , 32'h161DDF20 , 32'hCFDC0300 , 32'hFB5DB778} , 
{32'hC1F52C80 , 32'h1DEA6F40 , 32'h4D8EBB00 , 32'h0083C7ED , 32'h3D905180 , 32'h1CD52160 , 32'hDD80B200 , 32'h6C8B2780 , 32'h202B43C0 , 32'hE3117A80} , 
{32'h50B27080 , 32'h2037D580 , 32'hBBA18D00 , 32'h02FD5098 , 32'h42A41580 , 32'hFE70F188 , 32'h09902E20 , 32'h1B4F8920 , 32'h679F5980 , 32'hE1359F80} , 
{32'h7FFFFFFF , 32'hFC369358 , 32'hF266EA70 , 32'h92ECF480 , 32'hD9E06AC0 , 32'h33A76740 , 32'h4C822580 , 32'hA854C080 , 32'hFF803CD0 , 32'hF2C5D800} , 
{32'hC1765240 , 32'h03613C40 , 32'hD58A5800 , 32'hA5390180 , 32'hA4DB7180 , 32'hED50F220 , 32'h1CC65760 , 32'hF82BA478 , 32'hFFFAB0EE , 32'hDC950580} , 
{32'h000079EE , 32'h0001E8A1 , 32'h0001B78C , 32'h0004D352 , 32'h00014300 , 32'h000153BF , 32'h0002F3CF , 32'h000942A0 , 32'h000081A6 , 32'h00015E78} , 
{32'h489EA280 , 32'h07000118 , 32'h123BCEE0 , 32'hE1236440 , 32'h2CCF2000 , 32'h94E14600 , 32'hE30C55C0 , 32'hFB63BC58 , 32'h10C0CF80 , 32'hF3E25610} , 
{32'hFBE425E0 , 32'h1CEB1280 , 32'h151A53A0 , 32'h01BC89C8 , 32'h0CE29150 , 32'h01B60B40 , 32'h06692F90 , 32'h26436E00 , 32'h18E95440 , 32'h0EB55E70} , 
{32'h21938E80 , 32'h5B2F0D80 , 32'h0BFB8340 , 32'h06867F50 , 32'h04BF6F48 , 32'h1A748840 , 32'hFB547210 , 32'hEA935E60 , 32'hB7F33100 , 32'hFC52D7FC} , 
{32'h61AFD680 , 32'h4A6DA800 , 32'h00DECB2C , 32'hB0BCE700 , 32'hF063AA10 , 32'hAA7DD980 , 32'hEB65D520 , 32'hEB19BC40 , 32'h11FCD980 , 32'hD897BBC0} , 
{32'hFFFC720B , 32'hFFF8AD5C , 32'h00011B72 , 32'hFFFAC9AC , 32'h00046B4A , 32'h00038095 , 32'h00055B8A , 32'hFFFA03FC , 32'h000585C0 , 32'hFFF65EEB} , 
{32'hF854CFF0 , 32'hADE45000 , 32'hCC5A1280 , 32'h52A0CD00 , 32'h24D280C0 , 32'hD30E75C0 , 32'hED4F46C0 , 32'hE40FF8C0 , 32'hF6A4B9F0 , 32'hBE6D7180} , 
{32'hBFDDC500 , 32'h96542280 , 32'h0D59B690 , 32'h359688C0 , 32'hE4101740 , 32'h2A52A400 , 32'h006CAF88 , 32'hD6325CC0 , 32'h64BDB700 , 32'h0887C6B0} , 
{32'hEBB924A0 , 32'h7FFFFFFF , 32'h46F94C80 , 32'hFC8ED744 , 32'hD28D6BC0 , 32'h6F74E780 , 32'h0E2ECF50 , 32'h10EE3900 , 32'hD4713280 , 32'hC52F2100} , 
{32'hD5ACD140 , 32'h3C796880 , 32'hCF91D000 , 32'hDD5FB5C0 , 32'hF0E7FB80 , 32'h06E21F30 , 32'hDA783240 , 32'h0FF79900 , 32'h1E6C6820 , 32'hD6F57780} , 
{32'h6DF49980 , 32'hE773FD00 , 32'h16F71260 , 32'hEE78A5A0 , 32'hC0CA0480 , 32'hD56AFF00 , 32'hFF0084D3 , 32'h281C0640 , 32'h33BF58C0 , 32'h1C572F60}
};
logic signed [31:0] bias_0[37] = '{32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000 , 32'h00000000};
logic signed [31:0] bias_1[300] = '{32'hDD9F58C0 , 32'h0EEA81D0 , 32'hFAFB1C50 , 32'h2B412D00 , 32'hF1A4E860 , 32'hF982BBA8 , 32'hFDFC118C , 32'hF5D3AE00 , 32'hFA029140 , 32'hEE426660 , 32'hEA1B6AA0 , 32'h0E8487F0 , 32'h2561F9C0 , 32'hFE169E8C , 32'hEF38FEE0 , 32'h01F22654 , 32'hFDC36034 , 32'h06E20628 , 32'hD4A3EB80 , 32'hFECAD3B0 , 32'hFDEE950C , 32'hF52267E0 , 32'h2B608440 , 32'h073D0A70 , 32'h18B48D80 , 32'hFEB2F7F0 , 32'hFBC6C508 , 32'h02C39A08 , 32'hFE90E88C , 32'h3510FB40 , 32'hFD5EF710 , 32'h0CC2C810 , 32'hE58AED60 , 32'hF6DA5E60 , 32'hFEE76A10 , 32'h0368F5E0 , 32'h19363F00 , 32'hE4317A80 , 32'hF65CC1D0 , 32'h00B27F8E , 32'hE7A25C40 , 32'hF6F1F670 , 32'hFDDF1AE8 , 32'h05E0B128 , 32'h28D5C5C0 , 32'h2E90B2C0 , 32'hFF87CCA0 , 32'hFEF17DBC , 32'h0B14C910 , 32'hF7319A00 , 32'hFA0A72B8 , 32'hFC4FE16C , 32'hF351B280 , 32'h1454C2E0 , 32'hF7C20DC0 , 32'hFF16935A , 32'hFBE0DAB0 , 32'hFA4372A0 , 32'hFED441EC , 32'hBF388D80 , 32'hFBE1B2C8 , 32'hFCC043AC , 32'hFA2C3150 , 32'hFE794F40 , 32'h1443A360 , 32'hFA87C040 , 32'hF21B2710 , 32'h0370A80C , 32'hFDF5ED08 , 32'hD9863980 , 32'hF563EB30 , 32'hE034E4C0 , 32'hFCA16AA4 , 32'hFEB68834 , 32'hFDB00BE8 , 32'hD5496B80 , 32'hF3ED0D90 , 32'hFE2D59C0 , 32'h176D7D20 , 32'hEC8AEE00 , 32'hF3277240 , 32'h20201040 , 32'hF6CC5A20 , 32'hFBA8FE98 , 32'hD4AEF640 , 32'h1704C740 , 32'hCCB08940 , 32'hEDB300A0 , 32'hE8319300 , 32'hDE387E80 , 32'hFE362084 , 32'h1EF1F600 , 32'hFD35420C , 32'hDA703200 , 32'hEAC79C20 , 32'hFDFAABAC , 32'hFEA9DDE4 , 32'hFCE0B638 , 32'hF4BA7800 , 32'h09DDD560 , 32'h235A0600 , 32'hFDAB46BC , 32'hD2A51A40 , 32'h089CEA20 , 32'h356CBF40 , 32'hFE29BCA8 , 32'hE0C14060 , 32'hFE7849CC , 32'h13276740 , 32'h2E660840 , 32'hFBD93F38 , 32'h35964500 , 32'hF23810C0 , 32'hF8C45360 , 32'hD528DE80 , 32'h0DD4DE20 , 32'hDBF025C0 , 32'hFEB9CA58 , 32'h0A46D4F0 , 32'hFC4FF2E0 , 32'hECC99100 , 32'hF9402528 , 32'hEAA12D80 , 32'hEEC9F7A0 , 32'h1132B6E0 , 32'hF8DA7008 , 32'hFC5F7564 , 32'hFDAA67F8 , 32'hFEDAF234 , 32'hFB5426C8 , 32'hFC729C64 , 32'hFCA82D84 , 32'h0CB091B0 , 32'hF89F4230 , 32'hFC9A8374 , 32'h306AB140 , 32'h0F5EFD30 , 32'hFE3822C0 , 32'hFE382744 , 32'hE9B4A420 , 32'hF661A910 , 32'hFDDA94C4 , 32'hFA976E68 , 32'h1BED7C00 , 32'h20D86200 , 32'hF2ED8010 , 32'hEF0F73A0 , 32'hFEE8EDCC , 32'hEBC91360 , 32'hF889FD10 , 32'hF5ECBD30 , 32'hE652E660 , 32'hFEA6B848 , 32'hF7005EE0 , 32'hF1FE25E0 , 32'hFD650E34 , 32'h0A73BF10 , 32'hCC7D9600 , 32'hEDB35040 , 32'hF914DDF0 , 32'hFDA24124 , 32'hD0858080 , 32'hF89FBF90 , 32'h0EF39E50 , 32'h11005F40 , 32'hFDD362F8 , 32'h14DECB80 , 32'hF9E64CC0 , 32'hFB2407A0 , 32'hF0D23030 , 32'hE5487980 , 32'hF3242E40 , 32'hFE8092C0 , 32'hF5815D40 , 32'hEA7099A0 , 32'hE6A6B060 , 32'h1C681740 , 32'hEC53DD40 , 32'h07894258 , 32'hEE75B920 , 32'hE5184120 , 32'hFD643750 , 32'hF8EF6068 , 32'hFE492C20 , 32'hF2E73590 , 32'h1E7A8400 , 32'hE9DA14A0 , 32'hF8697590 , 32'h31ABEEC0 , 32'h17488CC0 , 32'hFDE9EEA8 , 32'hE640C940 , 32'h13983800 , 32'hF5CE0B90 , 32'hF9D7A978 , 32'hFE867998 , 32'hE488F040 , 32'hE731ADE0 , 32'hE3C20040 , 32'hFC7475A0 , 32'hFB177480 , 32'hFEE23A30 , 32'hFE45CD14 , 32'hFE16C110 , 32'hF1E40B40 , 32'hED9740C0 , 32'h067E0148 , 32'hFFD577F4 , 32'hEC82F1C0 , 32'h040919B8 , 32'hFEFB00F8 , 32'hFE41A068 , 32'hFEC1BC90 , 32'hF74BCBC0 , 32'hFCFF8E18 , 32'hE9CE41A0 , 32'h03909120 , 32'h100FEA80 , 32'hFD433B50 , 32'hFEBE73E8 , 32'hFC6872F0 , 32'hFCA53870 , 32'h0B818C10 , 32'hF2BD2470 , 32'hFBE86E88 , 32'hFB401818 , 32'hFCBDBB20 , 32'hEFAC0EE0 , 32'h13D640A0 , 32'hEBF8A2C0 , 32'hFE875344 , 32'hFF09DA66 , 32'hFF0130B5 , 32'hDEE68400 , 32'h0A714680 , 32'hFE84F434 , 32'hFE639D50 , 32'hF305E210 , 32'hFDC3A484 , 32'hCA6D7240 , 32'hFD412440 , 32'h2C3DEB40 , 32'hFE2DD230 , 32'hFFC680B8 , 32'hF0DA3B80 , 32'hEDCDA300 , 32'h30662E80 , 32'hF7BE1810 , 32'hECEA6A60 , 32'hE196B440 , 32'hFE92B234 , 32'h34A07140 , 32'hF3A91090 , 32'h01C4EB00 , 32'h0CE88CC0 , 32'h1F339880 , 32'hEFD822A0 , 32'hFC6AF148 , 32'hF8FFF070 , 32'hF2BE2010 , 32'h15E9DF20 , 32'hE6EB6DE0 , 32'hDB73F980 , 32'hFCC8EE5C , 32'hFCD409F4 , 32'hFE8A419C , 32'hF4ED09A0 , 32'hF922AAA0 , 32'hDD52CB00 , 32'h0BA2CDD0 , 32'hFCEFB5F0 , 32'hFD3E6554 , 32'hFF1BACB2 , 32'hED937E00 , 32'h24456980 , 32'h019A361C , 32'hFC06F8F8 , 32'h007C9AE5 , 32'hCDF48300 , 32'hFCE9AF04 , 32'hFDC6CFFC , 32'hF0AFC570 , 32'hFB3842D8 , 32'hF6814650 , 32'hFC1866DC , 32'hEC296120 , 32'hC2E3C380 , 32'hF5E23630 , 32'h07D5E568 , 32'hDA6446C0 , 32'hD66A0900 , 32'hFDB0F744 , 32'hFE620124 , 32'hF36BAC10 , 32'h1960DC40 , 32'hE1F05660 , 32'hF48F8E70 , 32'h0A63E5C0 , 32'hF6AA2B60 , 32'hFA6F8808};
logic signed [31:0] bias_2[100] = '{32'h0852FB80 , 32'hFCC8B83C , 32'h05100CD8 , 32'hFF025B44 , 32'hD775C1C0 , 32'h59B8DC80 , 32'h21F4D480 , 32'h2FFE1100 , 32'hFD05A24C , 32'hDA311880 , 32'h1AD43FE0 , 32'h06A8AB18 , 32'hCC0D0580 , 32'h430CB480 , 32'h08076840 , 32'h1BABB640 , 32'h04EF9BD8 , 32'h27E4FA40 , 32'h2884C280 , 32'hFC1D58EC , 32'h07777308 , 32'h2CDE2580 , 32'hE6451300 , 32'hFC6D7494 , 32'hF8705D70 , 32'h1D52C8C0 , 32'h02C99358 , 32'h32816D40 , 32'h11DF0200 , 32'h18252E80 , 32'hF6A13960 , 32'hEA7B20C0 , 32'hE210C600 , 32'h00F3628D , 32'hFF018954 , 32'hE00C7420 , 32'hDC9C4000 , 32'hC8F33900 , 32'hE932B6C0 , 32'hE3C2D880 , 32'hFC3B5CC8 , 32'hCF42EF80 , 32'h2A455440 , 32'hECF6BAE0 , 32'h4CF27D00 , 32'h0F209D40 , 32'hDAC05680 , 32'h30E2D700 , 32'h25587A00 , 32'h2E000FC0 , 32'hFAEF63F8 , 32'hF02C02B0 , 32'h0859DF40 , 32'h34565F00 , 32'h18A8D2E0 , 32'h519B0D00 , 32'h43B5A180 , 32'h4CCC3780 , 32'h1673A880 , 32'h49FE5E00 , 32'hEE67EB20 , 32'hF45367C0 , 32'hCD403480 , 32'h04DACFA0 , 32'h115B6F40 , 32'h0318C5AC , 32'hEA2B4620 , 32'h02670394 , 32'hEB6FF080 , 32'h02BAA6F4 , 32'hD422B5C0 , 32'h0D8386F0 , 32'hFBAD7EC0 , 32'h09209F60 , 32'hE27A5D00 , 32'h063E66C0 , 32'hEAF0EAE0 , 32'h0B74A8F0 , 32'h0D4A91F0 , 32'hF83EDE30 , 32'h3AC30C40 , 32'h19414680 , 32'h2F07D240 , 32'hF8564DE8 , 32'h11FD4480 , 32'h19C3BE00 , 32'hF1ABC070 , 32'h023EA840 , 32'h08CCB140 , 32'hFB606560 , 32'h2CCCCC80 , 32'hFE7F04C0 , 32'h3562FD40 , 32'h434CC680 , 32'hFD6FA1F8 , 32'hFA120B50 , 32'h10405B40 , 32'hE260DC80 , 32'h3E9EA2C0 , 32'h2671FB40};
logic signed [31:0] bias_3[10] = '{32'hF9F86C40 , 32'hD9CE1BC0 , 32'hFA273BF0 , 32'hFF377075 , 32'h06B7FB80 , 32'hE0A5AD60 , 32'h045D06E8 , 32'hD44CAC80 , 32'h52426B00 , 32'h0AF82900};


endpackage
